module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 ;
  assign n256 = ( ~x20 & x151 ) | ( ~x20 & x229 ) | ( x151 & x229 ) ;
  assign n257 = x236 ^ x106 ^ x21 ;
  assign n258 = ( x31 & x219 ) | ( x31 & ~x234 ) | ( x219 & ~x234 ) ;
  assign n259 = x236 ^ x224 ^ 1'b0 ;
  assign n260 = x238 & n259 ;
  assign n261 = ( x67 & x155 ) | ( x67 & ~x196 ) | ( x155 & ~x196 ) ;
  assign n262 = ( ~x234 & x239 ) | ( ~x234 & x247 ) | ( x239 & x247 ) ;
  assign n263 = x103 ^ x94 ^ 1'b0 ;
  assign n264 = x179 & n263 ;
  assign n265 = ( x63 & x126 ) | ( x63 & ~x227 ) | ( x126 & ~x227 ) ;
  assign n266 = ( x60 & ~x207 ) | ( x60 & x233 ) | ( ~x207 & x233 ) ;
  assign n270 = x230 ^ x179 ^ x173 ;
  assign n267 = x194 ^ x149 ^ x65 ;
  assign n268 = n267 ^ n257 ^ x192 ;
  assign n269 = x156 & ~n268 ;
  assign n271 = n270 ^ n269 ^ 1'b0 ;
  assign n272 = x136 & x199 ;
  assign n273 = ~x206 & n272 ;
  assign n274 = x76 & x153 ;
  assign n275 = n274 ^ x31 ^ 1'b0 ;
  assign n276 = ( x79 & ~x251 ) | ( x79 & n275 ) | ( ~x251 & n275 ) ;
  assign n277 = x213 ^ x187 ^ x76 ;
  assign n278 = x218 & ~n277 ;
  assign n279 = n278 ^ x178 ^ 1'b0 ;
  assign n280 = x252 ^ x158 ^ x138 ;
  assign n281 = n279 | n280 ;
  assign n282 = x11 | n281 ;
  assign n283 = n258 ^ x82 ^ x54 ;
  assign n284 = x196 & x201 ;
  assign n285 = n283 & n284 ;
  assign n286 = x227 ^ x183 ^ x20 ;
  assign n287 = x115 & x166 ;
  assign n288 = n287 ^ x68 ^ 1'b0 ;
  assign n289 = x250 & n288 ;
  assign n290 = n266 ^ x143 ^ x21 ;
  assign n291 = ( ~x24 & x139 ) | ( ~x24 & n287 ) | ( x139 & n287 ) ;
  assign n292 = x46 & x64 ;
  assign n293 = n292 ^ x110 ^ 1'b0 ;
  assign n294 = x189 & ~n293 ;
  assign n295 = ~x112 & n294 ;
  assign n296 = n295 ^ n279 ^ x28 ;
  assign n297 = x34 ^ x1 ^ 1'b0 ;
  assign n298 = ( x229 & n262 ) | ( x229 & n268 ) | ( n262 & n268 ) ;
  assign n299 = x99 & ~n268 ;
  assign n300 = ~x53 & n299 ;
  assign n301 = ( x0 & ~x21 ) | ( x0 & x57 ) | ( ~x21 & x57 ) ;
  assign n302 = x44 & ~n276 ;
  assign n303 = ~x141 & n302 ;
  assign n304 = n262 ^ x117 ^ x112 ;
  assign n305 = ( x131 & ~x152 ) | ( x131 & n304 ) | ( ~x152 & n304 ) ;
  assign n306 = n305 ^ x89 ^ x36 ;
  assign n307 = ( ~x58 & x70 ) | ( ~x58 & x164 ) | ( x70 & x164 ) ;
  assign n308 = ( ~x249 & n276 ) | ( ~x249 & n307 ) | ( n276 & n307 ) ;
  assign n309 = ( ~x165 & n306 ) | ( ~x165 & n308 ) | ( n306 & n308 ) ;
  assign n310 = n273 ^ x173 ^ x82 ;
  assign n311 = n310 ^ x242 ^ x195 ;
  assign n312 = x37 & ~n311 ;
  assign n313 = n261 ^ x159 ^ 1'b0 ;
  assign n314 = n313 ^ x231 ^ x193 ;
  assign n315 = ( x169 & ~x184 ) | ( x169 & n303 ) | ( ~x184 & n303 ) ;
  assign n316 = x114 & x173 ;
  assign n317 = ~x196 & n316 ;
  assign n318 = n317 ^ x209 ^ x128 ;
  assign n319 = x97 ^ x74 ^ 1'b0 ;
  assign n320 = x64 & n319 ;
  assign n321 = x179 & x219 ;
  assign n322 = ~n320 & n321 ;
  assign n323 = n322 ^ x253 ^ x69 ;
  assign n324 = ( ~x226 & n282 ) | ( ~x226 & n323 ) | ( n282 & n323 ) ;
  assign n325 = x185 ^ x76 ^ x48 ;
  assign n326 = ( ~x95 & x115 ) | ( ~x95 & n310 ) | ( x115 & n310 ) ;
  assign n327 = ( x96 & ~x190 ) | ( x96 & n293 ) | ( ~x190 & n293 ) ;
  assign n328 = x38 & ~n276 ;
  assign n329 = ~x150 & n328 ;
  assign n330 = x228 ^ x12 ^ 1'b0 ;
  assign n331 = x240 & n330 ;
  assign n332 = ( x92 & x132 ) | ( x92 & ~n331 ) | ( x132 & ~n331 ) ;
  assign n333 = ( n327 & ~n329 ) | ( n327 & n332 ) | ( ~n329 & n332 ) ;
  assign n334 = x37 & x49 ;
  assign n335 = n334 ^ x37 ^ 1'b0 ;
  assign n336 = x100 & x215 ;
  assign n337 = n336 ^ x179 ^ 1'b0 ;
  assign n338 = n337 ^ x116 ^ 1'b0 ;
  assign n339 = x188 & ~n338 ;
  assign n340 = x145 & x180 ;
  assign n341 = ~n339 & n340 ;
  assign n342 = x32 | n268 ;
  assign n343 = ( x27 & ~x164 ) | ( x27 & x245 ) | ( ~x164 & x245 ) ;
  assign n344 = ( ~x15 & x90 ) | ( ~x15 & n343 ) | ( x90 & n343 ) ;
  assign n345 = ( x171 & n342 ) | ( x171 & n344 ) | ( n342 & n344 ) ;
  assign n346 = ( x159 & ~x233 ) | ( x159 & n326 ) | ( ~x233 & n326 ) ;
  assign n347 = ( ~x5 & x127 ) | ( ~x5 & x248 ) | ( x127 & x248 ) ;
  assign n348 = x182 & n262 ;
  assign n349 = ~x140 & n348 ;
  assign n350 = ( n262 & n347 ) | ( n262 & n349 ) | ( n347 & n349 ) ;
  assign n351 = x238 ^ x162 ^ x137 ;
  assign n352 = ( ~x162 & x190 ) | ( ~x162 & x250 ) | ( x190 & x250 ) ;
  assign n353 = n352 ^ x148 ^ x66 ;
  assign n354 = x137 & ~n353 ;
  assign n355 = n351 & n354 ;
  assign n356 = n355 ^ x253 ^ x225 ;
  assign n357 = n350 & n356 ;
  assign n358 = ~x57 & n357 ;
  assign n359 = x231 ^ x61 ^ 1'b0 ;
  assign n360 = x47 & n359 ;
  assign n361 = n360 ^ n353 ^ 1'b0 ;
  assign n362 = n293 | n361 ;
  assign n363 = n332 ^ n280 ^ x38 ;
  assign n364 = x219 ^ x111 ^ x3 ;
  assign n365 = x1 & x240 ;
  assign n366 = ~x143 & n365 ;
  assign n367 = n277 ^ x190 ^ 1'b0 ;
  assign n368 = x245 & ~n367 ;
  assign n369 = ~n366 & n368 ;
  assign n370 = n369 ^ x26 ^ 1'b0 ;
  assign n371 = n364 | n370 ;
  assign n372 = x24 | n371 ;
  assign n373 = x112 ^ x44 ^ 1'b0 ;
  assign n374 = x199 & n373 ;
  assign n375 = x194 & n374 ;
  assign n376 = ~x124 & n375 ;
  assign n377 = x182 & x193 ;
  assign n378 = ~x49 & n377 ;
  assign n383 = x72 & x127 ;
  assign n384 = n383 ^ x20 ^ 1'b0 ;
  assign n381 = n307 ^ x204 ^ x151 ;
  assign n382 = x22 & ~n381 ;
  assign n385 = n384 ^ n382 ^ 1'b0 ;
  assign n386 = ( x228 & x231 ) | ( x228 & ~n385 ) | ( x231 & ~n385 ) ;
  assign n379 = x8 & x87 ;
  assign n380 = n379 ^ n337 ^ 1'b0 ;
  assign n387 = n386 ^ n380 ^ x175 ;
  assign n388 = x144 ^ x134 ^ 1'b0 ;
  assign n389 = ( n353 & ~n387 ) | ( n353 & n388 ) | ( ~n387 & n388 ) ;
  assign n390 = ~n378 & n389 ;
  assign n391 = n390 ^ x88 ^ 1'b0 ;
  assign n392 = n368 ^ n324 ^ 1'b0 ;
  assign n393 = x13 & n363 ;
  assign n394 = ( x206 & n304 ) | ( x206 & ~n352 ) | ( n304 & ~n352 ) ;
  assign n395 = ( ~x135 & x165 ) | ( ~x135 & x200 ) | ( x165 & x200 ) ;
  assign n396 = x212 & n395 ;
  assign n397 = n293 & n396 ;
  assign n398 = x2 & ~n397 ;
  assign n399 = n398 ^ x134 ^ 1'b0 ;
  assign n400 = ( x152 & n394 ) | ( x152 & ~n399 ) | ( n394 & ~n399 ) ;
  assign n401 = ( x60 & ~x184 ) | ( x60 & n397 ) | ( ~x184 & n397 ) ;
  assign n402 = n270 ^ x21 ^ 1'b0 ;
  assign n403 = x166 & ~n402 ;
  assign n404 = x177 & n403 ;
  assign n405 = n404 ^ n380 ^ 1'b0 ;
  assign n406 = x234 ^ x68 ^ 1'b0 ;
  assign n407 = x251 & n406 ;
  assign n408 = n405 & n407 ;
  assign n409 = n297 | n408 ;
  assign n410 = n409 ^ n360 ^ 1'b0 ;
  assign n411 = x231 ^ x216 ^ 1'b0 ;
  assign n412 = x233 & n411 ;
  assign n413 = n275 ^ x101 ^ 1'b0 ;
  assign n414 = n412 & ~n413 ;
  assign n415 = x162 ^ x123 ^ 1'b0 ;
  assign n416 = n414 & n415 ;
  assign n417 = x225 & n416 ;
  assign n418 = n417 ^ n374 ^ 1'b0 ;
  assign n419 = ( ~x39 & x131 ) | ( ~x39 & x169 ) | ( x131 & x169 ) ;
  assign n420 = x151 & n260 ;
  assign n421 = ~n419 & n420 ;
  assign n422 = n407 ^ n389 ^ x189 ;
  assign n423 = ( x22 & ~x32 ) | ( x22 & x49 ) | ( ~x32 & x49 ) ;
  assign n424 = n418 ^ x28 ^ 1'b0 ;
  assign n425 = n423 & ~n424 ;
  assign n426 = ( x16 & ~x24 ) | ( x16 & x249 ) | ( ~x24 & x249 ) ;
  assign n427 = ( ~x15 & n362 ) | ( ~x15 & n426 ) | ( n362 & n426 ) ;
  assign n428 = n346 & ~n427 ;
  assign n429 = n343 ^ x191 ^ x4 ;
  assign n430 = n426 & ~n429 ;
  assign n431 = n430 ^ x118 ^ 1'b0 ;
  assign n432 = ( x35 & x171 ) | ( x35 & n362 ) | ( x171 & n362 ) ;
  assign n433 = ( ~x49 & x54 ) | ( ~x49 & x208 ) | ( x54 & x208 ) ;
  assign n434 = n384 ^ x213 ^ x204 ;
  assign n435 = ( ~x0 & x153 ) | ( ~x0 & n265 ) | ( x153 & n265 ) ;
  assign n436 = ( x161 & ~x210 ) | ( x161 & n435 ) | ( ~x210 & n435 ) ;
  assign n437 = ~n434 & n436 ;
  assign n438 = n394 ^ x233 ^ x148 ;
  assign n439 = ( ~x127 & x150 ) | ( ~x127 & x251 ) | ( x150 & x251 ) ;
  assign n440 = ( x117 & ~n438 ) | ( x117 & n439 ) | ( ~n438 & n439 ) ;
  assign n441 = ( ~x9 & x204 ) | ( ~x9 & n310 ) | ( x204 & n310 ) ;
  assign n442 = x119 & n345 ;
  assign n443 = ~x125 & n442 ;
  assign n444 = x190 ^ x20 ^ 1'b0 ;
  assign n445 = x64 & n444 ;
  assign n446 = n445 ^ n360 ^ x219 ;
  assign n447 = ( ~x79 & x132 ) | ( ~x79 & n446 ) | ( x132 & n446 ) ;
  assign n448 = ( x19 & ~x224 ) | ( x19 & n399 ) | ( ~x224 & n399 ) ;
  assign n449 = x16 & x166 ;
  assign n450 = ~x13 & n449 ;
  assign n451 = x204 ^ x168 ^ x113 ;
  assign n452 = n450 | n451 ;
  assign n453 = n286 & ~n452 ;
  assign n454 = n453 ^ x227 ^ 1'b0 ;
  assign n459 = ( x130 & x155 ) | ( x130 & ~x209 ) | ( x155 & ~x209 ) ;
  assign n460 = ( x72 & n384 ) | ( x72 & n459 ) | ( n384 & n459 ) ;
  assign n456 = x88 ^ x62 ^ x30 ;
  assign n457 = x219 & ~n456 ;
  assign n458 = n457 ^ n258 ^ 1'b0 ;
  assign n461 = n460 ^ n458 ^ n322 ;
  assign n455 = n426 & ~n437 ;
  assign n462 = n461 ^ n455 ^ 1'b0 ;
  assign n463 = ~x90 & x122 ;
  assign n464 = ( x205 & n342 ) | ( x205 & n463 ) | ( n342 & n463 ) ;
  assign n465 = ( x64 & x191 ) | ( x64 & n351 ) | ( x191 & n351 ) ;
  assign n466 = n465 ^ x122 ^ x109 ;
  assign n467 = x55 & n403 ;
  assign n468 = n467 ^ x235 ^ 1'b0 ;
  assign n469 = n343 & n468 ;
  assign n470 = x171 & ~n469 ;
  assign n471 = n470 ^ n438 ^ x193 ;
  assign n472 = n471 ^ x147 ^ 1'b0 ;
  assign n473 = n307 ^ x108 ^ 1'b0 ;
  assign n474 = ( ~x30 & x44 ) | ( ~x30 & x206 ) | ( x44 & x206 ) ;
  assign n475 = ( x85 & n258 ) | ( x85 & n279 ) | ( n258 & n279 ) ;
  assign n476 = n475 ^ n279 ^ x144 ;
  assign n477 = n296 ^ x236 ^ x178 ;
  assign n478 = ( n287 & ~n476 ) | ( n287 & n477 ) | ( ~n476 & n477 ) ;
  assign n479 = x126 & n478 ;
  assign n480 = ~n474 & n479 ;
  assign n481 = n279 ^ x129 ^ x68 ;
  assign n482 = x145 ^ x107 ^ 1'b0 ;
  assign n483 = x96 & n482 ;
  assign n484 = n483 ^ x140 ^ 1'b0 ;
  assign n485 = n481 & n484 ;
  assign n489 = x205 & ~n364 ;
  assign n490 = n489 ^ x202 ^ x66 ;
  assign n491 = n469 & n490 ;
  assign n486 = x16 & x194 ;
  assign n487 = n486 ^ x33 ^ 1'b0 ;
  assign n488 = n487 ^ n266 ^ 1'b0 ;
  assign n492 = n491 ^ n488 ^ x218 ;
  assign n494 = x49 & ~x161 ;
  assign n493 = x108 ^ x76 ^ x6 ;
  assign n495 = n494 ^ n493 ^ n416 ;
  assign n496 = n397 | n495 ;
  assign n497 = n476 | n496 ;
  assign n498 = ( x61 & x160 ) | ( x61 & ~n392 ) | ( x160 & ~n392 ) ;
  assign n499 = ( x43 & x56 ) | ( x43 & ~x104 ) | ( x56 & ~x104 ) ;
  assign n500 = ( x100 & ~n374 ) | ( x100 & n499 ) | ( ~n374 & n499 ) ;
  assign n513 = x184 ^ x68 ^ 1'b0 ;
  assign n512 = ( x82 & ~x125 ) | ( x82 & n324 ) | ( ~x125 & n324 ) ;
  assign n503 = x45 & x86 ;
  assign n504 = ~x42 & n503 ;
  assign n505 = n504 ^ x78 ^ x49 ;
  assign n508 = ( x15 & x162 ) | ( x15 & ~n426 ) | ( x162 & ~n426 ) ;
  assign n506 = x156 ^ x105 ^ 1'b0 ;
  assign n507 = n306 & n506 ;
  assign n509 = n508 ^ n507 ^ 1'b0 ;
  assign n510 = ( ~x225 & n505 ) | ( ~x225 & n509 ) | ( n505 & n509 ) ;
  assign n501 = x213 ^ x145 ^ x34 ;
  assign n502 = ( x85 & n315 ) | ( x85 & n501 ) | ( n315 & n501 ) ;
  assign n511 = n510 ^ n502 ^ 1'b0 ;
  assign n514 = n513 ^ n512 ^ n511 ;
  assign n515 = x191 & x216 ;
  assign n516 = ~n260 & n515 ;
  assign n517 = ( x162 & ~n362 ) | ( x162 & n516 ) | ( ~n362 & n516 ) ;
  assign n518 = n517 ^ x39 ^ 1'b0 ;
  assign n519 = n304 ^ x168 ^ x155 ;
  assign n520 = n519 ^ n426 ^ x170 ;
  assign n521 = n520 ^ x17 ^ 1'b0 ;
  assign n522 = x160 & n521 ;
  assign n523 = n522 ^ x59 ^ 1'b0 ;
  assign n525 = x171 & n358 ;
  assign n524 = x65 & ~n520 ;
  assign n526 = n525 ^ n524 ^ 1'b0 ;
  assign n527 = n504 ^ n262 ^ 1'b0 ;
  assign n528 = x48 & ~n527 ;
  assign n529 = n528 ^ x187 ^ x65 ;
  assign n530 = ( x185 & ~n368 ) | ( x185 & n426 ) | ( ~n368 & n426 ) ;
  assign n531 = ( ~x28 & n529 ) | ( ~x28 & n530 ) | ( n529 & n530 ) ;
  assign n532 = x105 & x230 ;
  assign n533 = n532 ^ x87 ^ 1'b0 ;
  assign n534 = x201 ^ x170 ^ x50 ;
  assign n535 = x200 & ~n534 ;
  assign n536 = n535 ^ x182 ^ 1'b0 ;
  assign n537 = x89 & x231 ;
  assign n538 = ~x175 & n537 ;
  assign n539 = ( n533 & ~n536 ) | ( n533 & n538 ) | ( ~n536 & n538 ) ;
  assign n540 = ( ~x59 & n266 ) | ( ~x59 & n289 ) | ( n266 & n289 ) ;
  assign n542 = n434 ^ x232 ^ x143 ;
  assign n543 = n467 & ~n542 ;
  assign n544 = ~x142 & n543 ;
  assign n545 = x38 | n544 ;
  assign n546 = n545 ^ n478 ^ 1'b0 ;
  assign n541 = x213 & n308 ;
  assign n547 = n546 ^ n541 ^ n475 ;
  assign n548 = n540 & ~n547 ;
  assign n549 = n273 & n548 ;
  assign n550 = n433 ^ x63 ^ 1'b0 ;
  assign n551 = n550 ^ x85 ^ 1'b0 ;
  assign n552 = n322 ^ x212 ^ 1'b0 ;
  assign n553 = n551 | n552 ;
  assign n554 = x76 & n553 ;
  assign n555 = x250 ^ x225 ^ x144 ;
  assign n556 = n341 | n555 ;
  assign n557 = n556 ^ x115 ^ 1'b0 ;
  assign n558 = n545 ^ n477 ^ n300 ;
  assign n559 = x72 & ~x217 ;
  assign n560 = x140 & n559 ;
  assign n561 = ( x50 & x219 ) | ( x50 & ~x220 ) | ( x219 & ~x220 ) ;
  assign n562 = n561 ^ n414 ^ 1'b0 ;
  assign n563 = x146 ^ x98 ^ x89 ;
  assign n564 = n563 ^ n456 ^ x9 ;
  assign n565 = n499 ^ x92 ^ x2 ;
  assign n566 = n565 ^ n326 ^ n257 ;
  assign n567 = ( x231 & ~n387 ) | ( x231 & n566 ) | ( ~n387 & n566 ) ;
  assign n569 = ( x156 & ~x210 ) | ( x156 & n419 ) | ( ~x210 & n419 ) ;
  assign n568 = n290 | n376 ;
  assign n570 = n569 ^ n568 ^ 1'b0 ;
  assign n571 = x153 ^ x71 ^ 1'b0 ;
  assign n572 = x167 & n571 ;
  assign n573 = n572 ^ x209 ^ x148 ;
  assign n574 = n516 | n573 ;
  assign n575 = n563 & ~n574 ;
  assign n576 = x226 ^ x186 ^ x155 ;
  assign n577 = ( ~x42 & x85 ) | ( ~x42 & n576 ) | ( x85 & n576 ) ;
  assign n578 = n403 ^ x78 ^ 1'b0 ;
  assign n579 = x212 & n578 ;
  assign n580 = x151 & ~n579 ;
  assign n581 = n580 ^ x243 ^ 1'b0 ;
  assign n582 = n577 | n581 ;
  assign n583 = x78 & ~n582 ;
  assign n584 = n583 ^ n257 ^ 1'b0 ;
  assign n586 = x171 ^ x134 ^ x93 ;
  assign n587 = ( ~x27 & x148 ) | ( ~x27 & x154 ) | ( x148 & x154 ) ;
  assign n588 = ( ~x113 & n586 ) | ( ~x113 & n587 ) | ( n586 & n587 ) ;
  assign n589 = ( ~x211 & x234 ) | ( ~x211 & n588 ) | ( x234 & n588 ) ;
  assign n585 = ( x190 & x204 ) | ( x190 & ~n372 ) | ( x204 & ~n372 ) ;
  assign n590 = n589 ^ n585 ^ 1'b0 ;
  assign n591 = n332 & ~n590 ;
  assign n592 = n591 ^ n547 ^ n320 ;
  assign n593 = n592 ^ n314 ^ x114 ;
  assign n594 = n492 ^ x174 ^ 1'b0 ;
  assign n595 = n594 ^ n570 ^ x63 ;
  assign n596 = x199 ^ x172 ^ x115 ;
  assign n597 = x42 & x109 ;
  assign n598 = n596 & n597 ;
  assign n599 = n432 ^ x171 ^ 1'b0 ;
  assign n600 = ( n276 & n332 ) | ( n276 & ~n599 ) | ( n332 & ~n599 ) ;
  assign n601 = x175 ^ x29 ^ 1'b0 ;
  assign n602 = n601 ^ x124 ^ x97 ;
  assign n603 = ( n342 & n573 ) | ( n342 & n602 ) | ( n573 & n602 ) ;
  assign n604 = ( ~n598 & n600 ) | ( ~n598 & n603 ) | ( n600 & n603 ) ;
  assign n605 = n346 & ~n565 ;
  assign n606 = n451 & n605 ;
  assign n607 = n376 ^ x254 ^ x89 ;
  assign n608 = ( n324 & n606 ) | ( n324 & n607 ) | ( n606 & n607 ) ;
  assign n613 = ( x63 & ~x250 ) | ( x63 & n337 ) | ( ~x250 & n337 ) ;
  assign n612 = x224 & n380 ;
  assign n614 = n613 ^ n612 ^ 1'b0 ;
  assign n609 = x149 & ~n307 ;
  assign n610 = n609 ^ n501 ^ x103 ;
  assign n611 = x77 & ~n610 ;
  assign n615 = n614 ^ n611 ^ 1'b0 ;
  assign n620 = ( n306 & n516 ) | ( n306 & n519 ) | ( n516 & n519 ) ;
  assign n621 = n547 ^ n490 ^ 1'b0 ;
  assign n622 = n620 & n621 ;
  assign n616 = x91 & x137 ;
  assign n617 = n616 ^ n586 ^ 1'b0 ;
  assign n618 = n617 ^ x22 ^ 1'b0 ;
  assign n619 = n454 | n618 ;
  assign n623 = n622 ^ n619 ^ 1'b0 ;
  assign n624 = x245 ^ x131 ^ x37 ;
  assign n625 = n624 ^ n312 ^ 1'b0 ;
  assign n626 = ( x212 & n495 ) | ( x212 & n625 ) | ( n495 & n625 ) ;
  assign n627 = ( ~x217 & x251 ) | ( ~x217 & n626 ) | ( x251 & n626 ) ;
  assign n628 = n339 ^ x253 ^ 1'b0 ;
  assign n632 = x236 & n326 ;
  assign n629 = x50 & x71 ;
  assign n630 = ~x203 & n629 ;
  assign n631 = ( x89 & ~n606 ) | ( x89 & n630 ) | ( ~n606 & n630 ) ;
  assign n633 = n632 ^ n631 ^ 1'b0 ;
  assign n634 = ~x54 & x57 ;
  assign n635 = x77 & x157 ;
  assign n636 = ~x231 & n635 ;
  assign n637 = x120 & x184 ;
  assign n638 = ~x219 & n637 ;
  assign n639 = n335 | n638 ;
  assign n640 = ( n634 & ~n636 ) | ( n634 & n639 ) | ( ~n636 & n639 ) ;
  assign n641 = x29 & x110 ;
  assign n642 = ~x204 & n641 ;
  assign n643 = n642 ^ x60 ^ 1'b0 ;
  assign n644 = ( n483 & ~n640 ) | ( n483 & n643 ) | ( ~n640 & n643 ) ;
  assign n645 = x254 ^ x134 ^ x107 ;
  assign n646 = x61 ^ x56 ^ x13 ;
  assign n647 = n646 ^ n463 ^ 1'b0 ;
  assign n648 = ~x162 & n339 ;
  assign n649 = n296 | n648 ;
  assign n650 = n649 ^ n450 ^ 1'b0 ;
  assign n651 = n313 & ~n472 ;
  assign n652 = ~x227 & n651 ;
  assign n653 = x66 & x105 ;
  assign n654 = n653 ^ x43 ^ 1'b0 ;
  assign n655 = ~n349 & n654 ;
  assign n656 = n655 ^ n279 ^ 1'b0 ;
  assign n657 = n656 ^ n508 ^ x204 ;
  assign n658 = x214 ^ x41 ^ x22 ;
  assign n659 = n421 | n658 ;
  assign n660 = n657 & ~n659 ;
  assign n661 = n540 ^ n297 ^ x39 ;
  assign n662 = ( x128 & n587 ) | ( x128 & ~n661 ) | ( n587 & ~n661 ) ;
  assign n663 = x50 ^ x15 ^ 1'b0 ;
  assign n664 = x245 & ~n663 ;
  assign n665 = n664 ^ n466 ^ x117 ;
  assign n666 = n662 & ~n665 ;
  assign n668 = n475 ^ x181 ^ 1'b0 ;
  assign n667 = ~n283 & n389 ;
  assign n669 = n668 ^ n667 ^ n586 ;
  assign n670 = n669 ^ n643 ^ x246 ;
  assign n671 = ( x149 & x157 ) | ( x149 & ~x249 ) | ( x157 & ~x249 ) ;
  assign n672 = n671 ^ x144 ^ x14 ;
  assign n673 = ( n261 & n666 ) | ( n261 & n672 ) | ( n666 & n672 ) ;
  assign n674 = x134 ^ x71 ^ 1'b0 ;
  assign n675 = n303 ^ x237 ^ x166 ;
  assign n677 = x148 & x183 ;
  assign n678 = ~x124 & n677 ;
  assign n676 = x24 & x210 ;
  assign n679 = n678 ^ n676 ^ n451 ;
  assign n680 = n675 & ~n679 ;
  assign n681 = ~n674 & n680 ;
  assign n682 = ( ~n306 & n478 ) | ( ~n306 & n661 ) | ( n478 & n661 ) ;
  assign n683 = ( x66 & n437 ) | ( x66 & ~n682 ) | ( n437 & ~n682 ) ;
  assign n684 = ( n266 & ~n303 ) | ( n266 & n634 ) | ( ~n303 & n634 ) ;
  assign n685 = x242 ^ x225 ^ x45 ;
  assign n686 = x139 & ~n469 ;
  assign n687 = ( n355 & n685 ) | ( n355 & ~n686 ) | ( n685 & ~n686 ) ;
  assign n688 = ( n410 & n684 ) | ( n410 & n687 ) | ( n684 & n687 ) ;
  assign n689 = x205 ^ x164 ^ x32 ;
  assign n690 = n689 ^ x60 ^ x22 ;
  assign n691 = x244 & ~n293 ;
  assign n692 = n691 ^ n257 ^ 1'b0 ;
  assign n693 = ( x53 & x142 ) | ( x53 & ~n692 ) | ( x142 & ~n692 ) ;
  assign n694 = n693 ^ x235 ^ 1'b0 ;
  assign n695 = n690 & n694 ;
  assign n697 = x52 & ~x244 ;
  assign n698 = x253 ^ x159 ^ 1'b0 ;
  assign n699 = ~n560 & n698 ;
  assign n700 = n697 & n699 ;
  assign n696 = n335 ^ x1 ^ 1'b0 ;
  assign n701 = n700 ^ n696 ^ 1'b0 ;
  assign n702 = n701 ^ x246 ^ x13 ;
  assign n707 = ( x127 & x210 ) | ( x127 & ~n684 ) | ( x210 & ~n684 ) ;
  assign n708 = n598 ^ n569 ^ x144 ;
  assign n709 = x113 & n708 ;
  assign n710 = n709 ^ n576 ^ 1'b0 ;
  assign n711 = ( ~n587 & n707 ) | ( ~n587 & n710 ) | ( n707 & n710 ) ;
  assign n703 = x116 & n596 ;
  assign n704 = x205 | n703 ;
  assign n705 = n285 ^ x154 ^ x45 ;
  assign n706 = ( ~x82 & n704 ) | ( ~x82 & n705 ) | ( n704 & n705 ) ;
  assign n712 = n711 ^ n706 ^ 1'b0 ;
  assign n717 = n561 ^ n493 ^ x38 ;
  assign n716 = n545 ^ x164 ^ x38 ;
  assign n718 = n717 ^ n716 ^ n290 ;
  assign n714 = x39 & x165 ;
  assign n715 = n714 ^ x219 ^ 1'b0 ;
  assign n719 = n718 ^ n715 ^ n531 ;
  assign n713 = n553 ^ x166 ^ 1'b0 ;
  assign n720 = n719 ^ n713 ^ x59 ;
  assign n721 = ( n362 & n395 ) | ( n362 & n720 ) | ( n395 & n720 ) ;
  assign n722 = ( x71 & ~x126 ) | ( x71 & x211 ) | ( ~x126 & x211 ) ;
  assign n723 = n722 ^ n351 ^ x86 ;
  assign n724 = n723 ^ n432 ^ 1'b0 ;
  assign n725 = ( x160 & n435 ) | ( x160 & n504 ) | ( n435 & n504 ) ;
  assign n726 = x152 & x161 ;
  assign n727 = ~n725 & n726 ;
  assign n737 = ( x111 & n264 ) | ( x111 & n596 ) | ( n264 & n596 ) ;
  assign n739 = x218 ^ x134 ^ x38 ;
  assign n740 = ( x20 & ~n737 ) | ( x20 & n739 ) | ( ~n737 & n739 ) ;
  assign n736 = ( x31 & x125 ) | ( x31 & ~n368 ) | ( x125 & ~n368 ) ;
  assign n738 = ( ~n298 & n736 ) | ( ~n298 & n737 ) | ( n736 & n737 ) ;
  assign n731 = x67 & x109 ;
  assign n732 = n731 ^ x80 ^ 1'b0 ;
  assign n733 = n732 ^ n451 ^ x171 ;
  assign n734 = ( x28 & n636 ) | ( x28 & ~n733 ) | ( n636 & ~n733 ) ;
  assign n728 = x108 & x254 ;
  assign n729 = ~x122 & n728 ;
  assign n730 = n729 ^ n636 ^ x58 ;
  assign n735 = n734 ^ n730 ^ x97 ;
  assign n741 = n740 ^ n738 ^ n735 ;
  assign n742 = n523 ^ n458 ^ n440 ;
  assign n743 = n414 & ~n739 ;
  assign n744 = ~x18 & n743 ;
  assign n745 = n423 & ~n474 ;
  assign n746 = n745 ^ n363 ^ 1'b0 ;
  assign n747 = x204 ^ x37 ^ 1'b0 ;
  assign n748 = x93 & n747 ;
  assign n749 = n734 & n748 ;
  assign n750 = ~n393 & n749 ;
  assign n751 = ( n508 & ~n577 ) | ( n508 & n750 ) | ( ~n577 & n750 ) ;
  assign n752 = n710 ^ n646 ^ x10 ;
  assign n753 = ( x80 & ~n511 ) | ( x80 & n752 ) | ( ~n511 & n752 ) ;
  assign n757 = n558 ^ x167 ^ 1'b0 ;
  assign n758 = ~n283 & n757 ;
  assign n759 = ( ~x68 & n608 ) | ( ~x68 & n758 ) | ( n608 & n758 ) ;
  assign n760 = x21 & x198 ;
  assign n761 = n760 ^ x233 ^ 1'b0 ;
  assign n762 = n761 ^ x186 ^ 1'b0 ;
  assign n763 = n736 & ~n762 ;
  assign n764 = x64 & n763 ;
  assign n765 = ~n759 & n764 ;
  assign n754 = n618 ^ n384 ^ 1'b0 ;
  assign n755 = ~n520 & n754 ;
  assign n756 = n462 & n755 ;
  assign n766 = n765 ^ n756 ^ 1'b0 ;
  assign n767 = ( x28 & ~x129 ) | ( x28 & n320 ) | ( ~x129 & n320 ) ;
  assign n775 = n767 ^ n282 ^ x29 ;
  assign n768 = n767 ^ x91 ^ 1'b0 ;
  assign n769 = x249 ^ x79 ^ 1'b0 ;
  assign n770 = n426 & n769 ;
  assign n771 = ( x59 & ~n256 ) | ( x59 & n579 ) | ( ~n256 & n579 ) ;
  assign n772 = ( n563 & n770 ) | ( n563 & ~n771 ) | ( n770 & ~n771 ) ;
  assign n773 = ( x159 & ~n768 ) | ( x159 & n772 ) | ( ~n768 & n772 ) ;
  assign n774 = n773 ^ n431 ^ 1'b0 ;
  assign n776 = n775 ^ n774 ^ n471 ;
  assign n777 = n315 | n458 ;
  assign n778 = n777 ^ n381 ^ 1'b0 ;
  assign n779 = ( x123 & ~n558 ) | ( x123 & n778 ) | ( ~n558 & n778 ) ;
  assign n780 = ( ~x160 & n276 ) | ( ~x160 & n440 ) | ( n276 & n440 ) ;
  assign n781 = n609 ^ n341 ^ x12 ;
  assign n782 = x34 & x78 ;
  assign n783 = ~x238 & n782 ;
  assign n784 = n675 & n783 ;
  assign n785 = ( n780 & n781 ) | ( n780 & ~n784 ) | ( n781 & ~n784 ) ;
  assign n786 = ( x9 & ~x138 ) | ( x9 & n499 ) | ( ~x138 & n499 ) ;
  assign n800 = ~n327 & n767 ;
  assign n795 = n499 ^ n270 ^ x226 ;
  assign n796 = n795 ^ n412 ^ n343 ;
  assign n797 = n796 ^ n300 ^ x136 ;
  assign n794 = x76 & n414 ;
  assign n798 = n797 ^ n794 ^ 1'b0 ;
  assign n789 = n323 ^ x254 ^ x237 ;
  assign n790 = n789 ^ n775 ^ 1'b0 ;
  assign n791 = n530 & n790 ;
  assign n788 = n329 ^ n285 ^ 1'b0 ;
  assign n792 = n791 ^ n788 ^ x201 ;
  assign n793 = n792 ^ x231 ^ x140 ;
  assign n799 = n798 ^ n793 ^ 1'b0 ;
  assign n787 = x169 ^ x120 ^ 1'b0 ;
  assign n801 = n800 ^ n799 ^ n787 ;
  assign n802 = n778 ^ n483 ^ x196 ;
  assign n803 = n646 ^ n560 ^ n433 ;
  assign n804 = n644 & ~n715 ;
  assign n805 = n600 & n804 ;
  assign n806 = ( x97 & ~n332 ) | ( x97 & n423 ) | ( ~n332 & n423 ) ;
  assign n807 = n806 ^ n463 ^ x128 ;
  assign n808 = n807 ^ x254 ^ x124 ;
  assign n809 = x194 & ~n534 ;
  assign n810 = n809 ^ n393 ^ 1'b0 ;
  assign n811 = n810 ^ n690 ^ 1'b0 ;
  assign n818 = ( x211 & n257 ) | ( x211 & ~n267 ) | ( n257 & ~n267 ) ;
  assign n815 = x22 ^ x15 ^ 1'b0 ;
  assign n816 = n815 ^ x120 ^ 1'b0 ;
  assign n812 = ( ~x61 & n262 ) | ( ~x61 & n366 ) | ( n262 & n366 ) ;
  assign n813 = n812 ^ x200 ^ x73 ;
  assign n814 = x117 & n813 ;
  assign n817 = n816 ^ n814 ^ 1'b0 ;
  assign n819 = n818 ^ n817 ^ 1'b0 ;
  assign n820 = x92 ^ x2 ^ 1'b0 ;
  assign n821 = x233 & n820 ;
  assign n822 = n821 ^ n601 ^ n510 ;
  assign n823 = n587 ^ n460 ^ 1'b0 ;
  assign n824 = x164 & n823 ;
  assign n825 = x205 & n824 ;
  assign n826 = n822 & n825 ;
  assign n827 = n475 & ~n689 ;
  assign n828 = ~x239 & n827 ;
  assign n829 = n685 ^ n499 ^ x171 ;
  assign n830 = ( ~x199 & n333 ) | ( ~x199 & n441 ) | ( n333 & n441 ) ;
  assign n831 = ( n828 & n829 ) | ( n828 & n830 ) | ( n829 & n830 ) ;
  assign n832 = ~n826 & n831 ;
  assign n833 = n832 ^ x147 ^ 1'b0 ;
  assign n834 = n267 | n833 ;
  assign n835 = x139 & n822 ;
  assign n836 = n835 ^ n679 ^ n339 ;
  assign n837 = x59 & x114 ;
  assign n838 = n837 ^ n304 ^ 1'b0 ;
  assign n839 = n838 ^ x84 ^ 1'b0 ;
  assign n840 = x237 & n839 ;
  assign n841 = n840 ^ n604 ^ n585 ;
  assign n842 = n501 ^ x232 ^ x68 ;
  assign n843 = n842 ^ n697 ^ x164 ;
  assign n846 = x67 & n261 ;
  assign n847 = n846 ^ n307 ^ 1'b0 ;
  assign n848 = ( ~x68 & n380 ) | ( ~x68 & n847 ) | ( n380 & n847 ) ;
  assign n844 = n308 | n582 ;
  assign n845 = n506 & ~n844 ;
  assign n849 = n848 ^ n845 ^ 1'b0 ;
  assign n850 = x6 & n849 ;
  assign n851 = ~x147 & n850 ;
  assign n852 = n682 & ~n722 ;
  assign n853 = n852 ^ n512 ^ x12 ;
  assign n854 = n487 ^ x199 ^ x192 ;
  assign n855 = n795 ^ x138 ^ 1'b0 ;
  assign n856 = n854 & n855 ;
  assign n857 = ( x254 & n582 ) | ( x254 & n789 ) | ( n582 & n789 ) ;
  assign n858 = x52 & x220 ;
  assign n859 = n858 ^ n395 ^ 1'b0 ;
  assign n860 = n859 ^ n428 ^ n370 ;
  assign n861 = ( ~x244 & n351 ) | ( ~x244 & n860 ) | ( n351 & n860 ) ;
  assign n862 = ( n856 & n857 ) | ( n856 & ~n861 ) | ( n857 & ~n861 ) ;
  assign n863 = x76 & ~n518 ;
  assign n864 = n647 & n863 ;
  assign n865 = x75 & ~n587 ;
  assign n866 = ( x19 & x23 ) | ( x19 & n865 ) | ( x23 & n865 ) ;
  assign n867 = n866 ^ n751 ^ 1'b0 ;
  assign n868 = ~n504 & n867 ;
  assign n869 = n498 ^ n394 ^ 1'b0 ;
  assign n870 = n303 | n869 ;
  assign n871 = n696 ^ x231 ^ x45 ;
  assign n872 = n857 & ~n871 ;
  assign n873 = n538 & n755 ;
  assign n874 = n830 ^ n582 ^ n488 ;
  assign n875 = n646 ^ x7 ^ 1'b0 ;
  assign n876 = n874 | n875 ;
  assign n877 = ( x218 & n873 ) | ( x218 & n876 ) | ( n873 & n876 ) ;
  assign n880 = x252 ^ x181 ^ x166 ;
  assign n878 = x176 ^ x22 ^ 1'b0 ;
  assign n879 = x179 & n878 ;
  assign n881 = n880 ^ n879 ^ 1'b0 ;
  assign n882 = x114 & ~n881 ;
  assign n883 = ( n277 & ~n740 ) | ( n277 & n882 ) | ( ~n740 & n882 ) ;
  assign n884 = ( x203 & n865 ) | ( x203 & ~n883 ) | ( n865 & ~n883 ) ;
  assign n885 = ( x38 & ~x68 ) | ( x38 & n600 ) | ( ~x68 & n600 ) ;
  assign n886 = n446 | n885 ;
  assign n887 = n886 ^ x158 ^ 1'b0 ;
  assign n888 = ( ~x133 & n405 ) | ( ~x133 & n887 ) | ( n405 & n887 ) ;
  assign n889 = x70 & ~n539 ;
  assign n890 = ~x79 & n889 ;
  assign n891 = ( x62 & ~n671 ) | ( x62 & n733 ) | ( ~n671 & n733 ) ;
  assign n892 = ( n318 & ~n890 ) | ( n318 & n891 ) | ( ~n890 & n891 ) ;
  assign n893 = n892 ^ n765 ^ n564 ;
  assign n894 = ( x106 & x229 ) | ( x106 & n796 ) | ( x229 & n796 ) ;
  assign n899 = n422 ^ x95 ^ x94 ;
  assign n896 = x232 ^ x197 ^ x155 ;
  assign n897 = ( ~x78 & x218 ) | ( ~x78 & n896 ) | ( x218 & n896 ) ;
  assign n895 = n797 ^ n638 ^ 1'b0 ;
  assign n898 = n897 ^ n895 ^ n643 ;
  assign n900 = n899 ^ n898 ^ 1'b0 ;
  assign n901 = ~x161 & n393 ;
  assign n902 = ( ~n407 & n483 ) | ( ~n407 & n901 ) | ( n483 & n901 ) ;
  assign n903 = n880 & n899 ;
  assign n906 = x199 & ~n358 ;
  assign n907 = n906 ^ n339 ^ 1'b0 ;
  assign n904 = x209 & ~n358 ;
  assign n905 = ~n505 & n904 ;
  assign n908 = n907 ^ n905 ^ 1'b0 ;
  assign n909 = n462 & n908 ;
  assign n910 = n261 ^ x133 ^ 1'b0 ;
  assign n911 = ( ~x243 & n655 ) | ( ~x243 & n910 ) | ( n655 & n910 ) ;
  assign n912 = ( x189 & ~n435 ) | ( x189 & n911 ) | ( ~n435 & n911 ) ;
  assign n913 = n275 ^ x124 ^ x68 ;
  assign n914 = ( x167 & x225 ) | ( x167 & n305 ) | ( x225 & n305 ) ;
  assign n915 = ~n349 & n771 ;
  assign n916 = n915 ^ x194 ^ 1'b0 ;
  assign n917 = n520 | n686 ;
  assign n918 = ( x52 & n916 ) | ( x52 & ~n917 ) | ( n916 & ~n917 ) ;
  assign n919 = n914 & n918 ;
  assign n920 = ~x63 & n919 ;
  assign n922 = x120 ^ x24 ^ x3 ;
  assign n921 = x189 & x217 ;
  assign n923 = n922 ^ n921 ^ 1'b0 ;
  assign n924 = n923 ^ x234 ^ x80 ;
  assign n925 = ( x16 & x158 ) | ( x16 & n924 ) | ( x158 & n924 ) ;
  assign n926 = x163 ^ x149 ^ x55 ;
  assign n927 = n926 ^ n559 ^ 1'b0 ;
  assign n928 = x214 & n927 ;
  assign n929 = x224 & ~n368 ;
  assign n930 = ( x42 & x95 ) | ( x42 & ~x143 ) | ( x95 & ~x143 ) ;
  assign n931 = n633 & n930 ;
  assign n932 = n931 ^ n646 ^ 1'b0 ;
  assign n933 = n771 ^ x139 ^ x31 ;
  assign n934 = ( ~x142 & x250 ) | ( ~x142 & n636 ) | ( x250 & n636 ) ;
  assign n935 = n860 & ~n934 ;
  assign n936 = n707 ^ x20 ^ 1'b0 ;
  assign n937 = ( n933 & ~n935 ) | ( n933 & n936 ) | ( ~n935 & n936 ) ;
  assign n938 = n513 ^ x93 ^ 1'b0 ;
  assign n939 = n346 & ~n378 ;
  assign n940 = x202 ^ x178 ^ x101 ;
  assign n941 = n940 ^ n860 ^ x74 ;
  assign n942 = n939 & n941 ;
  assign n943 = n773 & n942 ;
  assign n944 = n366 | n943 ;
  assign n945 = n576 & ~n944 ;
  assign n946 = n364 ^ n310 ^ x54 ;
  assign n947 = n946 ^ n337 ^ x101 ;
  assign n948 = ( x125 & x250 ) | ( x125 & ~n947 ) | ( x250 & ~n947 ) ;
  assign n949 = ( n654 & n670 ) | ( n654 & n729 ) | ( n670 & n729 ) ;
  assign n950 = ( ~x38 & x169 ) | ( ~x38 & n826 ) | ( x169 & n826 ) ;
  assign n951 = n646 | n950 ;
  assign n952 = n951 ^ n561 ^ 1'b0 ;
  assign n953 = ( n466 & n556 ) | ( n466 & n670 ) | ( n556 & n670 ) ;
  assign n954 = n953 ^ x218 ^ x138 ;
  assign n955 = ( x114 & ~x198 ) | ( x114 & n954 ) | ( ~x198 & n954 ) ;
  assign n956 = x4 & ~n295 ;
  assign n957 = n775 & n956 ;
  assign n958 = n591 ^ x113 ^ 1'b0 ;
  assign n959 = ~n957 & n958 ;
  assign n960 = n672 & ~n727 ;
  assign n961 = ( n692 & n959 ) | ( n692 & n960 ) | ( n959 & n960 ) ;
  assign n962 = n961 ^ x165 ^ 1'b0 ;
  assign n964 = x179 & n824 ;
  assign n965 = ~x243 & n964 ;
  assign n963 = n591 & n752 ;
  assign n966 = n965 ^ n963 ^ x31 ;
  assign n967 = n966 ^ n761 ^ 1'b0 ;
  assign n968 = n879 ^ x82 ^ 1'b0 ;
  assign n969 = ~n257 & n968 ;
  assign n970 = n538 | n689 ;
  assign n971 = x95 | n970 ;
  assign n972 = ( n399 & n969 ) | ( n399 & n971 ) | ( n969 & n971 ) ;
  assign n973 = x208 ^ x165 ^ x117 ;
  assign n974 = n301 | n394 ;
  assign n975 = ( n342 & n973 ) | ( n342 & ~n974 ) | ( n973 & ~n974 ) ;
  assign n976 = n821 ^ n358 ^ 1'b0 ;
  assign n977 = n674 & ~n976 ;
  assign n978 = n890 ^ n366 ^ x141 ;
  assign n979 = ( x70 & n678 ) | ( x70 & n978 ) | ( n678 & n978 ) ;
  assign n980 = ( n899 & n965 ) | ( n899 & ~n979 ) | ( n965 & ~n979 ) ;
  assign n981 = ~x137 & n287 ;
  assign n982 = ( ~n705 & n838 ) | ( ~n705 & n981 ) | ( n838 & n981 ) ;
  assign n983 = ( ~n324 & n477 ) | ( ~n324 & n494 ) | ( n477 & n494 ) ;
  assign n984 = n983 ^ n265 ^ x80 ;
  assign n985 = n298 & n497 ;
  assign n986 = n985 ^ x201 ^ 1'b0 ;
  assign n987 = n986 ^ n971 ^ 1'b0 ;
  assign n988 = x42 & ~n987 ;
  assign n989 = n988 ^ n806 ^ 1'b0 ;
  assign n990 = x89 & n587 ;
  assign n991 = n950 ^ n610 ^ x214 ;
  assign n992 = x172 ^ x65 ^ 1'b0 ;
  assign n993 = x22 & n992 ;
  assign n994 = n491 & n993 ;
  assign n995 = ~n991 & n994 ;
  assign n996 = n922 ^ n812 ^ 1'b0 ;
  assign n997 = x38 & n996 ;
  assign n998 = ( ~x152 & n859 ) | ( ~x152 & n997 ) | ( n859 & n997 ) ;
  assign n999 = n998 ^ n283 ^ x153 ;
  assign n1000 = ~n711 & n954 ;
  assign n1001 = n840 ^ x116 ^ 1'b0 ;
  assign n1002 = n607 & n1001 ;
  assign n1003 = n711 ^ n355 ^ x85 ;
  assign n1004 = n1003 ^ n953 ^ n389 ;
  assign n1005 = x251 ^ x187 ^ x33 ;
  assign n1009 = x155 & ~n342 ;
  assign n1010 = n1009 ^ n737 ^ 1'b0 ;
  assign n1008 = x247 & ~n624 ;
  assign n1011 = n1010 ^ n1008 ^ 1'b0 ;
  assign n1006 = x233 & n307 ;
  assign n1007 = ~x38 & n1006 ;
  assign n1012 = n1011 ^ n1007 ^ n428 ;
  assign n1013 = n1012 ^ x129 ^ 1'b0 ;
  assign n1014 = ~n1005 & n1013 ;
  assign n1015 = n1014 ^ n395 ^ x11 ;
  assign n1016 = n1004 | n1015 ;
  assign n1017 = x86 & ~n280 ;
  assign n1018 = n1017 ^ x44 ^ 1'b0 ;
  assign n1019 = ( n293 & n374 ) | ( n293 & n481 ) | ( n374 & n481 ) ;
  assign n1020 = ( ~x28 & n1018 ) | ( ~x28 & n1019 ) | ( n1018 & n1019 ) ;
  assign n1021 = x5 & ~n429 ;
  assign n1022 = n1020 & n1021 ;
  assign n1023 = n1022 ^ n494 ^ n301 ;
  assign n1024 = ~n538 & n752 ;
  assign n1025 = n1024 ^ x239 ^ 1'b0 ;
  assign n1027 = x211 ^ x54 ^ 1'b0 ;
  assign n1028 = n477 & n1027 ;
  assign n1029 = n1028 ^ x178 ^ 1'b0 ;
  assign n1030 = x124 & n1029 ;
  assign n1026 = x204 ^ x192 ^ 1'b0 ;
  assign n1031 = n1030 ^ n1026 ^ 1'b0 ;
  assign n1032 = ( n427 & n1025 ) | ( n427 & ~n1031 ) | ( n1025 & ~n1031 ) ;
  assign n1033 = n291 & n440 ;
  assign n1034 = n1033 ^ n341 ^ 1'b0 ;
  assign n1035 = n478 & n1034 ;
  assign n1036 = n1035 ^ n556 ^ 1'b0 ;
  assign n1037 = n1032 | n1036 ;
  assign n1038 = n350 & ~n1020 ;
  assign n1039 = n704 & n1038 ;
  assign n1040 = ( n488 & n1005 ) | ( n488 & ~n1039 ) | ( n1005 & ~n1039 ) ;
  assign n1041 = ( ~n592 & n852 ) | ( ~n592 & n939 ) | ( n852 & n939 ) ;
  assign n1042 = ( x190 & ~n687 ) | ( x190 & n1041 ) | ( ~n687 & n1041 ) ;
  assign n1044 = ( x69 & ~x151 ) | ( x69 & x204 ) | ( ~x151 & x204 ) ;
  assign n1045 = x168 & n1044 ;
  assign n1043 = n399 ^ n326 ^ n291 ;
  assign n1046 = n1045 ^ n1043 ^ n500 ;
  assign n1047 = n1046 ^ x98 ^ 1'b0 ;
  assign n1048 = ( n287 & n472 ) | ( n287 & n562 ) | ( n472 & n562 ) ;
  assign n1049 = x127 & n1048 ;
  assign n1050 = n733 ^ n337 ^ x85 ;
  assign n1051 = n1050 ^ n466 ^ 1'b0 ;
  assign n1052 = n266 & n1051 ;
  assign n1053 = x174 ^ x30 ^ 1'b0 ;
  assign n1054 = x40 & n1053 ;
  assign n1055 = x202 | n828 ;
  assign n1056 = n1055 ^ n730 ^ n345 ;
  assign n1057 = x27 & n1056 ;
  assign n1058 = ~n530 & n1057 ;
  assign n1061 = n934 ^ n564 ^ 1'b0 ;
  assign n1059 = x188 ^ x150 ^ x6 ;
  assign n1060 = x153 & ~n1059 ;
  assign n1062 = n1061 ^ n1060 ^ 1'b0 ;
  assign n1063 = ( ~n277 & n655 ) | ( ~n277 & n1062 ) | ( n655 & n1062 ) ;
  assign n1064 = ( x32 & ~x174 ) | ( x32 & x206 ) | ( ~x174 & x206 ) ;
  assign n1065 = ( ~n830 & n1034 ) | ( ~n830 & n1064 ) | ( n1034 & n1064 ) ;
  assign n1066 = x243 & n1065 ;
  assign n1067 = n687 & n1066 ;
  assign n1070 = n339 & ~n732 ;
  assign n1071 = n1070 ^ n399 ^ 1'b0 ;
  assign n1072 = n1071 ^ n432 ^ x0 ;
  assign n1068 = n658 ^ n572 ^ n289 ;
  assign n1069 = ( ~x22 & n887 ) | ( ~x22 & n1068 ) | ( n887 & n1068 ) ;
  assign n1073 = n1072 ^ n1069 ^ n776 ;
  assign n1074 = n891 ^ n693 ^ 1'b0 ;
  assign n1075 = x68 & ~n1074 ;
  assign n1076 = n1075 ^ x232 ^ 1'b0 ;
  assign n1077 = ( n521 & n588 ) | ( n521 & ~n1076 ) | ( n588 & ~n1076 ) ;
  assign n1078 = ( x57 & n490 ) | ( x57 & n824 ) | ( n490 & n824 ) ;
  assign n1079 = n501 ^ n412 ^ x178 ;
  assign n1080 = x189 & n1079 ;
  assign n1081 = n1080 ^ n329 ^ 1'b0 ;
  assign n1082 = ~n848 & n1081 ;
  assign n1083 = ~n813 & n1082 ;
  assign n1084 = ( x144 & n456 ) | ( x144 & n617 ) | ( n456 & n617 ) ;
  assign n1085 = n1084 ^ n733 ^ 1'b0 ;
  assign n1086 = x192 & ~n1085 ;
  assign n1087 = n1086 ^ n384 ^ x97 ;
  assign n1088 = ( x113 & n1083 ) | ( x113 & ~n1087 ) | ( n1083 & ~n1087 ) ;
  assign n1089 = ( x78 & ~n973 ) | ( x78 & n1088 ) | ( ~n973 & n1088 ) ;
  assign n1090 = ~n1040 & n1089 ;
  assign n1091 = n1088 & n1090 ;
  assign n1092 = n556 ^ x87 ^ 1'b0 ;
  assign n1093 = n540 & ~n1092 ;
  assign n1096 = n882 ^ n740 ^ x115 ;
  assign n1094 = n307 ^ x95 ^ 1'b0 ;
  assign n1095 = ~n495 & n1094 ;
  assign n1097 = n1096 ^ n1095 ^ x133 ;
  assign n1098 = ( x217 & ~n1093 ) | ( x217 & n1097 ) | ( ~n1093 & n1097 ) ;
  assign n1099 = n301 ^ n285 ^ x224 ;
  assign n1100 = n1099 ^ n1015 ^ x150 ;
  assign n1101 = n704 ^ n296 ^ x172 ;
  assign n1102 = n1101 ^ n460 ^ n295 ;
  assign n1103 = n1102 ^ n391 ^ n283 ;
  assign n1111 = ( x85 & n267 ) | ( x85 & ~n476 ) | ( n267 & ~n476 ) ;
  assign n1112 = n1111 ^ n864 ^ x164 ;
  assign n1113 = ( x130 & n606 ) | ( x130 & ~n1112 ) | ( n606 & ~n1112 ) ;
  assign n1104 = ( n343 & n1003 ) | ( n343 & ~n1012 ) | ( n1003 & ~n1012 ) ;
  assign n1105 = n833 ^ x245 ^ 1'b0 ;
  assign n1106 = n722 ^ x195 ^ 1'b0 ;
  assign n1107 = x95 & n1106 ;
  assign n1108 = n291 & n1107 ;
  assign n1109 = ( ~n364 & n450 ) | ( ~n364 & n1108 ) | ( n450 & n1108 ) ;
  assign n1110 = ( n1104 & n1105 ) | ( n1104 & n1109 ) | ( n1105 & n1109 ) ;
  assign n1114 = n1113 ^ n1110 ^ x124 ;
  assign n1124 = x153 ^ x65 ^ x49 ;
  assign n1117 = x79 & n883 ;
  assign n1118 = n1117 ^ x127 ^ 1'b0 ;
  assign n1120 = n289 & ~n828 ;
  assign n1121 = n1120 ^ n587 ^ 1'b0 ;
  assign n1119 = x79 & ~n280 ;
  assign n1122 = n1121 ^ n1119 ^ 1'b0 ;
  assign n1123 = ( ~x246 & n1118 ) | ( ~x246 & n1122 ) | ( n1118 & n1122 ) ;
  assign n1115 = x105 & n901 ;
  assign n1116 = n1115 ^ n808 ^ 1'b0 ;
  assign n1125 = n1124 ^ n1123 ^ n1116 ;
  assign n1127 = n313 ^ x53 ^ 1'b0 ;
  assign n1128 = n682 & n1127 ;
  assign n1126 = n363 & n1083 ;
  assign n1129 = n1128 ^ n1126 ^ n596 ;
  assign n1130 = ( x142 & ~n358 ) | ( x142 & n566 ) | ( ~n358 & n566 ) ;
  assign n1131 = ( ~n326 & n622 ) | ( ~n326 & n1130 ) | ( n622 & n1130 ) ;
  assign n1132 = ~n1129 & n1131 ;
  assign n1133 = n1132 ^ n412 ^ 1'b0 ;
  assign n1136 = n895 ^ n466 ^ x151 ;
  assign n1137 = ( x44 & ~n1034 ) | ( x44 & n1136 ) | ( ~n1034 & n1136 ) ;
  assign n1134 = n748 ^ n441 ^ 1'b0 ;
  assign n1135 = x89 & n1134 ;
  assign n1138 = n1137 ^ n1135 ^ 1'b0 ;
  assign n1139 = ( ~x126 & n561 ) | ( ~x126 & n716 ) | ( n561 & n716 ) ;
  assign n1140 = n1139 ^ n384 ^ 1'b0 ;
  assign n1141 = n775 ^ n363 ^ n275 ;
  assign n1142 = n1141 ^ x249 ^ 1'b0 ;
  assign n1143 = n297 | n1142 ;
  assign n1144 = n350 & ~n1075 ;
  assign n1145 = ( n297 & ~n1143 ) | ( n297 & n1144 ) | ( ~n1143 & n1144 ) ;
  assign n1146 = n1140 & n1145 ;
  assign n1147 = n617 ^ x95 ^ 1'b0 ;
  assign n1148 = ~n553 & n1147 ;
  assign n1149 = ~n745 & n1148 ;
  assign n1150 = n556 & n1149 ;
  assign n1151 = n1146 & ~n1150 ;
  assign n1152 = ~n1138 & n1151 ;
  assign n1157 = x94 & ~n1079 ;
  assign n1155 = ( x82 & ~x119 ) | ( x82 & x214 ) | ( ~x119 & x214 ) ;
  assign n1153 = n304 ^ x180 ^ x153 ;
  assign n1154 = ( ~x17 & n282 ) | ( ~x17 & n1153 ) | ( n282 & n1153 ) ;
  assign n1156 = n1155 ^ n1154 ^ 1'b0 ;
  assign n1158 = n1157 ^ n1156 ^ n551 ;
  assign n1161 = x142 ^ x1 ^ 1'b0 ;
  assign n1159 = n678 ^ n391 ^ 1'b0 ;
  assign n1160 = ~n1121 & n1159 ;
  assign n1162 = n1161 ^ n1160 ^ n636 ;
  assign n1164 = ( x36 & n429 ) | ( x36 & n1011 ) | ( n429 & n1011 ) ;
  assign n1163 = x174 ^ x132 ^ x34 ;
  assign n1165 = n1164 ^ n1163 ^ n265 ;
  assign n1166 = n819 & ~n1165 ;
  assign n1174 = n614 ^ n499 ^ 1'b0 ;
  assign n1175 = n591 & n1174 ;
  assign n1176 = n1175 ^ n350 ^ x251 ;
  assign n1177 = n1176 ^ n664 ^ x93 ;
  assign n1171 = ( x77 & n258 ) | ( x77 & ~n1064 ) | ( n258 & ~n1064 ) ;
  assign n1172 = ( n1022 & ~n1118 ) | ( n1022 & n1171 ) | ( ~n1118 & n1171 ) ;
  assign n1167 = n504 ^ x149 ^ 1'b0 ;
  assign n1168 = x213 & ~n1139 ;
  assign n1169 = n1167 & n1168 ;
  assign n1170 = x113 & ~n1169 ;
  assign n1173 = n1172 ^ n1170 ^ 1'b0 ;
  assign n1178 = n1177 ^ n1173 ^ 1'b0 ;
  assign n1179 = n441 & n1178 ;
  assign n1180 = n1087 ^ n830 ^ x51 ;
  assign n1182 = x78 & x120 ;
  assign n1183 = ( ~n684 & n1140 ) | ( ~n684 & n1182 ) | ( n1140 & n1182 ) ;
  assign n1181 = x62 & n1014 ;
  assign n1184 = n1183 ^ n1181 ^ 1'b0 ;
  assign n1185 = n438 & n563 ;
  assign n1186 = n748 | n1185 ;
  assign n1187 = ( n681 & n740 ) | ( n681 & ~n810 ) | ( n740 & ~n810 ) ;
  assign n1188 = x122 & n339 ;
  assign n1189 = ( n308 & ~n1187 ) | ( n308 & n1188 ) | ( ~n1187 & n1188 ) ;
  assign n1190 = ( n1184 & ~n1186 ) | ( n1184 & n1189 ) | ( ~n1186 & n1189 ) ;
  assign n1191 = n273 & ~n1180 ;
  assign n1194 = x5 & x41 ;
  assign n1195 = ~n508 & n1194 ;
  assign n1196 = ~n469 & n818 ;
  assign n1197 = ~n1195 & n1196 ;
  assign n1192 = n660 ^ n530 ^ n485 ;
  assign n1193 = n1192 ^ n1036 ^ n662 ;
  assign n1198 = n1197 ^ n1193 ^ n948 ;
  assign n1199 = ( x127 & ~n879 ) | ( x127 & n1198 ) | ( ~n879 & n1198 ) ;
  assign n1202 = n946 ^ n828 ^ 1'b0 ;
  assign n1201 = n1161 ^ x117 ^ 1'b0 ;
  assign n1200 = ( x51 & x100 ) | ( x51 & ~n929 ) | ( x100 & ~n929 ) ;
  assign n1203 = n1202 ^ n1201 ^ n1200 ;
  assign n1204 = n745 ^ x55 ^ 1'b0 ;
  assign n1205 = n264 & ~n1204 ;
  assign n1206 = n618 & n1205 ;
  assign n1207 = x246 & ~n589 ;
  assign n1208 = ~x54 & n1207 ;
  assign n1210 = ~x153 & x214 ;
  assign n1209 = n795 ^ n707 ^ 1'b0 ;
  assign n1211 = n1210 ^ n1209 ^ n428 ;
  assign n1212 = n1010 ^ n435 ^ 1'b0 ;
  assign n1213 = n1211 | n1212 ;
  assign n1214 = ( ~x52 & x157 ) | ( ~x52 & x237 ) | ( x157 & x237 ) ;
  assign n1215 = n1162 ^ x197 ^ 1'b0 ;
  assign n1216 = n1214 & n1215 ;
  assign n1217 = ( x112 & ~n296 ) | ( x112 & n739 ) | ( ~n296 & n739 ) ;
  assign n1218 = ~n1020 & n1217 ;
  assign n1219 = ~x181 & n1218 ;
  assign n1223 = n632 & ~n761 ;
  assign n1224 = n1223 ^ n434 ^ 1'b0 ;
  assign n1221 = n270 & ~n525 ;
  assign n1220 = n337 ^ x252 ^ x189 ;
  assign n1222 = n1221 ^ n1220 ^ x86 ;
  assign n1225 = n1224 ^ n1222 ^ n622 ;
  assign n1226 = n1225 ^ n773 ^ 1'b0 ;
  assign n1227 = ( n638 & ~n876 ) | ( n638 & n896 ) | ( ~n876 & n896 ) ;
  assign n1233 = n260 ^ x237 ^ x63 ;
  assign n1234 = x216 ^ x196 ^ 1'b0 ;
  assign n1235 = n887 & n1234 ;
  assign n1236 = ( x250 & n1233 ) | ( x250 & n1235 ) | ( n1233 & n1235 ) ;
  assign n1230 = n910 ^ x141 ^ x27 ;
  assign n1231 = ( x53 & n344 ) | ( x53 & n1230 ) | ( n344 & n1230 ) ;
  assign n1232 = ( n410 & ~n579 ) | ( n410 & n1231 ) | ( ~n579 & n1231 ) ;
  assign n1228 = n1210 ^ n778 ^ 1'b0 ;
  assign n1229 = n1228 ^ n962 ^ x136 ;
  assign n1237 = n1236 ^ n1232 ^ n1229 ;
  assign n1238 = n352 & ~n1163 ;
  assign n1239 = n1238 ^ n350 ^ 1'b0 ;
  assign n1240 = n903 | n1239 ;
  assign n1241 = n997 | n1240 ;
  assign n1242 = n475 ^ x179 ^ 1'b0 ;
  assign n1243 = x119 & n1242 ;
  assign n1244 = x118 & ~n559 ;
  assign n1245 = ~n724 & n1244 ;
  assign n1246 = ( n632 & n1243 ) | ( n632 & n1245 ) | ( n1243 & n1245 ) ;
  assign n1247 = n614 ^ n504 ^ 1'b0 ;
  assign n1248 = n1153 & ~n1247 ;
  assign n1249 = n1248 ^ n745 ^ n399 ;
  assign n1250 = n1249 ^ n891 ^ x36 ;
  assign n1255 = n643 | n1056 ;
  assign n1256 = x76 ^ x41 ^ 1'b0 ;
  assign n1257 = x27 & n1256 ;
  assign n1258 = n630 ^ n353 ^ x167 ;
  assign n1259 = n286 ^ x103 ^ 1'b0 ;
  assign n1260 = n1258 | n1259 ;
  assign n1261 = n882 & ~n1260 ;
  assign n1262 = ( n439 & n561 ) | ( n439 & ~n1261 ) | ( n561 & ~n1261 ) ;
  assign n1263 = n1262 ^ x81 ^ 1'b0 ;
  assign n1264 = x169 & n1263 ;
  assign n1268 = ( x234 & ~n739 ) | ( x234 & n896 ) | ( ~n739 & n896 ) ;
  assign n1265 = n460 & n707 ;
  assign n1266 = ~x183 & n1265 ;
  assign n1267 = ( x247 & ~n890 ) | ( x247 & n1266 ) | ( ~n890 & n1266 ) ;
  assign n1269 = n1268 ^ n1267 ^ 1'b0 ;
  assign n1270 = ~n957 & n1269 ;
  assign n1271 = ( n1257 & ~n1264 ) | ( n1257 & n1270 ) | ( ~n1264 & n1270 ) ;
  assign n1272 = ( n807 & ~n1255 ) | ( n807 & n1271 ) | ( ~n1255 & n1271 ) ;
  assign n1251 = ( ~x36 & x45 ) | ( ~x36 & n293 ) | ( x45 & n293 ) ;
  assign n1252 = n840 & ~n1251 ;
  assign n1253 = ~x196 & n1252 ;
  assign n1254 = ( x168 & n984 ) | ( x168 & n1253 ) | ( n984 & n1253 ) ;
  assign n1273 = n1272 ^ n1254 ^ 1'b0 ;
  assign n1274 = n1250 | n1273 ;
  assign n1275 = ( n615 & n1103 ) | ( n615 & n1107 ) | ( n1103 & n1107 ) ;
  assign n1276 = x183 & n941 ;
  assign n1277 = ( n684 & n885 ) | ( n684 & n1276 ) | ( n885 & n1276 ) ;
  assign n1279 = n516 ^ n291 ^ n256 ;
  assign n1278 = ( ~x245 & n978 ) | ( ~x245 & n1164 ) | ( n978 & n1164 ) ;
  assign n1280 = n1279 ^ n1278 ^ 1'b0 ;
  assign n1281 = n624 ^ n410 ^ x70 ;
  assign n1282 = ( n834 & n1197 ) | ( n834 & ~n1281 ) | ( n1197 & ~n1281 ) ;
  assign n1283 = n570 & ~n1282 ;
  assign n1284 = n1283 ^ n662 ^ 1'b0 ;
  assign n1285 = x201 & ~n642 ;
  assign n1286 = n1285 ^ x50 ^ 1'b0 ;
  assign n1287 = n1110 & ~n1286 ;
  assign n1288 = n1287 ^ n490 ^ 1'b0 ;
  assign n1292 = x167 & x224 ;
  assign n1293 = n1292 ^ x124 ^ 1'b0 ;
  assign n1289 = ( x114 & ~n287 ) | ( x114 & n596 ) | ( ~n287 & n596 ) ;
  assign n1290 = x64 & ~n1289 ;
  assign n1291 = n1290 ^ x193 ^ 1'b0 ;
  assign n1294 = n1293 ^ n1291 ^ x44 ;
  assign n1295 = n587 | n1294 ;
  assign n1296 = ( ~x166 & n533 ) | ( ~x166 & n1295 ) | ( n533 & n1295 ) ;
  assign n1297 = n1296 ^ n1213 ^ n489 ;
  assign n1298 = ~x99 & n1140 ;
  assign n1299 = n1298 ^ x140 ^ 1'b0 ;
  assign n1300 = x65 | n1299 ;
  assign n1301 = n412 & n501 ;
  assign n1303 = n1268 ^ n1018 ^ n770 ;
  assign n1302 = n305 | n323 ;
  assign n1304 = n1303 ^ n1302 ^ n711 ;
  assign n1306 = ( ~x157 & x242 ) | ( ~x157 & n275 ) | ( x242 & n275 ) ;
  assign n1307 = ( n428 & ~n788 ) | ( n428 & n1306 ) | ( ~n788 & n1306 ) ;
  assign n1305 = ( x223 & n384 ) | ( x223 & ~n1270 ) | ( n384 & ~n1270 ) ;
  assign n1308 = n1307 ^ n1305 ^ 1'b0 ;
  assign n1309 = ( n393 & ~n472 ) | ( n393 & n981 ) | ( ~n472 & n981 ) ;
  assign n1310 = ~x64 & n693 ;
  assign n1311 = ( x252 & n770 ) | ( x252 & ~n1310 ) | ( n770 & ~n1310 ) ;
  assign n1312 = n1309 & n1311 ;
  assign n1313 = n555 | n692 ;
  assign n1314 = ~n894 & n1313 ;
  assign n1315 = n1314 ^ n1197 ^ 1'b0 ;
  assign n1316 = x155 & n1315 ;
  assign n1317 = n1316 ^ n562 ^ 1'b0 ;
  assign n1318 = n657 ^ x127 ^ 1'b0 ;
  assign n1319 = n662 ^ n647 ^ n428 ;
  assign n1320 = x135 & ~n1319 ;
  assign n1321 = n999 & n1320 ;
  assign n1322 = n1318 & n1321 ;
  assign n1323 = ( x5 & x151 ) | ( x5 & ~n882 ) | ( x151 & ~n882 ) ;
  assign n1324 = n403 & n1323 ;
  assign n1325 = n1324 ^ n573 ^ 1'b0 ;
  assign n1326 = n1122 ^ n796 ^ 1'b0 ;
  assign n1327 = n802 & n1326 ;
  assign n1328 = ~x6 & n1327 ;
  assign n1329 = ( ~x178 & n817 ) | ( ~x178 & n1328 ) | ( n817 & n1328 ) ;
  assign n1330 = ~n335 & n1329 ;
  assign n1331 = ( x57 & ~x207 ) | ( x57 & n1128 ) | ( ~x207 & n1128 ) ;
  assign n1332 = x176 & x227 ;
  assign n1333 = n1332 ^ x149 ^ 1'b0 ;
  assign n1334 = ( x73 & n767 ) | ( x73 & n1333 ) | ( n767 & n1333 ) ;
  assign n1335 = ~n678 & n1334 ;
  assign n1336 = ~n1281 & n1335 ;
  assign n1337 = x161 ^ x82 ^ 1'b0 ;
  assign n1338 = n725 & ~n1337 ;
  assign n1339 = ~x149 & n1338 ;
  assign n1340 = ( n297 & ~n1336 ) | ( n297 & n1339 ) | ( ~n1336 & n1339 ) ;
  assign n1341 = ( ~n738 & n1331 ) | ( ~n738 & n1340 ) | ( n1331 & n1340 ) ;
  assign n1350 = n539 ^ n488 ^ 1'b0 ;
  assign n1351 = ~n745 & n1350 ;
  assign n1349 = x175 & ~n368 ;
  assign n1352 = n1351 ^ n1349 ^ n742 ;
  assign n1344 = ( x121 & n308 ) | ( x121 & ~n333 ) | ( n308 & ~n333 ) ;
  assign n1345 = n344 & ~n1344 ;
  assign n1346 = ~x130 & n1345 ;
  assign n1342 = x126 & x129 ;
  assign n1343 = ~x65 & n1342 ;
  assign n1347 = n1346 ^ n1343 ^ n672 ;
  assign n1348 = ~n652 & n1347 ;
  assign n1353 = n1352 ^ n1348 ^ 1'b0 ;
  assign n1354 = ( x232 & n504 ) | ( x232 & ~n1353 ) | ( n504 & ~n1353 ) ;
  assign n1355 = n1135 ^ n313 ^ x234 ;
  assign n1356 = ( ~n742 & n754 ) | ( ~n742 & n1355 ) | ( n754 & n1355 ) ;
  assign n1357 = ~n933 & n1356 ;
  assign n1358 = ~n385 & n1357 ;
  assign n1359 = ( x222 & ~x244 ) | ( x222 & n370 ) | ( ~x244 & n370 ) ;
  assign n1360 = n673 & ~n1359 ;
  assign n1361 = ~n644 & n1360 ;
  assign n1362 = n1361 ^ n410 ^ 1'b0 ;
  assign n1363 = ( n862 & ~n1358 ) | ( n862 & n1362 ) | ( ~n1358 & n1362 ) ;
  assign n1364 = n1069 ^ n636 ^ n408 ;
  assign n1365 = n1364 ^ x3 ^ 1'b0 ;
  assign n1367 = n1289 ^ n266 ^ x214 ;
  assign n1366 = n1104 ^ n858 ^ n530 ;
  assign n1368 = n1367 ^ n1366 ^ n1036 ;
  assign n1369 = n403 & n426 ;
  assign n1370 = n1369 ^ n435 ^ 1'b0 ;
  assign n1371 = x5 & x83 ;
  assign n1372 = n1370 & n1371 ;
  assign n1373 = ( x191 & ~n914 ) | ( x191 & n1372 ) | ( ~n914 & n1372 ) ;
  assign n1374 = n1195 ^ x222 ^ x153 ;
  assign n1375 = n1374 ^ n783 ^ n617 ;
  assign n1376 = ( ~x99 & n752 ) | ( ~x99 & n1375 ) | ( n752 & n1375 ) ;
  assign n1377 = x76 & ~n270 ;
  assign n1378 = n447 & n1377 ;
  assign n1381 = ~n267 & n335 ;
  assign n1382 = ( ~n492 & n558 ) | ( ~n492 & n1381 ) | ( n558 & n1381 ) ;
  assign n1379 = n874 | n1164 ;
  assign n1380 = n1379 ^ n916 ^ 1'b0 ;
  assign n1383 = n1382 ^ n1380 ^ 1'b0 ;
  assign n1384 = n1378 | n1383 ;
  assign n1385 = n1384 ^ n1253 ^ n489 ;
  assign n1386 = n1183 & n1303 ;
  assign n1387 = n1386 ^ n400 ^ 1'b0 ;
  assign n1388 = n1387 ^ x70 ^ 1'b0 ;
  assign n1392 = n831 & ~n1251 ;
  assign n1393 = ~n620 & n1392 ;
  assign n1390 = n924 ^ x224 ^ x27 ;
  assign n1391 = ( ~x151 & x179 ) | ( ~x151 & n1390 ) | ( x179 & n1390 ) ;
  assign n1394 = n1393 ^ n1391 ^ x165 ;
  assign n1389 = n505 & n1319 ;
  assign n1395 = n1394 ^ n1389 ^ 1'b0 ;
  assign n1396 = ( n1193 & n1388 ) | ( n1193 & ~n1395 ) | ( n1388 & ~n1395 ) ;
  assign n1417 = n662 & ~n1210 ;
  assign n1418 = n1417 ^ n1268 ^ 1'b0 ;
  assign n1419 = ( x238 & n1050 ) | ( x238 & ~n1418 ) | ( n1050 & ~n1418 ) ;
  assign n1420 = ~n480 & n518 ;
  assign n1421 = ~n615 & n1420 ;
  assign n1422 = n1421 ^ n1048 ^ x186 ;
  assign n1423 = ( n1083 & n1419 ) | ( n1083 & n1422 ) | ( n1419 & n1422 ) ;
  assign n1424 = ( n1231 & n1336 ) | ( n1231 & ~n1423 ) | ( n1336 & ~n1423 ) ;
  assign n1406 = x246 ^ x192 ^ 1'b0 ;
  assign n1407 = n463 & n1406 ;
  assign n1411 = ( x18 & n473 ) | ( x18 & n510 ) | ( n473 & n510 ) ;
  assign n1412 = n642 ^ x67 ^ 1'b0 ;
  assign n1413 = n517 | n1412 ;
  assign n1414 = n1411 | n1413 ;
  assign n1408 = n1068 & ~n1183 ;
  assign n1409 = x139 & x243 ;
  assign n1410 = n1408 & n1409 ;
  assign n1415 = n1414 ^ n1410 ^ x49 ;
  assign n1416 = ( ~n913 & n1407 ) | ( ~n913 & n1415 ) | ( n1407 & n1415 ) ;
  assign n1398 = n716 ^ n337 ^ x38 ;
  assign n1399 = n1398 ^ n1171 ^ n349 ;
  assign n1397 = ~n1163 & n1164 ;
  assign n1400 = n1399 ^ n1397 ^ 1'b0 ;
  assign n1401 = n1279 ^ n1019 ^ n499 ;
  assign n1402 = n1401 ^ n438 ^ 1'b0 ;
  assign n1403 = n928 & ~n1402 ;
  assign n1404 = n370 | n1403 ;
  assign n1405 = ( n687 & ~n1400 ) | ( n687 & n1404 ) | ( ~n1400 & n1404 ) ;
  assign n1425 = n1424 ^ n1416 ^ n1405 ;
  assign n1426 = n440 & n895 ;
  assign n1427 = n1426 ^ n672 ^ 1'b0 ;
  assign n1428 = n517 | n1427 ;
  assign n1429 = ( x243 & ~n528 ) | ( x243 & n1233 ) | ( ~n528 & n1233 ) ;
  assign n1430 = ( ~x4 & x41 ) | ( ~x4 & n1429 ) | ( x41 & n1429 ) ;
  assign n1431 = ( x102 & n1407 ) | ( x102 & n1430 ) | ( n1407 & n1430 ) ;
  assign n1432 = ( n573 & ~n1291 ) | ( n573 & n1431 ) | ( ~n1291 & n1431 ) ;
  assign n1433 = ~x43 & n1432 ;
  assign n1434 = n1433 ^ n724 ^ 1'b0 ;
  assign n1435 = n1434 ^ n812 ^ 1'b0 ;
  assign n1436 = x176 & n1435 ;
  assign n1437 = x152 & x203 ;
  assign n1438 = n1437 ^ n885 ^ 1'b0 ;
  assign n1443 = n773 ^ x251 ^ 1'b0 ;
  assign n1444 = n573 | n1443 ;
  assign n1445 = n1444 ^ n587 ^ n466 ;
  assign n1439 = ( x147 & ~n512 ) | ( x147 & n828 ) | ( ~n512 & n828 ) ;
  assign n1440 = n1439 ^ n400 ^ x180 ;
  assign n1441 = x132 & n895 ;
  assign n1442 = ~n1440 & n1441 ;
  assign n1446 = n1445 ^ n1442 ^ x234 ;
  assign n1447 = n1446 ^ n374 ^ 1'b0 ;
  assign n1448 = n547 | n1447 ;
  assign n1449 = ~x169 & x254 ;
  assign n1458 = ( x150 & x196 ) | ( x150 & n414 ) | ( x196 & n414 ) ;
  assign n1452 = n435 & n739 ;
  assign n1459 = x165 & ~n1452 ;
  assign n1460 = ~n1458 & n1459 ;
  assign n1450 = ( x52 & n326 ) | ( x52 & ~n767 ) | ( n326 & ~n767 ) ;
  assign n1451 = n1450 ^ n702 ^ x170 ;
  assign n1453 = x181 & ~n1452 ;
  assign n1454 = n1453 ^ x54 ^ 1'b0 ;
  assign n1455 = ( x64 & n1451 ) | ( x64 & n1454 ) | ( n1451 & n1454 ) ;
  assign n1456 = ~n982 & n1455 ;
  assign n1457 = ~n959 & n1456 ;
  assign n1461 = n1460 ^ n1457 ^ x210 ;
  assign n1462 = ( x173 & n785 ) | ( x173 & ~n896 ) | ( n785 & ~n896 ) ;
  assign n1463 = ~x86 & n663 ;
  assign n1464 = n1463 ^ n647 ^ 1'b0 ;
  assign n1465 = n1462 & ~n1464 ;
  assign n1466 = n1465 ^ n1128 ^ n937 ;
  assign n1467 = n1466 ^ n561 ^ 1'b0 ;
  assign n1468 = n1416 & n1467 ;
  assign n1469 = n771 ^ n723 ^ n644 ;
  assign n1470 = ( ~x78 & n333 ) | ( ~x78 & n697 ) | ( n333 & n697 ) ;
  assign n1471 = n1470 ^ n343 ^ 1'b0 ;
  assign n1472 = n1046 | n1471 ;
  assign n1473 = n1014 & n1276 ;
  assign n1474 = n1137 ^ n327 ^ 1'b0 ;
  assign n1475 = ( n344 & n654 ) | ( n344 & n1039 ) | ( n654 & n1039 ) ;
  assign n1476 = n506 ^ x79 ^ x27 ;
  assign n1477 = n930 ^ n500 ^ 1'b0 ;
  assign n1478 = ~n1298 & n1477 ;
  assign n1479 = ~x71 & n256 ;
  assign n1480 = n1230 ^ x240 ^ 1'b0 ;
  assign n1481 = n1479 & ~n1480 ;
  assign n1482 = ( n312 & n1478 ) | ( n312 & ~n1481 ) | ( n1478 & ~n1481 ) ;
  assign n1483 = ~n1476 & n1482 ;
  assign n1484 = n1475 & n1483 ;
  assign n1485 = x248 ^ x154 ^ x120 ;
  assign n1486 = n1183 & n1378 ;
  assign n1487 = n1485 | n1486 ;
  assign n1488 = x61 & ~n1487 ;
  assign n1489 = n1488 ^ n701 ^ 1'b0 ;
  assign n1490 = n1258 | n1489 ;
  assign n1491 = n1490 ^ n422 ^ 1'b0 ;
  assign n1492 = x25 & n785 ;
  assign n1493 = n983 ^ x95 ^ 1'b0 ;
  assign n1494 = x40 & ~n1493 ;
  assign n1495 = n1494 ^ n1275 ^ n564 ;
  assign n1496 = n1495 ^ x251 ^ 1'b0 ;
  assign n1497 = x167 & n1496 ;
  assign n1498 = x223 & n385 ;
  assign n1499 = n1498 ^ n773 ^ 1'b0 ;
  assign n1500 = ( x210 & n1177 ) | ( x210 & ~n1499 ) | ( n1177 & ~n1499 ) ;
  assign n1501 = x157 & ~n1185 ;
  assign n1502 = ~n671 & n1501 ;
  assign n1504 = ~n324 & n1236 ;
  assign n1503 = x50 & ~n573 ;
  assign n1505 = n1504 ^ n1503 ^ 1'b0 ;
  assign n1506 = n1505 ^ n1254 ^ n1064 ;
  assign n1507 = ( n1500 & ~n1502 ) | ( n1500 & n1506 ) | ( ~n1502 & n1506 ) ;
  assign n1508 = n1257 ^ n772 ^ n735 ;
  assign n1509 = ~n573 & n1508 ;
  assign n1510 = ~x89 & n1509 ;
  assign n1511 = n1420 ^ n926 ^ x85 ;
  assign n1512 = n1065 ^ n469 ^ n304 ;
  assign n1513 = n1512 ^ n902 ^ 1'b0 ;
  assign n1514 = n910 & n1326 ;
  assign n1515 = ~x102 & n1514 ;
  assign n1516 = n1485 ^ n965 ^ 1'b0 ;
  assign n1517 = ~n1515 & n1516 ;
  assign n1518 = n1517 ^ n397 ^ 1'b0 ;
  assign n1524 = ( x96 & n940 ) | ( x96 & n1398 ) | ( n940 & n1398 ) ;
  assign n1525 = n1524 ^ n1137 ^ n551 ;
  assign n1519 = n346 & n1163 ;
  assign n1520 = n323 & n474 ;
  assign n1521 = n1519 & n1520 ;
  assign n1522 = n885 ^ x108 ^ 1'b0 ;
  assign n1523 = ~n1521 & n1522 ;
  assign n1526 = n1525 ^ n1523 ^ n882 ;
  assign n1527 = n1526 ^ n1011 ^ n304 ;
  assign n1528 = ( n267 & n772 ) | ( n267 & ~n1439 ) | ( n772 & ~n1439 ) ;
  assign n1530 = ( n929 & n1030 ) | ( n929 & ~n1311 ) | ( n1030 & ~n1311 ) ;
  assign n1529 = x81 & n961 ;
  assign n1531 = n1530 ^ n1529 ^ 1'b0 ;
  assign n1532 = n1275 ^ n510 ^ 1'b0 ;
  assign n1533 = n1075 & ~n1532 ;
  assign n1534 = n1533 ^ n1003 ^ 1'b0 ;
  assign n1539 = n351 | n1298 ;
  assign n1540 = n1071 | n1539 ;
  assign n1535 = n344 & ~n1230 ;
  assign n1536 = n1535 ^ n675 ^ 1'b0 ;
  assign n1537 = ( ~n615 & n675 ) | ( ~n615 & n1536 ) | ( n675 & n1536 ) ;
  assign n1538 = n1537 ^ x130 ^ x81 ;
  assign n1541 = n1540 ^ n1538 ^ 1'b0 ;
  assign n1542 = x178 & ~n1541 ;
  assign n1543 = n389 | n1072 ;
  assign n1544 = n458 ^ n368 ^ 1'b0 ;
  assign n1545 = ( x223 & n364 ) | ( x223 & n1544 ) | ( n364 & n1544 ) ;
  assign n1546 = n1543 | n1545 ;
  assign n1547 = n1352 ^ n751 ^ x186 ;
  assign n1548 = n1139 & n1547 ;
  assign n1549 = n1548 ^ n1166 ^ x186 ;
  assign n1550 = n1352 ^ n1036 ^ 1'b0 ;
  assign n1551 = ( x141 & n270 ) | ( x141 & ~n1550 ) | ( n270 & ~n1550 ) ;
  assign n1552 = n426 ^ x95 ^ 1'b0 ;
  assign n1553 = n1551 & n1552 ;
  assign n1554 = n678 ^ x64 ^ 1'b0 ;
  assign n1555 = n800 & ~n1554 ;
  assign n1556 = ( x125 & n497 ) | ( x125 & ~n1555 ) | ( n497 & ~n1555 ) ;
  assign n1557 = n1300 ^ n683 ^ 1'b0 ;
  assign n1560 = x115 & n582 ;
  assign n1561 = ( n276 & ~n481 ) | ( n276 & n1560 ) | ( ~n481 & n1560 ) ;
  assign n1558 = x51 & n1492 ;
  assign n1559 = n885 & ~n1558 ;
  assign n1562 = n1561 ^ n1559 ^ 1'b0 ;
  assign n1563 = n1296 ^ n569 ^ 1'b0 ;
  assign n1564 = ( n271 & ~n580 ) | ( n271 & n1563 ) | ( ~n580 & n1563 ) ;
  assign n1577 = n610 | n1177 ;
  assign n1578 = n1577 ^ n307 ^ 1'b0 ;
  assign n1579 = n849 & n1087 ;
  assign n1580 = ~n1578 & n1579 ;
  assign n1567 = ( x58 & n297 ) | ( x58 & n488 ) | ( n297 & n488 ) ;
  assign n1568 = x120 & ~n639 ;
  assign n1569 = n1568 ^ x40 ^ 1'b0 ;
  assign n1570 = ~n1567 & n1569 ;
  assign n1565 = ~n672 & n1064 ;
  assign n1566 = n1565 ^ n403 ^ 1'b0 ;
  assign n1571 = n1570 ^ n1566 ^ 1'b0 ;
  assign n1572 = ~n472 & n1571 ;
  assign n1573 = x21 & ~n1572 ;
  assign n1574 = ~x127 & x182 ;
  assign n1575 = ( ~x129 & n943 ) | ( ~x129 & n1574 ) | ( n943 & n1574 ) ;
  assign n1576 = n1573 | n1575 ;
  assign n1581 = n1580 ^ n1576 ^ 1'b0 ;
  assign n1582 = ( n1010 & ~n1180 ) | ( n1010 & n1581 ) | ( ~n1180 & n1581 ) ;
  assign n1583 = x16 & ~n954 ;
  assign n1587 = n1452 ^ n1124 ^ n494 ;
  assign n1584 = x124 & n897 ;
  assign n1585 = ( n911 & ~n1329 ) | ( n911 & n1584 ) | ( ~n1329 & n1584 ) ;
  assign n1586 = x133 & ~n1585 ;
  assign n1588 = n1587 ^ n1586 ^ 1'b0 ;
  assign n1589 = n822 ^ n483 ^ n271 ;
  assign n1590 = ( n511 & n758 ) | ( n511 & ~n1589 ) | ( n758 & ~n1589 ) ;
  assign n1603 = ( ~x2 & x18 ) | ( ~x2 & n297 ) | ( x18 & n297 ) ;
  assign n1602 = ( ~x169 & n882 ) | ( ~x169 & n946 ) | ( n882 & n946 ) ;
  assign n1604 = n1603 ^ n1602 ^ n1349 ;
  assign n1605 = n1228 & ~n1604 ;
  assign n1606 = ~x72 & n1605 ;
  assign n1607 = n1478 ^ x13 ^ 1'b0 ;
  assign n1608 = ~n1606 & n1607 ;
  assign n1591 = x166 & x194 ;
  assign n1592 = ~n930 & n1591 ;
  assign n1593 = ( x93 & ~n678 ) | ( x93 & n1592 ) | ( ~n678 & n1592 ) ;
  assign n1594 = ~n351 & n617 ;
  assign n1595 = n1594 ^ n1050 ^ 1'b0 ;
  assign n1596 = n866 & ~n1359 ;
  assign n1597 = ~n1595 & n1596 ;
  assign n1598 = x227 & ~n1481 ;
  assign n1599 = ( x243 & n1597 ) | ( x243 & ~n1598 ) | ( n1597 & ~n1598 ) ;
  assign n1600 = ( n766 & n1478 ) | ( n766 & ~n1599 ) | ( n1478 & ~n1599 ) ;
  assign n1601 = n1593 & n1600 ;
  assign n1609 = n1608 ^ n1601 ^ 1'b0 ;
  assign n1610 = ( x142 & ~n816 ) | ( x142 & n917 ) | ( ~n816 & n917 ) ;
  assign n1611 = x220 & n530 ;
  assign n1612 = ( n540 & n1282 ) | ( n540 & n1611 ) | ( n1282 & n1611 ) ;
  assign n1619 = n1430 ^ n1351 ^ 1'b0 ;
  assign n1620 = n363 & ~n1619 ;
  assign n1621 = ( ~n303 & n632 ) | ( ~n303 & n1343 ) | ( n632 & n1343 ) ;
  assign n1622 = ( n627 & n1620 ) | ( n627 & ~n1621 ) | ( n1620 & ~n1621 ) ;
  assign n1613 = x71 & x131 ;
  assign n1614 = n1613 ^ x195 ^ 1'b0 ;
  assign n1615 = x187 & ~n1614 ;
  assign n1616 = n317 & n1615 ;
  assign n1617 = ( x63 & n311 ) | ( x63 & ~n1616 ) | ( n311 & ~n1616 ) ;
  assign n1618 = n1617 ^ x34 ^ 1'b0 ;
  assign n1623 = n1622 ^ n1618 ^ 1'b0 ;
  assign n1624 = ( x17 & n303 ) | ( x17 & ~n573 ) | ( n303 & ~n573 ) ;
  assign n1625 = n1624 ^ n588 ^ n512 ;
  assign n1626 = n1625 ^ n1219 ^ n1213 ;
  assign n1627 = n1599 ^ n1534 ^ x216 ;
  assign n1628 = ( x246 & ~n770 ) | ( x246 & n1343 ) | ( ~n770 & n1343 ) ;
  assign n1630 = n1398 ^ n724 ^ n638 ;
  assign n1629 = ( n462 & ~n819 ) | ( n462 & n1308 ) | ( ~n819 & n1308 ) ;
  assign n1631 = n1630 ^ n1629 ^ n868 ;
  assign n1634 = n1364 ^ n851 ^ n511 ;
  assign n1632 = ( n673 & ~n735 ) | ( n673 & n938 ) | ( ~n735 & n938 ) ;
  assign n1633 = n1632 ^ n911 ^ x103 ;
  assign n1635 = n1634 ^ n1633 ^ n1280 ;
  assign n1636 = n988 ^ n891 ^ n632 ;
  assign n1637 = ( x194 & n856 ) | ( x194 & ~n1636 ) | ( n856 & ~n1636 ) ;
  assign n1638 = n1637 ^ n841 ^ n501 ;
  assign n1639 = n1638 ^ n384 ^ 1'b0 ;
  assign n1640 = n1267 ^ n1251 ^ x31 ;
  assign n1641 = x45 & n1640 ;
  assign n1642 = n1641 ^ x153 ^ 1'b0 ;
  assign n1643 = ( x86 & n981 ) | ( x86 & n1642 ) | ( n981 & n1642 ) ;
  assign n1646 = ( x128 & x153 ) | ( x128 & ~n331 ) | ( x153 & ~n331 ) ;
  assign n1644 = ( n353 & ~n589 ) | ( n353 & n1048 ) | ( ~n589 & n1048 ) ;
  assign n1645 = ( n386 & ~n567 ) | ( n386 & n1644 ) | ( ~n567 & n1644 ) ;
  assign n1647 = n1646 ^ n1645 ^ x163 ;
  assign n1649 = n573 ^ x131 ^ x26 ;
  assign n1650 = n745 | n1649 ;
  assign n1648 = n687 ^ n445 ^ n342 ;
  assign n1651 = n1650 ^ n1648 ^ x118 ;
  assign n1653 = ( n478 & n1044 ) | ( n478 & n1124 ) | ( n1044 & n1124 ) ;
  assign n1654 = n1653 ^ n526 ^ 1'b0 ;
  assign n1655 = n545 & n1654 ;
  assign n1652 = ( n1130 & ~n1430 ) | ( n1130 & n1548 ) | ( ~n1430 & n1548 ) ;
  assign n1656 = n1655 ^ n1652 ^ 1'b0 ;
  assign n1663 = x4 & ~n525 ;
  assign n1664 = n1343 & n1663 ;
  assign n1661 = n909 & ~n1445 ;
  assign n1662 = n1661 ^ x209 ^ 1'b0 ;
  assign n1665 = n1664 ^ n1662 ^ n499 ;
  assign n1657 = ( ~x40 & n530 ) | ( ~x40 & n636 ) | ( n530 & n636 ) ;
  assign n1658 = n1657 ^ n1544 ^ 1'b0 ;
  assign n1659 = x77 & n1658 ;
  assign n1660 = ~n697 & n1659 ;
  assign n1666 = n1665 ^ n1660 ^ 1'b0 ;
  assign n1667 = ( x26 & n778 ) | ( x26 & n1384 ) | ( n778 & n1384 ) ;
  assign n1668 = n1667 ^ n683 ^ n257 ;
  assign n1671 = n1390 ^ n1267 ^ n935 ;
  assign n1669 = ( x57 & ~x199 ) | ( x57 & n381 ) | ( ~x199 & n381 ) ;
  assign n1670 = n1669 ^ n498 ^ 1'b0 ;
  assign n1672 = n1671 ^ n1670 ^ n610 ;
  assign n1673 = n563 ^ x17 ^ 1'b0 ;
  assign n1674 = x36 & ~n1673 ;
  assign n1675 = n1306 & n1674 ;
  assign n1676 = n1672 & ~n1675 ;
  assign n1677 = ( ~n910 & n1011 ) | ( ~n910 & n1505 ) | ( n1011 & n1505 ) ;
  assign n1678 = x154 & n1677 ;
  assign n1682 = n759 ^ n489 ^ x218 ;
  assign n1679 = n487 | n716 ;
  assign n1680 = ( ~x164 & n840 ) | ( ~x164 & n1659 ) | ( n840 & n1659 ) ;
  assign n1681 = ( n483 & n1679 ) | ( n483 & ~n1680 ) | ( n1679 & ~n1680 ) ;
  assign n1683 = n1682 ^ n1681 ^ n262 ;
  assign n1684 = n719 & n835 ;
  assign n1685 = n1440 ^ n1429 ^ 1'b0 ;
  assign n1686 = n633 ^ n596 ^ 1'b0 ;
  assign n1687 = ~n1685 & n1686 ;
  assign n1688 = ~n1684 & n1687 ;
  assign n1689 = x150 & ~n768 ;
  assign n1690 = n983 | n1415 ;
  assign n1691 = n1087 ^ x254 ^ x96 ;
  assign n1692 = n1691 ^ n387 ^ n265 ;
  assign n1693 = n257 & ~n297 ;
  assign n1694 = ( n342 & n554 ) | ( n342 & ~n1693 ) | ( n554 & ~n1693 ) ;
  assign n1695 = n698 & n1694 ;
  assign n1696 = n1695 ^ n303 ^ 1'b0 ;
  assign n1697 = n1696 ^ n322 ^ 1'b0 ;
  assign n1698 = n483 ^ x142 ^ 1'b0 ;
  assign n1699 = ~n922 & n1698 ;
  assign n1700 = ( x150 & n380 ) | ( x150 & n1182 ) | ( n380 & n1182 ) ;
  assign n1701 = ( n778 & n1373 ) | ( n778 & n1700 ) | ( n1373 & n1700 ) ;
  assign n1702 = ( ~n716 & n1699 ) | ( ~n716 & n1701 ) | ( n1699 & n1701 ) ;
  assign n1706 = ~n306 & n1108 ;
  assign n1703 = n1420 ^ n1351 ^ 1'b0 ;
  assign n1704 = n1703 ^ n1302 ^ 1'b0 ;
  assign n1705 = n1403 & ~n1704 ;
  assign n1707 = n1706 ^ n1705 ^ 1'b0 ;
  assign n1708 = n1343 | n1707 ;
  assign n1709 = ( x120 & x209 ) | ( x120 & n610 ) | ( x209 & n610 ) ;
  assign n1710 = n1709 ^ x106 ^ 1'b0 ;
  assign n1711 = n933 & n1042 ;
  assign n1712 = n1711 ^ x159 ^ 1'b0 ;
  assign n1713 = n646 ^ x109 ^ 1'b0 ;
  assign n1714 = n1713 ^ n730 ^ x115 ;
  assign n1715 = n1401 ^ n512 ^ 1'b0 ;
  assign n1716 = n1714 | n1715 ;
  assign n1717 = ( n1710 & ~n1712 ) | ( n1710 & n1716 ) | ( ~n1712 & n1716 ) ;
  assign n1718 = n1169 | n1343 ;
  assign n1719 = n1718 ^ n1267 ^ 1'b0 ;
  assign n1720 = n1625 & ~n1719 ;
  assign n1721 = ~n1670 & n1720 ;
  assign n1722 = n1154 ^ n335 ^ x127 ;
  assign n1723 = n1722 ^ n831 ^ n627 ;
  assign n1724 = n1723 ^ n1016 ^ n589 ;
  assign n1725 = x254 & ~n304 ;
  assign n1726 = ~n555 & n1725 ;
  assign n1727 = n1726 ^ x20 ^ 1'b0 ;
  assign n1728 = n381 & ~n1727 ;
  assign n1729 = n1180 ^ n1010 ^ 1'b0 ;
  assign n1730 = ~n1728 & n1729 ;
  assign n1731 = n1279 ^ n1251 ^ n463 ;
  assign n1732 = n1731 ^ n1179 ^ n1133 ;
  assign n1733 = x118 & ~n937 ;
  assign n1734 = n1733 ^ n1370 ^ n1260 ;
  assign n1736 = x241 ^ x193 ^ x87 ;
  assign n1735 = x60 & ~n778 ;
  assign n1737 = n1736 ^ n1735 ^ 1'b0 ;
  assign n1738 = ( x221 & n1032 ) | ( x221 & ~n1737 ) | ( n1032 & ~n1737 ) ;
  assign n1739 = ( n885 & n1734 ) | ( n885 & n1738 ) | ( n1734 & n1738 ) ;
  assign n1743 = n1374 ^ n366 ^ x53 ;
  assign n1744 = n1679 ^ n585 ^ 1'b0 ;
  assign n1745 = n1743 & ~n1744 ;
  assign n1742 = x23 & ~n1101 ;
  assign n1746 = n1745 ^ n1742 ^ 1'b0 ;
  assign n1740 = n474 ^ n339 ^ n256 ;
  assign n1741 = n1141 | n1740 ;
  assign n1747 = n1746 ^ n1741 ^ 1'b0 ;
  assign n1748 = n438 ^ n345 ^ 1'b0 ;
  assign n1749 = ( ~n376 & n541 ) | ( ~n376 & n687 ) | ( n541 & n687 ) ;
  assign n1750 = n1107 & ~n1749 ;
  assign n1751 = ~n506 & n1750 ;
  assign n1752 = n1041 | n1751 ;
  assign n1753 = n1665 & ~n1752 ;
  assign n1754 = n513 | n1753 ;
  assign n1755 = n948 ^ n685 ^ n586 ;
  assign n1756 = ( ~x142 & x210 ) | ( ~x142 & n341 ) | ( x210 & n341 ) ;
  assign n1757 = n1280 ^ n1145 ^ 1'b0 ;
  assign n1758 = ~n1756 & n1757 ;
  assign n1759 = n1758 ^ n1182 ^ n551 ;
  assign n1760 = n1759 ^ n924 ^ 1'b0 ;
  assign n1761 = n1760 ^ n1393 ^ 1'b0 ;
  assign n1762 = ~n707 & n831 ;
  assign n1763 = n981 & n1762 ;
  assign n1767 = ~n600 & n934 ;
  assign n1764 = n1718 ^ n600 ^ 1'b0 ;
  assign n1765 = n670 & n1764 ;
  assign n1766 = n864 & n1765 ;
  assign n1768 = n1767 ^ n1766 ^ 1'b0 ;
  assign n1769 = ( x63 & ~n477 ) | ( x63 & n1401 ) | ( ~n477 & n1401 ) ;
  assign n1770 = n1769 ^ n1731 ^ n695 ;
  assign n1771 = ( n270 & ~n785 ) | ( n270 & n1528 ) | ( ~n785 & n1528 ) ;
  assign n1772 = n1770 & n1771 ;
  assign n1775 = n1657 ^ n1444 ^ n576 ;
  assign n1773 = n692 & n922 ;
  assign n1774 = n1505 & ~n1773 ;
  assign n1776 = n1775 ^ n1774 ^ 1'b0 ;
  assign n1777 = x218 | n732 ;
  assign n1778 = x8 & ~n1777 ;
  assign n1779 = n1778 ^ n1065 ^ 1'b0 ;
  assign n1788 = n768 ^ n325 ^ 1'b0 ;
  assign n1789 = n1202 | n1788 ;
  assign n1790 = n1789 ^ n732 ^ n525 ;
  assign n1782 = x190 & ~n549 ;
  assign n1783 = n678 & n1782 ;
  assign n1784 = n1783 ^ n887 ^ 1'b0 ;
  assign n1785 = n1784 ^ n871 ^ n474 ;
  assign n1780 = ( x68 & ~x85 ) | ( x68 & n297 ) | ( ~x85 & n297 ) ;
  assign n1781 = n1222 & ~n1780 ;
  assign n1786 = n1785 ^ n1781 ^ x28 ;
  assign n1787 = ( x254 & n606 ) | ( x254 & ~n1786 ) | ( n606 & ~n1786 ) ;
  assign n1791 = n1790 ^ n1787 ^ n946 ;
  assign n1792 = x169 ^ x102 ^ x59 ;
  assign n1793 = ( n630 & n1113 ) | ( n630 & ~n1792 ) | ( n1113 & ~n1792 ) ;
  assign n1794 = ( x180 & n640 ) | ( x180 & n696 ) | ( n640 & n696 ) ;
  assign n1795 = ~x13 & n326 ;
  assign n1796 = n1795 ^ x127 ^ 1'b0 ;
  assign n1797 = ( x71 & n1794 ) | ( x71 & n1796 ) | ( n1794 & n1796 ) ;
  assign n1798 = n1797 ^ n355 ^ x105 ;
  assign n1799 = ( n1136 & ~n1489 ) | ( n1136 & n1697 ) | ( ~n1489 & n1697 ) ;
  assign n1800 = n279 | n874 ;
  assign n1801 = x63 & n766 ;
  assign n1802 = ~n859 & n1801 ;
  assign n1803 = ( n335 & n561 ) | ( n335 & ~n1099 ) | ( n561 & ~n1099 ) ;
  assign n1804 = n1617 & ~n1803 ;
  assign n1805 = ~n1802 & n1804 ;
  assign n1806 = n1805 ^ n1531 ^ 1'b0 ;
  assign n1811 = x102 & ~n1359 ;
  assign n1812 = ~x253 & n1811 ;
  assign n1808 = x71 & n489 ;
  assign n1809 = n1808 ^ x18 ^ 1'b0 ;
  assign n1810 = ( n439 & ~n978 ) | ( n439 & n1809 ) | ( ~n978 & n1809 ) ;
  assign n1813 = n1812 ^ n1810 ^ n819 ;
  assign n1814 = ( x119 & ~x161 ) | ( x119 & n380 ) | ( ~x161 & n380 ) ;
  assign n1815 = ( n836 & ~n1451 ) | ( n836 & n1814 ) | ( ~n1451 & n1814 ) ;
  assign n1816 = ( n1311 & ~n1813 ) | ( n1311 & n1815 ) | ( ~n1813 & n1815 ) ;
  assign n1807 = ( n448 & n929 ) | ( n448 & n1044 ) | ( n929 & n1044 ) ;
  assign n1817 = n1816 ^ n1807 ^ 1'b0 ;
  assign n1818 = n1022 | n1817 ;
  assign n1822 = ( ~x219 & n632 ) | ( ~x219 & n1153 ) | ( n632 & n1153 ) ;
  assign n1823 = ~n1336 & n1822 ;
  assign n1821 = ( x199 & ~n511 ) | ( x199 & n1390 ) | ( ~n511 & n1390 ) ;
  assign n1819 = n471 & n664 ;
  assign n1820 = n1819 ^ n595 ^ n283 ;
  assign n1824 = n1823 ^ n1821 ^ n1820 ;
  assign n1825 = n798 ^ n360 ^ n326 ;
  assign n1826 = n1825 ^ n1003 ^ n960 ;
  assign n1827 = n866 & n1826 ;
  assign n1828 = n1213 ^ n422 ^ x90 ;
  assign n1829 = n1828 ^ n1272 ^ n697 ;
  assign n1830 = ( x141 & n1827 ) | ( x141 & ~n1829 ) | ( n1827 & ~n1829 ) ;
  assign n1838 = n1007 ^ n954 ^ x229 ;
  assign n1834 = ( x70 & x164 ) | ( x70 & ~x217 ) | ( x164 & ~x217 ) ;
  assign n1835 = n596 ^ n384 ^ 1'b0 ;
  assign n1836 = n1834 & n1835 ;
  assign n1831 = n1126 ^ n497 ^ n467 ;
  assign n1832 = ( n633 & ~n792 ) | ( n633 & n1831 ) | ( ~n792 & n1831 ) ;
  assign n1833 = ( n598 & n1306 ) | ( n598 & n1832 ) | ( n1306 & n1832 ) ;
  assign n1837 = n1836 ^ n1833 ^ n309 ;
  assign n1839 = n1838 ^ n1837 ^ 1'b0 ;
  assign n1840 = n1839 ^ n1447 ^ 1'b0 ;
  assign n1846 = ( x93 & n387 ) | ( x93 & ~n514 ) | ( n387 & ~n514 ) ;
  assign n1842 = n304 ^ x78 ^ x31 ;
  assign n1841 = ( ~x76 & n388 ) | ( ~x76 & n519 ) | ( n388 & n519 ) ;
  assign n1843 = n1842 ^ n1841 ^ n997 ;
  assign n1844 = n786 & ~n1843 ;
  assign n1845 = n327 & n1844 ;
  assign n1847 = n1846 ^ n1845 ^ 1'b0 ;
  assign n1848 = n797 | n1847 ;
  assign n1849 = ( n818 & n994 ) | ( n818 & n1848 ) | ( n994 & n1848 ) ;
  assign n1850 = n1289 ^ n435 ^ 1'b0 ;
  assign n1851 = n1850 ^ n1505 ^ n1275 ;
  assign n1852 = ~n1669 & n1851 ;
  assign n1853 = n1849 & n1852 ;
  assign n1854 = x170 & n476 ;
  assign n1855 = x143 & n1854 ;
  assign n1856 = ~n947 & n1855 ;
  assign n1860 = n788 ^ x190 ^ 1'b0 ;
  assign n1861 = n892 & ~n1860 ;
  assign n1857 = x69 & x192 ;
  assign n1858 = n780 & n1857 ;
  assign n1859 = ( n258 & ~n505 ) | ( n258 & n1858 ) | ( ~n505 & n1858 ) ;
  assign n1862 = n1861 ^ n1859 ^ n778 ;
  assign n1863 = n1611 ^ n799 ^ n531 ;
  assign n1864 = n671 | n1863 ;
  assign n1865 = ~x189 & n676 ;
  assign n1866 = n1865 ^ n724 ^ 1'b0 ;
  assign n1867 = n910 ^ n729 ^ 1'b0 ;
  assign n1868 = x187 & n1867 ;
  assign n1869 = n1866 & n1868 ;
  assign n1870 = n802 & n1148 ;
  assign n1871 = ~n437 & n1870 ;
  assign n1872 = ~n829 & n1871 ;
  assign n1873 = n1010 | n1872 ;
  assign n1874 = n1614 & ~n1873 ;
  assign n1875 = n1649 ^ x17 ^ 1'b0 ;
  assign n1876 = x69 & n1875 ;
  assign n1877 = ( x213 & x222 ) | ( x213 & n1340 ) | ( x222 & n1340 ) ;
  assign n1878 = n1877 ^ n617 ^ 1'b0 ;
  assign n1879 = ~n789 & n1878 ;
  assign n1880 = ( ~x15 & n448 ) | ( ~x15 & n1879 ) | ( n448 & n1879 ) ;
  assign n1881 = ( n439 & n1876 ) | ( n439 & n1880 ) | ( n1876 & n1880 ) ;
  assign n1882 = ~n732 & n1555 ;
  assign n1883 = n888 & n1882 ;
  assign n1884 = n1505 & ~n1883 ;
  assign n1885 = ( x248 & n1230 ) | ( x248 & n1302 ) | ( n1230 & n1302 ) ;
  assign n1886 = ( n314 & ~n713 ) | ( n314 & n1885 ) | ( ~n713 & n1885 ) ;
  assign n1887 = n1093 ^ n711 ^ n577 ;
  assign n1888 = n1887 ^ n1367 ^ 1'b0 ;
  assign n1889 = ( x42 & x235 ) | ( x42 & ~n1888 ) | ( x235 & ~n1888 ) ;
  assign n1894 = n275 ^ x149 ^ x84 ;
  assign n1893 = n380 & n1088 ;
  assign n1890 = ( x200 & ~x252 ) | ( x200 & n588 ) | ( ~x252 & n588 ) ;
  assign n1891 = ( n618 & n706 ) | ( n618 & ~n1890 ) | ( n706 & ~n1890 ) ;
  assign n1892 = ( n575 & ~n1833 ) | ( n575 & n1891 ) | ( ~n1833 & n1891 ) ;
  assign n1895 = n1894 ^ n1893 ^ n1892 ;
  assign n1896 = n1466 | n1895 ;
  assign n1897 = n1018 ^ x39 ^ 1'b0 ;
  assign n1898 = n1516 ^ n600 ^ 1'b0 ;
  assign n1899 = x89 & ~n1898 ;
  assign n1900 = n1899 ^ n1221 ^ n549 ;
  assign n1901 = n761 | n1485 ;
  assign n1902 = n940 ^ x59 ^ 1'b0 ;
  assign n1903 = n1901 | n1902 ;
  assign n1904 = n788 ^ n521 ^ x186 ;
  assign n1905 = ( n586 & ~n1903 ) | ( n586 & n1904 ) | ( ~n1903 & n1904 ) ;
  assign n1906 = ( n1200 & n1900 ) | ( n1200 & n1905 ) | ( n1900 & n1905 ) ;
  assign n1907 = n701 ^ n582 ^ 1'b0 ;
  assign n1908 = n717 & ~n1907 ;
  assign n1909 = n1153 ^ n528 ^ n300 ;
  assign n1910 = n1909 ^ x150 ^ 1'b0 ;
  assign n1911 = ~n358 & n1910 ;
  assign n1912 = ~x159 & n1911 ;
  assign n1913 = n1211 | n1912 ;
  assign n1914 = n1908 | n1913 ;
  assign n1915 = n1914 ^ n664 ^ n575 ;
  assign n1916 = n1075 & n1447 ;
  assign n1918 = n896 ^ n632 ^ 1'b0 ;
  assign n1917 = n830 & n1011 ;
  assign n1919 = n1918 ^ n1917 ^ 1'b0 ;
  assign n1920 = n1802 ^ n594 ^ x104 ;
  assign n1921 = ( n304 & n485 ) | ( n304 & n1920 ) | ( n485 & n1920 ) ;
  assign n1922 = ( ~n386 & n1466 ) | ( ~n386 & n1547 ) | ( n1466 & n1547 ) ;
  assign n1923 = ( x238 & ~n554 ) | ( x238 & n907 ) | ( ~n554 & n907 ) ;
  assign n1924 = ( n724 & n1164 ) | ( n724 & n1923 ) | ( n1164 & n1923 ) ;
  assign n1925 = x157 & ~n732 ;
  assign n1926 = ~n356 & n1925 ;
  assign n1927 = n464 & n1926 ;
  assign n1928 = n1924 | n1927 ;
  assign n1929 = n1928 ^ x236 ^ 1'b0 ;
  assign n1930 = ( n884 & n1592 ) | ( n884 & n1929 ) | ( n1592 & n1929 ) ;
  assign n1931 = n1930 ^ n351 ^ 1'b0 ;
  assign n1932 = ~n1630 & n1931 ;
  assign n1936 = n1185 ^ x157 ^ 1'b0 ;
  assign n1937 = n866 & ~n1936 ;
  assign n1933 = n1163 ^ n1019 ^ 1'b0 ;
  assign n1934 = n1446 | n1933 ;
  assign n1935 = ( n261 & n1713 ) | ( n261 & n1934 ) | ( n1713 & n1934 ) ;
  assign n1938 = n1937 ^ n1935 ^ n1632 ;
  assign n1939 = x87 & n895 ;
  assign n1940 = n1939 ^ n1567 ^ 1'b0 ;
  assign n1941 = n879 & ~n1940 ;
  assign n1942 = ( n285 & n735 ) | ( n285 & n750 ) | ( n735 & n750 ) ;
  assign n1943 = ( x226 & ~n1387 ) | ( x226 & n1942 ) | ( ~n1387 & n1942 ) ;
  assign n1944 = n1943 ^ n962 ^ 1'b0 ;
  assign n1945 = n1941 & ~n1944 ;
  assign n1946 = n331 & n910 ;
  assign n1947 = n866 & n1946 ;
  assign n1948 = n746 & n1947 ;
  assign n1949 = ( ~x180 & n1196 ) | ( ~x180 & n1318 ) | ( n1196 & n1318 ) ;
  assign n1950 = ( n1432 & ~n1948 ) | ( n1432 & n1949 ) | ( ~n1948 & n1949 ) ;
  assign n1951 = n633 ^ n623 ^ 1'b0 ;
  assign n1952 = ( x21 & ~n327 ) | ( x21 & n1650 ) | ( ~n327 & n1650 ) ;
  assign n1953 = n1910 ^ n513 ^ 1'b0 ;
  assign n1954 = x26 & n1953 ;
  assign n1955 = ~n554 & n1954 ;
  assign n1956 = n1848 ^ n471 ^ 1'b0 ;
  assign n1957 = n1955 | n1956 ;
  assign n1964 = n1743 ^ n1653 ^ 1'b0 ;
  assign n1965 = ~n594 & n1964 ;
  assign n1966 = n1965 ^ n1909 ^ n271 ;
  assign n1958 = ( ~x126 & n1126 ) | ( ~x126 & n1499 ) | ( n1126 & n1499 ) ;
  assign n1959 = n1206 | n1958 ;
  assign n1960 = n1959 ^ x164 ^ 1'b0 ;
  assign n1961 = ( ~x144 & n280 ) | ( ~x144 & n755 ) | ( n280 & n755 ) ;
  assign n1962 = n1237 & ~n1961 ;
  assign n1963 = n1960 & ~n1962 ;
  assign n1967 = n1966 ^ n1963 ^ 1'b0 ;
  assign n1968 = n1046 | n1967 ;
  assign n1971 = n789 ^ n666 ^ n358 ;
  assign n1972 = n1971 ^ n1164 ^ n634 ;
  assign n1969 = n258 ^ x246 ^ 1'b0 ;
  assign n1970 = n1969 ^ x254 ^ x0 ;
  assign n1973 = n1972 ^ n1970 ^ 1'b0 ;
  assign n1974 = ~n1091 & n1973 ;
  assign n1975 = n1946 ^ x114 ^ 1'b0 ;
  assign n1976 = x23 & ~n315 ;
  assign n1977 = n1976 ^ n1030 ^ 1'b0 ;
  assign n1978 = n1570 ^ n666 ^ 1'b0 ;
  assign n1979 = ( n289 & n1977 ) | ( n289 & n1978 ) | ( n1977 & n1978 ) ;
  assign n1980 = n1139 ^ x78 ^ 1'b0 ;
  assign n1981 = ~n828 & n1980 ;
  assign n1982 = ( n495 & n1407 ) | ( n495 & ~n1981 ) | ( n1407 & ~n1981 ) ;
  assign n1983 = x187 & ~n1385 ;
  assign n1984 = ~n1982 & n1983 ;
  assign n1985 = x199 & n1470 ;
  assign n1986 = n414 & ~n1985 ;
  assign n1987 = ~n1175 & n1986 ;
  assign n1988 = ( n617 & n1109 ) | ( n617 & n1987 ) | ( n1109 & n1987 ) ;
  assign n1989 = ( n346 & n1272 ) | ( n346 & ~n1988 ) | ( n1272 & ~n1988 ) ;
  assign n1990 = ( n264 & n950 ) | ( n264 & n955 ) | ( n950 & n955 ) ;
  assign n1991 = n1990 ^ n933 ^ n423 ;
  assign n1992 = n1564 ^ n306 ^ 1'b0 ;
  assign n1993 = ~n1991 & n1992 ;
  assign n1994 = ( x84 & x220 ) | ( x84 & n586 ) | ( x220 & n586 ) ;
  assign n1995 = n297 ^ n283 ^ 1'b0 ;
  assign n1996 = n256 & n1205 ;
  assign n1997 = n1996 ^ n1736 ^ 1'b0 ;
  assign n1998 = n1995 & ~n1997 ;
  assign n1999 = n1998 ^ n622 ^ 1'b0 ;
  assign n2000 = n1343 | n1999 ;
  assign n2001 = n2000 ^ n1300 ^ n1197 ;
  assign n2002 = ( ~n1479 & n1994 ) | ( ~n1479 & n2001 ) | ( n1994 & n2001 ) ;
  assign n2003 = ( x73 & x187 ) | ( x73 & n2002 ) | ( x187 & n2002 ) ;
  assign n2004 = ( n1164 & ~n1257 ) | ( n1164 & n1555 ) | ( ~n1257 & n1555 ) ;
  assign n2005 = n2004 ^ n1101 ^ 1'b0 ;
  assign n2006 = n1261 & n2005 ;
  assign n2007 = n2006 ^ n564 ^ 1'b0 ;
  assign n2008 = x243 ^ x162 ^ x119 ;
  assign n2009 = n959 ^ n268 ^ 1'b0 ;
  assign n2010 = ( n293 & n2008 ) | ( n293 & ~n2009 ) | ( n2008 & ~n2009 ) ;
  assign n2011 = n1011 & ~n1470 ;
  assign n2012 = n2010 & n2011 ;
  assign n2013 = n772 & ~n2012 ;
  assign n2014 = n2013 ^ n520 ^ 1'b0 ;
  assign n2015 = n2014 ^ n1854 ^ x222 ;
  assign n2016 = x58 & x203 ;
  assign n2017 = ~x122 & n2016 ;
  assign n2018 = ~n618 & n2017 ;
  assign n2019 = n2018 ^ n1331 ^ 1'b0 ;
  assign n2020 = n1812 | n2019 ;
  assign n2021 = n554 | n1037 ;
  assign n2022 = ( n1813 & n2020 ) | ( n1813 & n2021 ) | ( n2020 & n2021 ) ;
  assign n2023 = n273 | n488 ;
  assign n2024 = ( ~x253 & n1743 ) | ( ~x253 & n2023 ) | ( n1743 & n2023 ) ;
  assign n2025 = n1077 ^ n866 ^ 1'b0 ;
  assign n2026 = n1404 & ~n2025 ;
  assign n2027 = ( n1150 & n1394 ) | ( n1150 & n1926 ) | ( n1394 & n1926 ) ;
  assign n2029 = n1910 ^ n360 ^ x174 ;
  assign n2030 = ( n439 & n933 ) | ( n439 & ~n2029 ) | ( n933 & ~n2029 ) ;
  assign n2028 = ~n262 & n1610 ;
  assign n2031 = n2030 ^ n2028 ^ x49 ;
  assign n2032 = x176 & n260 ;
  assign n2033 = n2032 ^ x99 ^ 1'b0 ;
  assign n2034 = n752 ^ n742 ^ n257 ;
  assign n2035 = n2033 & ~n2034 ;
  assign n2036 = ( n656 & n1424 ) | ( n656 & n2035 ) | ( n1424 & n2035 ) ;
  assign n2037 = n2017 ^ n668 ^ 1'b0 ;
  assign n2038 = n403 & ~n2037 ;
  assign n2039 = n2038 ^ n1048 ^ n600 ;
  assign n2040 = n1241 & n2039 ;
  assign n2041 = n1528 ^ x229 ^ 1'b0 ;
  assign n2042 = n2040 | n2041 ;
  assign n2043 = ~n2036 & n2042 ;
  assign n2044 = n1213 | n1665 ;
  assign n2045 = n2044 ^ n445 ^ 1'b0 ;
  assign n2046 = ~n917 & n2045 ;
  assign n2047 = n314 ^ n289 ^ 1'b0 ;
  assign n2048 = n556 | n2047 ;
  assign n2049 = n2048 ^ x184 ^ x13 ;
  assign n2050 = n1812 ^ n627 ^ x41 ;
  assign n2051 = n1230 ^ n587 ^ x237 ;
  assign n2052 = n557 ^ n312 ^ x136 ;
  assign n2053 = ~n997 & n2052 ;
  assign n2054 = ( n582 & n2051 ) | ( n582 & ~n2053 ) | ( n2051 & ~n2053 ) ;
  assign n2055 = n419 ^ n268 ^ 1'b0 ;
  assign n2056 = n2055 ^ x174 ^ x97 ;
  assign n2057 = ( n2050 & ~n2054 ) | ( n2050 & n2056 ) | ( ~n2054 & n2056 ) ;
  assign n2058 = x183 & n471 ;
  assign n2059 = ~n400 & n2058 ;
  assign n2060 = n2059 ^ n682 ^ 1'b0 ;
  assign n2061 = ( ~x66 & n1854 ) | ( ~x66 & n2060 ) | ( n1854 & n2060 ) ;
  assign n2062 = ( x186 & n2017 ) | ( x186 & n2061 ) | ( n2017 & n2061 ) ;
  assign n2063 = n1049 | n2062 ;
  assign n2068 = ~n315 & n899 ;
  assign n2069 = n2068 ^ n676 ^ 1'b0 ;
  assign n2070 = ( n362 & n1995 ) | ( n362 & n2069 ) | ( n1995 & n2069 ) ;
  assign n2071 = ( x237 & n598 ) | ( x237 & ~n2070 ) | ( n598 & ~n2070 ) ;
  assign n2072 = ( x206 & ~n696 ) | ( x206 & n831 ) | ( ~n696 & n831 ) ;
  assign n2073 = ( ~n609 & n2071 ) | ( ~n609 & n2072 ) | ( n2071 & n2072 ) ;
  assign n2064 = n610 ^ x71 ^ 1'b0 ;
  assign n2065 = ( x202 & ~n625 ) | ( x202 & n2064 ) | ( ~n625 & n2064 ) ;
  assign n2066 = ( x23 & ~x40 ) | ( x23 & n732 ) | ( ~x40 & n732 ) ;
  assign n2067 = n2065 | n2066 ;
  assign n2074 = n2073 ^ n2067 ^ 1'b0 ;
  assign n2075 = x137 & ~n885 ;
  assign n2076 = n2075 ^ x44 ^ 1'b0 ;
  assign n2077 = n2076 ^ n1885 ^ 1'b0 ;
  assign n2082 = n1164 ^ n538 ^ 1'b0 ;
  assign n2083 = x238 & n2082 ;
  assign n2084 = ( n582 & n1326 ) | ( n582 & n2083 ) | ( n1326 & n2083 ) ;
  assign n2085 = ( ~n1103 & n1241 ) | ( ~n1103 & n1309 ) | ( n1241 & n1309 ) ;
  assign n2086 = ( n630 & n2084 ) | ( n630 & ~n2085 ) | ( n2084 & ~n2085 ) ;
  assign n2078 = n969 & n1217 ;
  assign n2079 = n297 & n2078 ;
  assign n2080 = n2079 ^ n982 ^ x68 ;
  assign n2081 = n589 | n2080 ;
  assign n2087 = n2086 ^ n2081 ^ 1'b0 ;
  assign n2088 = x22 & n1877 ;
  assign n2089 = n2088 ^ n1282 ^ 1'b0 ;
  assign n2090 = n407 | n861 ;
  assign n2091 = n2090 ^ n1156 ^ n708 ;
  assign n2092 = ( x6 & ~x162 ) | ( x6 & n1854 ) | ( ~x162 & n1854 ) ;
  assign n2093 = n1121 ^ n739 ^ 1'b0 ;
  assign n2094 = ~n702 & n2093 ;
  assign n2095 = ( n905 & n2092 ) | ( n905 & n2094 ) | ( n2092 & n2094 ) ;
  assign n2097 = ( n431 & n719 ) | ( n431 & n1709 ) | ( n719 & n1709 ) ;
  assign n2098 = n2097 ^ n1303 ^ n1069 ;
  assign n2096 = n1961 ^ n1798 ^ 1'b0 ;
  assign n2099 = n2098 ^ n2096 ^ x40 ;
  assign n2100 = n2055 ^ n835 ^ 1'b0 ;
  assign n2101 = n326 & n2100 ;
  assign n2102 = ~x8 & n2101 ;
  assign n2103 = n1282 ^ n986 ^ n384 ;
  assign n2104 = ( n798 & ~n969 ) | ( n798 & n2103 ) | ( ~n969 & n2103 ) ;
  assign n2105 = x192 & n433 ;
  assign n2106 = n2104 & ~n2105 ;
  assign n2107 = ( ~x112 & n802 ) | ( ~x112 & n1423 ) | ( n802 & n1423 ) ;
  assign n2108 = ~x41 & n2107 ;
  assign n2109 = n1474 ^ n734 ^ x143 ;
  assign n2110 = ( n849 & n1222 ) | ( n849 & ~n2109 ) | ( n1222 & ~n2109 ) ;
  assign n2113 = n1323 ^ n526 ^ x245 ;
  assign n2111 = n1814 ^ x216 ^ 1'b0 ;
  assign n2112 = ( n525 & n1291 ) | ( n525 & n2111 ) | ( n1291 & n2111 ) ;
  assign n2114 = n2113 ^ n2112 ^ n741 ;
  assign n2115 = n2114 ^ n971 ^ 1'b0 ;
  assign n2116 = n1072 ^ n835 ^ 1'b0 ;
  assign n2117 = ~n525 & n2116 ;
  assign n2118 = ( n418 & n606 ) | ( n418 & n2117 ) | ( n606 & n2117 ) ;
  assign n2119 = n387 | n2118 ;
  assign n2120 = n2115 & ~n2119 ;
  assign n2121 = n1853 | n2120 ;
  assign n2122 = n614 & n693 ;
  assign n2123 = n2122 ^ n586 ^ 1'b0 ;
  assign n2124 = ( x83 & ~x166 ) | ( x83 & n1468 ) | ( ~x166 & n1468 ) ;
  assign n2125 = n1243 ^ n887 ^ 1'b0 ;
  assign n2126 = n1095 & n2125 ;
  assign n2127 = n2126 ^ n575 ^ 1'b0 ;
  assign n2128 = n493 ^ x239 ^ 1'b0 ;
  assign n2129 = x81 & n464 ;
  assign n2130 = n1779 & n2129 ;
  assign n2131 = n337 ^ x152 ^ x81 ;
  assign n2132 = x160 & ~n2131 ;
  assign n2133 = x10 & ~n2008 ;
  assign n2134 = ~n345 & n2133 ;
  assign n2135 = n1683 & ~n2134 ;
  assign n2136 = ~n733 & n1394 ;
  assign n2137 = ~n1164 & n2136 ;
  assign n2138 = n2137 ^ n1644 ^ 1'b0 ;
  assign n2139 = n2138 ^ n1555 ^ n1097 ;
  assign n2140 = ~n1708 & n2139 ;
  assign n2141 = n923 ^ n493 ^ 1'b0 ;
  assign n2142 = ( n416 & n559 ) | ( n416 & ~n697 ) | ( n559 & ~n697 ) ;
  assign n2143 = ( n1648 & n2141 ) | ( n1648 & n2142 ) | ( n2141 & n2142 ) ;
  assign n2144 = n2117 ^ n1516 ^ x178 ;
  assign n2145 = ( x23 & n1705 ) | ( x23 & n2144 ) | ( n1705 & n2144 ) ;
  assign n2146 = n2145 ^ n2039 ^ 1'b0 ;
  assign n2147 = x191 | n565 ;
  assign n2148 = n2147 ^ n911 ^ n750 ;
  assign n2149 = n1969 ^ x107 ^ 1'b0 ;
  assign n2150 = ( n286 & n967 ) | ( n286 & n2149 ) | ( n967 & n2149 ) ;
  assign n2151 = n1979 ^ x76 ^ 1'b0 ;
  assign n2152 = x143 & n2151 ;
  assign n2153 = n718 | n810 ;
  assign n2154 = n2153 ^ n257 ^ 1'b0 ;
  assign n2155 = ( n333 & n706 ) | ( n333 & n933 ) | ( n706 & n933 ) ;
  assign n2156 = n1067 ^ n967 ^ 1'b0 ;
  assign n2157 = ~n2155 & n2156 ;
  assign n2158 = n2157 ^ n799 ^ x85 ;
  assign n2159 = n436 | n514 ;
  assign n2160 = n1634 & ~n2159 ;
  assign n2161 = n1341 | n2160 ;
  assign n2162 = n682 | n2161 ;
  assign n2163 = ( n2154 & n2158 ) | ( n2154 & ~n2162 ) | ( n2158 & ~n2162 ) ;
  assign n2164 = n392 & n1646 ;
  assign n2165 = n495 & n2164 ;
  assign n2166 = n2165 ^ x153 ^ x22 ;
  assign n2167 = n1076 ^ n840 ^ n787 ;
  assign n2168 = ~n313 & n1593 ;
  assign n2169 = ( n2166 & ~n2167 ) | ( n2166 & n2168 ) | ( ~n2167 & n2168 ) ;
  assign n2170 = n584 & n623 ;
  assign n2171 = ~n2051 & n2170 ;
  assign n2172 = ( ~n513 & n1602 ) | ( ~n513 & n2171 ) | ( n1602 & n2171 ) ;
  assign n2173 = n2172 ^ n999 ^ n887 ;
  assign n2174 = n602 | n833 ;
  assign n2175 = n542 ^ n326 ^ x66 ;
  assign n2176 = ( n285 & n426 ) | ( n285 & ~n803 ) | ( n426 & ~n803 ) ;
  assign n2177 = ( ~x186 & n257 ) | ( ~x186 & n2176 ) | ( n257 & n2176 ) ;
  assign n2178 = ( n822 & n1068 ) | ( n822 & n2177 ) | ( n1068 & n2177 ) ;
  assign n2179 = n483 & ~n1643 ;
  assign n2180 = n392 & ~n1064 ;
  assign n2181 = n1430 ^ n1112 ^ 1'b0 ;
  assign n2182 = ~n2180 & n2181 ;
  assign n2183 = ( x6 & ~x31 ) | ( x6 & x113 ) | ( ~x31 & x113 ) ;
  assign n2184 = ( n352 & ~n1095 ) | ( n352 & n2183 ) | ( ~n1095 & n2183 ) ;
  assign n2185 = n2184 ^ n603 ^ 1'b0 ;
  assign n2187 = n675 ^ n520 ^ x207 ;
  assign n2186 = n853 & n1419 ;
  assign n2188 = n2187 ^ n2186 ^ 1'b0 ;
  assign n2189 = ~n943 & n1078 ;
  assign n2190 = n2189 ^ n862 ^ 1'b0 ;
  assign n2191 = n2190 ^ n745 ^ 1'b0 ;
  assign n2192 = n2191 ^ n1612 ^ n493 ;
  assign n2193 = ( n1163 & n2188 ) | ( n1163 & ~n2192 ) | ( n2188 & ~n2192 ) ;
  assign n2194 = x133 | n740 ;
  assign n2195 = ( n261 & n1400 ) | ( n261 & ~n2194 ) | ( n1400 & ~n2194 ) ;
  assign n2203 = x116 & ~n828 ;
  assign n2204 = n1524 & n2203 ;
  assign n2196 = ( n643 & ~n1303 ) | ( n643 & n1997 ) | ( ~n1303 & n1997 ) ;
  assign n2199 = x194 & ~n575 ;
  assign n2197 = x81 & ~n1046 ;
  assign n2198 = n2197 ^ n682 ^ 1'b0 ;
  assign n2200 = n2199 ^ n2198 ^ 1'b0 ;
  assign n2201 = n2200 ^ n1492 ^ n376 ;
  assign n2202 = ~n2196 & n2201 ;
  assign n2205 = n2204 ^ n2202 ^ 1'b0 ;
  assign n2206 = n1611 ^ n1005 ^ n724 ;
  assign n2207 = n2206 ^ n1818 ^ n1789 ;
  assign n2208 = x191 & n873 ;
  assign n2209 = n2065 ^ n1997 ^ n1673 ;
  assign n2210 = ~n1543 & n1946 ;
  assign n2211 = x244 & n748 ;
  assign n2212 = ~n2210 & n2211 ;
  assign n2213 = ( x79 & n1067 ) | ( x79 & n2212 ) | ( n1067 & n2212 ) ;
  assign n2214 = n1526 ^ n1048 ^ 1'b0 ;
  assign n2215 = x89 & ~n873 ;
  assign n2216 = ~n851 & n2215 ;
  assign n2217 = ~n2131 & n2216 ;
  assign n2218 = n2086 ^ n1894 ^ n1563 ;
  assign n2229 = n1003 ^ n636 ^ 1'b0 ;
  assign n2230 = n2229 ^ n895 ^ x205 ;
  assign n2231 = n885 & n2230 ;
  assign n2232 = n2231 ^ n965 ^ 1'b0 ;
  assign n2233 = n724 & n2232 ;
  assign n2219 = n596 | n865 ;
  assign n2220 = n910 | n2219 ;
  assign n2221 = x167 & n1655 ;
  assign n2222 = n2221 ^ n313 ^ 1'b0 ;
  assign n2223 = n293 | n560 ;
  assign n2224 = n1336 & ~n2223 ;
  assign n2225 = n2224 ^ n2062 ^ 1'b0 ;
  assign n2226 = ~n2222 & n2225 ;
  assign n2227 = n2220 & n2226 ;
  assign n2228 = n2227 ^ n1940 ^ 1'b0 ;
  assign n2234 = n2233 ^ n2228 ^ 1'b0 ;
  assign n2236 = x104 & ~n1129 ;
  assign n2237 = n740 & n2236 ;
  assign n2235 = n1631 & n1988 ;
  assign n2238 = n2237 ^ n2235 ^ 1'b0 ;
  assign n2239 = x229 & n2238 ;
  assign n2240 = n2239 ^ x14 ^ 1'b0 ;
  assign n2241 = n1573 | n2240 ;
  assign n2242 = n848 & ~n2241 ;
  assign n2243 = n1451 ^ n910 ^ x204 ;
  assign n2249 = x180 & n930 ;
  assign n2250 = n896 & n2249 ;
  assign n2251 = ( x159 & n748 ) | ( x159 & n2250 ) | ( n748 & n2250 ) ;
  assign n2252 = ( n523 & n1096 ) | ( n523 & ~n1566 ) | ( n1096 & ~n1566 ) ;
  assign n2253 = n1073 ^ n1026 ^ 1'b0 ;
  assign n2254 = n2252 & n2253 ;
  assign n2255 = ( n2210 & ~n2251 ) | ( n2210 & n2254 ) | ( ~n2251 & n2254 ) ;
  assign n2244 = n475 ^ n356 ^ 1'b0 ;
  assign n2245 = n540 & ~n1485 ;
  assign n2246 = ~x198 & n2245 ;
  assign n2247 = ( n1076 & n1101 ) | ( n1076 & ~n2246 ) | ( n1101 & ~n2246 ) ;
  assign n2248 = ( ~n1385 & n2244 ) | ( ~n1385 & n2247 ) | ( n2244 & n2247 ) ;
  assign n2256 = n2255 ^ n2248 ^ n1974 ;
  assign n2257 = ( x78 & n2243 ) | ( x78 & n2256 ) | ( n2243 & n2256 ) ;
  assign n2258 = n713 | n1918 ;
  assign n2259 = n2258 ^ n1000 ^ 1'b0 ;
  assign n2270 = ( n841 & n1000 ) | ( n841 & ~n2025 ) | ( n1000 & ~n2025 ) ;
  assign n2266 = ( n397 & n672 ) | ( n397 & n1093 ) | ( n672 & n1093 ) ;
  assign n2267 = n2266 ^ n975 ^ n826 ;
  assign n2264 = n2010 ^ n1624 ^ 1'b0 ;
  assign n2265 = n434 & ~n2264 ;
  assign n2268 = n2267 ^ n2265 ^ 1'b0 ;
  assign n2269 = x172 & n2268 ;
  assign n2261 = n1176 ^ n717 ^ 1'b0 ;
  assign n2262 = n618 | n2261 ;
  assign n2263 = n797 & ~n2262 ;
  assign n2271 = n2270 ^ n2269 ^ n2263 ;
  assign n2260 = x70 & x172 ;
  assign n2272 = n2271 ^ n2260 ^ n857 ;
  assign n2273 = ( ~x243 & n499 ) | ( ~x243 & n997 ) | ( n499 & n997 ) ;
  assign n2274 = n2273 ^ n842 ^ 1'b0 ;
  assign n2275 = n1039 | n1567 ;
  assign n2276 = n2275 ^ n454 ^ 1'b0 ;
  assign n2277 = n924 ^ n663 ^ 1'b0 ;
  assign n2278 = n2276 | n2277 ;
  assign n2279 = n2278 ^ n386 ^ 1'b0 ;
  assign n2280 = n538 ^ n315 ^ 1'b0 ;
  assign n2281 = ~n1819 & n2280 ;
  assign n2282 = ~n1781 & n2281 ;
  assign n2283 = n1276 ^ n663 ^ n627 ;
  assign n2284 = n1836 & n2283 ;
  assign n2285 = n2284 ^ n2039 ^ 1'b0 ;
  assign n2286 = ( n2250 & ~n2282 ) | ( n2250 & n2285 ) | ( ~n2282 & n2285 ) ;
  assign n2287 = ~n502 & n572 ;
  assign n2288 = ~n2286 & n2287 ;
  assign n2289 = n2196 ^ n485 ^ 1'b0 ;
  assign n2290 = n1323 & ~n2289 ;
  assign n2291 = ~x3 & n2290 ;
  assign n2292 = ~n335 & n865 ;
  assign n2293 = n2292 ^ n539 ^ 1'b0 ;
  assign n2294 = n499 & n763 ;
  assign n2295 = n580 & n2294 ;
  assign n2296 = n2295 ^ n1563 ^ n745 ;
  assign n2297 = n1542 & n2296 ;
  assign n2298 = ~n2293 & n2297 ;
  assign n2299 = n711 ^ n257 ^ 1'b0 ;
  assign n2300 = n920 | n2299 ;
  assign n2301 = ( n748 & ~n1667 ) | ( n748 & n2300 ) | ( ~n1667 & n2300 ) ;
  assign n2302 = n894 ^ x194 ^ 1'b0 ;
  assign n2303 = x37 & n2302 ;
  assign n2304 = ~n2301 & n2303 ;
  assign n2314 = x32 | n1825 ;
  assign n2308 = n1276 ^ n847 ^ 1'b0 ;
  assign n2309 = n314 ^ x135 ^ 1'b0 ;
  assign n2310 = ( n2039 & ~n2308 ) | ( n2039 & n2309 ) | ( ~n2308 & n2309 ) ;
  assign n2307 = ~n495 & n695 ;
  assign n2311 = n2310 ^ n2307 ^ 1'b0 ;
  assign n2305 = ( n1164 & n1224 ) | ( n1164 & ~n1334 ) | ( n1224 & ~n1334 ) ;
  assign n2306 = n1436 & n2305 ;
  assign n2312 = n2311 ^ n2306 ^ 1'b0 ;
  assign n2313 = n2312 ^ n598 ^ n422 ;
  assign n2315 = n2314 ^ n2313 ^ n779 ;
  assign n2318 = x235 & n983 ;
  assign n2319 = ( n1039 & ~n1923 ) | ( n1039 & n2318 ) | ( ~n1923 & n2318 ) ;
  assign n2316 = n799 | n941 ;
  assign n2317 = n2316 ^ n1981 ^ n1724 ;
  assign n2320 = n2319 ^ n2317 ^ x123 ;
  assign n2331 = n2094 ^ n901 ^ n883 ;
  assign n2328 = x119 & ~n610 ;
  assign n2329 = ~x179 & n2328 ;
  assign n2330 = n2329 ^ n789 ^ n737 ;
  assign n2332 = n2331 ^ n2330 ^ n1839 ;
  assign n2326 = n2126 ^ n874 ^ n766 ;
  assign n2321 = n293 | n533 ;
  assign n2322 = n2321 ^ n1823 ^ 1'b0 ;
  assign n2323 = n467 & n2322 ;
  assign n2324 = n2323 ^ n410 ^ 1'b0 ;
  assign n2325 = n2324 ^ x147 ^ 1'b0 ;
  assign n2327 = n2326 ^ n2325 ^ n1838 ;
  assign n2333 = n2332 ^ n2327 ^ n437 ;
  assign n2334 = n2117 ^ n262 ^ 1'b0 ;
  assign n2335 = ~n1749 & n2334 ;
  assign n2336 = n1427 & n1440 ;
  assign n2337 = n2336 ^ x69 ^ 1'b0 ;
  assign n2338 = ( ~n509 & n2335 ) | ( ~n509 & n2337 ) | ( n2335 & n2337 ) ;
  assign n2339 = x104 & n829 ;
  assign n2340 = ~x20 & n2339 ;
  assign n2341 = n1236 ^ x30 ^ 1'b0 ;
  assign n2342 = ~n2340 & n2341 ;
  assign n2343 = n2342 ^ n1834 ^ x65 ;
  assign n2344 = n2343 ^ n835 ^ 1'b0 ;
  assign n2345 = n2338 & ~n2344 ;
  assign n2346 = ~n403 & n2345 ;
  assign n2347 = n2346 ^ n2166 ^ 1'b0 ;
  assign n2348 = n2347 ^ n1530 ^ n995 ;
  assign n2354 = ( ~n1563 & n2017 ) | ( ~n1563 & n2269 ) | ( n2017 & n2269 ) ;
  assign n2350 = ( ~n314 & n577 ) | ( ~n314 & n1306 ) | ( n577 & n1306 ) ;
  assign n2349 = ( n626 & n1653 ) | ( n626 & n1731 ) | ( n1653 & n1731 ) ;
  assign n2351 = n2350 ^ n2349 ^ n1278 ;
  assign n2352 = n2351 ^ n1469 ^ 1'b0 ;
  assign n2353 = n2352 ^ n883 ^ x235 ;
  assign n2355 = n2354 ^ n2353 ^ n1237 ;
  assign n2366 = n1058 ^ n434 ^ 1'b0 ;
  assign n2367 = n550 | n2366 ;
  assign n2368 = n2367 ^ n2062 ^ 1'b0 ;
  assign n2369 = ~n1766 & n2368 ;
  assign n2356 = n1908 ^ n1662 ^ n1466 ;
  assign n2357 = ( ~n528 & n1048 ) | ( ~n528 & n2356 ) | ( n1048 & n2356 ) ;
  assign n2360 = ( n572 & n934 ) | ( n572 & ~n1012 ) | ( n934 & ~n1012 ) ;
  assign n2358 = x123 & n425 ;
  assign n2359 = n1825 & n2358 ;
  assign n2361 = n2360 ^ n2359 ^ 1'b0 ;
  assign n2362 = ~n295 & n2361 ;
  assign n2363 = ~n2357 & n2362 ;
  assign n2364 = n785 & n2363 ;
  assign n2365 = n2364 ^ n1567 ^ n1284 ;
  assign n2370 = n2369 ^ n2365 ^ n2036 ;
  assign n2371 = ~n936 & n1200 ;
  assign n2372 = ( x189 & ~x236 ) | ( x189 & n2371 ) | ( ~x236 & n2371 ) ;
  assign n2373 = n481 & n1224 ;
  assign n2375 = n1264 ^ x21 ^ 1'b0 ;
  assign n2374 = n1595 ^ n1367 ^ 1'b0 ;
  assign n2376 = n2375 ^ n2374 ^ n570 ;
  assign n2377 = n1023 & ~n1297 ;
  assign n2378 = ( n1319 & n2376 ) | ( n1319 & ~n2377 ) | ( n2376 & ~n2377 ) ;
  assign n2379 = n1104 & ~n1740 ;
  assign n2380 = ~x14 & n2379 ;
  assign n2381 = n2380 ^ n2137 ^ n893 ;
  assign n2382 = n2381 ^ n265 ^ 1'b0 ;
  assign n2383 = n2382 ^ n1812 ^ 1'b0 ;
  assign n2384 = n1909 & ~n2383 ;
  assign n2385 = n2384 ^ n349 ^ 1'b0 ;
  assign n2386 = n999 & ~n2385 ;
  assign n2387 = n1388 ^ n1220 ^ n1044 ;
  assign n2391 = n834 ^ n775 ^ n671 ;
  assign n2392 = n2391 ^ n1236 ^ n997 ;
  assign n2388 = n1845 ^ n433 ^ n419 ;
  assign n2389 = n1153 & n2388 ;
  assign n2390 = ~n1315 & n2389 ;
  assign n2393 = n2392 ^ n2390 ^ 1'b0 ;
  assign n2394 = n1515 ^ n1363 ^ 1'b0 ;
  assign n2395 = n947 & ~n1163 ;
  assign n2396 = n2395 ^ n1196 ^ 1'b0 ;
  assign n2397 = ( n573 & n687 ) | ( n573 & ~n2396 ) | ( n687 & ~n2396 ) ;
  assign n2398 = n2397 ^ n840 ^ x229 ;
  assign n2399 = n645 ^ x231 ^ 1'b0 ;
  assign n2400 = x38 & ~n2399 ;
  assign n2401 = ( x248 & n343 ) | ( x248 & ~n2400 ) | ( n343 & ~n2400 ) ;
  assign n2402 = ( n2100 & ~n2398 ) | ( n2100 & n2401 ) | ( ~n2398 & n2401 ) ;
  assign n2403 = x159 & ~n1430 ;
  assign n2404 = ~x104 & n2403 ;
  assign n2405 = n1048 ^ n971 ^ n567 ;
  assign n2406 = ( n1096 & ~n1807 ) | ( n1096 & n2405 ) | ( ~n1807 & n2405 ) ;
  assign n2407 = n784 | n1727 ;
  assign n2408 = n2407 ^ n290 ^ 1'b0 ;
  assign n2409 = ~n1059 & n2408 ;
  assign n2410 = ( n2404 & ~n2406 ) | ( n2404 & n2409 ) | ( ~n2406 & n2409 ) ;
  assign n2411 = n1354 ^ n930 ^ 1'b0 ;
  assign n2412 = n1693 | n2038 ;
  assign n2413 = n2412 ^ n1731 ^ 1'b0 ;
  assign n2414 = n2413 ^ n1804 ^ 1'b0 ;
  assign n2415 = n2145 & n2414 ;
  assign n2416 = n868 ^ n861 ^ n669 ;
  assign n2417 = x78 & ~n564 ;
  assign n2418 = ( n523 & n815 ) | ( n523 & n2417 ) | ( n815 & n2417 ) ;
  assign n2419 = ( n1200 & n2042 ) | ( n1200 & ~n2418 ) | ( n2042 & ~n2418 ) ;
  assign n2426 = n1368 ^ n1226 ^ 1'b0 ;
  assign n2420 = n266 & n1508 ;
  assign n2421 = n2420 ^ n627 ^ 1'b0 ;
  assign n2422 = n2351 & n2421 ;
  assign n2423 = n1544 | n2422 ;
  assign n2424 = n660 & ~n2423 ;
  assign n2425 = ( n1957 & n1988 ) | ( n1957 & ~n2424 ) | ( n1988 & ~n2424 ) ;
  assign n2427 = n2426 ^ n2425 ^ n1491 ;
  assign n2428 = n1235 & ~n2424 ;
  assign n2429 = n2374 ^ n1876 ^ 1'b0 ;
  assign n2430 = n2059 ^ n2023 ^ 1'b0 ;
  assign n2431 = n2430 ^ n2392 ^ 1'b0 ;
  assign n2432 = ~n1314 & n2431 ;
  assign n2433 = n1270 ^ n1111 ^ n798 ;
  assign n2434 = n531 | n1195 ;
  assign n2435 = n853 ^ n516 ^ 1'b0 ;
  assign n2436 = n2434 | n2435 ;
  assign n2437 = n607 & ~n2436 ;
  assign n2438 = n1329 & n2437 ;
  assign n2439 = n1396 | n2438 ;
  assign n2440 = n2433 | n2439 ;
  assign n2441 = ( n1987 & n2432 ) | ( n1987 & ~n2440 ) | ( n2432 & ~n2440 ) ;
  assign n2442 = ( x5 & ~x251 ) | ( x5 & n718 ) | ( ~x251 & n718 ) ;
  assign n2443 = n2442 ^ n1962 ^ 1'b0 ;
  assign n2444 = n2443 ^ n1672 ^ n407 ;
  assign n2445 = n1297 ^ n1284 ^ 1'b0 ;
  assign n2446 = ( x198 & ~x206 ) | ( x198 & n601 ) | ( ~x206 & n601 ) ;
  assign n2455 = ( n792 & ~n843 ) | ( n792 & n1173 ) | ( ~n843 & n1173 ) ;
  assign n2456 = ( n351 & n502 ) | ( n351 & n2166 ) | ( n502 & n2166 ) ;
  assign n2457 = x166 & n662 ;
  assign n2458 = ~n258 & n2457 ;
  assign n2459 = ( n492 & n2405 ) | ( n492 & n2458 ) | ( n2405 & n2458 ) ;
  assign n2460 = ( n264 & n2456 ) | ( n264 & n2459 ) | ( n2456 & n2459 ) ;
  assign n2461 = n2455 | n2460 ;
  assign n2462 = n1404 ^ x2 ^ 1'b0 ;
  assign n2463 = ~n2461 & n2462 ;
  assign n2447 = n546 | n1504 ;
  assign n2448 = n2447 ^ x201 ^ 1'b0 ;
  assign n2449 = n707 & ~n2448 ;
  assign n2450 = ~n1016 & n2449 ;
  assign n2451 = n1261 ^ n1101 ^ n483 ;
  assign n2452 = n2451 ^ n1251 ^ n329 ;
  assign n2453 = n1404 & n2452 ;
  assign n2454 = ~n2450 & n2453 ;
  assign n2464 = n2463 ^ n2454 ^ 1'b0 ;
  assign n2465 = x64 & ~n370 ;
  assign n2466 = n2465 ^ n907 ^ 1'b0 ;
  assign n2467 = ( ~n656 & n758 ) | ( ~n656 & n2466 ) | ( n758 & n2466 ) ;
  assign n2468 = x25 & n2466 ;
  assign n2469 = n2468 ^ n991 ^ 1'b0 ;
  assign n2470 = ( n891 & ~n2467 ) | ( n891 & n2469 ) | ( ~n2467 & n2469 ) ;
  assign n2471 = x121 & ~n796 ;
  assign n2472 = n2471 ^ n1699 ^ n307 ;
  assign n2473 = n366 | n775 ;
  assign n2474 = x129 | n2473 ;
  assign n2475 = n1883 ^ n308 ^ x39 ;
  assign n2476 = n1146 ^ n916 ^ n551 ;
  assign n2477 = n1144 | n1734 ;
  assign n2478 = n2477 ^ n1980 ^ 1'b0 ;
  assign n2479 = x9 & ~n2478 ;
  assign n2480 = n2479 ^ n403 ^ 1'b0 ;
  assign n2488 = ~n910 & n1376 ;
  assign n2489 = n2488 ^ n368 ^ 1'b0 ;
  assign n2490 = ( ~n957 & n1126 ) | ( ~n957 & n2434 ) | ( n1126 & n2434 ) ;
  assign n2491 = x35 & ~n2490 ;
  assign n2492 = n2489 & n2491 ;
  assign n2481 = ( ~n555 & n965 ) | ( ~n555 & n1101 ) | ( n965 & n1101 ) ;
  assign n2482 = ( n349 & n1390 ) | ( n349 & n2481 ) | ( n1390 & n2481 ) ;
  assign n2483 = n320 ^ x91 ^ 1'b0 ;
  assign n2484 = n2483 ^ n983 ^ 1'b0 ;
  assign n2485 = n2482 | n2484 ;
  assign n2486 = n989 & n2072 ;
  assign n2487 = ( n1597 & n2485 ) | ( n1597 & n2486 ) | ( n2485 & n2486 ) ;
  assign n2493 = n2492 ^ n2487 ^ n994 ;
  assign n2494 = ( ~n372 & n2110 ) | ( ~n372 & n2493 ) | ( n2110 & n2493 ) ;
  assign n2495 = ( n873 & n1446 ) | ( n873 & n1993 ) | ( n1446 & n1993 ) ;
  assign n2497 = n2138 ^ n1320 ^ 1'b0 ;
  assign n2498 = n2497 ^ n965 ^ x245 ;
  assign n2499 = n1455 & ~n2137 ;
  assign n2500 = n2498 & n2499 ;
  assign n2496 = ~n991 & n1703 ;
  assign n2501 = n2500 ^ n2496 ^ 1'b0 ;
  assign n2502 = n2036 ^ n1525 ^ 1'b0 ;
  assign n2509 = n531 | n811 ;
  assign n2510 = n2509 ^ n627 ^ 1'b0 ;
  assign n2503 = n555 ^ n467 ^ 1'b0 ;
  assign n2504 = n1004 ^ n355 ^ x230 ;
  assign n2505 = n567 & ~n1097 ;
  assign n2506 = ~n2504 & n2505 ;
  assign n2507 = n2503 | n2506 ;
  assign n2508 = n2507 ^ n386 ^ 1'b0 ;
  assign n2511 = n2510 ^ n2508 ^ n1534 ;
  assign n2512 = x97 & ~n1336 ;
  assign n2513 = ( ~x129 & n1823 ) | ( ~x129 & n2512 ) | ( n1823 & n2512 ) ;
  assign n2514 = n1217 & n2513 ;
  assign n2515 = n426 | n1005 ;
  assign n2526 = n667 | n1250 ;
  assign n2527 = n2526 ^ n1584 ^ x70 ;
  assign n2528 = n2527 ^ n2086 ^ n772 ;
  assign n2523 = n1784 ^ n1188 ^ n982 ;
  assign n2524 = n2523 ^ x8 ^ 1'b0 ;
  assign n2522 = n2252 ^ n280 ^ x65 ;
  assign n2525 = n2524 ^ n2522 ^ 1'b0 ;
  assign n2519 = ~n335 & n2375 ;
  assign n2520 = n2519 ^ n1220 ^ 1'b0 ;
  assign n2516 = n625 ^ n293 ^ 1'b0 ;
  assign n2517 = ~n470 & n2516 ;
  assign n2518 = ~n286 & n2517 ;
  assign n2521 = n2520 ^ n2518 ^ 1'b0 ;
  assign n2529 = n2528 ^ n2525 ^ n2521 ;
  assign n2530 = n2529 ^ n1492 ^ 1'b0 ;
  assign n2531 = n591 ^ n469 ^ 1'b0 ;
  assign n2532 = ~n1370 & n2531 ;
  assign n2533 = ( n2100 & n2350 ) | ( n2100 & n2532 ) | ( n2350 & n2532 ) ;
  assign n2534 = ~n1739 & n2533 ;
  assign n2535 = n2534 ^ n980 ^ 1'b0 ;
  assign n2536 = n1614 ^ x171 ^ 1'b0 ;
  assign n2537 = n1276 ^ n1274 ^ n465 ;
  assign n2538 = n509 & n900 ;
  assign n2539 = n2537 & n2538 ;
  assign n2540 = n1412 | n1822 ;
  assign n2541 = ~n625 & n1226 ;
  assign n2542 = n2541 ^ x12 ^ 1'b0 ;
  assign n2543 = n2540 & ~n2542 ;
  assign n2544 = n2282 | n2305 ;
  assign n2545 = n2544 ^ n374 ^ 1'b0 ;
  assign n2546 = n1230 ^ n689 ^ x181 ;
  assign n2547 = n1570 ^ n1462 ^ 1'b0 ;
  assign n2548 = x103 & ~n765 ;
  assign n2549 = n335 & n2548 ;
  assign n2550 = n1714 & ~n2549 ;
  assign n2551 = ( n1893 & n2547 ) | ( n1893 & ~n2550 ) | ( n2547 & ~n2550 ) ;
  assign n2552 = ( x179 & n2546 ) | ( x179 & n2551 ) | ( n2546 & n2551 ) ;
  assign n2556 = n346 ^ x85 ^ 1'b0 ;
  assign n2557 = ( x78 & n566 ) | ( x78 & ~n2556 ) | ( n566 & ~n2556 ) ;
  assign n2558 = n2557 ^ n1980 ^ n1306 ;
  assign n2559 = n436 | n2558 ;
  assign n2560 = n664 & ~n2559 ;
  assign n2553 = ( ~x137 & n737 ) | ( ~x137 & n1610 ) | ( n737 & n1610 ) ;
  assign n2554 = n1703 & n2553 ;
  assign n2555 = n2554 ^ n1206 ^ 1'b0 ;
  assign n2561 = n2560 ^ n2555 ^ 1'b0 ;
  assign n2562 = n494 ^ n322 ^ x228 ;
  assign n2563 = ( x42 & ~n1432 ) | ( x42 & n2562 ) | ( ~n1432 & n2562 ) ;
  assign n2564 = x85 & ~n1955 ;
  assign n2565 = n536 & n2564 ;
  assign n2566 = n303 | n890 ;
  assign n2567 = n2565 & ~n2566 ;
  assign n2568 = n2563 | n2567 ;
  assign n2569 = n2568 ^ n2124 ^ 1'b0 ;
  assign n2570 = n2061 ^ n1758 ^ n1444 ;
  assign n2571 = x50 | n586 ;
  assign n2572 = n1257 ^ x140 ^ 1'b0 ;
  assign n2573 = x124 & ~n2305 ;
  assign n2574 = n2573 ^ n1899 ^ 1'b0 ;
  assign n2575 = n551 ^ x243 ^ 1'b0 ;
  assign n2576 = n2575 ^ n2471 ^ 1'b0 ;
  assign n2577 = ~n2574 & n2576 ;
  assign n2578 = ~n433 & n1894 ;
  assign n2579 = n2578 ^ x118 ^ 1'b0 ;
  assign n2580 = n2579 ^ n2461 ^ n410 ;
  assign n2581 = n857 | n2155 ;
  assign n2582 = x70 | n2581 ;
  assign n2583 = x230 & ~n1152 ;
  assign n2584 = n471 ^ x169 ^ 1'b0 ;
  assign n2585 = ( x229 & ~n506 ) | ( x229 & n1088 ) | ( ~n506 & n1088 ) ;
  assign n2586 = x40 & ~n539 ;
  assign n2587 = n2586 ^ n436 ^ 1'b0 ;
  assign n2588 = n2587 ^ n1653 ^ 1'b0 ;
  assign n2589 = n2154 & n2588 ;
  assign n2590 = n2541 ^ n1205 ^ n423 ;
  assign n2591 = n767 & ~n1382 ;
  assign n2592 = n977 ^ x162 ^ 1'b0 ;
  assign n2593 = n2591 | n2592 ;
  assign n2594 = n2593 ^ n1206 ^ 1'b0 ;
  assign n2597 = n1980 ^ n378 ^ x206 ;
  assign n2595 = ( x64 & x108 ) | ( x64 & ~n1842 ) | ( x108 & ~n1842 ) ;
  assign n2596 = n2595 ^ n1175 ^ n324 ;
  assign n2598 = n2597 ^ n2596 ^ n1083 ;
  assign n2599 = n2598 ^ n668 ^ 1'b0 ;
  assign n2600 = n2594 & ~n2599 ;
  assign n2601 = ( ~n1786 & n2590 ) | ( ~n1786 & n2600 ) | ( n2590 & n2600 ) ;
  assign n2602 = ~n565 & n1075 ;
  assign n2603 = ( x8 & n1300 ) | ( x8 & n2602 ) | ( n1300 & n2602 ) ;
  assign n2604 = ~n279 & n1639 ;
  assign n2605 = n1705 ^ n1691 ^ n523 ;
  assign n2606 = n2605 ^ n1077 ^ n508 ;
  assign n2607 = ~n356 & n2512 ;
  assign n2608 = n1670 ^ n1044 ^ 1'b0 ;
  assign n2609 = ( ~n480 & n2607 ) | ( ~n480 & n2608 ) | ( n2607 & n2608 ) ;
  assign n2610 = ( ~n333 & n2523 ) | ( ~n333 & n2609 ) | ( n2523 & n2609 ) ;
  assign n2611 = n822 ^ x73 ^ x1 ;
  assign n2612 = n1239 | n1970 ;
  assign n2613 = n2611 | n2612 ;
  assign n2625 = x160 & ~n646 ;
  assign n2614 = n1965 ^ n1362 ^ n1331 ;
  assign n2615 = ( n384 & ~n1630 ) | ( n384 & n1965 ) | ( ~n1630 & n1965 ) ;
  assign n2616 = n2615 ^ n1015 ^ 1'b0 ;
  assign n2617 = n613 | n2616 ;
  assign n2618 = n2617 ^ x233 ^ 1'b0 ;
  assign n2619 = x93 & ~n2618 ;
  assign n2620 = ~n1315 & n2619 ;
  assign n2621 = n2620 ^ n1620 ^ 1'b0 ;
  assign n2622 = n1734 ^ n349 ^ 1'b0 ;
  assign n2623 = n1876 & n2622 ;
  assign n2624 = ( ~n2614 & n2621 ) | ( ~n2614 & n2623 ) | ( n2621 & n2623 ) ;
  assign n2626 = n2625 ^ n2624 ^ 1'b0 ;
  assign n2627 = n2613 & n2626 ;
  assign n2628 = n1169 ^ n1079 ^ x72 ;
  assign n2629 = n2628 ^ n1099 ^ n632 ;
  assign n2630 = n530 ^ x248 ^ 1'b0 ;
  assign n2631 = n932 & n2630 ;
  assign n2633 = n1468 ^ n1188 ^ n332 ;
  assign n2632 = n816 ^ x196 ^ x49 ;
  assign n2634 = n2633 ^ n2632 ^ n1693 ;
  assign n2635 = n2631 & ~n2634 ;
  assign n2636 = ~n1405 & n2635 ;
  assign n2637 = n2636 ^ n1714 ^ 1'b0 ;
  assign n2640 = ( x10 & n370 ) | ( x10 & ~n648 ) | ( n370 & ~n648 ) ;
  assign n2641 = ( n646 & ~n1189 ) | ( n646 & n2640 ) | ( ~n1189 & n2640 ) ;
  assign n2638 = n2452 ^ n735 ^ n429 ;
  assign n2639 = ( ~x63 & n1620 ) | ( ~x63 & n2638 ) | ( n1620 & n2638 ) ;
  assign n2642 = n2641 ^ n2639 ^ n656 ;
  assign n2643 = ~n2171 & n2642 ;
  assign n2660 = n1210 ^ n978 ^ 1'b0 ;
  assign n2661 = n1220 & n2660 ;
  assign n2662 = n2661 ^ n1710 ^ n1209 ;
  assign n2657 = ( ~x64 & x215 ) | ( ~x64 & n2066 ) | ( x215 & n2066 ) ;
  assign n2656 = ~n1920 & n2342 ;
  assign n2658 = n2657 ^ n2656 ^ 1'b0 ;
  assign n2659 = n2658 ^ n1830 ^ 1'b0 ;
  assign n2663 = n2662 ^ n2659 ^ 1'b0 ;
  assign n2664 = n1054 & ~n2663 ;
  assign n2665 = x111 & n2664 ;
  assign n2666 = n2665 ^ n591 ^ 1'b0 ;
  assign n2644 = n1630 ^ n1126 ^ 1'b0 ;
  assign n2647 = n898 ^ n533 ^ 1'b0 ;
  assign n2648 = x26 & n2647 ;
  assign n2649 = n2648 ^ n1302 ^ n587 ;
  assign n2650 = n1071 & n1128 ;
  assign n2651 = n2649 & n2650 ;
  assign n2652 = ( ~n640 & n2000 ) | ( ~n640 & n2651 ) | ( n2000 & n2651 ) ;
  assign n2645 = n1604 ^ n1352 ^ n279 ;
  assign n2646 = n1666 & n2645 ;
  assign n2653 = n2652 ^ n2646 ^ 1'b0 ;
  assign n2654 = n2644 & n2653 ;
  assign n2655 = n974 & n2654 ;
  assign n2667 = n2666 ^ n2655 ^ n812 ;
  assign n2676 = n1203 ^ n1022 ^ 1'b0 ;
  assign n2668 = n1570 ^ n861 ^ 1'b0 ;
  assign n2669 = n2668 ^ n656 ^ n625 ;
  assign n2670 = n2669 ^ n2424 ^ n1153 ;
  assign n2671 = n950 ^ n561 ^ 1'b0 ;
  assign n2672 = ( n902 & n1494 ) | ( n902 & n2671 ) | ( n1494 & n2671 ) ;
  assign n2673 = n2672 ^ n2391 ^ n1054 ;
  assign n2674 = n2673 ^ n1423 ^ n1130 ;
  assign n2675 = n2670 & ~n2674 ;
  assign n2677 = n2676 ^ n2675 ^ 1'b0 ;
  assign n2678 = n1084 & ~n2057 ;
  assign n2679 = ~x209 & n2678 ;
  assign n2680 = n1347 ^ n1028 ^ 1'b0 ;
  assign n2681 = n2680 ^ n1537 ^ x222 ;
  assign n2682 = n2681 ^ n1738 ^ n400 ;
  assign n2683 = n2682 ^ n1593 ^ 1'b0 ;
  assign n2684 = n1442 | n2683 ;
  assign n2687 = n282 ^ x181 ^ 1'b0 ;
  assign n2688 = x5 & n2687 ;
  assign n2689 = n1062 | n2460 ;
  assign n2690 = n2688 | n2689 ;
  assign n2685 = ~n1145 & n2110 ;
  assign n2686 = n2685 ^ n1759 ^ 1'b0 ;
  assign n2691 = n2690 ^ n2686 ^ n385 ;
  assign n2692 = ( ~n604 & n1173 ) | ( ~n604 & n2162 ) | ( n1173 & n2162 ) ;
  assign n2693 = n1250 ^ x167 ^ x35 ;
  assign n2694 = ~n891 & n2440 ;
  assign n2695 = ~n2693 & n2694 ;
  assign n2696 = n2692 | n2695 ;
  assign n2697 = n1102 ^ x134 ^ x48 ;
  assign n2698 = ( n923 & n2391 ) | ( n923 & n2697 ) | ( n2391 & n2697 ) ;
  assign n2699 = n1065 & ~n1858 ;
  assign n2700 = n280 & n2699 ;
  assign n2701 = ~n1736 & n2700 ;
  assign n2702 = ( ~n508 & n1624 ) | ( ~n508 & n2701 ) | ( n1624 & n2701 ) ;
  assign n2703 = ~n916 & n2702 ;
  assign n2704 = n2703 ^ n685 ^ 1'b0 ;
  assign n2709 = n971 ^ n865 ^ x154 ;
  assign n2710 = n2709 ^ x179 ^ 1'b0 ;
  assign n2711 = ~n1510 & n2710 ;
  assign n2705 = ( n1110 & ~n1649 ) | ( n1110 & n1722 ) | ( ~n1649 & n1722 ) ;
  assign n2706 = ~n391 & n988 ;
  assign n2707 = ( n276 & n572 ) | ( n276 & n2706 ) | ( n572 & n2706 ) ;
  assign n2708 = ( ~n1797 & n2705 ) | ( ~n1797 & n2707 ) | ( n2705 & n2707 ) ;
  assign n2712 = n2711 ^ n2708 ^ x38 ;
  assign n2713 = n1064 ^ n498 ^ 1'b0 ;
  assign n2714 = x21 & n2713 ;
  assign n2715 = ( n2066 & n2661 ) | ( n2066 & ~n2714 ) | ( n2661 & ~n2714 ) ;
  assign n2716 = ( n1440 & n2562 ) | ( n1440 & ~n2715 ) | ( n2562 & ~n2715 ) ;
  assign n2717 = n2716 ^ n2697 ^ n2693 ;
  assign n2718 = n617 ^ x241 ^ x79 ;
  assign n2719 = n2503 ^ x49 ^ 1'b0 ;
  assign n2720 = n322 | n2719 ;
  assign n2721 = n2718 | n2720 ;
  assign n2722 = n2721 ^ n981 ^ 1'b0 ;
  assign n2723 = n2722 ^ n1642 ^ 1'b0 ;
  assign n2724 = ( n534 & ~n924 ) | ( n534 & n2723 ) | ( ~n924 & n2723 ) ;
  assign n2725 = x0 & ~n476 ;
  assign n2730 = n1081 ^ n778 ^ 1'b0 ;
  assign n2731 = n897 | n2730 ;
  assign n2732 = ( n1163 & n1645 ) | ( n1163 & ~n2731 ) | ( n1645 & ~n2731 ) ;
  assign n2728 = n1573 ^ n997 ^ n613 ;
  assign n2726 = n466 ^ x114 ^ 1'b0 ;
  assign n2727 = x119 | n2726 ;
  assign n2729 = n2728 ^ n2727 ^ 1'b0 ;
  assign n2733 = n2732 ^ n2729 ^ 1'b0 ;
  assign n2734 = ( x172 & ~n711 ) | ( x172 & n2187 ) | ( ~n711 & n2187 ) ;
  assign n2735 = n810 & n2734 ;
  assign n2736 = n1229 ^ n859 ^ n783 ;
  assign n2737 = ( n324 & ~n410 ) | ( n324 & n2736 ) | ( ~n410 & n2736 ) ;
  assign n2738 = n2644 & n2737 ;
  assign n2739 = n2735 & n2738 ;
  assign n2740 = n283 | n2739 ;
  assign n2742 = n273 | n2485 ;
  assign n2743 = n1819 & ~n2742 ;
  assign n2741 = x0 & n1699 ;
  assign n2744 = n2743 ^ n2741 ^ 1'b0 ;
  assign n2748 = n2330 ^ n1909 ^ 1'b0 ;
  assign n2749 = ~n1304 & n2206 ;
  assign n2750 = ( n883 & n2748 ) | ( n883 & n2749 ) | ( n2748 & n2749 ) ;
  assign n2751 = n2750 ^ n2701 ^ n2417 ;
  assign n2745 = ~n1444 & n1466 ;
  assign n2746 = n2745 ^ n549 ^ 1'b0 ;
  assign n2752 = n2751 ^ n2746 ^ n2481 ;
  assign n2747 = ~n627 & n2746 ;
  assign n2753 = n2752 ^ n2747 ^ 1'b0 ;
  assign n2754 = n1427 ^ x51 ^ 1'b0 ;
  assign n2755 = ( n702 & n1662 ) | ( n702 & ~n2391 ) | ( n1662 & ~n2391 ) ;
  assign n2756 = n2755 ^ n932 ^ x225 ;
  assign n2757 = ( n1643 & n2405 ) | ( n1643 & n2756 ) | ( n2405 & n2756 ) ;
  assign n2758 = n676 & n2757 ;
  assign n2759 = n2758 ^ n325 ^ 1'b0 ;
  assign n2760 = ( n427 & ~n595 ) | ( n427 & n1877 ) | ( ~n595 & n1877 ) ;
  assign n2761 = n2760 ^ n2511 ^ n1206 ;
  assign n2769 = x169 & n744 ;
  assign n2770 = ( n849 & ~n1481 ) | ( n849 & n2769 ) | ( ~n1481 & n2769 ) ;
  assign n2762 = n2083 ^ n1802 ^ 1'b0 ;
  assign n2763 = n852 | n2762 ;
  assign n2764 = n529 & ~n1722 ;
  assign n2765 = n2764 ^ n2640 ^ n434 ;
  assign n2766 = n2765 ^ n1310 ^ n1197 ;
  assign n2767 = n1387 | n2766 ;
  assign n2768 = n2763 & ~n2767 ;
  assign n2771 = n2770 ^ n2768 ^ n2594 ;
  assign n2772 = n1072 ^ x1 ^ 1'b0 ;
  assign n2773 = n851 | n2772 ;
  assign n2774 = n2126 & ~n2773 ;
  assign n2775 = ~n2089 & n2774 ;
  assign n2776 = ~x210 & n1909 ;
  assign n2777 = n1620 ^ n1121 ^ n480 ;
  assign n2778 = n880 & ~n2777 ;
  assign n2779 = ( n844 & n1162 ) | ( n844 & n2778 ) | ( n1162 & n2778 ) ;
  assign n2780 = n2779 ^ n2565 ^ n1673 ;
  assign n2781 = ~n2776 & n2780 ;
  assign n2782 = n2781 ^ n463 ^ 1'b0 ;
  assign n2783 = n2782 ^ n478 ^ 1'b0 ;
  assign n2784 = n1141 | n2783 ;
  assign n2785 = ( n771 & n1213 ) | ( n771 & ~n2263 ) | ( n1213 & ~n2263 ) ;
  assign n2786 = n462 & ~n2481 ;
  assign n2787 = ~n1518 & n2786 ;
  assign n2788 = ( n2020 & n2722 ) | ( n2020 & ~n2787 ) | ( n2722 & ~n2787 ) ;
  assign n2789 = n506 & n2038 ;
  assign n2790 = n2789 ^ n298 ^ 1'b0 ;
  assign n2791 = n450 & ~n2790 ;
  assign n2792 = x13 | n2791 ;
  assign n2793 = n884 & ~n2792 ;
  assign n2795 = n1555 ^ n573 ^ 1'b0 ;
  assign n2796 = n858 & ~n2795 ;
  assign n2794 = ( n979 & ~n1274 ) | ( n979 & n1651 ) | ( ~n1274 & n1651 ) ;
  assign n2797 = n2796 ^ n2794 ^ n1351 ;
  assign n2798 = ~n478 & n984 ;
  assign n2799 = n2798 ^ x103 ^ 1'b0 ;
  assign n2800 = n2799 ^ n2111 ^ n630 ;
  assign n2801 = n1407 ^ n923 ^ 1'b0 ;
  assign n2802 = x41 & n2801 ;
  assign n2803 = n2802 ^ n2168 ^ 1'b0 ;
  assign n2804 = ~n2661 & n2803 ;
  assign n2805 = n2804 ^ n303 ^ 1'b0 ;
  assign n2806 = ~n2800 & n2805 ;
  assign n2807 = n2237 ^ n1217 ^ 1'b0 ;
  assign n2808 = n787 & n1713 ;
  assign n2809 = n2780 & ~n2808 ;
  assign n2810 = n1268 ^ n1126 ^ n589 ;
  assign n2811 = n1157 ^ n534 ^ x224 ;
  assign n2812 = ( ~x31 & x195 ) | ( ~x31 & n559 ) | ( x195 & n559 ) ;
  assign n2813 = ~n973 & n2812 ;
  assign n2814 = n2813 ^ x69 ^ x1 ;
  assign n2815 = n1225 & n2814 ;
  assign n2816 = n2811 & n2815 ;
  assign n2817 = ( n416 & n2810 ) | ( n416 & ~n2816 ) | ( n2810 & ~n2816 ) ;
  assign n2818 = n1007 | n1445 ;
  assign n2819 = n2818 ^ n885 ^ 1'b0 ;
  assign n2820 = n2166 ^ n1714 ^ 1'b0 ;
  assign n2821 = n1486 | n2820 ;
  assign n2822 = n2819 & ~n2821 ;
  assign n2823 = n836 | n1121 ;
  assign n2824 = n556 & ~n2823 ;
  assign n2825 = n2675 & ~n2824 ;
  assign n2826 = n2822 & n2825 ;
  assign n2827 = n1673 ^ n257 ^ x137 ;
  assign n2828 = ( ~n673 & n1228 ) | ( ~n673 & n2827 ) | ( n1228 & n2827 ) ;
  assign n2829 = ( n981 & n1113 ) | ( n981 & n2828 ) | ( n1113 & n2828 ) ;
  assign n2830 = n1816 ^ x146 ^ 1'b0 ;
  assign n2831 = n2829 | n2830 ;
  assign n2832 = n658 ^ x233 ^ x158 ;
  assign n2833 = n1584 | n2250 ;
  assign n2834 = n2833 ^ n1814 ^ 1'b0 ;
  assign n2835 = ( n923 & n2832 ) | ( n923 & ~n2834 ) | ( n2832 & ~n2834 ) ;
  assign n2836 = x123 & n2835 ;
  assign n2837 = n387 & n2836 ;
  assign n2838 = ( n489 & n2831 ) | ( n489 & n2837 ) | ( n2831 & n2837 ) ;
  assign n2839 = n736 & ~n2838 ;
  assign n2840 = n2839 ^ n1790 ^ 1'b0 ;
  assign n2841 = n2050 ^ n1113 ^ 1'b0 ;
  assign n2842 = n936 ^ n362 ^ x221 ;
  assign n2843 = n1319 & n2045 ;
  assign n2844 = n1257 ^ n1111 ^ x125 ;
  assign n2845 = n2111 ^ n833 ^ 1'b0 ;
  assign n2846 = n2844 & ~n2845 ;
  assign n2847 = ~n1135 & n2846 ;
  assign n2849 = x200 & x250 ;
  assign n2850 = n2849 ^ n529 ^ 1'b0 ;
  assign n2848 = n1759 ^ n719 ^ n433 ;
  assign n2851 = n2850 ^ n2848 ^ n2524 ;
  assign n2853 = n802 ^ n676 ^ 1'b0 ;
  assign n2854 = n1399 ^ n800 ^ 1'b0 ;
  assign n2855 = n2853 & ~n2854 ;
  assign n2856 = n1858 | n2855 ;
  assign n2852 = n1694 & ~n2155 ;
  assign n2857 = n2856 ^ n2852 ^ 1'b0 ;
  assign n2858 = ( n935 & n1997 ) | ( n935 & n2017 ) | ( n1997 & n2017 ) ;
  assign n2859 = n2858 ^ n2331 ^ x123 ;
  assign n2861 = ~n628 & n1645 ;
  assign n2862 = n2861 ^ n1126 ^ 1'b0 ;
  assign n2863 = n1765 & n2862 ;
  assign n2860 = n967 ^ n389 ^ n291 ;
  assign n2864 = n2863 ^ n2860 ^ n2163 ;
  assign n2866 = n1751 & n2105 ;
  assign n2867 = n2866 ^ n1638 ^ 1'b0 ;
  assign n2868 = ~n1777 & n2167 ;
  assign n2869 = n2867 & n2868 ;
  assign n2870 = n2869 ^ n2734 ^ 1'b0 ;
  assign n2871 = n1632 & ~n2870 ;
  assign n2865 = n2651 ^ n1915 ^ x112 ;
  assign n2872 = n2871 ^ n2865 ^ 1'b0 ;
  assign n2873 = n2194 & ~n2872 ;
  assign n2875 = ( n822 & n1068 ) | ( n822 & n1366 ) | ( n1068 & n1366 ) ;
  assign n2876 = n2875 ^ n792 ^ 1'b0 ;
  assign n2877 = n1702 & ~n2876 ;
  assign n2874 = n2098 ^ n1388 ^ x92 ;
  assign n2878 = n2877 ^ n2874 ^ 1'b0 ;
  assign n2879 = x80 | n2878 ;
  assign n2880 = ( ~x10 & x197 ) | ( ~x10 & n485 ) | ( x197 & n485 ) ;
  assign n2881 = ( n1304 & n1722 ) | ( n1304 & ~n2880 ) | ( n1722 & ~n2880 ) ;
  assign n2882 = n834 ^ x232 ^ 1'b0 ;
  assign n2883 = n1648 ^ n322 ^ 1'b0 ;
  assign n2884 = n1519 ^ n1463 ^ n1217 ;
  assign n2885 = ( ~n547 & n2562 ) | ( ~n547 & n2884 ) | ( n2562 & n2884 ) ;
  assign n2886 = n2329 | n2810 ;
  assign n2887 = ( ~n1937 & n2885 ) | ( ~n1937 & n2886 ) | ( n2885 & n2886 ) ;
  assign n2888 = n2288 | n2887 ;
  assign n2889 = n2888 ^ n1862 ^ 1'b0 ;
  assign n2890 = n2889 ^ n2415 ^ 1'b0 ;
  assign n2891 = n2883 & ~n2890 ;
  assign n2894 = x33 & n966 ;
  assign n2895 = ~n1172 & n2894 ;
  assign n2892 = x120 & ~n1893 ;
  assign n2893 = ~n2001 & n2892 ;
  assign n2896 = n2895 ^ n2893 ^ 1'b0 ;
  assign n2899 = n697 ^ n327 ^ x243 ;
  assign n2900 = n2899 ^ n692 ^ x12 ;
  assign n2901 = n2184 ^ n559 ^ 1'b0 ;
  assign n2902 = n2901 ^ x207 ^ 1'b0 ;
  assign n2903 = n2734 & ~n2902 ;
  assign n2904 = ( n1224 & n2900 ) | ( n1224 & n2903 ) | ( n2900 & n2903 ) ;
  assign n2897 = n997 & ~n1949 ;
  assign n2898 = n1675 & n2897 ;
  assign n2905 = n2904 ^ n2898 ^ n454 ;
  assign n2906 = n1023 & ~n2905 ;
  assign n2907 = n2856 ^ n2343 ^ n852 ;
  assign n2908 = n2907 ^ n2583 ^ n1915 ;
  assign n2909 = n1694 ^ x90 ^ 1'b0 ;
  assign n2910 = n2909 ^ n1427 ^ n1291 ;
  assign n2911 = x197 & ~n2910 ;
  assign n2912 = ( n1202 & n2908 ) | ( n1202 & ~n2911 ) | ( n2908 & ~n2911 ) ;
  assign n2916 = x223 & n363 ;
  assign n2917 = n2916 ^ n1340 ^ 1'b0 ;
  assign n2915 = ( n570 & ~n988 ) | ( n570 & n2187 ) | ( ~n988 & n2187 ) ;
  assign n2913 = ( n1407 & n2099 ) | ( n1407 & n2230 ) | ( n2099 & n2230 ) ;
  assign n2914 = n2913 ^ n1356 ^ n892 ;
  assign n2918 = n2917 ^ n2915 ^ n2914 ;
  assign n2924 = n946 ^ n534 ^ 1'b0 ;
  assign n2925 = n2924 ^ n2014 ^ 1'b0 ;
  assign n2926 = x52 & ~n2925 ;
  assign n2920 = ( n1354 & n1696 ) | ( n1354 & ~n2690 ) | ( n1696 & ~n2690 ) ;
  assign n2921 = n899 & ~n2920 ;
  assign n2922 = ~n701 & n2921 ;
  assign n2919 = n2027 | n2452 ;
  assign n2923 = n2922 ^ n2919 ^ 1'b0 ;
  assign n2927 = n2926 ^ n2923 ^ x225 ;
  assign n2928 = ( ~x141 & x161 ) | ( ~x141 & n1346 ) | ( x161 & n1346 ) ;
  assign n2929 = ~n2461 & n2662 ;
  assign n2930 = n2929 ^ x212 ^ 1'b0 ;
  assign n2931 = ( n792 & ~n2928 ) | ( n792 & n2930 ) | ( ~n2928 & n2930 ) ;
  assign n2932 = n2931 ^ n570 ^ x126 ;
  assign n2933 = n954 & ~n2335 ;
  assign n2934 = ( ~n648 & n1157 ) | ( ~n648 & n2933 ) | ( n1157 & n2933 ) ;
  assign n2935 = n268 & n2094 ;
  assign n2936 = ( ~n461 & n2512 ) | ( ~n461 & n2935 ) | ( n2512 & n2935 ) ;
  assign n2937 = n428 & ~n2936 ;
  assign n2938 = n2937 ^ n1331 ^ 1'b0 ;
  assign n2939 = n2097 & ~n2938 ;
  assign n2940 = n1039 | n1932 ;
  assign n2941 = x56 & ~n1923 ;
  assign n2942 = n1359 & n2941 ;
  assign n2943 = n374 & ~n2942 ;
  assign n2944 = ( n746 & ~n1670 ) | ( n746 & n2943 ) | ( ~n1670 & n2943 ) ;
  assign n2945 = n1230 ^ x22 ^ 1'b0 ;
  assign n2946 = ( n1279 & ~n1475 ) | ( n1279 & n2945 ) | ( ~n1475 & n2945 ) ;
  assign n2947 = ( n2940 & n2944 ) | ( n2940 & ~n2946 ) | ( n2944 & ~n2946 ) ;
  assign n2948 = n2814 ^ n460 ^ n345 ;
  assign n2949 = n1728 ^ n1583 ^ x114 ;
  assign n2950 = n2949 ^ n2458 ^ n2111 ;
  assign n2951 = ( ~n510 & n1537 ) | ( ~n510 & n2950 ) | ( n1537 & n2950 ) ;
  assign n2953 = ( n865 & n946 ) | ( n865 & n2295 ) | ( n946 & n2295 ) ;
  assign n2952 = n965 ^ n745 ^ n499 ;
  assign n2954 = n2953 ^ n2952 ^ 1'b0 ;
  assign n2955 = n2147 & ~n2954 ;
  assign n2956 = n692 | n2955 ;
  assign n2957 = n2956 ^ n2664 ^ 1'b0 ;
  assign n2958 = n672 | n1834 ;
  assign n2959 = n2958 ^ n1604 ^ n1262 ;
  assign n2960 = ~n1484 & n2959 ;
  assign n2961 = n1865 ^ x92 ^ 1'b0 ;
  assign n2962 = n2302 & n2961 ;
  assign n2963 = n2962 ^ n509 ^ x31 ;
  assign n2964 = n2963 ^ n2504 ^ n774 ;
  assign n2965 = x119 & n1718 ;
  assign n2966 = n710 & n1730 ;
  assign n2967 = n2966 ^ n883 ^ 1'b0 ;
  assign n2968 = ( n1481 & n2965 ) | ( n1481 & ~n2967 ) | ( n2965 & ~n2967 ) ;
  assign n2974 = n1003 ^ x138 ^ 1'b0 ;
  assign n2975 = n1431 & n2974 ;
  assign n2976 = ( x246 & n2942 ) | ( x246 & n2975 ) | ( n2942 & n2975 ) ;
  assign n2977 = n2976 ^ n626 ^ 1'b0 ;
  assign n2970 = x184 & ~n737 ;
  assign n2969 = ~n601 & n2084 ;
  assign n2971 = n2970 ^ n2969 ^ 1'b0 ;
  assign n2972 = ~n1395 & n2230 ;
  assign n2973 = n2971 & n2972 ;
  assign n2978 = n2977 ^ n2973 ^ n1228 ;
  assign n2979 = ( n381 & n938 ) | ( n381 & n2187 ) | ( n938 & n2187 ) ;
  assign n2980 = n2060 ^ n876 ^ x230 ;
  assign n2981 = ( n932 & n1239 ) | ( n932 & ~n2980 ) | ( n1239 & ~n2980 ) ;
  assign n2982 = n2979 & n2981 ;
  assign n2983 = ~n256 & n2982 ;
  assign n2986 = n976 | n1923 ;
  assign n2987 = n2430 ^ n2084 ^ x28 ;
  assign n2988 = ( n333 & ~n2986 ) | ( n333 & n2987 ) | ( ~n2986 & n2987 ) ;
  assign n2989 = x226 & n1910 ;
  assign n2990 = ~n310 & n2989 ;
  assign n2991 = ( n275 & n817 ) | ( n275 & n2909 ) | ( n817 & n2909 ) ;
  assign n2992 = ( n2988 & ~n2990 ) | ( n2988 & n2991 ) | ( ~n2990 & n2991 ) ;
  assign n2984 = ( ~n264 & n1189 ) | ( ~n264 & n1486 ) | ( n1189 & n1486 ) ;
  assign n2985 = n305 & ~n2984 ;
  assign n2993 = n2992 ^ n2985 ^ n1712 ;
  assign n2994 = ( x212 & n1251 ) | ( x212 & ~n2993 ) | ( n1251 & ~n2993 ) ;
  assign n2995 = n992 ^ x227 ^ 1'b0 ;
  assign n2996 = ~n1800 & n2995 ;
  assign n2997 = n2996 ^ n1154 ^ n977 ;
  assign n3000 = n795 ^ x157 ^ x67 ;
  assign n2999 = n1616 ^ n631 ^ 1'b0 ;
  assign n3001 = n3000 ^ n2999 ^ 1'b0 ;
  assign n3002 = n2644 & n3001 ;
  assign n2998 = n1553 & n2367 ;
  assign n3003 = n3002 ^ n2998 ^ 1'b0 ;
  assign n3004 = n3003 ^ n473 ^ 1'b0 ;
  assign n3006 = ( n1129 & n1198 ) | ( n1129 & ~n2709 ) | ( n1198 & ~n2709 ) ;
  assign n3005 = ( n445 & n1696 ) | ( n445 & n2165 ) | ( n1696 & n2165 ) ;
  assign n3007 = n3006 ^ n3005 ^ n883 ;
  assign n3008 = n1685 ^ n1410 ^ n447 ;
  assign n3009 = x165 & n2934 ;
  assign n3010 = n2317 & n3009 ;
  assign n3011 = ( n599 & ~n655 ) | ( n599 & n986 ) | ( ~n655 & n986 ) ;
  assign n3012 = n1569 | n2886 ;
  assign n3013 = n3012 ^ n2212 ^ 1'b0 ;
  assign n3014 = ~n953 & n1632 ;
  assign n3015 = n3013 & n3014 ;
  assign n3016 = n990 ^ n836 ^ 1'b0 ;
  assign n3017 = n3016 ^ n1139 ^ 1'b0 ;
  assign n3018 = x29 & ~n2069 ;
  assign n3019 = n1840 ^ n275 ^ 1'b0 ;
  assign n3020 = n2878 | n3019 ;
  assign n3021 = n1076 & ~n3020 ;
  assign n3022 = ~n1172 & n2979 ;
  assign n3023 = n1155 & ~n3022 ;
  assign n3024 = n3021 & n3023 ;
  assign n3025 = ~n1314 & n2503 ;
  assign n3026 = ~n1916 & n2561 ;
  assign n3027 = n843 & n2349 ;
  assign n3028 = n544 & n3027 ;
  assign n3029 = n3028 ^ n1536 ^ n802 ;
  assign n3030 = n808 & ~n3029 ;
  assign n3031 = ~n1411 & n3030 ;
  assign n3032 = ( n1113 & n2820 ) | ( n1113 & ~n3031 ) | ( n2820 & ~n3031 ) ;
  assign n3033 = n3032 ^ n2633 ^ n1791 ;
  assign n3037 = ( n267 & n636 ) | ( n267 & n1946 ) | ( n636 & n1946 ) ;
  assign n3038 = n1566 | n3037 ;
  assign n3039 = n736 | n3038 ;
  assign n3034 = n1841 ^ n856 ^ x164 ;
  assign n3035 = n2004 | n3034 ;
  assign n3036 = n1599 | n3035 ;
  assign n3040 = n3039 ^ n3036 ^ 1'b0 ;
  assign n3041 = ~n1428 & n1680 ;
  assign n3042 = n3041 ^ x108 ^ 1'b0 ;
  assign n3043 = ( ~n1103 & n1722 ) | ( ~n1103 & n3042 ) | ( n1722 & n3042 ) ;
  assign n3044 = n2899 ^ n547 ^ 1'b0 ;
  assign n3045 = x224 & ~n1370 ;
  assign n3046 = ~n3044 & n3045 ;
  assign n3047 = n2084 & n3046 ;
  assign n3048 = n1815 | n1980 ;
  assign n3049 = n754 | n3048 ;
  assign n3050 = n3049 ^ n1905 ^ n972 ;
  assign n3051 = x50 & ~x223 ;
  assign n3052 = ( ~n1485 & n1937 ) | ( ~n1485 & n2829 ) | ( n1937 & n2829 ) ;
  assign n3053 = n3052 ^ n1384 ^ 1'b0 ;
  assign n3054 = n3051 | n3053 ;
  assign n3055 = ( n898 & ~n3050 ) | ( n898 & n3054 ) | ( ~n3050 & n3054 ) ;
  assign n3056 = n2858 ^ n2337 ^ n456 ;
  assign n3057 = ( ~n712 & n2139 ) | ( ~n712 & n3056 ) | ( n2139 & n3056 ) ;
  assign n3058 = n742 ^ n678 ^ n376 ;
  assign n3059 = n3058 ^ n885 ^ 1'b0 ;
  assign n3060 = n3059 ^ n1569 ^ 1'b0 ;
  assign n3061 = n977 ^ n296 ^ x249 ;
  assign n3063 = x200 & n1946 ;
  assign n3064 = ~n1241 & n3063 ;
  assign n3062 = ~n1150 & n1222 ;
  assign n3065 = n3064 ^ n3062 ^ 1'b0 ;
  assign n3066 = ( n874 & n3061 ) | ( n874 & n3065 ) | ( n3061 & n3065 ) ;
  assign n3067 = n2539 & n3066 ;
  assign n3068 = n3060 & ~n3067 ;
  assign n3069 = n1611 ^ n1482 ^ n1282 ;
  assign n3070 = n1205 & n1895 ;
  assign n3071 = ( ~n2659 & n3069 ) | ( ~n2659 & n3070 ) | ( n3069 & n3070 ) ;
  assign n3072 = n741 ^ x118 ^ 1'b0 ;
  assign n3073 = x113 & n3072 ;
  assign n3074 = ~n2360 & n3073 ;
  assign n3075 = n3074 ^ x222 ^ 1'b0 ;
  assign n3076 = n3075 ^ n2657 ^ n1950 ;
  assign n3077 = n3076 ^ n2587 ^ 1'b0 ;
  assign n3078 = n498 & ~n3077 ;
  assign n3079 = n879 & n3078 ;
  assign n3080 = ~n3071 & n3079 ;
  assign n3081 = n2087 ^ n1114 ^ 1'b0 ;
  assign n3082 = n3081 ^ n370 ^ 1'b0 ;
  assign n3083 = n739 | n3082 ;
  assign n3084 = ( n738 & ~n1049 ) | ( n738 & n2500 ) | ( ~n1049 & n2500 ) ;
  assign n3085 = ~x39 & n3084 ;
  assign n3086 = n939 & n3039 ;
  assign n3087 = n3086 ^ n1108 ^ 1'b0 ;
  assign n3088 = x127 & n2471 ;
  assign n3089 = ~n1794 & n3088 ;
  assign n3090 = n1400 | n3089 ;
  assign n3091 = n2013 ^ n711 ^ 1'b0 ;
  assign n3092 = n838 & ~n3091 ;
  assign n3093 = ( n2722 & n3090 ) | ( n2722 & n3092 ) | ( n3090 & n3092 ) ;
  assign n3094 = ( n802 & n1135 ) | ( n802 & n1164 ) | ( n1135 & n1164 ) ;
  assign n3095 = ( x223 & ~n688 ) | ( x223 & n3094 ) | ( ~n688 & n3094 ) ;
  assign n3096 = n1266 | n1833 ;
  assign n3097 = n3095 | n3096 ;
  assign n3098 = n3097 ^ n1523 ^ 1'b0 ;
  assign n3099 = n393 & n3098 ;
  assign n3100 = ~n781 & n1140 ;
  assign n3101 = ~n2090 & n3100 ;
  assign n3102 = n3101 ^ n499 ^ 1'b0 ;
  assign n3103 = n1131 & ~n3102 ;
  assign n3104 = n3103 ^ n890 ^ 1'b0 ;
  assign n3105 = n3099 & ~n3104 ;
  assign n3107 = n1545 ^ x107 ^ x9 ;
  assign n3106 = ( n1330 & n2107 ) | ( n1330 & n2803 ) | ( n2107 & n2803 ) ;
  assign n3108 = n3107 ^ n3106 ^ 1'b0 ;
  assign n3109 = n2757 & n3108 ;
  assign n3110 = n1644 ^ n1291 ^ n1187 ;
  assign n3111 = n2309 ^ n2191 ^ 1'b0 ;
  assign n3112 = ( n771 & n3110 ) | ( n771 & ~n3111 ) | ( n3110 & ~n3111 ) ;
  assign n3120 = n704 | n1123 ;
  assign n3121 = n1407 | n3120 ;
  assign n3122 = n3121 ^ n1647 ^ 1'b0 ;
  assign n3116 = ( x249 & ~n1685 ) | ( x249 & n2812 ) | ( ~n1685 & n2812 ) ;
  assign n3117 = n3116 ^ n1940 ^ n1584 ;
  assign n3118 = ~n268 & n3117 ;
  assign n3119 = n3118 ^ n439 ^ 1'b0 ;
  assign n3113 = n1909 ^ x127 ^ 1'b0 ;
  assign n3114 = n3113 ^ n3089 ^ n722 ;
  assign n3115 = n3114 ^ n1675 ^ n1187 ;
  assign n3123 = n3122 ^ n3119 ^ n3115 ;
  assign n3124 = n599 & ~n1813 ;
  assign n3125 = n3124 ^ n2278 ^ n2043 ;
  assign n3126 = n2308 ^ n311 ^ x54 ;
  assign n3127 = n3126 ^ n1356 ^ 1'b0 ;
  assign n3128 = n1344 | n3127 ;
  assign n3129 = ( n2118 & n2340 ) | ( n2118 & ~n2755 ) | ( n2340 & ~n2755 ) ;
  assign n3130 = ~n443 & n3129 ;
  assign n3131 = ~n3128 & n3130 ;
  assign n3132 = n2360 & n3131 ;
  assign n3133 = n3132 ^ n550 ^ 1'b0 ;
  assign n3134 = n453 ^ x89 ^ 1'b0 ;
  assign n3135 = n2918 & n3134 ;
  assign n3136 = ~n324 & n3135 ;
  assign n3137 = x247 & ~n2214 ;
  assign n3138 = n3137 ^ n1249 ^ 1'b0 ;
  assign n3139 = ( n1666 & ~n1821 ) | ( n1666 & n3138 ) | ( ~n1821 & n3138 ) ;
  assign n3140 = ( ~n1717 & n2238 ) | ( ~n1717 & n2247 ) | ( n2238 & n2247 ) ;
  assign n3141 = n3140 ^ n2701 ^ 1'b0 ;
  assign n3143 = ( n618 & n943 ) | ( n618 & ~n1025 ) | ( n943 & ~n1025 ) ;
  assign n3142 = n2812 ^ n1003 ^ n436 ;
  assign n3144 = n3143 ^ n3142 ^ n2095 ;
  assign n3145 = n1171 ^ n891 ^ n618 ;
  assign n3146 = ( n802 & n999 ) | ( n802 & n3145 ) | ( n999 & n3145 ) ;
  assign n3147 = n3146 ^ n2756 ^ n1408 ;
  assign n3148 = n1039 ^ n386 ^ 1'b0 ;
  assign n3149 = ( ~n550 & n662 ) | ( ~n550 & n3148 ) | ( n662 & n3148 ) ;
  assign n3153 = n1295 ^ n579 ^ 1'b0 ;
  assign n3154 = n1988 & n3153 ;
  assign n3150 = n750 ^ n332 ^ 1'b0 ;
  assign n3151 = n697 | n3150 ;
  assign n3152 = n669 & ~n3151 ;
  assign n3155 = n3154 ^ n3152 ^ n2999 ;
  assign n3156 = n2229 | n3017 ;
  assign n3157 = n1822 ^ n1156 ^ n857 ;
  assign n3158 = x158 & n511 ;
  assign n3159 = ~n1236 & n3158 ;
  assign n3160 = n3157 & ~n3159 ;
  assign n3161 = ( n282 & ~n1618 ) | ( n282 & n3037 ) | ( ~n1618 & n3037 ) ;
  assign n3162 = n3160 | n3161 ;
  assign n3163 = n853 & ~n2421 ;
  assign n3164 = ( ~n1923 & n2829 ) | ( ~n1923 & n3163 ) | ( n2829 & n3163 ) ;
  assign n3168 = n1156 & ~n2035 ;
  assign n3169 = n3168 ^ x201 ^ 1'b0 ;
  assign n3165 = n775 ^ x219 ^ 1'b0 ;
  assign n3166 = n654 | n3165 ;
  assign n3167 = n3166 ^ n1635 ^ 1'b0 ;
  assign n3170 = n3169 ^ n3167 ^ 1'b0 ;
  assign n3171 = n2354 & ~n3170 ;
  assign n3172 = n1634 ^ x132 ^ 1'b0 ;
  assign n3173 = n1627 ^ n1518 ^ 1'b0 ;
  assign n3174 = n2418 ^ x71 ^ 1'b0 ;
  assign n3175 = n544 | n3174 ;
  assign n3176 = n3175 ^ n1190 ^ 1'b0 ;
  assign n3177 = n2574 ^ n1245 ^ x90 ;
  assign n3180 = n719 ^ x213 ^ 1'b0 ;
  assign n3181 = x140 & n3180 ;
  assign n3182 = n1225 ^ n911 ^ n325 ;
  assign n3183 = n3182 ^ n1650 ^ 1'b0 ;
  assign n3184 = n3181 & n3183 ;
  assign n3185 = ( n974 & ~n995 ) | ( n974 & n3184 ) | ( ~n995 & n3184 ) ;
  assign n3186 = n3185 ^ n2327 ^ n324 ;
  assign n3178 = n1644 ^ n1043 ^ n512 ;
  assign n3179 = n3178 ^ n913 ^ 1'b0 ;
  assign n3187 = n3186 ^ n3179 ^ n2736 ;
  assign n3188 = ( n3176 & n3177 ) | ( n3176 & ~n3187 ) | ( n3177 & ~n3187 ) ;
  assign n3189 = ( n512 & n1099 ) | ( n512 & n1300 ) | ( n1099 & n1300 ) ;
  assign n3190 = ( x87 & n646 ) | ( x87 & n2204 ) | ( n646 & n2204 ) ;
  assign n3191 = n3190 ^ n1078 ^ n797 ;
  assign n3192 = n2799 ^ n1543 ^ 1'b0 ;
  assign n3193 = n1865 & ~n3192 ;
  assign n3194 = ~n639 & n3193 ;
  assign n3195 = n1344 & n3194 ;
  assign n3196 = n3195 ^ n3103 ^ n2034 ;
  assign n3197 = n2173 ^ n1731 ^ 1'b0 ;
  assign n3198 = ~n3196 & n3197 ;
  assign n3201 = ( n1069 & n1113 ) | ( n1069 & n1767 ) | ( n1113 & n1767 ) ;
  assign n3199 = n441 & n2450 ;
  assign n3200 = ~n1548 & n3199 ;
  assign n3202 = n3201 ^ n3200 ^ x252 ;
  assign n3203 = n784 & n1758 ;
  assign n3204 = n736 & n3203 ;
  assign n3205 = n1307 & ~n3204 ;
  assign n3206 = ~n1899 & n3205 ;
  assign n3207 = n561 & n668 ;
  assign n3208 = n3207 ^ x72 ^ 1'b0 ;
  assign n3209 = ( n689 & n1175 ) | ( n689 & n1910 ) | ( n1175 & n1910 ) ;
  assign n3210 = ( ~n425 & n945 ) | ( ~n425 & n3209 ) | ( n945 & n3209 ) ;
  assign n3213 = n2134 ^ n320 ^ x121 ;
  assign n3211 = n393 & ~n1261 ;
  assign n3212 = n3211 ^ n3178 ^ n1211 ;
  assign n3214 = n3213 ^ n3212 ^ n2828 ;
  assign n3215 = ( n3208 & ~n3210 ) | ( n3208 & n3214 ) | ( ~n3210 & n3214 ) ;
  assign n3216 = n1557 & n2076 ;
  assign n3217 = n2755 ^ n1164 ^ x2 ;
  assign n3218 = n3217 ^ n1424 ^ 1'b0 ;
  assign n3219 = ( ~n3121 & n3216 ) | ( ~n3121 & n3218 ) | ( n3216 & n3218 ) ;
  assign n3220 = n1381 ^ n290 ^ 1'b0 ;
  assign n3221 = ( x184 & n678 ) | ( x184 & ~n802 ) | ( n678 & ~n802 ) ;
  assign n3222 = n1460 ^ n1128 ^ 1'b0 ;
  assign n3223 = n3221 | n3222 ;
  assign n3225 = n1155 ^ n795 ^ n310 ;
  assign n3224 = n2562 ^ n1095 ^ 1'b0 ;
  assign n3226 = n3225 ^ n3224 ^ 1'b0 ;
  assign n3227 = n3226 ^ x130 ^ 1'b0 ;
  assign n3228 = x209 & ~n3227 ;
  assign n3229 = n3216 ^ n2180 ^ n2132 ;
  assign n3230 = ~n257 & n401 ;
  assign n3231 = n3230 ^ n3126 ^ n1336 ;
  assign n3232 = ( n378 & n558 ) | ( n378 & ~n3225 ) | ( n558 & ~n3225 ) ;
  assign n3233 = ( x61 & x247 ) | ( x61 & n742 ) | ( x247 & n742 ) ;
  assign n3234 = n3233 ^ n2308 ^ x150 ;
  assign n3235 = n3234 ^ n1787 ^ n1494 ;
  assign n3236 = ( n3119 & n3232 ) | ( n3119 & ~n3235 ) | ( n3232 & ~n3235 ) ;
  assign n3244 = n1943 ^ x126 ^ 1'b0 ;
  assign n3245 = ~n418 & n3244 ;
  assign n3239 = x1 & x16 ;
  assign n3240 = ~n414 & n3239 ;
  assign n3241 = ( x203 & ~n2117 ) | ( x203 & n3240 ) | ( ~n2117 & n3240 ) ;
  assign n3242 = n3241 ^ n1037 ^ x142 ;
  assign n3243 = ( n1067 & n1206 ) | ( n1067 & ~n3242 ) | ( n1206 & ~n3242 ) ;
  assign n3246 = n3245 ^ n3243 ^ n408 ;
  assign n3247 = n3246 ^ n617 ^ 1'b0 ;
  assign n3248 = n3247 ^ n833 ^ x161 ;
  assign n3237 = n547 | n939 ;
  assign n3238 = n3052 & ~n3237 ;
  assign n3249 = n3248 ^ n3238 ^ 1'b0 ;
  assign n3250 = n493 | n512 ;
  assign n3251 = x187 & ~n1370 ;
  assign n3252 = ~n530 & n3251 ;
  assign n3253 = ( n1050 & n3250 ) | ( n1050 & n3252 ) | ( n3250 & n3252 ) ;
  assign n3254 = n2413 & n3253 ;
  assign n3255 = ( n665 & n2701 ) | ( n665 & n2976 ) | ( n2701 & n2976 ) ;
  assign n3256 = n2924 ^ n362 ^ 1'b0 ;
  assign n3257 = n1003 | n2018 ;
  assign n3258 = ( n262 & n3256 ) | ( n262 & n3257 ) | ( n3256 & n3257 ) ;
  assign n3261 = ~n1157 & n1257 ;
  assign n3262 = n3261 ^ n1731 ^ n1217 ;
  assign n3259 = n1733 ^ n980 ^ 1'b0 ;
  assign n3260 = n2704 & n3259 ;
  assign n3263 = n3262 ^ n3260 ^ 1'b0 ;
  assign n3264 = ( n876 & ~n1370 ) | ( n876 & n2922 ) | ( ~n1370 & n2922 ) ;
  assign n3265 = n3264 ^ n512 ^ 1'b0 ;
  assign n3266 = n1629 & ~n3265 ;
  assign n3267 = n1734 ^ n1103 ^ 1'b0 ;
  assign n3268 = ( x150 & n453 ) | ( x150 & n2065 ) | ( n453 & n2065 ) ;
  assign n3269 = n3268 ^ n722 ^ 1'b0 ;
  assign n3270 = n556 ^ n276 ^ 1'b0 ;
  assign n3271 = n695 & n3270 ;
  assign n3272 = ( ~n663 & n3269 ) | ( ~n663 & n3271 ) | ( n3269 & n3271 ) ;
  assign n3274 = x54 & x249 ;
  assign n3275 = n3274 ^ n853 ^ 1'b0 ;
  assign n3276 = ~n1848 & n3275 ;
  assign n3273 = n2965 ^ n2680 ^ n326 ;
  assign n3277 = n3276 ^ n3273 ^ 1'b0 ;
  assign n3278 = ~n739 & n3277 ;
  assign n3282 = n1129 | n1361 ;
  assign n3283 = n1032 & ~n3282 ;
  assign n3284 = n1341 | n3283 ;
  assign n3285 = x108 & ~n3284 ;
  assign n3286 = n2031 ^ n1148 ^ 1'b0 ;
  assign n3287 = n3285 | n3286 ;
  assign n3279 = ( n280 & n332 ) | ( n280 & ~n901 ) | ( n332 & ~n901 ) ;
  assign n3280 = n3279 ^ n2563 ^ n1675 ;
  assign n3281 = n3280 ^ n1865 ^ n989 ;
  assign n3288 = n3287 ^ n3281 ^ n2422 ;
  assign n3289 = n3278 & n3288 ;
  assign n3290 = ~n843 & n3289 ;
  assign n3291 = n1025 ^ n368 ^ 1'b0 ;
  assign n3292 = n652 | n3291 ;
  assign n3293 = n3292 ^ n1766 ^ n1656 ;
  assign n3294 = n3293 ^ n2212 ^ n639 ;
  assign n3295 = n2932 ^ n2302 ^ 1'b0 ;
  assign n3296 = n1653 & n2668 ;
  assign n3297 = n3296 ^ n1546 ^ 1'b0 ;
  assign n3298 = n3297 ^ n2036 ^ n1422 ;
  assign n3299 = n3298 ^ x240 ^ 1'b0 ;
  assign n3300 = ~n502 & n3299 ;
  assign n3301 = n1463 ^ x227 ^ 1'b0 ;
  assign n3302 = n3202 & n3301 ;
  assign n3303 = n3302 ^ n1073 ^ 1'b0 ;
  assign n3304 = n1192 & ~n1300 ;
  assign n3305 = n3304 ^ n860 ^ 1'b0 ;
  assign n3306 = ( n696 & n3199 ) | ( n696 & n3305 ) | ( n3199 & n3305 ) ;
  assign n3307 = n3306 ^ n2097 ^ x144 ;
  assign n3314 = n2482 ^ n1712 ^ n1567 ;
  assign n3310 = n586 | n2349 ;
  assign n3308 = ( x166 & n333 ) | ( x166 & ~n1065 ) | ( n333 & ~n1065 ) ;
  assign n3309 = n3308 ^ n1504 ^ n560 ;
  assign n3311 = n3310 ^ n3309 ^ n2858 ;
  assign n3312 = n2952 ^ n1822 ^ 1'b0 ;
  assign n3313 = n3311 | n3312 ;
  assign n3315 = n3314 ^ n3313 ^ n879 ;
  assign n3317 = n896 ^ x62 ^ 1'b0 ;
  assign n3318 = n3317 ^ n1039 ^ 1'b0 ;
  assign n3319 = n528 & ~n3318 ;
  assign n3316 = n2469 & ~n3101 ;
  assign n3320 = n3319 ^ n3316 ^ 1'b0 ;
  assign n3321 = n425 & n1458 ;
  assign n3322 = n3321 ^ x72 ^ 1'b0 ;
  assign n3323 = n3322 ^ n2117 ^ n1353 ;
  assign n3324 = ( n652 & n2417 ) | ( n652 & n3323 ) | ( n2417 & n3323 ) ;
  assign n3325 = n3324 ^ n948 ^ 1'b0 ;
  assign n3326 = n1721 ^ n491 ^ 1'b0 ;
  assign n3327 = ( n1236 & ~n3243 ) | ( n1236 & n3326 ) | ( ~n3243 & n3326 ) ;
  assign n3328 = n1721 | n1957 ;
  assign n3329 = n2537 | n3328 ;
  assign n3330 = n2160 | n3329 ;
  assign n3331 = ( n834 & n935 ) | ( n834 & ~n1420 ) | ( n935 & ~n1420 ) ;
  assign n3332 = n304 | n3331 ;
  assign n3333 = n959 | n3332 ;
  assign n3334 = ~n2396 & n3333 ;
  assign n3335 = n523 & n3334 ;
  assign n3336 = n2740 | n3335 ;
  assign n3337 = n1644 & ~n3336 ;
  assign n3340 = n2215 ^ n1831 ^ n536 ;
  assign n3338 = n912 ^ x45 ^ 1'b0 ;
  assign n3339 = n465 & ~n3338 ;
  assign n3341 = n3340 ^ n3339 ^ 1'b0 ;
  assign n3342 = n2640 & n3341 ;
  assign n3348 = x36 | n280 ;
  assign n3345 = x91 & ~n1201 ;
  assign n3346 = n3345 ^ n1276 ^ 1'b0 ;
  assign n3347 = ( n767 & n2002 ) | ( n767 & ~n3346 ) | ( n2002 & ~n3346 ) ;
  assign n3349 = n3348 ^ n3347 ^ n1046 ;
  assign n3343 = n1450 ^ n1258 ^ n933 ;
  assign n3344 = ( n580 & n3065 ) | ( n580 & ~n3343 ) | ( n3065 & ~n3343 ) ;
  assign n3350 = n3349 ^ n3344 ^ n2194 ;
  assign n3351 = n2985 ^ n1856 ^ 1'b0 ;
  assign n3358 = n1513 & n2198 ;
  assign n3355 = ( x150 & n386 ) | ( x150 & ~n436 ) | ( n386 & ~n436 ) ;
  assign n3356 = ~n1433 & n3355 ;
  assign n3357 = ~x6 & n3356 ;
  assign n3352 = ~x25 & n2628 ;
  assign n3353 = n1289 ^ n750 ^ 1'b0 ;
  assign n3354 = ( n681 & n3352 ) | ( n681 & ~n3353 ) | ( n3352 & ~n3353 ) ;
  assign n3359 = n3358 ^ n3357 ^ n3354 ;
  assign n3360 = n391 ^ x126 ^ 1'b0 ;
  assign n3361 = n1041 | n1304 ;
  assign n3362 = n3360 & ~n3361 ;
  assign n3363 = n1018 ^ n506 ^ x248 ;
  assign n3364 = ( x103 & n277 ) | ( x103 & ~n3363 ) | ( n277 & ~n3363 ) ;
  assign n3365 = n3364 ^ n1209 ^ 1'b0 ;
  assign n3366 = n3365 ^ n526 ^ 1'b0 ;
  assign n3367 = n2892 ^ n1432 ^ 1'b0 ;
  assign n3368 = ( n2715 & ~n3366 ) | ( n2715 & n3367 ) | ( ~n3366 & n3367 ) ;
  assign n3369 = ( n1758 & n1924 ) | ( n1758 & ~n3368 ) | ( n1924 & ~n3368 ) ;
  assign n3370 = ( n347 & ~n1153 ) | ( n347 & n3369 ) | ( ~n1153 & n3369 ) ;
  assign n3371 = ( n2391 & n2697 ) | ( n2391 & ~n3370 ) | ( n2697 & ~n3370 ) ;
  assign n3373 = ( n775 & n1084 ) | ( n775 & n1924 ) | ( n1084 & n1924 ) ;
  assign n3372 = n774 & n2157 ;
  assign n3374 = n3373 ^ n3372 ^ 1'b0 ;
  assign n3375 = n3374 ^ n642 ^ 1'b0 ;
  assign n3379 = ( n374 & n1258 ) | ( n374 & ~n2928 ) | ( n1258 & ~n2928 ) ;
  assign n3380 = ( x228 & ~n467 ) | ( x228 & n3379 ) | ( ~n467 & n3379 ) ;
  assign n3381 = n3380 ^ n2727 ^ 1'b0 ;
  assign n3376 = n2718 ^ n485 ^ 1'b0 ;
  assign n3377 = n1172 & ~n3376 ;
  assign n3378 = ~n1802 & n3377 ;
  assign n3382 = n3381 ^ n3378 ^ 1'b0 ;
  assign n3383 = ( n1086 & ~n2436 ) | ( n1086 & n3382 ) | ( ~n2436 & n3382 ) ;
  assign n3384 = ~n1751 & n3383 ;
  assign n3385 = n290 & n3384 ;
  assign n3390 = x243 & n853 ;
  assign n3391 = ~n2117 & n3390 ;
  assign n3386 = ~n678 & n2532 ;
  assign n3387 = ~x7 & n3386 ;
  assign n3388 = n3387 ^ n1739 ^ x199 ;
  assign n3389 = n2791 | n3388 ;
  assign n3392 = n3391 ^ n3389 ^ 1'b0 ;
  assign n3397 = ( x88 & ~n2417 ) | ( x88 & n3121 ) | ( ~n2417 & n3121 ) ;
  assign n3396 = n1400 & ~n1773 ;
  assign n3398 = n3397 ^ n3396 ^ 1'b0 ;
  assign n3393 = n2393 | n2679 ;
  assign n3394 = n3393 ^ n2915 ^ 1'b0 ;
  assign n3395 = ~n2775 & n3394 ;
  assign n3399 = n3398 ^ n3395 ^ 1'b0 ;
  assign n3400 = ( n1294 & n1915 ) | ( n1294 & n3273 ) | ( n1915 & n3273 ) ;
  assign n3401 = n3400 ^ n603 ^ 1'b0 ;
  assign n3405 = ( ~x54 & n538 ) | ( ~x54 & n569 ) | ( n538 & n569 ) ;
  assign n3406 = n1677 | n3405 ;
  assign n3402 = n1096 ^ n448 ^ n364 ;
  assign n3403 = ~n950 & n3402 ;
  assign n3404 = n3403 ^ n1610 ^ n1012 ;
  assign n3407 = n3406 ^ n3404 ^ n1352 ;
  assign n3408 = n3134 ^ n2451 ^ n778 ;
  assign n3409 = n1329 ^ n1010 ^ 1'b0 ;
  assign n3410 = n3408 & n3409 ;
  assign n3411 = ( n1487 & n3397 ) | ( n1487 & ~n3410 ) | ( n3397 & ~n3410 ) ;
  assign n3412 = n879 ^ n431 ^ n399 ;
  assign n3413 = n3412 ^ x45 ^ 1'b0 ;
  assign n3414 = n1220 & ~n2102 ;
  assign n3415 = n3414 ^ n3193 ^ 1'b0 ;
  assign n3416 = ~n1364 & n1919 ;
  assign n3417 = n3416 ^ n2582 ^ n1255 ;
  assign n3418 = ~n1359 & n2814 ;
  assign n3419 = n3418 ^ n721 ^ 1'b0 ;
  assign n3420 = n3417 | n3419 ;
  assign n3421 = n1649 & n2295 ;
  assign n3425 = n1429 ^ n1261 ^ n880 ;
  assign n3424 = n894 & n1107 ;
  assign n3426 = n3425 ^ n3424 ^ 1'b0 ;
  assign n3427 = n3426 ^ n1670 ^ 1'b0 ;
  assign n3422 = x148 & n559 ;
  assign n3423 = ~n429 & n3422 ;
  assign n3428 = n3427 ^ n3423 ^ 1'b0 ;
  assign n3429 = n1466 ^ n708 ^ 1'b0 ;
  assign n3430 = n489 & n3429 ;
  assign n3431 = n2325 ^ n1979 ^ 1'b0 ;
  assign n3432 = ( ~x19 & n256 ) | ( ~x19 & n350 ) | ( n256 & n350 ) ;
  assign n3433 = ( n787 & n2204 ) | ( n787 & ~n3432 ) | ( n2204 & ~n3432 ) ;
  assign n3435 = n962 | n2992 ;
  assign n3434 = n1836 & n3198 ;
  assign n3436 = n3435 ^ n3434 ^ 1'b0 ;
  assign n3437 = n3246 ^ n476 ^ 1'b0 ;
  assign n3438 = n439 ^ x63 ^ 1'b0 ;
  assign n3439 = x206 & n3438 ;
  assign n3440 = ( ~n602 & n1020 ) | ( ~n602 & n3439 ) | ( n1020 & n3439 ) ;
  assign n3441 = ( x125 & n529 ) | ( x125 & ~n3382 ) | ( n529 & ~n3382 ) ;
  assign n3442 = ~n3440 & n3441 ;
  assign n3443 = n3437 & n3442 ;
  assign n3444 = n3443 ^ n3067 ^ n2188 ;
  assign n3445 = n2845 ^ n1404 ^ 1'b0 ;
  assign n3447 = n1523 & n2421 ;
  assign n3448 = n2069 & n3447 ;
  assign n3446 = ( n752 & ~n1662 ) | ( n752 & n2562 ) | ( ~n1662 & n2562 ) ;
  assign n3449 = n3448 ^ n3446 ^ n2158 ;
  assign n3450 = n3445 | n3449 ;
  assign n3451 = n2570 ^ n488 ^ 1'b0 ;
  assign n3452 = n3263 & n3451 ;
  assign n3453 = x159 & ~n2224 ;
  assign n3454 = ( ~n345 & n2185 ) | ( ~n345 & n3453 ) | ( n2185 & n3453 ) ;
  assign n3455 = x172 & n916 ;
  assign n3456 = ( n2889 & n2967 ) | ( n2889 & ~n3455 ) | ( n2967 & ~n3455 ) ;
  assign n3463 = x184 & n1172 ;
  assign n3464 = n1385 & n3463 ;
  assign n3465 = ( x213 & n1966 ) | ( x213 & n3464 ) | ( n1966 & n3464 ) ;
  assign n3466 = n3465 ^ n856 ^ n800 ;
  assign n3457 = n2790 ^ n879 ^ 1'b0 ;
  assign n3458 = ( ~n531 & n542 ) | ( ~n531 & n935 ) | ( n542 & n935 ) ;
  assign n3459 = n3458 ^ n1548 ^ n797 ;
  assign n3460 = ( x99 & ~n3457 ) | ( x99 & n3459 ) | ( ~n3457 & n3459 ) ;
  assign n3461 = n796 | n2127 ;
  assign n3462 = n3460 & ~n3461 ;
  assign n3467 = n3466 ^ n3462 ^ n1621 ;
  assign n3468 = ~x214 & n1165 ;
  assign n3469 = x78 & ~n3468 ;
  assign n3470 = n3469 ^ x97 ^ 1'b0 ;
  assign n3471 = n759 ^ n754 ^ 1'b0 ;
  assign n3478 = n1182 & n2644 ;
  assign n3479 = ~n331 & n3478 ;
  assign n3480 = ( ~n565 & n1588 ) | ( ~n565 & n3479 ) | ( n1588 & n3479 ) ;
  assign n3481 = n3056 ^ n416 ^ 1'b0 ;
  assign n3482 = ( n770 & n3480 ) | ( n770 & n3481 ) | ( n3480 & n3481 ) ;
  assign n3472 = ( x192 & ~n423 ) | ( x192 & n1281 ) | ( ~n423 & n1281 ) ;
  assign n3473 = ~n811 & n3472 ;
  assign n3474 = n3473 ^ n1089 ^ 1'b0 ;
  assign n3475 = ~n342 & n1320 ;
  assign n3476 = n3475 ^ n2118 ^ n1748 ;
  assign n3477 = ~n3474 & n3476 ;
  assign n3483 = n3482 ^ n3477 ^ 1'b0 ;
  assign n3494 = n1736 ^ n911 ^ x91 ;
  assign n3495 = n3494 ^ x146 ^ 1'b0 ;
  assign n3496 = n1890 ^ x225 ^ 1'b0 ;
  assign n3497 = x14 & ~n3496 ;
  assign n3498 = n3495 & n3497 ;
  assign n3493 = ( n676 & n1507 ) | ( n676 & n1556 ) | ( n1507 & n1556 ) ;
  assign n3499 = n3498 ^ n3493 ^ n2453 ;
  assign n3487 = n1981 ^ n1073 ^ n562 ;
  assign n3488 = n1286 ^ n257 ^ 1'b0 ;
  assign n3489 = ~n3487 & n3488 ;
  assign n3490 = ~n2546 & n3489 ;
  assign n3484 = n738 ^ x112 ^ 1'b0 ;
  assign n3485 = n2524 ^ n1669 ^ 1'b0 ;
  assign n3486 = ( n3402 & n3484 ) | ( n3402 & n3485 ) | ( n3484 & n3485 ) ;
  assign n3491 = n3490 ^ n3486 ^ x221 ;
  assign n3492 = n3491 ^ n2695 ^ n2214 ;
  assign n3500 = n3499 ^ n3492 ^ n2009 ;
  assign n3501 = n1583 ^ n526 ^ 1'b0 ;
  assign n3502 = n3501 ^ n3385 ^ 1'b0 ;
  assign n3503 = ~x72 & n508 ;
  assign n3506 = n748 & n1288 ;
  assign n3507 = n3506 ^ n1971 ^ 1'b0 ;
  assign n3504 = n2398 ^ n2098 ^ n1620 ;
  assign n3505 = n3504 ^ n984 ^ x230 ;
  assign n3508 = n3507 ^ n3505 ^ 1'b0 ;
  assign n3509 = n3503 | n3508 ;
  assign n3510 = n698 & ~n3216 ;
  assign n3514 = n1499 & ~n1722 ;
  assign n3515 = n2770 | n3514 ;
  assign n3511 = x15 & n410 ;
  assign n3512 = n2681 ^ n464 ^ 1'b0 ;
  assign n3513 = ~n3511 & n3512 ;
  assign n3516 = n3515 ^ n3513 ^ 1'b0 ;
  assign n3517 = n610 ^ n606 ^ 1'b0 ;
  assign n3518 = n329 & ~n1766 ;
  assign n3519 = n1720 & n2316 ;
  assign n3520 = n1449 & n3519 ;
  assign n3521 = n3518 | n3520 ;
  assign n3522 = n3517 & ~n3521 ;
  assign n3523 = n3522 ^ n1784 ^ x198 ;
  assign n3524 = ~n582 & n3481 ;
  assign n3525 = n3524 ^ n1786 ^ 1'b0 ;
  assign n3526 = n3525 ^ n1162 ^ 1'b0 ;
  assign n3527 = ( n556 & n2706 ) | ( n556 & ~n3526 ) | ( n2706 & ~n3526 ) ;
  assign n3528 = n2187 ^ x90 ^ 1'b0 ;
  assign n3529 = x185 & n3528 ;
  assign n3530 = n275 & n1313 ;
  assign n3531 = x194 ^ x113 ^ 1'b0 ;
  assign n3532 = n3531 ^ n2295 ^ n594 ;
  assign n3533 = n295 | n1924 ;
  assign n3534 = n920 & ~n3533 ;
  assign n3535 = ( ~n1573 & n3532 ) | ( ~n1573 & n3534 ) | ( n3532 & n3534 ) ;
  assign n3536 = ( n2953 & n3530 ) | ( n2953 & n3535 ) | ( n3530 & n3535 ) ;
  assign n3537 = ( n1055 & n1401 ) | ( n1055 & n3536 ) | ( n1401 & n3536 ) ;
  assign n3539 = n1993 ^ n1832 ^ 1'b0 ;
  assign n3540 = n2714 & n3539 ;
  assign n3538 = n2638 ^ n1268 ^ 1'b0 ;
  assign n3541 = n3540 ^ n3538 ^ 1'b0 ;
  assign n3542 = n2784 | n3541 ;
  assign n3546 = n684 ^ n356 ^ 1'b0 ;
  assign n3543 = n2450 ^ x94 ^ 1'b0 ;
  assign n3544 = ( x209 & ~n474 ) | ( x209 & n1179 ) | ( ~n474 & n1179 ) ;
  assign n3545 = ( ~n1771 & n3543 ) | ( ~n1771 & n3544 ) | ( n3543 & n3544 ) ;
  assign n3547 = n3546 ^ n3545 ^ n2527 ;
  assign n3548 = ~x53 & n3547 ;
  assign n3549 = n2112 ^ n1536 ^ n1333 ;
  assign n3554 = ~x199 & n802 ;
  assign n3550 = ( n1101 & ~n1373 ) | ( n1101 & n1588 ) | ( ~n1373 & n1588 ) ;
  assign n3551 = ~n730 & n1865 ;
  assign n3552 = ~x41 & n3551 ;
  assign n3553 = n3550 | n3552 ;
  assign n3555 = n3554 ^ n3553 ^ 1'b0 ;
  assign n3556 = n3555 ^ n1575 ^ 1'b0 ;
  assign n3557 = n3122 | n3556 ;
  assign n3558 = n1593 & n2814 ;
  assign n3559 = n582 & n3558 ;
  assign n3560 = ( n585 & n3557 ) | ( n585 & n3559 ) | ( n3557 & n3559 ) ;
  assign n3561 = ( x40 & n2292 ) | ( x40 & n2513 ) | ( n2292 & n2513 ) ;
  assign n3562 = n3561 ^ n1179 ^ n412 ;
  assign n3563 = ~n687 & n742 ;
  assign n3564 = n3563 ^ n2605 ^ n1432 ;
  assign n3568 = n1012 ^ n717 ^ 1'b0 ;
  assign n3566 = n1928 ^ n1662 ^ n887 ;
  assign n3567 = n3566 ^ n1390 ^ n1002 ;
  assign n3565 = n1977 ^ n401 ^ n307 ;
  assign n3569 = n3568 ^ n3567 ^ n3565 ;
  assign n3570 = n3146 & ~n3569 ;
  assign n3571 = ~n2097 & n3570 ;
  assign n3572 = n1333 | n1531 ;
  assign n3573 = n3201 | n3572 ;
  assign n3574 = x37 & n3573 ;
  assign n3575 = n3574 ^ n2450 ^ 1'b0 ;
  assign n3577 = n1866 ^ n1834 ^ n337 ;
  assign n3578 = n3577 ^ n1325 ^ 1'b0 ;
  assign n3579 = n2727 & ~n3578 ;
  assign n3576 = ~n275 & n1649 ;
  assign n3580 = n3579 ^ n3576 ^ 1'b0 ;
  assign n3581 = n2017 | n3580 ;
  assign n3582 = n3575 | n3581 ;
  assign n3583 = n3457 ^ n2867 ^ x11 ;
  assign n3584 = n3536 ^ n2583 ^ n560 ;
  assign n3585 = n633 ^ x76 ^ 1'b0 ;
  assign n3586 = ( x103 & ~x130 ) | ( x103 & n473 ) | ( ~x130 & n473 ) ;
  assign n3587 = ( n1671 & n3585 ) | ( n1671 & ~n3586 ) | ( n3585 & ~n3586 ) ;
  assign n3588 = ~n351 & n3587 ;
  assign n3589 = n1364 ^ n508 ^ 1'b0 ;
  assign n3590 = ( x75 & n2199 ) | ( x75 & n2558 ) | ( n2199 & n2558 ) ;
  assign n3591 = n3452 ^ n3437 ^ n1250 ;
  assign n3593 = x8 & ~n1442 ;
  assign n3594 = n3593 ^ n1669 ^ 1'b0 ;
  assign n3595 = n2934 & ~n3594 ;
  assign n3592 = n960 & n1984 ;
  assign n3596 = n3595 ^ n3592 ^ 1'b0 ;
  assign n3597 = n721 & ~n3531 ;
  assign n3598 = ~n984 & n3597 ;
  assign n3599 = n3598 ^ n1089 ^ 1'b0 ;
  assign n3600 = n1516 & ~n3599 ;
  assign n3601 = n2407 ^ n712 ^ n566 ;
  assign n3602 = n3601 ^ n796 ^ 1'b0 ;
  assign n3603 = n513 & ~n3602 ;
  assign n3604 = n3439 ^ n2895 ^ n1518 ;
  assign n3605 = n2992 ^ n2605 ^ 1'b0 ;
  assign n3606 = n2380 & n3605 ;
  assign n3607 = n2003 & ~n3606 ;
  assign n3608 = n2099 & n3607 ;
  assign n3609 = n1171 & ~n1799 ;
  assign n3610 = ~n3187 & n3609 ;
  assign n3611 = n3610 ^ n2609 ^ 1'b0 ;
  assign n3612 = n2813 ^ n2700 ^ n780 ;
  assign n3613 = n3612 ^ n3255 ^ n2807 ;
  assign n3614 = ~n317 & n705 ;
  assign n3615 = ~n692 & n3614 ;
  assign n3616 = ( ~n314 & n708 ) | ( ~n314 & n3615 ) | ( n708 & n3615 ) ;
  assign n3617 = x195 & ~n1025 ;
  assign n3618 = n3617 ^ n2677 ^ 1'b0 ;
  assign n3619 = n3616 & ~n3618 ;
  assign n3620 = ~n3107 & n3619 ;
  assign n3621 = ~n381 & n1683 ;
  assign n3622 = n681 ^ n257 ^ 1'b0 ;
  assign n3623 = ~n3621 & n3622 ;
  assign n3624 = n2748 ^ n1688 ^ n1550 ;
  assign n3625 = ( n324 & ~n3623 ) | ( n324 & n3624 ) | ( ~n3623 & n3624 ) ;
  assign n3628 = x213 & ~n1581 ;
  assign n3629 = n1966 & n3628 ;
  assign n3626 = n708 ^ x77 ^ 1'b0 ;
  assign n3627 = n3626 ^ n1581 ^ x210 ;
  assign n3630 = n3629 ^ n3627 ^ n711 ;
  assign n3636 = n2506 ^ n2397 ^ n1862 ;
  assign n3633 = x218 ^ x38 ^ x29 ;
  assign n3634 = x71 | n3633 ;
  assign n3631 = ~n1366 & n1400 ;
  assign n3632 = n2069 & n3631 ;
  assign n3635 = n3634 ^ n3632 ^ 1'b0 ;
  assign n3637 = n3636 ^ n3635 ^ x56 ;
  assign n3638 = n2154 ^ n333 ^ x38 ;
  assign n3639 = n3638 ^ n972 ^ 1'b0 ;
  assign n3640 = n2419 & n3639 ;
  assign n3641 = n546 ^ x88 ^ 1'b0 ;
  assign n3642 = n2672 & n3641 ;
  assign n3643 = n3450 ^ n1950 ^ x234 ;
  assign n3644 = n3476 ^ n3380 ^ n1474 ;
  assign n3645 = n3644 ^ n2673 ^ n2344 ;
  assign n3646 = ( n1461 & n2451 ) | ( n1461 & ~n3245 ) | ( n2451 & ~n3245 ) ;
  assign n3647 = n1096 | n3646 ;
  assign n3648 = ( x138 & n852 ) | ( x138 & ~n1560 ) | ( n852 & ~n1560 ) ;
  assign n3649 = n3648 ^ n531 ^ x38 ;
  assign n3650 = x143 & n3649 ;
  assign n3651 = ( ~n1713 & n2357 ) | ( ~n1713 & n3650 ) | ( n2357 & n3650 ) ;
  assign n3652 = n3651 ^ n1516 ^ 1'b0 ;
  assign n3653 = n866 & ~n3652 ;
  assign n3654 = n595 & ~n1987 ;
  assign n3655 = n3654 ^ n1650 ^ n817 ;
  assign n3656 = n2106 ^ n868 ^ 1'b0 ;
  assign n3657 = n3655 & n3656 ;
  assign n3658 = n2344 & n3657 ;
  assign n3660 = ( x82 & n1152 ) | ( x82 & ~n1308 ) | ( n1152 & ~n1308 ) ;
  assign n3659 = n979 ^ n713 ^ n471 ;
  assign n3661 = n3660 ^ n3659 ^ n3008 ;
  assign n3662 = n1920 ^ n1824 ^ n950 ;
  assign n3664 = n2448 ^ n1295 ^ x13 ;
  assign n3663 = n2042 ^ n828 ^ n308 ;
  assign n3665 = n3664 ^ n3663 ^ 1'b0 ;
  assign n3666 = n3662 | n3665 ;
  assign n3667 = n2392 | n3666 ;
  assign n3668 = ( n345 & n606 ) | ( n345 & n1260 ) | ( n606 & n1260 ) ;
  assign n3669 = n1544 & ~n3029 ;
  assign n3670 = n2357 & n3669 ;
  assign n3671 = ( n1627 & ~n3668 ) | ( n1627 & n3670 ) | ( ~n3668 & n3670 ) ;
  assign n3674 = n1892 ^ n549 ^ 1'b0 ;
  assign n3675 = n3674 ^ n3211 ^ n508 ;
  assign n3676 = x4 & n2038 ;
  assign n3677 = ~n339 & n3676 ;
  assign n3678 = ( ~x5 & n3675 ) | ( ~x5 & n3677 ) | ( n3675 & n3677 ) ;
  assign n3672 = n3498 ^ n2597 ^ n891 ;
  assign n3673 = ~x155 & n3672 ;
  assign n3679 = n3678 ^ n3673 ^ n741 ;
  assign n3680 = n1540 & ~n3679 ;
  assign n3681 = n3680 ^ n2958 ^ 1'b0 ;
  assign n3682 = n1135 & n2858 ;
  assign n3683 = x233 & n1790 ;
  assign n3684 = ~n3682 & n3683 ;
  assign n3685 = n586 | n3684 ;
  assign n3686 = n2145 | n3685 ;
  assign n3687 = n1686 ^ n1186 ^ 1'b0 ;
  assign n3688 = n1549 ^ n260 ^ 1'b0 ;
  assign n3689 = n3687 & ~n3688 ;
  assign n3690 = n3689 ^ n2546 ^ n1550 ;
  assign n3691 = n3690 ^ n1897 ^ 1'b0 ;
  assign n3692 = n3686 & n3691 ;
  assign n3695 = ~n1998 & n3232 ;
  assign n3696 = n3166 & n3695 ;
  assign n3693 = n1806 & n2152 ;
  assign n3694 = n3693 ^ n1982 ^ 1'b0 ;
  assign n3697 = n3696 ^ n3694 ^ 1'b0 ;
  assign n3698 = n460 & n2672 ;
  assign n3699 = n429 & n3698 ;
  assign n3700 = ~n2597 & n2801 ;
  assign n3701 = ~n2765 & n3700 ;
  assign n3702 = n3701 ^ n2892 ^ 1'b0 ;
  assign n3703 = n3699 | n3702 ;
  assign n3704 = n1843 ^ n1164 ^ 1'b0 ;
  assign n3707 = ( ~n891 & n1955 ) | ( ~n891 & n3044 ) | ( n1955 & n3044 ) ;
  assign n3708 = n3707 ^ n639 ^ 1'b0 ;
  assign n3709 = n2051 & ~n3708 ;
  assign n3705 = ~n310 & n3355 ;
  assign n3706 = ( n1935 & n3134 ) | ( n1935 & n3705 ) | ( n3134 & n3705 ) ;
  assign n3710 = n3709 ^ n3706 ^ n1946 ;
  assign n3711 = n441 & n1382 ;
  assign n3712 = n3677 & n3711 ;
  assign n3713 = n3054 & ~n3712 ;
  assign n3714 = n323 & ~n3000 ;
  assign n3715 = ~n602 & n3714 ;
  assign n3716 = n3715 ^ n577 ^ n489 ;
  assign n3717 = n2098 ^ n1723 ^ n556 ;
  assign n3718 = ( n885 & n1814 ) | ( n885 & ~n3717 ) | ( n1814 & ~n3717 ) ;
  assign n3719 = n801 & ~n3718 ;
  assign n3720 = n3716 & n3719 ;
  assign n3721 = n3720 ^ n1423 ^ n1365 ;
  assign n3722 = ( x18 & ~n3713 ) | ( x18 & n3721 ) | ( ~n3713 & n3721 ) ;
  assign n3723 = n3262 ^ n3160 ^ n613 ;
  assign n3724 = n3439 & ~n3723 ;
  assign n3725 = ~n3201 & n3724 ;
  assign n3726 = n2998 ^ n2149 ^ n1623 ;
  assign n3727 = x177 & ~n1901 ;
  assign n3728 = n3727 ^ n2963 ^ 1'b0 ;
  assign n3729 = n2943 & ~n3728 ;
  assign n3730 = ( n1300 & ~n3726 ) | ( n1300 & n3729 ) | ( ~n3726 & n3729 ) ;
  assign n3734 = ~n594 & n1846 ;
  assign n3735 = ~n786 & n3734 ;
  assign n3736 = n3735 ^ n1783 ^ 1'b0 ;
  assign n3731 = ( n588 & n831 ) | ( n588 & ~n2591 ) | ( n831 & ~n2591 ) ;
  assign n3732 = n3731 ^ n1454 ^ n689 ;
  assign n3733 = n3732 ^ n1043 ^ 1'b0 ;
  assign n3737 = n3736 ^ n3733 ^ x212 ;
  assign n3738 = ( n1229 & n1442 ) | ( n1229 & n2278 ) | ( n1442 & n2278 ) ;
  assign n3739 = ( n325 & n799 ) | ( n325 & ~n2396 ) | ( n799 & ~n2396 ) ;
  assign n3740 = n3739 ^ n1961 ^ n1599 ;
  assign n3741 = ( x174 & n1675 ) | ( x174 & ~n3740 ) | ( n1675 & ~n3740 ) ;
  assign n3742 = n3738 | n3741 ;
  assign n3743 = n3742 ^ n1450 ^ 1'b0 ;
  assign n3744 = ~n2529 & n3743 ;
  assign n3745 = x62 & n1638 ;
  assign n3746 = n1429 & n3745 ;
  assign n3747 = ( n481 & n561 ) | ( n481 & n1010 ) | ( n561 & n1010 ) ;
  assign n3748 = n3747 ^ n3080 ^ 1'b0 ;
  assign n3749 = n3346 ^ n859 ^ 1'b0 ;
  assign n3752 = ~n1306 & n1985 ;
  assign n3753 = n1465 & n3752 ;
  assign n3750 = ~x193 & n1717 ;
  assign n3751 = n3750 ^ n2976 ^ n433 ;
  assign n3754 = n3753 ^ n3751 ^ n2623 ;
  assign n3755 = n3754 ^ n3008 ^ x249 ;
  assign n3756 = n3749 & ~n3755 ;
  assign n3764 = n3752 ^ n658 ^ n617 ;
  assign n3762 = n1337 & n2448 ;
  assign n3757 = n271 & ~n1163 ;
  assign n3758 = n3757 ^ n353 ^ 1'b0 ;
  assign n3759 = ~n2853 & n3234 ;
  assign n3760 = ( n1796 & n3758 ) | ( n1796 & ~n3759 ) | ( n3758 & ~n3759 ) ;
  assign n3761 = n3760 ^ n1510 ^ 1'b0 ;
  assign n3763 = n3762 ^ n3761 ^ n683 ;
  assign n3765 = n3764 ^ n3763 ^ n287 ;
  assign n3766 = n1608 & ~n3174 ;
  assign n3767 = n3765 & n3766 ;
  assign n3769 = ~n509 & n2517 ;
  assign n3770 = n3769 ^ n374 ^ 1'b0 ;
  assign n3771 = ( ~x125 & n266 ) | ( ~x125 & n3770 ) | ( n266 & n3770 ) ;
  assign n3768 = n895 & ~n2167 ;
  assign n3772 = n3771 ^ n3768 ^ 1'b0 ;
  assign n3773 = n3772 ^ n913 ^ 1'b0 ;
  assign n3774 = ( ~n387 & n3767 ) | ( ~n387 & n3773 ) | ( n3767 & n3773 ) ;
  assign n3775 = n1834 | n1839 ;
  assign n3776 = n3775 ^ n1258 ^ 1'b0 ;
  assign n3777 = n3776 ^ n2798 ^ x177 ;
  assign n3778 = ~n1005 & n1347 ;
  assign n3779 = ~x28 & n3778 ;
  assign n3780 = n3777 & ~n3779 ;
  assign n3781 = n2756 ^ n874 ^ x5 ;
  assign n3782 = ~n740 & n1512 ;
  assign n3783 = n3782 ^ n566 ^ 1'b0 ;
  assign n3784 = ( n1950 & n2867 ) | ( n1950 & n3783 ) | ( n2867 & n3783 ) ;
  assign n3785 = n3784 ^ n3103 ^ n2885 ;
  assign n3786 = n3489 ^ n681 ^ 1'b0 ;
  assign n3787 = ~x98 & n1473 ;
  assign n3788 = n1200 & n1254 ;
  assign n3789 = ~n1137 & n3788 ;
  assign n3790 = ( n521 & n1566 ) | ( n521 & n2706 ) | ( n1566 & n2706 ) ;
  assign n3791 = ~n3789 & n3790 ;
  assign n3792 = n3787 | n3791 ;
  assign n3793 = n3792 ^ n2187 ^ n1962 ;
  assign n3794 = ~x21 & n1232 ;
  assign n3795 = x219 & ~n3794 ;
  assign n3796 = n3795 ^ n1210 ^ 1'b0 ;
  assign n3797 = n2224 ^ x112 ^ 1'b0 ;
  assign n3798 = n410 & ~n3797 ;
  assign n3799 = n3798 ^ n3435 ^ 1'b0 ;
  assign n3800 = n498 & n3799 ;
  assign n3801 = n2460 & n3800 ;
  assign n3802 = n3796 & ~n3801 ;
  assign n3803 = ~n1876 & n3802 ;
  assign n3804 = n1122 ^ n998 ^ n586 ;
  assign n3805 = n2191 ^ n1408 ^ 1'b0 ;
  assign n3806 = n3146 & n3805 ;
  assign n3807 = x109 & ~n3806 ;
  assign n3808 = ( n386 & ~n3804 ) | ( n386 & n3807 ) | ( ~n3804 & n3807 ) ;
  assign n3809 = n1062 | n3808 ;
  assign n3810 = ( x156 & n437 ) | ( x156 & n598 ) | ( n437 & n598 ) ;
  assign n3811 = n3810 ^ n2777 ^ n2433 ;
  assign n3812 = n511 ^ x208 ^ 1'b0 ;
  assign n3813 = ~n3811 & n3812 ;
  assign n3814 = ( n1177 & n2667 ) | ( n1177 & n3813 ) | ( n2667 & n3813 ) ;
  assign n3815 = ( n758 & ~n1107 ) | ( n758 & n1620 ) | ( ~n1107 & n1620 ) ;
  assign n3816 = ~n3285 & n3815 ;
  assign n3817 = ~n667 & n3816 ;
  assign n3818 = n3817 ^ n1787 ^ x17 ;
  assign n3819 = n1042 & n3818 ;
  assign n3820 = ( n892 & n1258 ) | ( n892 & n2562 ) | ( n1258 & n2562 ) ;
  assign n3823 = ( n458 & ~n1036 ) | ( n458 & n2677 ) | ( ~n1036 & n2677 ) ;
  assign n3821 = n1279 | n2312 ;
  assign n3822 = ~n1485 & n3821 ;
  assign n3824 = n3823 ^ n3822 ^ 1'b0 ;
  assign n3825 = n613 ^ x158 ^ 1'b0 ;
  assign n3826 = ( n1881 & ~n2755 ) | ( n1881 & n3825 ) | ( ~n2755 & n3825 ) ;
  assign n3827 = ( n1372 & n3709 ) | ( n1372 & n3826 ) | ( n3709 & n3826 ) ;
  assign n3832 = ( n585 & ~n1849 ) | ( n585 & n3706 ) | ( ~n1849 & n3706 ) ;
  assign n3829 = n2391 ^ x37 ^ 1'b0 ;
  assign n3830 = n2470 | n3829 ;
  assign n3831 = n1067 & ~n3830 ;
  assign n3828 = n753 & n3011 ;
  assign n3833 = n3832 ^ n3831 ^ n3828 ;
  assign n3836 = ~n1445 & n1516 ;
  assign n3837 = n3836 ^ n761 ^ 1'b0 ;
  assign n3834 = ( x187 & x242 ) | ( x187 & n329 ) | ( x242 & n329 ) ;
  assign n3835 = ~n1807 & n3834 ;
  assign n3838 = n3837 ^ n3835 ^ x145 ;
  assign n3839 = ( n1015 & n3605 ) | ( n1015 & ~n3838 ) | ( n3605 & ~n3838 ) ;
  assign n3840 = n1697 | n3453 ;
  assign n3841 = ( n1697 & n3494 ) | ( n1697 & n3840 ) | ( n3494 & n3840 ) ;
  assign n3842 = n704 | n3841 ;
  assign n3843 = n3839 | n3842 ;
  assign n3844 = n2952 ^ n1440 ^ 1'b0 ;
  assign n3845 = ( x83 & n439 ) | ( x83 & ~n2319 ) | ( n439 & ~n2319 ) ;
  assign n3846 = n859 & ~n3845 ;
  assign n3847 = ( n626 & n1497 ) | ( n626 & n3163 ) | ( n1497 & n3163 ) ;
  assign n3848 = ( x59 & n781 ) | ( x59 & n1186 ) | ( n781 & n1186 ) ;
  assign n3849 = ( x132 & n448 ) | ( x132 & ~n1084 ) | ( n448 & ~n1084 ) ;
  assign n3850 = n1221 | n1253 ;
  assign n3851 = n3849 & ~n3850 ;
  assign n3852 = n3851 ^ n2700 ^ 1'b0 ;
  assign n3853 = n3848 & ~n3852 ;
  assign n3854 = ( n829 & n3847 ) | ( n829 & n3853 ) | ( n3847 & n3853 ) ;
  assign n3855 = n1508 & ~n1820 ;
  assign n3856 = ~n2711 & n3855 ;
  assign n3857 = n3856 ^ n1152 ^ 1'b0 ;
  assign n3858 = n2233 ^ n1961 ^ n741 ;
  assign n3865 = n1463 ^ x185 ^ 1'b0 ;
  assign n3866 = n708 & n3865 ;
  assign n3867 = n3866 ^ n831 ^ 1'b0 ;
  assign n3868 = n1683 ^ x100 ^ 1'b0 ;
  assign n3869 = n1163 | n3868 ;
  assign n3870 = ( n2538 & n3867 ) | ( n2538 & ~n3869 ) | ( n3867 & ~n3869 ) ;
  assign n3862 = n345 & ~n384 ;
  assign n3863 = n3862 ^ n401 ^ 1'b0 ;
  assign n3861 = n1870 ^ n1077 ^ 1'b0 ;
  assign n3864 = n3863 ^ n3861 ^ n1347 ;
  assign n3859 = ~n502 & n2936 ;
  assign n3860 = ~n3157 & n3859 ;
  assign n3871 = n3870 ^ n3864 ^ n3860 ;
  assign n3872 = n283 | n3177 ;
  assign n3873 = n2746 | n3872 ;
  assign n3874 = n2183 ^ n2066 ^ x243 ;
  assign n3875 = ( ~x205 & n1830 ) | ( ~x205 & n2162 ) | ( n1830 & n2162 ) ;
  assign n3876 = n3259 & n3875 ;
  assign n3877 = n3876 ^ n1216 ^ 1'b0 ;
  assign n3880 = ( x89 & n453 ) | ( x89 & ~n3113 ) | ( n453 & ~n3113 ) ;
  assign n3878 = ( ~n290 & n924 ) | ( ~n290 & n2057 ) | ( n924 & n2057 ) ;
  assign n3879 = ( n1606 & n1665 ) | ( n1606 & ~n3878 ) | ( n1665 & ~n3878 ) ;
  assign n3881 = n3880 ^ n3879 ^ 1'b0 ;
  assign n3888 = n1412 ^ n618 ^ 1'b0 ;
  assign n3889 = n363 & n3888 ;
  assign n3890 = n738 & n3889 ;
  assign n3891 = ~x159 & n3890 ;
  assign n3892 = ( n1067 & n1474 ) | ( n1067 & ~n3891 ) | ( n1474 & ~n3891 ) ;
  assign n3893 = n3655 ^ n465 ^ 1'b0 ;
  assign n3894 = ~n3892 & n3893 ;
  assign n3884 = n1394 ^ x190 ^ 1'b0 ;
  assign n3885 = n3884 ^ n3264 ^ n1872 ;
  assign n3886 = ( ~n1588 & n1905 ) | ( ~n1588 & n3885 ) | ( n1905 & n3885 ) ;
  assign n3882 = n2589 ^ n1186 ^ 1'b0 ;
  assign n3883 = n838 & ~n3882 ;
  assign n3887 = n3886 ^ n3883 ^ n1291 ;
  assign n3895 = n3894 ^ n3887 ^ n2520 ;
  assign n3896 = n1101 | n1440 ;
  assign n3897 = n932 & ~n3752 ;
  assign n3898 = n3897 ^ n2057 ^ n1023 ;
  assign n3899 = n2196 ^ x60 ^ 1'b0 ;
  assign n3900 = ( n1065 & ~n1284 ) | ( n1065 & n3899 ) | ( ~n1284 & n3899 ) ;
  assign n3901 = n1910 & n3900 ;
  assign n3902 = n3898 & n3901 ;
  assign n3903 = n3902 ^ n2625 ^ 1'b0 ;
  assign n3904 = n3896 & ~n3903 ;
  assign n3905 = n3904 ^ n2945 ^ 1'b0 ;
  assign n3906 = n2744 ^ n788 ^ x30 ;
  assign n3907 = n1311 ^ n672 ^ 1'b0 ;
  assign n3908 = n2229 | n3907 ;
  assign n3909 = n3908 ^ n2794 ^ n1295 ;
  assign n3910 = ( n901 & n1163 ) | ( n901 & n1227 ) | ( n1163 & n1227 ) ;
  assign n3911 = n3910 ^ n1411 ^ 1'b0 ;
  assign n3912 = ( n1391 & ~n1468 ) | ( n1391 & n3516 ) | ( ~n1468 & n3516 ) ;
  assign n3913 = n346 & ~n2308 ;
  assign n3914 = n3913 ^ x123 ^ 1'b0 ;
  assign n3917 = n1291 ^ n947 ^ x70 ;
  assign n3915 = x136 & n770 ;
  assign n3916 = n3915 ^ x246 ^ 1'b0 ;
  assign n3918 = n3917 ^ n3916 ^ n1075 ;
  assign n3919 = ( n3486 & ~n3914 ) | ( n3486 & n3918 ) | ( ~n3914 & n3918 ) ;
  assign n3920 = ( n1344 & n1385 ) | ( n1344 & ~n3919 ) | ( n1385 & ~n3919 ) ;
  assign n3922 = n1129 ^ n325 ^ x237 ;
  assign n3923 = ( n384 & n3446 ) | ( n384 & ~n3922 ) | ( n3446 & ~n3922 ) ;
  assign n3921 = ( x131 & x227 ) | ( x131 & ~n1684 ) | ( x227 & ~n1684 ) ;
  assign n3924 = n3923 ^ n3921 ^ n1820 ;
  assign n3925 = ( x57 & ~n395 ) | ( x57 & n1135 ) | ( ~n395 & n1135 ) ;
  assign n3926 = n3925 ^ n436 ^ 1'b0 ;
  assign n3927 = n2958 & ~n3926 ;
  assign n3928 = n3671 & n3927 ;
  assign n3929 = n3928 ^ x168 ^ 1'b0 ;
  assign n3930 = n3740 | n3929 ;
  assign n3931 = n3930 ^ n1997 ^ 1'b0 ;
  assign n3932 = ~x88 & n1914 ;
  assign n3933 = n1839 & n3932 ;
  assign n3934 = ( n622 & n2092 ) | ( n622 & n3933 ) | ( n2092 & n3933 ) ;
  assign n3935 = n2915 ^ x27 ^ 1'b0 ;
  assign n3936 = x147 & n1710 ;
  assign n3937 = n2034 & n3936 ;
  assign n3939 = n1002 & ~n2482 ;
  assign n3940 = n3939 ^ x72 ^ 1'b0 ;
  assign n3938 = n3115 ^ n2981 ^ 1'b0 ;
  assign n3941 = n3940 ^ n3938 ^ n2859 ;
  assign n3942 = n2157 ^ n2029 ^ 1'b0 ;
  assign n3943 = ( n1049 & n2409 ) | ( n1049 & ~n3942 ) | ( n2409 & ~n3942 ) ;
  assign n3955 = x89 | n539 ;
  assign n3954 = n2613 ^ n1773 ^ 1'b0 ;
  assign n3956 = n3955 ^ n3954 ^ n2956 ;
  assign n3944 = n622 & n2433 ;
  assign n3945 = n3944 ^ n674 ^ 1'b0 ;
  assign n3946 = n3945 ^ n1447 ^ 1'b0 ;
  assign n3947 = n1010 ^ n538 ^ x31 ;
  assign n3948 = n1709 | n3947 ;
  assign n3949 = n2206 ^ n1274 ^ 1'b0 ;
  assign n3950 = n3949 ^ n3749 ^ n1827 ;
  assign n3951 = ( n2910 & n3948 ) | ( n2910 & n3950 ) | ( n3948 & n3950 ) ;
  assign n3952 = n3951 ^ n2049 ^ n872 ;
  assign n3953 = ( ~n1928 & n3946 ) | ( ~n1928 & n3952 ) | ( n3946 & n3952 ) ;
  assign n3957 = n3956 ^ n3953 ^ 1'b0 ;
  assign n3958 = n3140 | n3957 ;
  assign n3959 = ( n733 & n1220 ) | ( n733 & ~n1301 ) | ( n1220 & ~n1301 ) ;
  assign n3960 = n3959 ^ n385 ^ 1'b0 ;
  assign n3961 = ~n1434 & n3960 ;
  assign n3962 = n1138 & n2495 ;
  assign n3963 = x149 ^ x8 ^ 1'b0 ;
  assign n3964 = ~n2906 & n3946 ;
  assign n3965 = ~n3963 & n3964 ;
  assign n3966 = n2357 | n3712 ;
  assign n3967 = n2145 | n3966 ;
  assign n3968 = x6 | n2563 ;
  assign n3969 = ( n1815 & ~n1864 ) | ( n1815 & n3968 ) | ( ~n1864 & n3968 ) ;
  assign n3970 = n2517 ^ n1233 ^ n704 ;
  assign n3971 = ( ~n261 & n464 ) | ( ~n261 & n824 ) | ( n464 & n824 ) ;
  assign n3972 = ( n298 & n401 ) | ( n298 & ~n3971 ) | ( n401 & ~n3971 ) ;
  assign n3973 = n3972 ^ n559 ^ 1'b0 ;
  assign n3974 = n995 & n3973 ;
  assign n3975 = n3974 ^ x236 ^ 1'b0 ;
  assign n3976 = ~n3970 & n3975 ;
  assign n3977 = ~n1671 & n2820 ;
  assign n3978 = x21 & ~n3977 ;
  assign n3979 = n1667 & ~n3479 ;
  assign n3980 = n3979 ^ n3146 ^ 1'b0 ;
  assign n3981 = n3978 & ~n3980 ;
  assign n3982 = n1288 ^ n1014 ^ n474 ;
  assign n3983 = ( ~n938 & n3981 ) | ( ~n938 & n3982 ) | ( n3981 & n3982 ) ;
  assign n3984 = n3983 ^ n1176 ^ 1'b0 ;
  assign n3985 = n3984 ^ n3465 ^ n1430 ;
  assign n3986 = n3753 ^ n1982 ^ 1'b0 ;
  assign n3987 = ~x177 & n3986 ;
  assign n3988 = ( n2932 & n3696 ) | ( n2932 & ~n3987 ) | ( n3696 & ~n3987 ) ;
  assign n3989 = n3988 ^ n3801 ^ n1504 ;
  assign n3991 = x123 & ~n509 ;
  assign n3990 = ~n654 & n682 ;
  assign n3992 = n3991 ^ n3990 ^ 1'b0 ;
  assign n3993 = ( n1385 & n1587 ) | ( n1385 & n3992 ) | ( n1587 & n3992 ) ;
  assign n3994 = n3993 ^ n378 ^ 1'b0 ;
  assign n3995 = ~n1692 & n3994 ;
  assign n3996 = n3995 ^ n689 ^ 1'b0 ;
  assign n4000 = ( n513 & ~n1935 ) | ( n513 & n3230 ) | ( ~n1935 & n3230 ) ;
  assign n4001 = n4000 ^ n1466 ^ n668 ;
  assign n4002 = n928 & ~n4001 ;
  assign n4003 = n4002 ^ x144 ^ 1'b0 ;
  assign n4004 = n4003 ^ n1376 ^ n1343 ;
  assign n4005 = ( ~n2108 & n3626 ) | ( ~n2108 & n4004 ) | ( n3626 & n4004 ) ;
  assign n3997 = n362 ^ x189 ^ 1'b0 ;
  assign n3998 = n3997 ^ n1545 ^ 1'b0 ;
  assign n3999 = n429 | n3998 ;
  assign n4006 = n4005 ^ n3999 ^ n3580 ;
  assign n4007 = ( ~n554 & n1261 ) | ( ~n554 & n2141 ) | ( n1261 & n2141 ) ;
  assign n4008 = n4007 ^ x155 ^ 1'b0 ;
  assign n4009 = n3704 & ~n4008 ;
  assign n4010 = n1894 ^ n1725 ^ n374 ;
  assign n4011 = ~n1862 & n4010 ;
  assign n4018 = ( n1317 & ~n1937 ) | ( n1317 & n3422 ) | ( ~n1937 & n3422 ) ;
  assign n4019 = n1197 & n4018 ;
  assign n4020 = n4019 ^ n1032 ^ 1'b0 ;
  assign n4013 = n1422 ^ n771 ^ 1'b0 ;
  assign n4014 = x180 & n4013 ;
  assign n4015 = n4014 ^ n1206 ^ n609 ;
  assign n4016 = n1611 ^ x27 ^ 1'b0 ;
  assign n4017 = ~n4015 & n4016 ;
  assign n4012 = n1850 ^ n711 ^ x89 ;
  assign n4021 = n4020 ^ n4017 ^ n4012 ;
  assign n4022 = ( n1072 & n2065 ) | ( n1072 & ~n2523 ) | ( n2065 & ~n2523 ) ;
  assign n4023 = ( n401 & ~n1073 ) | ( n401 & n4022 ) | ( ~n1073 & n4022 ) ;
  assign n4024 = x172 & ~n2777 ;
  assign n4025 = n4024 ^ n2464 ^ 1'b0 ;
  assign n4026 = x199 & n1310 ;
  assign n4027 = n4026 ^ n2330 ^ 1'b0 ;
  assign n4028 = ( x125 & n300 ) | ( x125 & n4027 ) | ( n300 & n4027 ) ;
  assign n4029 = n2844 & ~n3364 ;
  assign n4030 = ~n4028 & n4029 ;
  assign n4031 = n4004 ^ n1275 ^ 1'b0 ;
  assign n4032 = n2094 & ~n4031 ;
  assign n4042 = n1430 ^ n704 ^ 1'b0 ;
  assign n4037 = n1137 ^ n1069 ^ 1'b0 ;
  assign n4038 = ~n1294 & n4037 ;
  assign n4039 = x51 & n474 ;
  assign n4040 = n4039 ^ n1229 ^ 1'b0 ;
  assign n4041 = ( ~n1308 & n4038 ) | ( ~n1308 & n4040 ) | ( n4038 & n4040 ) ;
  assign n4043 = n4042 ^ n4041 ^ 1'b0 ;
  assign n4033 = ( n1012 & n1440 ) | ( n1012 & n2359 ) | ( n1440 & n2359 ) ;
  assign n4034 = ~n432 & n1236 ;
  assign n4035 = ( n2798 & n3765 ) | ( n2798 & ~n4034 ) | ( n3765 & ~n4034 ) ;
  assign n4036 = n4033 & ~n4035 ;
  assign n4044 = n4043 ^ n4036 ^ 1'b0 ;
  assign n4045 = n3655 ^ n2061 ^ 1'b0 ;
  assign n4046 = n1827 ^ n801 ^ n461 ;
  assign n4047 = n4046 ^ n1317 ^ n614 ;
  assign n4048 = n4047 ^ n1838 ^ 1'b0 ;
  assign n4049 = n1962 | n4048 ;
  assign n4050 = n3970 ^ n687 ^ 1'b0 ;
  assign n4051 = n895 & n4050 ;
  assign n4052 = n4051 ^ n2102 ^ 1'b0 ;
  assign n4053 = ( ~n840 & n946 ) | ( ~n840 & n2072 ) | ( n946 & n2072 ) ;
  assign n4054 = n561 & n4053 ;
  assign n4055 = ( n660 & ~n991 ) | ( n660 & n1484 ) | ( ~n991 & n1484 ) ;
  assign n4056 = ( n2596 & n4054 ) | ( n2596 & n4055 ) | ( n4054 & n4055 ) ;
  assign n4057 = ( n716 & n2495 ) | ( n716 & n4017 ) | ( n2495 & n4017 ) ;
  assign n4059 = ~n349 & n2714 ;
  assign n4060 = n4059 ^ n607 ^ 1'b0 ;
  assign n4058 = ( n741 & n1361 ) | ( n741 & n2979 ) | ( n1361 & n2979 ) ;
  assign n4061 = n4060 ^ n4058 ^ 1'b0 ;
  assign n4062 = n1991 ^ n640 ^ x90 ;
  assign n4063 = n4062 ^ n3568 ^ n2859 ;
  assign n4064 = ( ~n3437 & n4061 ) | ( ~n3437 & n4063 ) | ( n4061 & n4063 ) ;
  assign n4068 = ( x120 & n1139 ) | ( x120 & n1398 ) | ( n1139 & n1398 ) ;
  assign n4065 = n3834 ^ n3472 ^ 1'b0 ;
  assign n4066 = n2899 | n4065 ;
  assign n4067 = n4066 ^ n2835 ^ n752 ;
  assign n4069 = n4068 ^ n4067 ^ 1'b0 ;
  assign n4070 = n4064 & n4069 ;
  assign n4071 = ( n337 & ~n972 ) | ( n337 & n1458 ) | ( ~n972 & n1458 ) ;
  assign n4072 = n4071 ^ n2668 ^ 1'b0 ;
  assign n4073 = n1260 | n4072 ;
  assign n4074 = n4073 ^ n2392 ^ n1393 ;
  assign n4075 = ~n3124 & n4074 ;
  assign n4076 = ( n1448 & n4042 ) | ( n1448 & ~n4075 ) | ( n4042 & ~n4075 ) ;
  assign n4077 = ( n585 & ~n1994 ) | ( n585 & n4076 ) | ( ~n1994 & n4076 ) ;
  assign n4083 = n718 & ~n975 ;
  assign n4084 = ( n1690 & ~n3662 ) | ( n1690 & n4083 ) | ( ~n3662 & n4083 ) ;
  assign n4078 = n3301 ^ n797 ^ 1'b0 ;
  assign n4085 = n4084 ^ n4078 ^ n2426 ;
  assign n4079 = ( ~n679 & n1602 ) | ( ~n679 & n3208 ) | ( n1602 & n3208 ) ;
  assign n4080 = ( n599 & ~n3216 ) | ( n599 & n4079 ) | ( ~n3216 & n4079 ) ;
  assign n4081 = n1155 & n4080 ;
  assign n4082 = n4078 & n4081 ;
  assign n4086 = n4085 ^ n4082 ^ n3064 ;
  assign n4087 = n853 & ~n1821 ;
  assign n4088 = n1736 | n4087 ;
  assign n4089 = n4088 ^ n2348 ^ 1'b0 ;
  assign n4090 = ( n470 & n540 ) | ( n470 & n1894 ) | ( n540 & n1894 ) ;
  assign n4091 = n4090 ^ n670 ^ 1'b0 ;
  assign n4092 = ~n4089 & n4091 ;
  assign n4093 = ~n4086 & n4092 ;
  assign n4094 = n4028 ^ n3122 ^ 1'b0 ;
  assign n4100 = x171 & n1245 ;
  assign n4101 = n313 & n807 ;
  assign n4102 = n761 | n4101 ;
  assign n4103 = x220 | n4102 ;
  assign n4104 = ~n4100 & n4103 ;
  assign n4105 = x229 & ~n502 ;
  assign n4106 = ~n4104 & n4105 ;
  assign n4095 = n3146 ^ n1323 ^ n638 ;
  assign n4096 = n4095 ^ x171 ^ 1'b0 ;
  assign n4097 = ~n704 & n4096 ;
  assign n4098 = n4097 ^ n1793 ^ 1'b0 ;
  assign n4099 = n1995 & n4098 ;
  assign n4107 = n4106 ^ n4099 ^ n962 ;
  assign n4108 = n347 ^ x158 ^ 1'b0 ;
  assign n4109 = x202 & n4108 ;
  assign n4110 = n4109 ^ n2217 ^ 1'b0 ;
  assign n4111 = n1361 | n4110 ;
  assign n4112 = n2330 | n4111 ;
  assign n4113 = n2029 | n4112 ;
  assign n4114 = ~n458 & n4113 ;
  assign n4115 = n4114 ^ n529 ^ 1'b0 ;
  assign n4116 = x187 & ~n3148 ;
  assign n4117 = ~n3308 & n4116 ;
  assign n4118 = n1272 ^ x188 ^ 1'b0 ;
  assign n4119 = n497 & ~n3298 ;
  assign n4120 = n4119 ^ n3161 ^ n2344 ;
  assign n4121 = ( n983 & n4118 ) | ( n983 & n4120 ) | ( n4118 & n4120 ) ;
  assign n4122 = n2634 ^ n872 ^ n587 ;
  assign n4123 = ( ~n1192 & n1233 ) | ( ~n1192 & n4122 ) | ( n1233 & n4122 ) ;
  assign n4131 = n1398 ^ n613 ^ x198 ;
  assign n4130 = ( x186 & n1403 ) | ( x186 & ~n4066 ) | ( n1403 & ~n4066 ) ;
  assign n4124 = n2853 ^ n1245 ^ 1'b0 ;
  assign n4125 = n2558 ^ x89 ^ 1'b0 ;
  assign n4126 = n4124 | n4125 ;
  assign n4127 = x133 & n2883 ;
  assign n4128 = n4126 & n4127 ;
  assign n4129 = n4128 ^ n2644 ^ n2108 ;
  assign n4132 = n4131 ^ n4130 ^ n4129 ;
  assign n4133 = n969 ^ x237 ^ 1'b0 ;
  assign n4134 = x176 & ~n4133 ;
  assign n4135 = n2844 & ~n4010 ;
  assign n4136 = n4135 ^ n876 ^ 1'b0 ;
  assign n4137 = n2595 ^ x70 ^ 1'b0 ;
  assign n4138 = ( n1089 & n4136 ) | ( n1089 & n4137 ) | ( n4136 & n4137 ) ;
  assign n4139 = n797 & n4138 ;
  assign n4150 = x50 & n733 ;
  assign n4147 = n1050 & ~n1341 ;
  assign n4148 = n624 | n1143 ;
  assign n4149 = n4147 & ~n4148 ;
  assign n4140 = x202 & ~n598 ;
  assign n4141 = n945 & n4140 ;
  assign n4142 = n3849 ^ n1904 ^ n395 ;
  assign n4143 = n2021 ^ n704 ^ 1'b0 ;
  assign n4144 = n1303 & n4143 ;
  assign n4145 = ( n3309 & n4142 ) | ( n3309 & n4144 ) | ( n4142 & n4144 ) ;
  assign n4146 = ( n2317 & ~n4141 ) | ( n2317 & n4145 ) | ( ~n4141 & n4145 ) ;
  assign n4151 = n4150 ^ n4149 ^ n4146 ;
  assign n4155 = n912 & ~n1025 ;
  assign n4152 = n1688 ^ n903 ^ n899 ;
  assign n4153 = ( n686 & n3257 ) | ( n686 & n4152 ) | ( n3257 & n4152 ) ;
  assign n4154 = n2812 | n4153 ;
  assign n4156 = n4155 ^ n4154 ^ 1'b0 ;
  assign n4157 = n3106 ^ n601 ^ 1'b0 ;
  assign n4158 = ( x138 & n4156 ) | ( x138 & n4157 ) | ( n4156 & n4157 ) ;
  assign n4159 = n3471 & ~n4158 ;
  assign n4160 = n3577 & n4159 ;
  assign n4163 = n3129 ^ n523 ^ 1'b0 ;
  assign n4164 = ~n2597 & n4163 ;
  assign n4161 = ( n287 & n1261 ) | ( n287 & n1306 ) | ( n1261 & n1306 ) ;
  assign n4162 = n1268 & ~n4161 ;
  assign n4165 = n4164 ^ n4162 ^ 1'b0 ;
  assign n4166 = n4165 ^ n3801 ^ x9 ;
  assign n4167 = ~n3471 & n3813 ;
  assign n4168 = n697 ^ n267 ^ 1'b0 ;
  assign n4169 = ~n650 & n4168 ;
  assign n4170 = n4169 ^ x204 ^ 1'b0 ;
  assign n4171 = ~n2099 & n4170 ;
  assign n4172 = ~n1399 & n4171 ;
  assign n4173 = ~n1462 & n4172 ;
  assign n4174 = n4173 ^ n3276 ^ 1'b0 ;
  assign n4175 = n4167 & ~n4174 ;
  assign n4176 = ( x130 & n304 ) | ( x130 & n3013 ) | ( n304 & n3013 ) ;
  assign n4177 = x129 & ~n4176 ;
  assign n4178 = n4177 ^ n3262 ^ 1'b0 ;
  assign n4179 = ( ~n801 & n1162 ) | ( ~n801 & n1998 ) | ( n1162 & n1998 ) ;
  assign n4180 = ( n570 & n1123 ) | ( n570 & n2596 ) | ( n1123 & n2596 ) ;
  assign n4181 = ~n1884 & n4180 ;
  assign n4182 = ~x176 & n4181 ;
  assign n4183 = n4182 ^ n916 ^ 1'b0 ;
  assign n4184 = ~n4179 & n4183 ;
  assign n4185 = n4184 ^ n2733 ^ n1229 ;
  assign n4186 = n4185 ^ n1789 ^ 1'b0 ;
  assign n4187 = n4178 & n4186 ;
  assign n4188 = ~n1524 & n4187 ;
  assign n4189 = n4188 ^ n924 ^ 1'b0 ;
  assign n4193 = n1306 & ~n1561 ;
  assign n4194 = n4193 ^ n1784 ^ n1010 ;
  assign n4190 = x127 & n318 ;
  assign n4191 = ~n2106 & n4190 ;
  assign n4192 = ( n652 & ~n1010 ) | ( n652 & n4191 ) | ( ~n1010 & n4191 ) ;
  assign n4195 = n4194 ^ n4192 ^ x85 ;
  assign n4200 = ( x226 & n1706 ) | ( x226 & n2109 ) | ( n1706 & n2109 ) ;
  assign n4198 = ( ~x74 & x131 ) | ( ~x74 & n1099 ) | ( x131 & n1099 ) ;
  assign n4197 = n672 ^ n364 ^ x209 ;
  assign n4196 = n897 & ~n1998 ;
  assign n4199 = n4198 ^ n4197 ^ n4196 ;
  assign n4201 = n4200 ^ n4199 ^ n4052 ;
  assign n4202 = x30 & n2676 ;
  assign n4203 = n4202 ^ n1141 ^ 1'b0 ;
  assign n4204 = n4203 ^ n3200 ^ n1308 ;
  assign n4205 = n608 ^ x26 ^ 1'b0 ;
  assign n4206 = n4204 & n4205 ;
  assign n4207 = ~n514 & n1649 ;
  assign n4208 = ~n498 & n4207 ;
  assign n4209 = ( n1506 & n3426 ) | ( n1506 & ~n4208 ) | ( n3426 & ~n4208 ) ;
  assign n4210 = n4209 ^ n1039 ^ x222 ;
  assign n4218 = n633 & n1012 ;
  assign n4219 = ~x194 & n4218 ;
  assign n4217 = ( n306 & n807 ) | ( n306 & ~n2517 ) | ( n807 & ~n2517 ) ;
  assign n4220 = n4219 ^ n4217 ^ x215 ;
  assign n4215 = n910 & n3269 ;
  assign n4216 = n4215 ^ n1019 ^ 1'b0 ;
  assign n4221 = n4220 ^ n4216 ^ n715 ;
  assign n4222 = n3271 & n4221 ;
  assign n4211 = n2340 ^ n275 ^ 1'b0 ;
  assign n4212 = ~n1626 & n4211 ;
  assign n4213 = ~n2917 & n4212 ;
  assign n4214 = n4213 ^ n3392 ^ n2344 ;
  assign n4223 = n4222 ^ n4214 ^ n3178 ;
  assign n4224 = n2983 & ~n3877 ;
  assign n4225 = ( n1089 & ~n1420 ) | ( n1089 & n3256 ) | ( ~n1420 & n3256 ) ;
  assign n4226 = ( n674 & n4106 ) | ( n674 & ~n4225 ) | ( n4106 & ~n4225 ) ;
  assign n4227 = n3981 ^ n2951 ^ n1848 ;
  assign n4228 = n2594 ^ n2229 ^ 1'b0 ;
  assign n4229 = n2436 ^ n1226 ^ n687 ;
  assign n4230 = n541 & n4229 ;
  assign n4231 = n4230 ^ n3160 ^ 1'b0 ;
  assign n4232 = n1720 ^ x54 ^ 1'b0 ;
  assign n4233 = ~n557 & n2286 ;
  assign n4234 = n4233 ^ n4124 ^ 1'b0 ;
  assign n4235 = ~n1977 & n4234 ;
  assign n4236 = n4235 ^ n2048 ^ 1'b0 ;
  assign n4237 = ( x134 & ~n1382 ) | ( x134 & n2165 ) | ( ~n1382 & n2165 ) ;
  assign n4238 = n3016 | n4237 ;
  assign n4239 = n4236 | n4238 ;
  assign n4240 = n2597 ^ n2063 ^ n1728 ;
  assign n4241 = n4240 ^ n775 ^ x68 ;
  assign n4242 = ~n370 & n4241 ;
  assign n4243 = n4242 ^ n1897 ^ 1'b0 ;
  assign n4244 = ( n4106 & ~n4239 ) | ( n4106 & n4243 ) | ( ~n4239 & n4243 ) ;
  assign n4245 = n356 & n3176 ;
  assign n4246 = x242 & n2850 ;
  assign n4247 = n4246 ^ n3720 ^ 1'b0 ;
  assign n4248 = ( n623 & n4245 ) | ( n623 & ~n4247 ) | ( n4245 & ~n4247 ) ;
  assign n4249 = n436 ^ x215 ^ 1'b0 ;
  assign n4250 = n3128 ^ n453 ^ 1'b0 ;
  assign n4251 = n4249 & n4250 ;
  assign n4252 = x206 & n671 ;
  assign n4253 = n4252 ^ n3664 ^ 1'b0 ;
  assign n4254 = ( n1291 & n4043 ) | ( n1291 & n4253 ) | ( n4043 & n4253 ) ;
  assign n4255 = ~n748 & n1834 ;
  assign n4256 = n436 | n3497 ;
  assign n4257 = ( n3892 & ~n4255 ) | ( n3892 & n4256 ) | ( ~n4255 & n4256 ) ;
  assign n4258 = n1640 & n3179 ;
  assign n4259 = n1185 & n4258 ;
  assign n4260 = n2162 & ~n4259 ;
  assign n4261 = ~n4257 & n4260 ;
  assign n4262 = ~n2845 & n4261 ;
  assign n4263 = n258 & n1598 ;
  assign n4264 = x79 & ~n1253 ;
  assign n4265 = n4264 ^ x96 ^ 1'b0 ;
  assign n4266 = ( n268 & n1636 ) | ( n268 & ~n4265 ) | ( n1636 & ~n4265 ) ;
  assign n4267 = n4266 ^ n2344 ^ 1'b0 ;
  assign n4268 = n565 | n4267 ;
  assign n4270 = n1079 ^ x254 ^ 1'b0 ;
  assign n4271 = n475 & n4270 ;
  assign n4269 = n868 & ~n1926 ;
  assign n4272 = n4271 ^ n4269 ^ 1'b0 ;
  assign n4273 = x124 & ~n4272 ;
  assign n4274 = ~n2384 & n4273 ;
  assign n4275 = n4274 ^ n3110 ^ n2279 ;
  assign n4276 = n935 & ~n1783 ;
  assign n4277 = ~x137 & n4276 ;
  assign n4278 = n4277 ^ n2707 ^ 1'b0 ;
  assign n4279 = n4256 & ~n4278 ;
  assign n4280 = ( n588 & n2329 ) | ( n588 & n4279 ) | ( n2329 & n4279 ) ;
  assign n4282 = n3218 ^ n971 ^ x121 ;
  assign n4281 = n1460 | n1904 ;
  assign n4283 = n4282 ^ n4281 ^ n308 ;
  assign n4284 = ( n556 & n1146 ) | ( n556 & ~n2810 ) | ( n1146 & ~n2810 ) ;
  assign n4285 = n4284 ^ n916 ^ 1'b0 ;
  assign n4286 = n3545 ^ n1680 ^ 1'b0 ;
  assign n4287 = ~n3744 & n4286 ;
  assign n4288 = n4287 ^ x215 ^ 1'b0 ;
  assign n4289 = n4288 ^ n885 ^ 1'b0 ;
  assign n4290 = n2698 & n4289 ;
  assign n4291 = ( n466 & n585 ) | ( n466 & ~n891 ) | ( n585 & ~n891 ) ;
  assign n4292 = n1465 & n3317 ;
  assign n4293 = ~n1836 & n4292 ;
  assign n4294 = ~n586 & n4293 ;
  assign n4295 = ( n1228 & ~n2367 ) | ( n1228 & n4294 ) | ( ~n2367 & n4294 ) ;
  assign n4296 = ~n3770 & n4295 ;
  assign n4297 = ~n623 & n4296 ;
  assign n4298 = ~n2259 & n2958 ;
  assign n4299 = ~n4297 & n4298 ;
  assign n4300 = n4299 ^ n3992 ^ 1'b0 ;
  assign n4301 = ~n1578 & n4300 ;
  assign n4302 = ( ~n3443 & n4291 ) | ( ~n3443 & n4301 ) | ( n4291 & n4301 ) ;
  assign n4303 = n1829 ^ n623 ^ 1'b0 ;
  assign n4304 = n3686 & n4303 ;
  assign n4305 = n4304 ^ n1048 ^ 1'b0 ;
  assign n4306 = n257 ^ x131 ^ 1'b0 ;
  assign n4307 = n705 & ~n4306 ;
  assign n4308 = n1649 & n4307 ;
  assign n4309 = n4308 ^ n3103 ^ 1'b0 ;
  assign n4310 = n992 ^ n874 ^ n873 ;
  assign n4311 = n4310 ^ n2114 ^ x110 ;
  assign n4312 = n1714 ^ n853 ^ 1'b0 ;
  assign n4313 = n347 & ~n4312 ;
  assign n4314 = n1229 & n2448 ;
  assign n4315 = ~n1069 & n4314 ;
  assign n4316 = n1251 ^ n445 ^ n289 ;
  assign n4317 = ( ~n3497 & n3968 ) | ( ~n3497 & n4316 ) | ( n3968 & n4316 ) ;
  assign n4318 = n973 | n2346 ;
  assign n4319 = n4318 ^ n2627 ^ 1'b0 ;
  assign n4320 = ( n4315 & n4317 ) | ( n4315 & ~n4319 ) | ( n4317 & ~n4319 ) ;
  assign n4321 = n4313 | n4320 ;
  assign n4322 = n4321 ^ n1182 ^ 1'b0 ;
  assign n4324 = n2750 ^ n1760 ^ n1516 ;
  assign n4325 = n4324 ^ n1745 ^ 1'b0 ;
  assign n4326 = n1419 ^ n325 ^ x151 ;
  assign n4327 = n4326 ^ n2574 ^ 1'b0 ;
  assign n4328 = ( n3248 & ~n4325 ) | ( n3248 & n4327 ) | ( ~n4325 & n4327 ) ;
  assign n4323 = ~n2460 & n2615 ;
  assign n4329 = n4328 ^ n4323 ^ 1'b0 ;
  assign n4330 = n3512 & n3575 ;
  assign n4331 = ~n1267 & n4330 ;
  assign n4332 = n439 & ~n1331 ;
  assign n4333 = n4042 ^ n3593 ^ 1'b0 ;
  assign n4334 = n4333 ^ n1783 ^ n829 ;
  assign n4335 = n4334 ^ n974 ^ 1'b0 ;
  assign n4336 = n343 & n4335 ;
  assign n4337 = n4336 ^ n2644 ^ 1'b0 ;
  assign n4338 = ( n380 & n4332 ) | ( n380 & n4337 ) | ( n4332 & n4337 ) ;
  assign n4339 = n4189 ^ n2185 ^ n1532 ;
  assign n4342 = n3731 ^ n347 ^ 1'b0 ;
  assign n4340 = n3997 ^ n561 ^ n350 ;
  assign n4341 = n2233 & ~n4340 ;
  assign n4343 = n4342 ^ n4341 ^ 1'b0 ;
  assign n4344 = n2096 ^ n1703 ^ 1'b0 ;
  assign n4345 = ( n2778 & n3502 ) | ( n2778 & n4344 ) | ( n3502 & n4344 ) ;
  assign n4346 = n1504 ^ n666 ^ 1'b0 ;
  assign n4349 = n2246 ^ n822 ^ 1'b0 ;
  assign n4347 = n3199 ^ n773 ^ 1'b0 ;
  assign n4348 = n3919 & n4347 ;
  assign n4350 = n4349 ^ n4348 ^ n3707 ;
  assign n4351 = n2254 ^ n273 ^ 1'b0 ;
  assign n4352 = n818 & n3147 ;
  assign n4353 = n4351 & n4352 ;
  assign n4354 = n1473 ^ n1368 ^ 1'b0 ;
  assign n4355 = n1363 & ~n3651 ;
  assign n4356 = ~n4354 & n4355 ;
  assign n4357 = n4067 ^ n2400 ^ n2322 ;
  assign n4362 = n3000 ^ n1225 ^ n317 ;
  assign n4359 = n1444 ^ n655 ^ 1'b0 ;
  assign n4360 = ( ~n1040 & n1994 ) | ( ~n1040 & n3050 ) | ( n1994 & n3050 ) ;
  assign n4361 = n4359 & n4360 ;
  assign n4363 = n4362 ^ n4361 ^ 1'b0 ;
  assign n4358 = n2707 ^ n1891 ^ n596 ;
  assign n4364 = n4363 ^ n4358 ^ 1'b0 ;
  assign n4365 = n287 & ~n4364 ;
  assign n4366 = n3860 ^ n701 ^ 1'b0 ;
  assign n4370 = x229 | n1849 ;
  assign n4367 = n693 ^ n504 ^ n492 ;
  assign n4368 = n4367 ^ n3899 ^ n322 ;
  assign n4369 = n3475 & n4368 ;
  assign n4371 = n4370 ^ n4369 ^ 1'b0 ;
  assign n4372 = n1842 ^ n1798 ^ 1'b0 ;
  assign n4373 = ~n4371 & n4372 ;
  assign n4374 = n1308 & ~n4373 ;
  assign n4375 = n1831 ^ n817 ^ x92 ;
  assign n4376 = ( ~x141 & n1189 ) | ( ~x141 & n1818 ) | ( n1189 & n1818 ) ;
  assign n4377 = n1305 | n4376 ;
  assign n4378 = n451 & ~n4377 ;
  assign n4379 = ( n2276 & n4375 ) | ( n2276 & ~n4378 ) | ( n4375 & ~n4378 ) ;
  assign n4380 = n2312 ^ n1516 ^ 1'b0 ;
  assign n4381 = x15 & ~n4380 ;
  assign n4382 = ( n4374 & ~n4379 ) | ( n4374 & n4381 ) | ( ~n4379 & n4381 ) ;
  assign n4383 = n2700 ^ x114 ^ 1'b0 ;
  assign n4384 = n1325 & ~n4383 ;
  assign n4385 = ( n1751 & ~n1984 ) | ( n1751 & n4384 ) | ( ~n1984 & n4384 ) ;
  assign n4386 = ( n487 & n587 ) | ( n487 & ~n4385 ) | ( n587 & ~n4385 ) ;
  assign n4387 = ( ~n841 & n2187 ) | ( ~n841 & n2878 ) | ( n2187 & n2878 ) ;
  assign n4388 = n3873 ^ n310 ^ 1'b0 ;
  assign n4389 = ~n4387 & n4388 ;
  assign n4390 = n2625 ^ n1845 ^ n447 ;
  assign n4391 = x230 & n1103 ;
  assign n4392 = n4391 ^ x81 ^ 1'b0 ;
  assign n4393 = n1030 & n4392 ;
  assign n4394 = ( n1288 & n4173 ) | ( n1288 & n4393 ) | ( n4173 & n4393 ) ;
  assign n4397 = ( n1179 & n1703 ) | ( n1179 & ~n4137 ) | ( n1703 & ~n4137 ) ;
  assign n4396 = n3403 ^ n1837 ^ n594 ;
  assign n4395 = n3904 ^ n3046 ^ n1982 ;
  assign n4398 = n4397 ^ n4396 ^ n4395 ;
  assign n4399 = n4398 ^ n3873 ^ 1'b0 ;
  assign n4402 = ( ~n324 & n512 ) | ( ~n324 & n3054 ) | ( n512 & n3054 ) ;
  assign n4403 = ( n1665 & n3075 ) | ( n1665 & ~n4402 ) | ( n3075 & ~n4402 ) ;
  assign n4400 = ~n1489 & n2968 ;
  assign n4401 = ~n1623 & n4400 ;
  assign n4404 = n4403 ^ n4401 ^ 1'b0 ;
  assign n4405 = n2676 ^ n1382 ^ 1'b0 ;
  assign n4406 = n2471 & ~n4061 ;
  assign n4407 = n3587 & n4406 ;
  assign n4408 = x140 | n874 ;
  assign n4409 = ( ~n322 & n1298 ) | ( ~n322 & n4408 ) | ( n1298 & n4408 ) ;
  assign n4413 = n666 ^ x231 ^ x191 ;
  assign n4410 = n1777 ^ n436 ^ x236 ;
  assign n4411 = n4410 ^ n2841 ^ 1'b0 ;
  assign n4412 = ~n3738 & n4411 ;
  assign n4414 = n4413 ^ n4412 ^ n1709 ;
  assign n4415 = n4409 & n4414 ;
  assign n4416 = n4079 ^ n2732 ^ n1015 ;
  assign n4419 = n1047 ^ n892 ^ 1'b0 ;
  assign n4420 = n1967 & ~n4419 ;
  assign n4421 = ( x129 & ~n3224 ) | ( x129 & n4420 ) | ( ~n3224 & n4420 ) ;
  assign n4417 = n3036 & ~n3203 ;
  assign n4418 = n1384 & n4417 ;
  assign n4422 = n4421 ^ n4418 ^ 1'b0 ;
  assign n4423 = n4422 ^ n2679 ^ 1'b0 ;
  assign n4424 = n4416 & n4423 ;
  assign n4425 = n4076 ^ n775 ^ n275 ;
  assign n4430 = ( x13 & ~n446 ) | ( x13 & n531 ) | ( ~n446 & n531 ) ;
  assign n4431 = ~n3097 & n4027 ;
  assign n4432 = n4430 & ~n4431 ;
  assign n4433 = n836 & n4432 ;
  assign n4426 = x126 & n1832 ;
  assign n4427 = n4336 ^ n3773 ^ 1'b0 ;
  assign n4428 = n883 & ~n4427 ;
  assign n4429 = n4426 & n4428 ;
  assign n4434 = n4433 ^ n4429 ^ 1'b0 ;
  assign n4436 = n408 | n1293 ;
  assign n4437 = n4436 ^ n2187 ^ 1'b0 ;
  assign n4435 = ~n692 & n1990 ;
  assign n4438 = n4437 ^ n4435 ^ n768 ;
  assign n4439 = ( n1197 & ~n1849 ) | ( n1197 & n3849 ) | ( ~n1849 & n3849 ) ;
  assign n4440 = n967 & n4439 ;
  assign n4441 = n3177 ^ n988 ^ n778 ;
  assign n4442 = ( n2215 & n4440 ) | ( n2215 & n4441 ) | ( n4440 & n4441 ) ;
  assign n4443 = ~n3703 & n4442 ;
  assign n4444 = n2040 ^ x202 ^ 1'b0 ;
  assign n4445 = n3094 & ~n4444 ;
  assign n4446 = n1689 ^ n792 ^ n341 ;
  assign n4447 = ~n3124 & n4446 ;
  assign n4448 = ~n4445 & n4447 ;
  assign n4449 = n4448 ^ n1940 ^ n1423 ;
  assign n4450 = n3870 ^ n2592 ^ n848 ;
  assign n4451 = x65 & n4450 ;
  assign n4452 = ( n844 & n2316 ) | ( n844 & n4451 ) | ( n2316 & n4451 ) ;
  assign n4453 = n3221 ^ x12 ^ 1'b0 ;
  assign n4454 = n4453 ^ n3130 ^ n2752 ;
  assign n4465 = ( x5 & ~n591 ) | ( x5 & n1440 ) | ( ~n591 & n1440 ) ;
  assign n4464 = x48 & ~n279 ;
  assign n4455 = ~n1398 & n1997 ;
  assign n4456 = n4455 ^ n916 ^ 1'b0 ;
  assign n4457 = ~n660 & n1414 ;
  assign n4458 = ~n4456 & n4457 ;
  assign n4459 = ~n466 & n2608 ;
  assign n4460 = ~n3530 & n4459 ;
  assign n4461 = n1302 & n1790 ;
  assign n4462 = n4461 ^ n2166 ^ 1'b0 ;
  assign n4463 = ( ~n4458 & n4460 ) | ( ~n4458 & n4462 ) | ( n4460 & n4462 ) ;
  assign n4466 = n4465 ^ n4464 ^ n4463 ;
  assign n4467 = n3156 ^ n1396 ^ 1'b0 ;
  assign n4468 = ( ~n1616 & n1893 ) | ( ~n1616 & n2071 ) | ( n1893 & n2071 ) ;
  assign n4469 = n4468 ^ x250 ^ 1'b0 ;
  assign n4470 = ( ~n3061 & n4266 ) | ( ~n3061 & n4469 ) | ( n4266 & n4469 ) ;
  assign n4471 = n2359 ^ n1311 ^ 1'b0 ;
  assign n4472 = x16 & n1135 ;
  assign n4473 = ~n4471 & n4472 ;
  assign n4474 = n4473 ^ x125 ^ 1'b0 ;
  assign n4481 = ( ~n1355 & n1780 ) | ( ~n1355 & n1970 ) | ( n1780 & n1970 ) ;
  assign n4478 = ( ~x35 & n2356 ) | ( ~x35 & n3261 ) | ( n2356 & n3261 ) ;
  assign n4479 = ( ~n675 & n1105 ) | ( ~n675 & n4478 ) | ( n1105 & n4478 ) ;
  assign n4475 = n4359 ^ n2295 ^ n2079 ;
  assign n4476 = ( n438 & n742 ) | ( n438 & ~n4475 ) | ( n742 & ~n4475 ) ;
  assign n4477 = n917 | n4476 ;
  assign n4480 = n4479 ^ n4477 ^ n1888 ;
  assign n4482 = n4481 ^ n4480 ^ 1'b0 ;
  assign n4483 = ~n4474 & n4482 ;
  assign n4484 = ~n3178 & n3692 ;
  assign n4485 = n871 | n1138 ;
  assign n4486 = x196 | n4485 ;
  assign n4487 = n4484 | n4486 ;
  assign n4488 = ( n1262 & n2510 ) | ( n1262 & ~n4375 ) | ( n2510 & ~n4375 ) ;
  assign n4489 = n799 & n2051 ;
  assign n4490 = n1047 | n4489 ;
  assign n4491 = n4490 ^ n3710 ^ n3417 ;
  assign n4492 = n4491 ^ n3487 ^ n1962 ;
  assign n4493 = n3987 ^ n2928 ^ n897 ;
  assign n4494 = ( n1418 & ~n3177 ) | ( n1418 & n4493 ) | ( ~n3177 & n4493 ) ;
  assign n4495 = n3476 ^ n1786 ^ n1144 ;
  assign n4496 = ~n490 & n4495 ;
  assign n4497 = n4496 ^ n1367 ^ 1'b0 ;
  assign n4498 = n4497 ^ n4466 ^ n3458 ;
  assign n4499 = n4307 ^ n2810 ^ n421 ;
  assign n4503 = n601 | n3503 ;
  assign n4504 = n778 & ~n4503 ;
  assign n4505 = n4504 ^ n2176 ^ n500 ;
  assign n4501 = n3331 ^ n1558 ^ n1340 ;
  assign n4502 = ~n2755 & n4501 ;
  assign n4506 = n4505 ^ n4502 ^ n4022 ;
  assign n4500 = n4178 ^ n1145 ^ 1'b0 ;
  assign n4507 = n4506 ^ n4500 ^ n3723 ;
  assign n4508 = n1100 ^ n573 ^ x75 ;
  assign n4509 = n4508 ^ n3681 ^ 1'b0 ;
  assign n4510 = ~n885 & n4509 ;
  assign n4511 = ~n1783 & n2504 ;
  assign n4512 = ~n4510 & n4511 ;
  assign n4513 = n4512 ^ n3254 ^ 1'b0 ;
  assign n4514 = n3113 & n4513 ;
  assign n4515 = n401 | n871 ;
  assign n4516 = n1129 & ~n4515 ;
  assign n4517 = n4516 ^ n2312 ^ 1'b0 ;
  assign n4521 = ( n681 & n925 ) | ( n681 & ~n1370 ) | ( n925 & ~n1370 ) ;
  assign n4522 = ( x199 & n1395 ) | ( x199 & n4521 ) | ( n1395 & n4521 ) ;
  assign n4518 = ( n724 & n912 ) | ( n724 & n3505 ) | ( n912 & n3505 ) ;
  assign n4519 = ( n1644 & ~n2530 ) | ( n1644 & n4518 ) | ( ~n2530 & n4518 ) ;
  assign n4520 = n4519 ^ n3878 ^ n3368 ;
  assign n4523 = n4522 ^ n4520 ^ n1508 ;
  assign n4524 = ( x54 & ~x75 ) | ( x54 & n911 ) | ( ~x75 & n911 ) ;
  assign n4525 = ( ~n803 & n1144 ) | ( ~n803 & n4524 ) | ( n1144 & n4524 ) ;
  assign n4526 = n746 & ~n3412 ;
  assign n4527 = ( n1977 & n2094 ) | ( n1977 & n4526 ) | ( n2094 & n4526 ) ;
  assign n4528 = n4527 ^ n3991 ^ n2526 ;
  assign n4529 = ( ~n877 & n1703 ) | ( ~n877 & n4528 ) | ( n1703 & n4528 ) ;
  assign n4530 = ( n2739 & n4525 ) | ( n2739 & ~n4529 ) | ( n4525 & ~n4529 ) ;
  assign n4531 = x125 & ~n4530 ;
  assign n4532 = ~n2495 & n4531 ;
  assign n4533 = n3185 ^ n977 ^ n819 ;
  assign n4534 = n2212 & n4533 ;
  assign n4535 = ( n4106 & n4532 ) | ( n4106 & ~n4534 ) | ( n4532 & ~n4534 ) ;
  assign n4536 = ( n3753 & n4523 ) | ( n3753 & n4535 ) | ( n4523 & n4535 ) ;
  assign n4537 = ( n4017 & ~n4517 ) | ( n4017 & n4536 ) | ( ~n4517 & n4536 ) ;
  assign n4538 = n939 & ~n2183 ;
  assign n4539 = ( x87 & n1458 ) | ( x87 & n2804 ) | ( n1458 & n2804 ) ;
  assign n4540 = n4538 & n4539 ;
  assign n4541 = n4540 ^ n1224 ^ 1'b0 ;
  assign n4542 = ~x105 & n1125 ;
  assign n4543 = n4542 ^ n268 ^ 1'b0 ;
  assign n4544 = x227 & n4543 ;
  assign n4545 = ~n2212 & n4544 ;
  assign n4546 = ~n842 & n4545 ;
  assign n4547 = n3542 ^ n3259 ^ 1'b0 ;
  assign n4553 = ( ~n1669 & n2210 ) | ( ~n1669 & n3143 ) | ( n2210 & n3143 ) ;
  assign n4548 = x140 & n705 ;
  assign n4549 = ~n1079 & n4548 ;
  assign n4550 = n4549 ^ n1108 ^ 1'b0 ;
  assign n4551 = n2113 | n4550 ;
  assign n4552 = n4551 ^ n2392 ^ n1089 ;
  assign n4554 = n4553 ^ n4552 ^ x64 ;
  assign n4555 = n4554 ^ n3431 ^ 1'b0 ;
  assign n4556 = ( n923 & n2556 ) | ( n923 & n3073 ) | ( n2556 & n3073 ) ;
  assign n4557 = n4083 ^ n3425 ^ 1'b0 ;
  assign n4558 = x78 & n4557 ;
  assign n4559 = ~n690 & n2957 ;
  assign n4560 = ( ~n4556 & n4558 ) | ( ~n4556 & n4559 ) | ( n4558 & n4559 ) ;
  assign n4561 = n1141 | n1158 ;
  assign n4562 = n517 & ~n4561 ;
  assign n4563 = n1555 ^ x22 ^ 1'b0 ;
  assign n4568 = n1592 ^ n1479 ^ 1'b0 ;
  assign n4569 = n4568 ^ n2295 ^ 1'b0 ;
  assign n4570 = ( n696 & n2700 ) | ( n696 & ~n4569 ) | ( n2700 & ~n4569 ) ;
  assign n4571 = n840 & n4570 ;
  assign n4564 = n998 ^ n286 ^ 1'b0 ;
  assign n4565 = x110 & ~n4564 ;
  assign n4566 = n1575 & n4565 ;
  assign n4567 = n727 | n4566 ;
  assign n4572 = n4571 ^ n4567 ^ 1'b0 ;
  assign n4573 = n4563 & ~n4572 ;
  assign n4574 = n4573 ^ n1772 ^ 1'b0 ;
  assign n4575 = ( n1078 & n1524 ) | ( n1078 & n2515 ) | ( n1524 & n2515 ) ;
  assign n4576 = n3406 ^ n1195 ^ 1'b0 ;
  assign n4577 = n3666 & ~n4576 ;
  assign n4578 = n4577 ^ n3460 ^ 1'b0 ;
  assign n4579 = ~n4575 & n4578 ;
  assign n4580 = n3116 ^ n806 ^ n418 ;
  assign n4581 = n4580 ^ n2407 ^ 1'b0 ;
  assign n4584 = n2080 ^ n563 ^ 1'b0 ;
  assign n4582 = n603 ^ n307 ^ 1'b0 ;
  assign n4583 = n4582 ^ n2102 ^ n301 ;
  assign n4585 = n4584 ^ n4583 ^ n2384 ;
  assign n4586 = n4208 ^ n1148 ^ n734 ;
  assign n4587 = n4586 ^ n3273 ^ n2114 ;
  assign n4588 = n2352 & n2661 ;
  assign n4589 = n3177 & n4588 ;
  assign n4592 = n3056 ^ n2107 ^ 1'b0 ;
  assign n4593 = n4556 ^ n622 ^ n305 ;
  assign n4594 = n4593 ^ n920 ^ n654 ;
  assign n4595 = n718 ^ x212 ^ x139 ;
  assign n4596 = n608 & n4595 ;
  assign n4597 = n4241 ^ n526 ^ 1'b0 ;
  assign n4598 = n4596 & n4597 ;
  assign n4599 = ( ~n4592 & n4594 ) | ( ~n4592 & n4598 ) | ( n4594 & n4598 ) ;
  assign n4600 = ~n2556 & n4599 ;
  assign n4601 = n4600 ^ n4075 ^ 1'b0 ;
  assign n4590 = n550 | n2556 ;
  assign n4591 = n4590 ^ n1644 ^ 1'b0 ;
  assign n4602 = n4601 ^ n4591 ^ 1'b0 ;
  assign n4603 = n1235 ^ n1220 ^ 1'b0 ;
  assign n4604 = ( n1837 & ~n1863 ) | ( n1837 & n4603 ) | ( ~n1863 & n4603 ) ;
  assign n4605 = n4604 ^ n2549 ^ n836 ;
  assign n4612 = n3186 ^ n920 ^ n722 ;
  assign n4613 = n4612 ^ n2135 ^ n1197 ;
  assign n4609 = n2076 ^ n999 ^ 1'b0 ;
  assign n4606 = n1646 ^ x161 ^ 1'b0 ;
  assign n4607 = n4606 ^ n4316 ^ 1'b0 ;
  assign n4608 = n394 & n4607 ;
  assign n4610 = n4609 ^ n4608 ^ n1267 ;
  assign n4611 = n4610 ^ n408 ^ x27 ;
  assign n4614 = n4613 ^ n4611 ^ 1'b0 ;
  assign n4615 = n2686 | n4614 ;
  assign n4616 = n1126 | n4615 ;
  assign n4617 = n1089 | n4616 ;
  assign n4618 = n2528 ^ n1071 ^ n954 ;
  assign n4619 = n4618 ^ n3152 ^ n1918 ;
  assign n4620 = x27 & ~n2448 ;
  assign n4621 = n4620 ^ x19 ^ 1'b0 ;
  assign n4622 = n4621 ^ n4499 ^ n604 ;
  assign n4623 = n4195 ^ n2623 ^ n2048 ;
  assign n4624 = ~n3593 & n3600 ;
  assign n4630 = ( ~n1249 & n2106 ) | ( ~n1249 & n2222 ) | ( n2106 & n2222 ) ;
  assign n4631 = ~n454 & n4630 ;
  assign n4632 = n4631 ^ n2529 ^ 1'b0 ;
  assign n4626 = ( n1058 & n1315 ) | ( n1058 & ~n4234 ) | ( n1315 & ~n4234 ) ;
  assign n4627 = n2962 ^ n627 ^ 1'b0 ;
  assign n4628 = n4627 ^ x72 ^ 1'b0 ;
  assign n4629 = ~n4626 & n4628 ;
  assign n4625 = n2066 ^ n963 ^ x29 ;
  assign n4633 = n4632 ^ n4629 ^ n4625 ;
  assign n4634 = ( x86 & n586 ) | ( x86 & ~n1251 ) | ( n586 & ~n1251 ) ;
  assign n4635 = n4634 ^ n2406 ^ n1909 ;
  assign n4636 = ( n2917 & ~n4311 ) | ( n2917 & n4635 ) | ( ~n4311 & n4635 ) ;
  assign n4637 = ~n549 & n1732 ;
  assign n4638 = ~n2388 & n4637 ;
  assign n4639 = n4638 ^ n3984 ^ n2829 ;
  assign n4640 = n974 | n3543 ;
  assign n4641 = ( n1191 & n2256 ) | ( n1191 & ~n4640 ) | ( n2256 & ~n4640 ) ;
  assign n4645 = n2210 ^ n2204 ^ n557 ;
  assign n4646 = n4645 ^ n1895 ^ n464 ;
  assign n4642 = n640 ^ n531 ^ x76 ;
  assign n4643 = n4642 ^ n3184 ^ 1'b0 ;
  assign n4644 = n1798 & ~n4643 ;
  assign n4647 = n4646 ^ n4644 ^ n2332 ;
  assign n4648 = n4641 & n4647 ;
  assign n4649 = n4648 ^ n4155 ^ 1'b0 ;
  assign n4653 = n3947 ^ n625 ^ x226 ;
  assign n4652 = ( n1193 & n2187 ) | ( n1193 & n4295 ) | ( n2187 & n4295 ) ;
  assign n4650 = n1694 ^ n1621 ^ 1'b0 ;
  assign n4651 = ( ~n1786 & n3203 ) | ( ~n1786 & n4650 ) | ( n3203 & n4650 ) ;
  assign n4654 = n4653 ^ n4652 ^ n4651 ;
  assign n4655 = ~n2558 & n4654 ;
  assign n4656 = n2804 & n4655 ;
  assign n4657 = n685 | n1145 ;
  assign n4658 = n2639 & ~n4657 ;
  assign n4659 = n4658 ^ n648 ^ x130 ;
  assign n4660 = n4659 ^ n3982 ^ 1'b0 ;
  assign n4661 = n4660 ^ n2370 ^ 1'b0 ;
  assign n4662 = n1585 & n4133 ;
  assign n4663 = n3403 ^ n1450 ^ 1'b0 ;
  assign n4664 = n1485 | n4663 ;
  assign n4665 = n1777 ^ n656 ^ 1'b0 ;
  assign n4666 = n282 & ~n4665 ;
  assign n4667 = n4666 ^ n2899 ^ 1'b0 ;
  assign n4668 = n4664 | n4667 ;
  assign n4669 = n1373 | n2373 ;
  assign n4670 = n4669 ^ n1073 ^ 1'b0 ;
  assign n4671 = n2382 ^ x167 ^ 1'b0 ;
  assign n4672 = ( ~x147 & n1122 ) | ( ~x147 & n2885 ) | ( n1122 & n2885 ) ;
  assign n4673 = ( n2666 & ~n3959 ) | ( n2666 & n4672 ) | ( ~n3959 & n4672 ) ;
  assign n4674 = n3317 ^ n1281 ^ n778 ;
  assign n4675 = n2175 & ~n4674 ;
  assign n4676 = n4675 ^ n3919 ^ 1'b0 ;
  assign n4677 = n1460 | n4676 ;
  assign n4678 = n1639 & ~n4677 ;
  assign n4679 = n763 & ~n1657 ;
  assign n4680 = n4679 ^ n1278 ^ 1'b0 ;
  assign n4681 = n1621 & ~n2746 ;
  assign n4682 = n2100 ^ n1863 ^ n1323 ;
  assign n4683 = n4682 ^ n271 ^ 1'b0 ;
  assign n4684 = ~n4681 & n4683 ;
  assign n4685 = ~n4680 & n4684 ;
  assign n4686 = ( n2495 & ~n4237 ) | ( n2495 & n4685 ) | ( ~n4237 & n4685 ) ;
  assign n4687 = ~n1921 & n4090 ;
  assign n4688 = ( n1816 & ~n4686 ) | ( n1816 & n4687 ) | ( ~n4686 & n4687 ) ;
  assign n4690 = ~n810 & n1220 ;
  assign n4691 = ~n584 & n4690 ;
  assign n4692 = n4691 ^ n2000 ^ n1219 ;
  assign n4693 = n4692 ^ n2695 ^ 1'b0 ;
  assign n4689 = n3370 & ~n4086 ;
  assign n4694 = n4693 ^ n4689 ^ 1'b0 ;
  assign n4697 = ( ~n505 & n2248 ) | ( ~n505 & n3621 ) | ( n2248 & n3621 ) ;
  assign n4695 = n4090 & ~n4674 ;
  assign n4696 = n4695 ^ n2091 ^ 1'b0 ;
  assign n4698 = n4697 ^ n4696 ^ n2260 ;
  assign n4699 = n4294 ^ n3370 ^ 1'b0 ;
  assign n4700 = n3050 | n4699 ;
  assign n4702 = x117 & n879 ;
  assign n4701 = n3826 ^ n3493 ^ n1054 ;
  assign n4703 = n4702 ^ n4701 ^ n3369 ;
  assign n4704 = ~n870 & n4326 ;
  assign n4705 = n4704 ^ n433 ^ 1'b0 ;
  assign n4706 = ( x194 & n2777 ) | ( x194 & n3522 ) | ( n2777 & n3522 ) ;
  assign n4707 = ( n3288 & ~n4705 ) | ( n3288 & n4706 ) | ( ~n4705 & n4706 ) ;
  assign n4714 = x228 & n374 ;
  assign n4708 = x230 & x236 ;
  assign n4709 = ~n410 & n4708 ;
  assign n4710 = n2551 & ~n4709 ;
  assign n4711 = n301 & ~n2601 ;
  assign n4712 = n4711 ^ n822 ^ 1'b0 ;
  assign n4713 = n4710 & n4712 ;
  assign n4715 = n4714 ^ n4713 ^ 1'b0 ;
  assign n4716 = ~n4707 & n4715 ;
  assign n4717 = n4716 ^ n4480 ^ n2384 ;
  assign n4721 = n3638 ^ n429 ^ x41 ;
  assign n4722 = n4721 ^ n1359 ^ n1258 ;
  assign n4720 = ( ~n952 & n1945 ) | ( ~n952 & n2071 ) | ( n1945 & n2071 ) ;
  assign n4723 = n4722 ^ n4720 ^ 1'b0 ;
  assign n4719 = n2923 | n3128 ;
  assign n4724 = n4723 ^ n4719 ^ 1'b0 ;
  assign n4725 = n4724 ^ n2996 ^ n2283 ;
  assign n4718 = n1479 & n3407 ;
  assign n4726 = n4725 ^ n4718 ^ 1'b0 ;
  assign n4727 = n423 & ~n2697 ;
  assign n4728 = ( ~x236 & n1616 ) | ( ~x236 & n4727 ) | ( n1616 & n4727 ) ;
  assign n4729 = ~n1998 & n4728 ;
  assign n4730 = n1888 ^ n1804 ^ n1047 ;
  assign n4731 = ~n4047 & n4730 ;
  assign n4732 = n4074 & n4731 ;
  assign n4733 = n4732 ^ n2097 ^ 1'b0 ;
  assign n4734 = n3252 ^ n326 ^ 1'b0 ;
  assign n4735 = ( n1997 & n2576 ) | ( n1997 & n4674 ) | ( n2576 & n4674 ) ;
  assign n4736 = n478 & ~n4735 ;
  assign n4737 = n4736 ^ n1538 ^ 1'b0 ;
  assign n4738 = n4734 & n4737 ;
  assign n4739 = n1179 & ~n3861 ;
  assign n4740 = n745 & n4739 ;
  assign n4741 = ( n2214 & ~n3902 ) | ( n2214 & n4740 ) | ( ~n3902 & n4740 ) ;
  assign n4744 = n1351 & ~n2475 ;
  assign n4745 = n1978 & ~n4744 ;
  assign n4742 = n1311 & n1793 ;
  assign n4743 = n1460 & n4742 ;
  assign n4746 = n4745 ^ n4743 ^ n2889 ;
  assign n4747 = ( n3313 & n4741 ) | ( n3313 & n4746 ) | ( n4741 & n4746 ) ;
  assign n4748 = x213 & n4747 ;
  assign n4749 = ~n1023 & n2951 ;
  assign n4750 = ~n800 & n4749 ;
  assign n4751 = n1710 & ~n2061 ;
  assign n4752 = n1622 & n4751 ;
  assign n4753 = n786 & n4752 ;
  assign n4754 = ( ~n643 & n2867 ) | ( ~n643 & n4630 ) | ( n2867 & n4630 ) ;
  assign n4755 = ~n1432 & n4754 ;
  assign n4756 = n3991 ^ n1833 ^ n859 ;
  assign n4757 = ( x90 & ~n1447 ) | ( x90 & n2076 ) | ( ~n1447 & n2076 ) ;
  assign n4758 = n3474 | n3767 ;
  assign n4759 = n4758 ^ n3670 ^ 1'b0 ;
  assign n4760 = ( ~n1504 & n4757 ) | ( ~n1504 & n4759 ) | ( n4757 & n4759 ) ;
  assign n4761 = ( n2928 & n3173 ) | ( n2928 & n4760 ) | ( n3173 & n4760 ) ;
  assign n4762 = ( ~n2319 & n3212 ) | ( ~n2319 & n4761 ) | ( n3212 & n4761 ) ;
  assign n4763 = ( ~n939 & n4756 ) | ( ~n939 & n4762 ) | ( n4756 & n4762 ) ;
  assign n4764 = n2325 & ~n3985 ;
  assign n4765 = n587 | n4764 ;
  assign n4766 = n3981 ^ n3971 ^ n520 ;
  assign n4767 = n2430 ^ x28 ^ 1'b0 ;
  assign n4768 = n4767 ^ n4301 ^ n610 ;
  assign n4769 = n1416 & ~n4768 ;
  assign n4770 = n1545 & ~n3945 ;
  assign n4771 = ( x245 & ~n900 ) | ( x245 & n4770 ) | ( ~n900 & n4770 ) ;
  assign n4772 = n4771 ^ n3211 ^ n1713 ;
  assign n4773 = n4772 ^ n3945 ^ 1'b0 ;
  assign n4774 = ( x106 & ~n428 ) | ( x106 & n2079 ) | ( ~n428 & n2079 ) ;
  assign n4775 = n2128 | n4774 ;
  assign n4776 = n4775 ^ n1458 ^ n399 ;
  assign n4777 = n4776 ^ n2065 ^ n363 ;
  assign n4778 = n418 & ~n1230 ;
  assign n4779 = ( n2152 & n2230 ) | ( n2152 & ~n4778 ) | ( n2230 & ~n4778 ) ;
  assign n4780 = n4095 ^ n3475 ^ 1'b0 ;
  assign n4781 = n1274 | n4780 ;
  assign n4783 = n4090 ^ n776 ^ 1'b0 ;
  assign n4784 = ( x22 & n765 ) | ( x22 & ~n4783 ) | ( n765 & ~n4783 ) ;
  assign n4782 = n1164 & ~n1401 ;
  assign n4785 = n4784 ^ n4782 ^ n4528 ;
  assign n4786 = ~n256 & n3697 ;
  assign n4787 = n1198 | n4117 ;
  assign n4790 = n902 & n954 ;
  assign n4791 = ~x147 & n4790 ;
  assign n4788 = n3155 ^ n2466 ^ n2160 ;
  assign n4789 = n4788 ^ n4169 ^ 1'b0 ;
  assign n4792 = n4791 ^ n4789 ^ 1'b0 ;
  assign n4793 = ~n3673 & n4792 ;
  assign n4794 = n3582 ^ n2662 ^ n2246 ;
  assign n4795 = ( x218 & n2810 ) | ( x218 & n4395 ) | ( n2810 & n4395 ) ;
  assign n4796 = n1938 ^ n700 ^ 1'b0 ;
  assign n4797 = n3167 & ~n4796 ;
  assign n4798 = n4797 ^ n3556 ^ 1'b0 ;
  assign n4799 = n2193 | n2820 ;
  assign n4800 = n1846 | n4799 ;
  assign n4801 = n4691 ^ n2374 ^ x247 ;
  assign n4802 = n4801 ^ n3013 ^ n791 ;
  assign n4803 = n4802 ^ n2905 ^ 1'b0 ;
  assign n4804 = n3317 & ~n4803 ;
  assign n4805 = x232 & ~n2028 ;
  assign n4806 = n1299 & n4805 ;
  assign n4807 = n1593 ^ n1525 ^ x205 ;
  assign n4808 = ( ~n1544 & n3445 ) | ( ~n1544 & n4807 ) | ( n3445 & n4807 ) ;
  assign n4809 = n4808 ^ n4653 ^ 1'b0 ;
  assign n4810 = ~n4806 & n4809 ;
  assign n4811 = n1020 & n4810 ;
  assign n4814 = ( n1108 & n1837 ) | ( n1108 & n2652 ) | ( n1837 & n2652 ) ;
  assign n4812 = n2053 ^ n1694 ^ 1'b0 ;
  assign n4813 = n2736 & ~n4812 ;
  assign n4815 = n4814 ^ n4813 ^ n4478 ;
  assign n4816 = n416 | n2049 ;
  assign n4817 = n556 | n1424 ;
  assign n4818 = n957 & n1830 ;
  assign n4819 = n2315 & ~n4818 ;
  assign n4820 = ~x105 & n3544 ;
  assign n4821 = n1513 & n3315 ;
  assign n4822 = n553 ^ n364 ^ 1'b0 ;
  assign n4823 = n1299 | n4571 ;
  assign n4824 = n2933 | n4823 ;
  assign n4825 = ( ~n565 & n4822 ) | ( ~n565 & n4824 ) | ( n4822 & n4824 ) ;
  assign n4828 = n2196 ^ n784 ^ x117 ;
  assign n4826 = ( ~x12 & n2008 ) | ( ~x12 & n3507 ) | ( n2008 & n3507 ) ;
  assign n4827 = n4826 ^ n1083 ^ n688 ;
  assign n4829 = n4828 ^ n4827 ^ n1118 ;
  assign n4830 = ( n329 & n1201 ) | ( n329 & ~n3398 ) | ( n1201 & ~n3398 ) ;
  assign n4831 = n4830 ^ n2208 ^ x198 ;
  assign n4832 = n4831 ^ n1838 ^ 1'b0 ;
  assign n4833 = n4829 & ~n4832 ;
  assign n4834 = ( x100 & n293 ) | ( x100 & ~n567 ) | ( n293 & ~n567 ) ;
  assign n4835 = n761 | n4834 ;
  assign n4836 = n4835 ^ n2092 ^ 1'b0 ;
  assign n4839 = x141 & ~n1587 ;
  assign n4837 = n4692 ^ n3439 ^ n2240 ;
  assign n4838 = n395 & n4837 ;
  assign n4840 = n4839 ^ n4838 ^ 1'b0 ;
  assign n4841 = ( n360 & ~n4836 ) | ( n360 & n4840 ) | ( ~n4836 & n4840 ) ;
  assign n4842 = n368 | n1266 ;
  assign n4843 = n1475 ^ n1118 ^ 1'b0 ;
  assign n4844 = ~n2031 & n4843 ;
  assign n4845 = n3130 & ~n3287 ;
  assign n4846 = ~n4844 & n4845 ;
  assign n4847 = ( n2571 & n4248 ) | ( n2571 & n4846 ) | ( n4248 & n4846 ) ;
  assign n4848 = n1408 ^ n287 ^ 1'b0 ;
  assign n4849 = ~n778 & n2095 ;
  assign n4850 = n4848 & n4849 ;
  assign n4851 = ( n4735 & n4847 ) | ( n4735 & ~n4850 ) | ( n4847 & ~n4850 ) ;
  assign n4860 = n2602 ^ x119 ^ 1'b0 ;
  assign n4861 = x207 & n4860 ;
  assign n4852 = n2898 ^ n995 ^ 1'b0 ;
  assign n4853 = n2072 & ~n4852 ;
  assign n4854 = ~n3498 & n4853 ;
  assign n4855 = n2847 & n4854 ;
  assign n4856 = n4855 ^ n3710 ^ 1'b0 ;
  assign n4857 = n1012 & ~n4856 ;
  assign n4858 = n4857 ^ n2632 ^ 1'b0 ;
  assign n4859 = n4858 ^ n1702 ^ 1'b0 ;
  assign n4862 = n4861 ^ n4859 ^ n3515 ;
  assign n4863 = ( n789 & n1746 ) | ( n789 & n4672 ) | ( n1746 & n4672 ) ;
  assign n4864 = ( n526 & ~n1894 ) | ( n526 & n4863 ) | ( ~n1894 & n4863 ) ;
  assign n4865 = ( ~x229 & n1545 ) | ( ~x229 & n2422 ) | ( n1545 & n2422 ) ;
  assign n4866 = x53 | n3391 ;
  assign n4867 = n4865 | n4866 ;
  assign n4868 = n4867 ^ n4011 ^ 1'b0 ;
  assign n4869 = n4868 ^ n4592 ^ n2806 ;
  assign n4870 = n1876 & ~n4869 ;
  assign n4871 = n4864 & n4870 ;
  assign n4872 = n3343 ^ n1989 ^ 1'b0 ;
  assign n4873 = ~n957 & n4633 ;
  assign n4874 = ( n805 & n1789 ) | ( n805 & ~n3124 ) | ( n1789 & ~n3124 ) ;
  assign n4875 = n4874 ^ n3479 ^ n763 ;
  assign n4876 = n2137 & ~n3696 ;
  assign n4877 = n4876 ^ n1331 ^ n516 ;
  assign n4878 = n4877 ^ n3779 ^ n3257 ;
  assign n4881 = n1789 ^ n1010 ^ 1'b0 ;
  assign n4879 = n929 & n4412 ;
  assign n4880 = ~n690 & n4879 ;
  assign n4882 = n4881 ^ n4880 ^ 1'b0 ;
  assign n4883 = n4878 | n4882 ;
  assign n4884 = n1177 | n4723 ;
  assign n4885 = n4384 ^ n1587 ^ n1084 ;
  assign n4886 = n4885 ^ n2537 ^ x197 ;
  assign n4891 = ~n1097 & n2701 ;
  assign n4892 = n1948 & n4891 ;
  assign n4887 = n1463 & n2117 ;
  assign n4888 = n4887 ^ n1538 ^ 1'b0 ;
  assign n4889 = n2271 ^ n389 ^ 1'b0 ;
  assign n4890 = n4888 & ~n4889 ;
  assign n4893 = n4892 ^ n4890 ^ 1'b0 ;
  assign n4894 = n4554 ^ n638 ^ 1'b0 ;
  assign n4895 = n4893 & ~n4894 ;
  assign n4896 = ( ~n3097 & n4886 ) | ( ~n3097 & n4895 ) | ( n4886 & n4895 ) ;
  assign n4897 = n4896 ^ n4165 ^ n3851 ;
  assign n4898 = n2481 | n3156 ;
  assign n4899 = n4898 ^ n759 ^ 1'b0 ;
  assign n4900 = n3090 & n4256 ;
  assign n4901 = n2550 | n2889 ;
  assign n4902 = n1276 | n4901 ;
  assign n4903 = n4209 & ~n4902 ;
  assign n4904 = n4900 & n4903 ;
  assign n4905 = n2756 ^ n2676 ^ n1072 ;
  assign n4906 = n4905 ^ x247 ^ 1'b0 ;
  assign n4907 = x199 & ~n3749 ;
  assign n4908 = ~n892 & n4907 ;
  assign n4909 = n2475 | n4908 ;
  assign n4910 = n3034 & ~n4909 ;
  assign n4911 = n4906 & ~n4910 ;
  assign n4912 = n4911 ^ n3191 ^ 1'b0 ;
  assign n4913 = ( n2309 & n4815 ) | ( n2309 & ~n4912 ) | ( n4815 & ~n4912 ) ;
  assign n4914 = n2061 ^ n1732 ^ 1'b0 ;
  assign n4919 = n4396 ^ n2238 ^ 1'b0 ;
  assign n4920 = ~n2372 & n4919 ;
  assign n4916 = n4066 ^ n1098 ^ 1'b0 ;
  assign n4917 = n4333 | n4916 ;
  assign n4918 = n1109 & ~n4917 ;
  assign n4921 = n4920 ^ n4918 ^ 1'b0 ;
  assign n4915 = n317 & n2054 ;
  assign n4922 = n4921 ^ n4915 ^ 1'b0 ;
  assign n4923 = n898 | n4521 ;
  assign n4924 = n843 & n1414 ;
  assign n4925 = n4924 ^ n2254 ^ n2036 ;
  assign n4926 = n4925 ^ n4042 ^ n2806 ;
  assign n4927 = n3703 ^ n1140 ^ 1'b0 ;
  assign n4928 = n283 | n1352 ;
  assign n4929 = n4928 ^ n1699 ^ 1'b0 ;
  assign n4930 = ( n582 & n1846 ) | ( n582 & n4929 ) | ( n1846 & n4929 ) ;
  assign n4931 = n4640 & n4930 ;
  assign n4932 = ~n2524 & n4931 ;
  assign n4938 = n3758 ^ n3005 ^ n1457 ;
  assign n4933 = n1485 ^ n700 ^ 1'b0 ;
  assign n4934 = n2641 | n4933 ;
  assign n4935 = n983 ^ n335 ^ 1'b0 ;
  assign n4936 = ~n4934 & n4935 ;
  assign n4937 = n894 & ~n4936 ;
  assign n4939 = n4938 ^ n4937 ^ n4231 ;
  assign n4940 = n3187 | n4346 ;
  assign n4941 = n2557 | n4940 ;
  assign n4942 = ( ~n722 & n1924 ) | ( ~n722 & n2917 ) | ( n1924 & n2917 ) ;
  assign n4943 = n4942 ^ n3323 ^ n1924 ;
  assign n4944 = n4885 | n4943 ;
  assign n4945 = n2288 & ~n4944 ;
  assign n4946 = n2160 ^ n587 ^ 1'b0 ;
  assign n4947 = n4779 & n4941 ;
  assign n4948 = n2114 & n4947 ;
  assign n4949 = n4376 ^ n1224 ^ 1'b0 ;
  assign n4950 = ( ~n1059 & n1294 ) | ( ~n1059 & n2895 ) | ( n1294 & n2895 ) ;
  assign n4951 = ( n2412 & n4001 ) | ( n2412 & ~n4950 ) | ( n4001 & ~n4950 ) ;
  assign n4952 = n3656 ^ n1700 ^ n1508 ;
  assign n4953 = n2382 ^ n1274 ^ 1'b0 ;
  assign n4954 = n4650 | n4953 ;
  assign n4955 = n332 & n1770 ;
  assign n4956 = n4955 ^ n854 ^ 1'b0 ;
  assign n4957 = n4956 ^ n2896 ^ 1'b0 ;
  assign n4958 = n4173 | n4957 ;
  assign n4960 = x136 & ~n287 ;
  assign n4961 = n4960 ^ n1525 ^ x240 ;
  assign n4962 = ( ~n562 & n4371 ) | ( ~n562 & n4961 ) | ( n4371 & n4961 ) ;
  assign n4959 = n685 | n3474 ;
  assign n4963 = n4962 ^ n4959 ^ 1'b0 ;
  assign n4964 = n2945 ^ n1500 ^ 1'b0 ;
  assign n4965 = n3717 & n4964 ;
  assign n4966 = n4965 ^ n2224 ^ n1666 ;
  assign n4967 = n4966 ^ n4291 ^ n2694 ;
  assign n4968 = n4626 | n4967 ;
  assign n4969 = n2052 | n4968 ;
  assign n4970 = n4615 ^ n1310 ^ 1'b0 ;
  assign n4971 = n312 & ~n4970 ;
  assign n4972 = ( ~n1375 & n2486 ) | ( ~n1375 & n3648 ) | ( n2486 & n3648 ) ;
  assign n4973 = n1655 & ~n4972 ;
  assign n4974 = n4973 ^ x226 ^ 1'b0 ;
  assign n4975 = ( n1730 & ~n4173 ) | ( n1730 & n4974 ) | ( ~n4173 & n4974 ) ;
  assign n4976 = n4975 ^ n3798 ^ n2706 ;
  assign n4977 = ( ~n421 & n4532 ) | ( ~n421 & n4618 ) | ( n4532 & n4618 ) ;
  assign n4978 = n625 | n2315 ;
  assign n4979 = n1948 ^ n1830 ^ 1'b0 ;
  assign n4980 = n710 & ~n4979 ;
  assign n4981 = n4978 | n4980 ;
  assign n4982 = n4781 ^ n2780 ^ x129 ;
  assign n4983 = n1803 | n2720 ;
  assign n4984 = n4983 ^ n2848 ^ n2121 ;
  assign n4988 = ( ~n1079 & n2067 ) | ( ~n1079 & n4974 ) | ( n2067 & n4974 ) ;
  assign n4989 = ( n1998 & ~n2965 ) | ( n1998 & n4988 ) | ( ~n2965 & n4988 ) ;
  assign n4985 = n2269 ^ n2042 ^ n1962 ;
  assign n4986 = n3626 & ~n4985 ;
  assign n4987 = n1201 & n4986 ;
  assign n4990 = n4989 ^ n4987 ^ x199 ;
  assign n4991 = ( ~x194 & n817 ) | ( ~x194 & n1279 ) | ( n817 & n1279 ) ;
  assign n4992 = ~n640 & n2392 ;
  assign n4993 = n4992 ^ n2077 ^ 1'b0 ;
  assign n4994 = n4993 ^ n934 ^ 1'b0 ;
  assign n4995 = ( n925 & ~n4991 ) | ( n925 & n4994 ) | ( ~n4991 & n4994 ) ;
  assign n4996 = n2624 & ~n2780 ;
  assign n4997 = ( n351 & ~n3242 ) | ( n351 & n4996 ) | ( ~n3242 & n4996 ) ;
  assign n4999 = n2562 ^ n561 ^ n530 ;
  assign n5000 = n4999 ^ n3331 ^ 1'b0 ;
  assign n5001 = n533 | n5000 ;
  assign n4998 = ( n502 & n1550 ) | ( n502 & n2797 ) | ( n1550 & n2797 ) ;
  assign n5002 = n5001 ^ n4998 ^ 1'b0 ;
  assign n5003 = ( x85 & n385 ) | ( x85 & n1018 ) | ( n385 & n1018 ) ;
  assign n5004 = n5003 ^ n1055 ^ n610 ;
  assign n5005 = n5004 ^ n1393 ^ x219 ;
  assign n5006 = n5005 ^ n3896 ^ 1'b0 ;
  assign n5007 = n3061 ^ n2230 ^ n2160 ;
  assign n5008 = n3497 ^ n2382 ^ n1953 ;
  assign n5009 = n3646 | n5008 ;
  assign n5010 = n529 & ~n5009 ;
  assign n5011 = n5007 & ~n5010 ;
  assign n5012 = ~n4705 & n5011 ;
  assign n5013 = ~n356 & n1530 ;
  assign n5014 = ~n1007 & n3912 ;
  assign n5015 = ( ~n2014 & n2620 ) | ( ~n2014 & n3510 ) | ( n2620 & n3510 ) ;
  assign n5016 = n466 | n1858 ;
  assign n5017 = n706 & ~n5016 ;
  assign n5018 = n3806 ^ n1628 ^ n770 ;
  assign n5019 = n5018 ^ n2614 ^ 1'b0 ;
  assign n5020 = ~n2978 & n5019 ;
  assign n5021 = n5020 ^ n3779 ^ 1'b0 ;
  assign n5022 = n5017 | n5021 ;
  assign n5023 = n1720 & n1945 ;
  assign n5024 = n2920 & n5023 ;
  assign n5025 = ( x211 & n2313 ) | ( x211 & n5024 ) | ( n2313 & n5024 ) ;
  assign n5026 = ( x75 & n647 ) | ( x75 & n923 ) | ( n647 & n923 ) ;
  assign n5027 = ( n4740 & n4926 ) | ( n4740 & n5026 ) | ( n4926 & n5026 ) ;
  assign n5028 = n4486 ^ n690 ^ 1'b0 ;
  assign n5029 = ( n304 & n2393 ) | ( n304 & n3092 ) | ( n2393 & n3092 ) ;
  assign n5030 = x227 | n5029 ;
  assign n5031 = n5030 ^ n723 ^ 1'b0 ;
  assign n5032 = n5028 & n5031 ;
  assign n5033 = n606 | n5032 ;
  assign n5034 = n3237 ^ n3225 ^ n1086 ;
  assign n5035 = n1684 & ~n5034 ;
  assign n5036 = n5035 ^ n1401 ^ 1'b0 ;
  assign n5037 = ( ~n1978 & n2947 ) | ( ~n1978 & n5036 ) | ( n2947 & n5036 ) ;
  assign n5038 = x94 | n5001 ;
  assign n5039 = n4645 ^ n1797 ^ x220 ;
  assign n5040 = n5039 ^ n3634 ^ n1302 ;
  assign n5043 = n3532 ^ n737 ^ n505 ;
  assign n5041 = ( x177 & n531 ) | ( x177 & ~n798 ) | ( n531 & ~n798 ) ;
  assign n5042 = ( n2267 & n3412 ) | ( n2267 & ~n5041 ) | ( n3412 & ~n5041 ) ;
  assign n5044 = n5043 ^ n5042 ^ n2675 ;
  assign n5045 = n2077 | n3019 ;
  assign n5046 = n5044 | n5045 ;
  assign n5052 = n4930 ^ n1198 ^ x144 ;
  assign n5049 = n3279 ^ n1573 ^ n273 ;
  assign n5050 = n861 | n5049 ;
  assign n5047 = ~n565 & n4638 ;
  assign n5048 = ( n1233 & ~n1971 ) | ( n1233 & n5047 ) | ( ~n1971 & n5047 ) ;
  assign n5051 = n5050 ^ n5048 ^ n4651 ;
  assign n5053 = n5052 ^ n5051 ^ 1'b0 ;
  assign n5054 = ( ~n4007 & n4674 ) | ( ~n4007 & n5053 ) | ( n4674 & n5053 ) ;
  assign n5055 = n774 & ~n2080 ;
  assign n5056 = ~n423 & n5055 ;
  assign n5057 = ( ~n2182 & n2692 ) | ( ~n2182 & n5056 ) | ( n2692 & n5056 ) ;
  assign n5058 = n445 & ~n2751 ;
  assign n5059 = ~n3808 & n5058 ;
  assign n5060 = n2779 ^ n1374 ^ 1'b0 ;
  assign n5061 = n5060 ^ n1416 ^ x150 ;
  assign n5062 = n301 & ~n5061 ;
  assign n5063 = n1724 & n5062 ;
  assign n5064 = n2582 ^ n2562 ^ n1193 ;
  assign n5065 = n5064 ^ n2234 ^ n852 ;
  assign n5066 = ( n2907 & n5063 ) | ( n2907 & n5065 ) | ( n5063 & n5065 ) ;
  assign n5086 = ( n1211 & ~n1701 ) | ( n1211 & n2076 ) | ( ~n1701 & n2076 ) ;
  assign n5082 = n1164 ^ n830 ^ n563 ;
  assign n5083 = n5082 ^ n3849 ^ 1'b0 ;
  assign n5084 = n1776 | n5083 ;
  assign n5080 = n4653 ^ n551 ^ 1'b0 ;
  assign n5081 = ~n3870 & n5080 ;
  assign n5076 = n3245 ^ n2887 ^ n1169 ;
  assign n5075 = n499 & n1230 ;
  assign n5077 = n5076 ^ n5075 ^ n394 ;
  assign n5078 = n2404 | n5077 ;
  assign n5079 = n5078 ^ n2102 ^ 1'b0 ;
  assign n5085 = n5084 ^ n5081 ^ n5079 ;
  assign n5067 = x16 & n312 ;
  assign n5068 = n5067 ^ x252 ^ 1'b0 ;
  assign n5069 = ( ~n1358 & n2063 ) | ( ~n1358 & n5068 ) | ( n2063 & n5068 ) ;
  assign n5070 = n2651 | n5069 ;
  assign n5071 = n5070 ^ n3058 ^ 1'b0 ;
  assign n5072 = ( n851 & n2205 ) | ( n851 & ~n2259 ) | ( n2205 & ~n2259 ) ;
  assign n5073 = ~n740 & n5072 ;
  assign n5074 = ~n5071 & n5073 ;
  assign n5087 = n5086 ^ n5085 ^ n5074 ;
  assign n5088 = ( n2574 & n3963 ) | ( n2574 & n4208 ) | ( n3963 & n4208 ) ;
  assign n5089 = n5088 ^ n2602 ^ 1'b0 ;
  assign n5090 = n453 | n5089 ;
  assign n5091 = n5090 ^ n2803 ^ n494 ;
  assign n5092 = n1892 ^ x200 ^ x11 ;
  assign n5093 = n2246 & n5092 ;
  assign n5094 = ( ~n2538 & n3549 ) | ( ~n2538 & n5093 ) | ( n3549 & n5093 ) ;
  assign n5095 = n1423 ^ n785 ^ 1'b0 ;
  assign n5096 = n1717 & ~n5095 ;
  assign n5097 = n5096 ^ n2538 ^ 1'b0 ;
  assign n5098 = n5097 ^ n4523 ^ n3046 ;
  assign n5099 = n1664 ^ n994 ^ x180 ;
  assign n5100 = x92 & ~n5099 ;
  assign n5101 = n2329 & n5100 ;
  assign n5105 = n3216 ^ x114 ^ 1'b0 ;
  assign n5106 = ~n1779 & n5105 ;
  assign n5102 = n4085 ^ n1743 ^ x125 ;
  assign n5103 = n5072 ^ x82 ^ 1'b0 ;
  assign n5104 = ~n5102 & n5103 ;
  assign n5107 = n5106 ^ n5104 ^ 1'b0 ;
  assign n5108 = n1827 & n5107 ;
  assign n5109 = x56 & ~n3256 ;
  assign n5110 = n5109 ^ n1370 ^ 1'b0 ;
  assign n5111 = n5110 ^ n3310 ^ n2525 ;
  assign n5112 = n5111 ^ n1198 ^ n408 ;
  assign n5113 = n1351 & ~n2810 ;
  assign n5114 = n5113 ^ n695 ^ 1'b0 ;
  assign n5115 = n5114 ^ n3783 ^ n3505 ;
  assign n5116 = n5115 ^ n4844 ^ n487 ;
  assign n5117 = ~n257 & n701 ;
  assign n5118 = ~n1643 & n5117 ;
  assign n5119 = n3841 ^ n3415 ^ 1'b0 ;
  assign n5120 = n1129 | n3237 ;
  assign n5121 = n1682 & ~n5120 ;
  assign n5122 = n5119 | n5121 ;
  assign n5123 = n1031 & ~n5122 ;
  assign n5124 = n1440 & ~n2482 ;
  assign n5125 = ~n1160 & n5124 ;
  assign n5126 = n5125 ^ n681 ^ x236 ;
  assign n5127 = n5126 ^ n1646 ^ 1'b0 ;
  assign n5128 = n2866 ^ n1772 ^ n662 ;
  assign n5129 = n2217 ^ n1793 ^ n1054 ;
  assign n5130 = n279 | n5129 ;
  assign n5131 = n5128 | n5130 ;
  assign n5132 = n3587 ^ n686 ^ 1'b0 ;
  assign n5133 = ~n962 & n2008 ;
  assign n5134 = ( ~n3787 & n5132 ) | ( ~n3787 & n5133 ) | ( n5132 & n5133 ) ;
  assign n5135 = n4404 & n4589 ;
  assign n5136 = n1095 ^ n286 ^ 1'b0 ;
  assign n5137 = n1071 & ~n5136 ;
  assign n5138 = n4510 ^ n980 ^ 1'b0 ;
  assign n5139 = n2131 & n5138 ;
  assign n5140 = n306 & n5086 ;
  assign n5141 = n3600 ^ n1896 ^ n1331 ;
  assign n5142 = n5141 ^ n2887 ^ x251 ;
  assign n5144 = n864 | n1305 ;
  assign n5145 = n600 & ~n5144 ;
  assign n5143 = x129 & ~n1981 ;
  assign n5146 = n5145 ^ n5143 ^ 1'b0 ;
  assign n5152 = n3479 ^ n471 ^ 1'b0 ;
  assign n5153 = ( n732 & n1376 ) | ( n732 & ~n2958 ) | ( n1376 & ~n2958 ) ;
  assign n5154 = n5152 | n5153 ;
  assign n5155 = n5154 ^ x57 ^ 1'b0 ;
  assign n5147 = n3672 ^ n1138 ^ n1086 ;
  assign n5148 = n1465 ^ x88 ^ 1'b0 ;
  assign n5149 = ~n5147 & n5148 ;
  assign n5150 = ( n1022 & n2860 ) | ( n1022 & ~n5149 ) | ( n2860 & ~n5149 ) ;
  assign n5151 = n2012 | n5150 ;
  assign n5156 = n5155 ^ n5151 ^ 1'b0 ;
  assign n5157 = n5146 & n5156 ;
  assign n5158 = n2812 & n5157 ;
  assign n5159 = ~n1155 & n4373 ;
  assign n5163 = n1798 ^ n1691 ^ n997 ;
  assign n5161 = n1241 & ~n4568 ;
  assign n5162 = n5161 ^ n2640 ^ 1'b0 ;
  assign n5160 = n320 | n4255 ;
  assign n5164 = n5163 ^ n5162 ^ n5160 ;
  assign n5165 = n5164 ^ n3358 ^ n1040 ;
  assign n5166 = n3370 ^ n1428 ^ x168 ;
  assign n5167 = n1730 & ~n4988 ;
  assign n5168 = n5167 ^ n1623 ^ 1'b0 ;
  assign n5169 = x207 & n2615 ;
  assign n5170 = n5169 ^ n3070 ^ 1'b0 ;
  assign n5171 = n3704 & ~n5170 ;
  assign n5172 = ( n2639 & n5092 ) | ( n2639 & ~n5171 ) | ( n5092 & ~n5171 ) ;
  assign n5173 = ( x83 & n5168 ) | ( x83 & n5172 ) | ( n5168 & n5172 ) ;
  assign n5174 = n1525 | n2986 ;
  assign n5175 = x51 | n5174 ;
  assign n5176 = n721 & n2928 ;
  assign n5177 = ( n1050 & n3095 ) | ( n1050 & ~n5176 ) | ( n3095 & ~n5176 ) ;
  assign n5178 = n3889 & n5177 ;
  assign n5179 = n2351 & n5178 ;
  assign n5180 = n1473 | n5179 ;
  assign n5181 = ~n3440 & n5180 ;
  assign n5182 = n5181 ^ n2474 ^ 1'b0 ;
  assign n5183 = ( n1193 & n4937 ) | ( n1193 & ~n5182 ) | ( n4937 & ~n5182 ) ;
  assign n5184 = ( n1431 & n3252 ) | ( n1431 & ~n5183 ) | ( n3252 & ~n5183 ) ;
  assign n5187 = n1825 ^ n1462 ^ 1'b0 ;
  assign n5188 = x147 & ~n5187 ;
  assign n5185 = x232 & ~n1961 ;
  assign n5186 = n1926 & n5185 ;
  assign n5189 = n5188 ^ n5186 ^ n4681 ;
  assign n5190 = n5189 ^ n2185 ^ 1'b0 ;
  assign n5191 = ~x36 & n5190 ;
  assign n5192 = n5191 ^ n2348 ^ 1'b0 ;
  assign n5193 = ( n1136 & ~n1288 ) | ( n1136 & n1614 ) | ( ~n1288 & n1614 ) ;
  assign n5194 = n5193 ^ n3509 ^ n2889 ;
  assign n5195 = n4586 ^ n3335 ^ n1968 ;
  assign n5196 = n1849 ^ n1756 ^ 1'b0 ;
  assign n5197 = n2981 ^ n2662 ^ 1'b0 ;
  assign n5198 = ~n1202 & n3425 ;
  assign n5199 = n5198 ^ n2400 ^ 1'b0 ;
  assign n5200 = n2009 | n5199 ;
  assign n5201 = ~n1783 & n4612 ;
  assign n5202 = n5200 & n5201 ;
  assign n5205 = n1014 ^ x111 ^ x107 ;
  assign n5203 = n768 & ~n3037 ;
  assign n5204 = n5203 ^ n1340 ^ 1'b0 ;
  assign n5206 = n5205 ^ n5204 ^ n3986 ;
  assign n5208 = x147 & ~n1005 ;
  assign n5207 = ~n1346 & n5065 ;
  assign n5209 = n5208 ^ n5207 ^ 1'b0 ;
  assign n5210 = n3716 | n4062 ;
  assign n5211 = n5210 ^ n3151 ^ 1'b0 ;
  assign n5212 = n5211 ^ n489 ^ 1'b0 ;
  assign n5213 = n2121 ^ n1280 ^ n351 ;
  assign n5214 = ( ~n4606 & n5212 ) | ( ~n4606 & n5213 ) | ( n5212 & n5213 ) ;
  assign n5215 = n5214 ^ n1842 ^ 1'b0 ;
  assign n5216 = n5215 ^ n4933 ^ 1'b0 ;
  assign n5217 = n2271 ^ n2121 ^ 1'b0 ;
  assign n5218 = ~n595 & n5217 ;
  assign n5219 = ~n443 & n471 ;
  assign n5220 = ~x133 & n5219 ;
  assign n5221 = n3092 | n5220 ;
  assign n5222 = n2545 & n5221 ;
  assign n5223 = x137 & ~n1025 ;
  assign n5224 = n5223 ^ n3163 ^ n2569 ;
  assign n5225 = n5224 ^ n4500 ^ n3195 ;
  assign n5226 = n5042 ^ n4348 ^ n2848 ;
  assign n5230 = ~n2120 & n3403 ;
  assign n5228 = n2372 ^ n1440 ^ n1408 ;
  assign n5227 = ( ~n681 & n1657 ) | ( ~n681 & n3103 ) | ( n1657 & n3103 ) ;
  assign n5229 = n5228 ^ n5227 ^ n291 ;
  assign n5231 = n5230 ^ n5229 ^ n1743 ;
  assign n5232 = ( ~n859 & n2413 ) | ( ~n859 & n5177 ) | ( n2413 & n5177 ) ;
  assign n5233 = n2803 ^ n1834 ^ 1'b0 ;
  assign n5234 = n5232 & n5233 ;
  assign n5235 = n5234 ^ n4950 ^ n1879 ;
  assign n5236 = n3042 ^ n1448 ^ n784 ;
  assign n5237 = n5236 ^ n4576 ^ n4003 ;
  assign n5238 = n3792 ^ n475 ^ 1'b0 ;
  assign n5239 = ( n911 & ~n5237 ) | ( n911 & n5238 ) | ( ~n5237 & n5238 ) ;
  assign n5240 = ~n739 & n3709 ;
  assign n5241 = n5240 ^ n1640 ^ 1'b0 ;
  assign n5250 = n608 & ~n1304 ;
  assign n5251 = n5250 ^ n1432 ^ 1'b0 ;
  assign n5252 = ( n403 & n1837 ) | ( n403 & n5251 ) | ( n1837 & n5251 ) ;
  assign n5253 = ( ~n286 & n3456 ) | ( ~n286 & n5252 ) | ( n3456 & n5252 ) ;
  assign n5245 = ( ~x227 & n1346 ) | ( ~x227 & n2434 ) | ( n1346 & n2434 ) ;
  assign n5246 = ( ~n401 & n1845 ) | ( ~n401 & n5245 ) | ( n1845 & n5245 ) ;
  assign n5247 = n425 & ~n5246 ;
  assign n5248 = ~n2326 & n5247 ;
  assign n5242 = n1826 ^ n1820 ^ n738 ;
  assign n5243 = n865 | n5242 ;
  assign n5244 = n5243 ^ n893 ^ 1'b0 ;
  assign n5249 = n5248 ^ n5244 ^ n2261 ;
  assign n5254 = n5253 ^ n5249 ^ n776 ;
  assign n5255 = n5254 ^ n4090 ^ 1'b0 ;
  assign n5256 = ~n5241 & n5255 ;
  assign n5261 = n1317 & n2210 ;
  assign n5262 = n5261 ^ n4003 ^ 1'b0 ;
  assign n5260 = ~n2708 & n4028 ;
  assign n5258 = ~n3358 & n4293 ;
  assign n5257 = n3968 ^ n1341 ^ 1'b0 ;
  assign n5259 = n5258 ^ n5257 ^ n2627 ;
  assign n5263 = n5262 ^ n5260 ^ n5259 ;
  assign n5264 = ( n4759 & n5256 ) | ( n4759 & ~n5263 ) | ( n5256 & ~n5263 ) ;
  assign n5265 = ( n401 & n550 ) | ( n401 & ~n1352 ) | ( n550 & ~n1352 ) ;
  assign n5266 = n5265 ^ n2631 ^ n1102 ;
  assign n5267 = n5266 ^ n4757 ^ x79 ;
  assign n5268 = ( n1387 & n2157 ) | ( n1387 & n5267 ) | ( n2157 & n5267 ) ;
  assign n5269 = n1743 ^ n1323 ^ 1'b0 ;
  assign n5270 = ( n1481 & n2588 ) | ( n1481 & ~n5269 ) | ( n2588 & ~n5269 ) ;
  assign n5271 = n2856 & ~n5270 ;
  assign n5272 = ( n3495 & n5268 ) | ( n3495 & ~n5271 ) | ( n5268 & ~n5271 ) ;
  assign n5273 = n2720 ^ n1982 ^ 1'b0 ;
  assign n5274 = x186 & n506 ;
  assign n5275 = n5273 & n5274 ;
  assign n5276 = n2148 ^ x56 ^ 1'b0 ;
  assign n5277 = n266 & ~n648 ;
  assign n5278 = n5277 ^ n2597 ^ n737 ;
  assign n5279 = n4138 ^ n1920 ^ 1'b0 ;
  assign n5280 = n5279 ^ x150 ^ 1'b0 ;
  assign n5281 = ~n1354 & n5280 ;
  assign n5282 = ( n2788 & ~n3626 ) | ( n2788 & n5281 ) | ( ~n3626 & n5281 ) ;
  assign n5283 = ( n1989 & n2142 ) | ( n1989 & ~n3844 ) | ( n2142 & ~n3844 ) ;
  assign n5284 = ( ~n2018 & n2753 ) | ( ~n2018 & n2886 ) | ( n2753 & n2886 ) ;
  assign n5285 = n3377 ^ n2920 ^ 1'b0 ;
  assign n5286 = n2606 & ~n5285 ;
  assign n5287 = ~n5284 & n5286 ;
  assign n5288 = n3010 & ~n5287 ;
  assign n5293 = n1972 ^ x33 ^ 1'b0 ;
  assign n5292 = n1614 | n3283 ;
  assign n5294 = n5293 ^ n5292 ^ 1'b0 ;
  assign n5289 = n3967 & ~n4917 ;
  assign n5290 = n1769 & n5289 ;
  assign n5291 = n2773 | n5290 ;
  assign n5295 = n5294 ^ n5291 ^ 1'b0 ;
  assign n5298 = n3701 ^ n1193 ^ n737 ;
  assign n5296 = n2595 | n3125 ;
  assign n5297 = n5296 ^ n1340 ^ 1'b0 ;
  assign n5299 = n5298 ^ n5297 ^ n857 ;
  assign n5300 = n3246 ^ n1419 ^ 1'b0 ;
  assign n5301 = n5300 ^ n2168 ^ n1045 ;
  assign n5302 = n1235 ^ n918 ^ n401 ;
  assign n5303 = n5302 ^ n4602 ^ n2283 ;
  assign n5304 = ~n296 & n2176 ;
  assign n5305 = n5304 ^ x22 ^ 1'b0 ;
  assign n5306 = n1303 & ~n5305 ;
  assign n5307 = n5306 ^ n1901 ^ 1'b0 ;
  assign n5308 = ~n453 & n1382 ;
  assign n5309 = ~n5307 & n5308 ;
  assign n5310 = n5309 ^ n3791 ^ n2898 ;
  assign n5315 = n2865 ^ n884 ^ 1'b0 ;
  assign n5316 = x46 & n5315 ;
  assign n5317 = n5316 ^ n4169 ^ x185 ;
  assign n5312 = n5163 ^ n4426 ^ n1186 ;
  assign n5311 = ( n718 & n1905 ) | ( n718 & n4802 ) | ( n1905 & n4802 ) ;
  assign n5313 = n5312 ^ n5311 ^ n2882 ;
  assign n5314 = ~n4830 & n5313 ;
  assign n5318 = n5317 ^ n5314 ^ 1'b0 ;
  assign n5319 = n798 & n5318 ;
  assign n5320 = n4484 & n5319 ;
  assign n5321 = n4956 ^ n3340 ^ n673 ;
  assign n5322 = n3314 & n5321 ;
  assign n5323 = n5322 ^ n4293 ^ n3523 ;
  assign n5324 = n436 & ~n3825 ;
  assign n5325 = n5324 ^ n1366 ^ 1'b0 ;
  assign n5326 = n5325 ^ n4841 ^ n1545 ;
  assign n5327 = n4993 ^ n4668 ^ n721 ;
  assign n5328 = n3458 ^ n1909 ^ n1358 ;
  assign n5329 = n5328 ^ n3636 ^ n1609 ;
  assign n5330 = n4740 ^ n4101 ^ 1'b0 ;
  assign n5331 = n755 & n2707 ;
  assign n5332 = ~n5330 & n5331 ;
  assign n5337 = n1156 ^ n569 ^ 1'b0 ;
  assign n5336 = n4864 ^ n1967 ^ n618 ;
  assign n5333 = n831 & n847 ;
  assign n5334 = n1664 | n5333 ;
  assign n5335 = n5334 ^ n980 ^ 1'b0 ;
  assign n5338 = n5337 ^ n5336 ^ n5335 ;
  assign n5339 = ( n5329 & n5332 ) | ( n5329 & n5338 ) | ( n5332 & n5338 ) ;
  assign n5341 = n1131 ^ n840 ^ n796 ;
  assign n5340 = n3111 | n5034 ;
  assign n5342 = n5341 ^ n5340 ^ 1'b0 ;
  assign n5343 = n5342 ^ n4338 ^ n2443 ;
  assign n5344 = ( n1358 & n2608 ) | ( n1358 & n4211 ) | ( n2608 & n4211 ) ;
  assign n5345 = n5344 ^ n2541 ^ 1'b0 ;
  assign n5346 = n2776 ^ n2652 ^ n2200 ;
  assign n5347 = ( ~x88 & x208 ) | ( ~x88 & n5346 ) | ( x208 & n5346 ) ;
  assign n5348 = n2965 & n4608 ;
  assign n5349 = ( ~n394 & n842 ) | ( ~n394 & n1524 ) | ( n842 & n1524 ) ;
  assign n5350 = n5349 ^ n2583 ^ x179 ;
  assign n5352 = n2737 ^ n739 ^ x174 ;
  assign n5351 = ( n1302 & n2478 ) | ( n1302 & n4362 ) | ( n2478 & n4362 ) ;
  assign n5353 = n5352 ^ n5351 ^ 1'b0 ;
  assign n5354 = ( n2421 & n3735 ) | ( n2421 & ~n5353 ) | ( n3735 & ~n5353 ) ;
  assign n5355 = x60 & ~n3234 ;
  assign n5356 = n5355 ^ x71 ^ 1'b0 ;
  assign n5357 = n5354 & n5356 ;
  assign n5358 = ~n3000 & n5357 ;
  assign n5359 = ~n5350 & n5358 ;
  assign n5360 = x27 & n2194 ;
  assign n5361 = ~n2644 & n5360 ;
  assign n5362 = n4342 & ~n5361 ;
  assign n5365 = n1940 & ~n3626 ;
  assign n5363 = ( n341 & n2592 ) | ( n341 & ~n3811 ) | ( n2592 & ~n3811 ) ;
  assign n5364 = n5363 ^ n3314 ^ n3111 ;
  assign n5366 = n5365 ^ n5364 ^ 1'b0 ;
  assign n5367 = ~n3437 & n5366 ;
  assign n5368 = ( n893 & n1448 ) | ( n893 & ~n2487 ) | ( n1448 & ~n2487 ) ;
  assign n5369 = x237 | n3034 ;
  assign n5370 = ( ~n2571 & n3491 ) | ( ~n2571 & n5364 ) | ( n3491 & n5364 ) ;
  assign n5371 = n4066 & ~n5370 ;
  assign n5372 = n5371 ^ n1205 ^ 1'b0 ;
  assign n5373 = n3297 ^ n2273 ^ n2076 ;
  assign n5374 = n3276 & n5373 ;
  assign n5375 = n436 | n5374 ;
  assign n5376 = n2602 & ~n5375 ;
  assign n5377 = n466 | n3413 ;
  assign n5384 = n1854 ^ n1457 ^ 1'b0 ;
  assign n5385 = n2726 | n5384 ;
  assign n5386 = n647 | n5385 ;
  assign n5387 = n4608 | n5386 ;
  assign n5379 = n751 & n3458 ;
  assign n5380 = n399 & n5379 ;
  assign n5381 = n5380 ^ n2087 ^ 1'b0 ;
  assign n5382 = ~n1672 & n5381 ;
  assign n5378 = n3629 ^ n2076 ^ 1'b0 ;
  assign n5383 = n5382 ^ n5378 ^ n4483 ;
  assign n5388 = n5387 ^ n5383 ^ 1'b0 ;
  assign n5389 = ~n1985 & n1993 ;
  assign n5390 = ~n3601 & n5389 ;
  assign n5391 = n5390 ^ n2583 ^ 1'b0 ;
  assign n5392 = ~n454 & n471 ;
  assign n5393 = n2332 ^ n1980 ^ n1388 ;
  assign n5394 = n5393 ^ n2829 ^ 1'b0 ;
  assign n5399 = n2247 ^ x190 ^ 1'b0 ;
  assign n5395 = ( ~n2305 & n2895 ) | ( ~n2305 & n4828 ) | ( n2895 & n4828 ) ;
  assign n5396 = ( n1141 & n1470 ) | ( n1141 & ~n5395 ) | ( n1470 & ~n5395 ) ;
  assign n5397 = ( x254 & n1193 ) | ( x254 & ~n5396 ) | ( n1193 & ~n5396 ) ;
  assign n5398 = ~n5251 & n5397 ;
  assign n5400 = n5399 ^ n5398 ^ 1'b0 ;
  assign n5401 = ( ~n5392 & n5394 ) | ( ~n5392 & n5400 ) | ( n5394 & n5400 ) ;
  assign n5402 = n771 ^ n695 ^ 1'b0 ;
  assign n5403 = n5402 ^ n5052 ^ n4787 ;
  assign n5404 = ~n572 & n1191 ;
  assign n5407 = n1930 & ~n4791 ;
  assign n5405 = ( n1304 & n2097 ) | ( n1304 & n2401 ) | ( n2097 & n2401 ) ;
  assign n5406 = ~n3668 & n5405 ;
  assign n5408 = n5407 ^ n5406 ^ 1'b0 ;
  assign n5409 = ( n2132 & n3060 ) | ( n2132 & n5408 ) | ( n3060 & n5408 ) ;
  assign n5410 = ( n4241 & n5404 ) | ( n4241 & ~n5409 ) | ( n5404 & ~n5409 ) ;
  assign n5411 = n5410 ^ n3200 ^ n1214 ;
  assign n5412 = ( ~x78 & n1171 ) | ( ~x78 & n1196 ) | ( n1171 & n1196 ) ;
  assign n5413 = ~n5133 & n5412 ;
  assign n5414 = n4283 & n5413 ;
  assign n5415 = ( n2060 & n2100 ) | ( n2060 & n2694 ) | ( n2100 & n2694 ) ;
  assign n5416 = ~n2026 & n5415 ;
  assign n5417 = n3764 ^ n3261 ^ 1'b0 ;
  assign n5420 = n2374 ^ n1985 ^ 1'b0 ;
  assign n5418 = ~n707 & n2187 ;
  assign n5419 = n5418 ^ n2043 ^ 1'b0 ;
  assign n5421 = n5420 ^ n5419 ^ n3730 ;
  assign n5422 = x17 & ~n689 ;
  assign n5423 = ~n3297 & n5422 ;
  assign n5424 = ( n534 & ~n683 ) | ( n534 & n4217 ) | ( ~n683 & n4217 ) ;
  assign n5425 = n593 & ~n5424 ;
  assign n5426 = n5425 ^ n5055 ^ 1'b0 ;
  assign n5427 = n3283 ^ n2063 ^ 1'b0 ;
  assign n5428 = n5426 & n5427 ;
  assign n5429 = ( ~n1706 & n3564 ) | ( ~n1706 & n5428 ) | ( n3564 & n5428 ) ;
  assign n5430 = n3264 ^ n1125 ^ 1'b0 ;
  assign n5431 = n5430 ^ n4627 ^ n3675 ;
  assign n5432 = n1030 ^ x90 ^ x59 ;
  assign n5433 = n2282 ^ n1423 ^ x91 ;
  assign n5434 = n5433 ^ n5317 ^ 1'b0 ;
  assign n5435 = n5432 | n5434 ;
  assign n5436 = n3076 ^ n1475 ^ 1'b0 ;
  assign n5437 = n721 & n5436 ;
  assign n5438 = n5437 ^ n1851 ^ 1'b0 ;
  assign n5439 = n3616 & n5438 ;
  assign n5440 = n2146 | n5368 ;
  assign n5441 = ~n758 & n2469 ;
  assign n5442 = x178 & ~n3226 ;
  assign n5443 = n3360 & n5442 ;
  assign n5444 = ( n3656 & ~n5441 ) | ( n3656 & n5443 ) | ( ~n5441 & n5443 ) ;
  assign n5445 = ~n1603 & n5270 ;
  assign n5446 = n5445 ^ n1848 ^ 1'b0 ;
  assign n5447 = x15 & n1656 ;
  assign n5448 = n1102 & n5447 ;
  assign n5449 = ( n604 & n4342 ) | ( n604 & n4974 ) | ( n4342 & n4974 ) ;
  assign n5450 = n5448 & ~n5449 ;
  assign n5451 = ( n766 & n1582 ) | ( n766 & n3240 ) | ( n1582 & n3240 ) ;
  assign n5452 = n2757 & n5451 ;
  assign n5453 = ~n2778 & n2844 ;
  assign n5454 = n5453 ^ n2185 ^ 1'b0 ;
  assign n5455 = ( n1544 & n5028 ) | ( n1544 & ~n5454 ) | ( n5028 & ~n5454 ) ;
  assign n5456 = n1232 & n1856 ;
  assign n5457 = n1225 & ~n5456 ;
  assign n5458 = ~n5455 & n5457 ;
  assign n5459 = ~n692 & n819 ;
  assign n5460 = n5459 ^ n4988 ^ 1'b0 ;
  assign n5461 = n5460 ^ n3004 ^ x189 ;
  assign n5462 = n3340 ^ n2192 ^ 1'b0 ;
  assign n5463 = n2820 | n5462 ;
  assign n5464 = n1165 & n5463 ;
  assign n5465 = ( n1046 & n2541 ) | ( n1046 & ~n5464 ) | ( n2541 & ~n5464 ) ;
  assign n5468 = ( ~x107 & n462 ) | ( ~x107 & n1745 ) | ( n462 & n1745 ) ;
  assign n5466 = ~n1583 & n3308 ;
  assign n5467 = x227 & n5466 ;
  assign n5469 = n5468 ^ n5467 ^ 1'b0 ;
  assign n5470 = n5469 ^ n4532 ^ 1'b0 ;
  assign n5471 = n1020 | n3339 ;
  assign n5472 = n4771 & n5471 ;
  assign n5473 = n5472 ^ n3025 ^ 1'b0 ;
  assign n5474 = n5470 & ~n5473 ;
  assign n5475 = n2466 ^ x112 ^ 1'b0 ;
  assign n5476 = n1759 & n5036 ;
  assign n5477 = n5476 ^ n3743 ^ 1'b0 ;
  assign n5478 = ( n2416 & n5475 ) | ( n2416 & n5477 ) | ( n5475 & n5477 ) ;
  assign n5488 = ~n408 & n3707 ;
  assign n5489 = n5488 ^ n1553 ^ 1'b0 ;
  assign n5483 = x160 & x229 ;
  assign n5484 = n626 & n5483 ;
  assign n5485 = n5484 ^ n1981 ^ 1'b0 ;
  assign n5486 = n519 & n5485 ;
  assign n5479 = n1390 & n2885 ;
  assign n5480 = n1429 & n5479 ;
  assign n5481 = n3064 | n5480 ;
  assign n5482 = n5481 ^ n1978 ^ 1'b0 ;
  assign n5487 = n5486 ^ n5482 ^ n2960 ;
  assign n5490 = n5489 ^ n5487 ^ n1877 ;
  assign n5491 = n1195 | n5490 ;
  assign n5492 = n1948 & ~n5491 ;
  assign n5493 = n2563 ^ n685 ^ 1'b0 ;
  assign n5494 = n1625 & n5493 ;
  assign n5495 = n5494 ^ n3435 ^ n1076 ;
  assign n5496 = n4572 ^ n1664 ^ 1'b0 ;
  assign n5497 = ~n4490 & n5496 ;
  assign n5498 = n3187 ^ n840 ^ x238 ;
  assign n5499 = ( x13 & n911 ) | ( x13 & ~n1429 ) | ( n911 & ~n1429 ) ;
  assign n5500 = n5499 ^ n2811 ^ 1'b0 ;
  assign n5501 = n5500 ^ n1103 ^ x242 ;
  assign n5502 = n4756 ^ n1693 ^ n1362 ;
  assign n5503 = n2084 & ~n3200 ;
  assign n5504 = ~x226 & n5503 ;
  assign n5505 = n5502 | n5504 ;
  assign n5506 = n5505 ^ x76 ^ 1'b0 ;
  assign n5507 = n5501 | n5506 ;
  assign n5508 = n3382 | n4241 ;
  assign n5509 = n1264 & n5508 ;
  assign n5510 = n2754 & n4464 ;
  assign n5511 = n5510 ^ n3661 ^ 1'b0 ;
  assign n5512 = n5511 ^ n3067 ^ 1'b0 ;
  assign n5513 = ( n4280 & n5509 ) | ( n4280 & n5512 ) | ( n5509 & n5512 ) ;
  assign n5514 = ( n466 & ~n4529 ) | ( n466 & n5513 ) | ( ~n4529 & n5513 ) ;
  assign n5520 = n550 & ~n1139 ;
  assign n5515 = n5232 ^ n5111 ^ n3942 ;
  assign n5516 = n1738 ^ n1037 ^ n912 ;
  assign n5517 = n5516 ^ n2230 ^ 1'b0 ;
  assign n5518 = n816 | n5517 ;
  assign n5519 = ( n2106 & ~n5515 ) | ( n2106 & n5518 ) | ( ~n5515 & n5518 ) ;
  assign n5521 = n5520 ^ n5519 ^ 1'b0 ;
  assign n5522 = n791 ^ n673 ^ 1'b0 ;
  assign n5523 = n5522 ^ n3324 ^ n2448 ;
  assign n5524 = n5523 ^ n2375 ^ n394 ;
  assign n5525 = n798 & n5524 ;
  assign n5526 = n2510 & n5525 ;
  assign n5527 = x29 & n1129 ;
  assign n5528 = n271 & ~n5527 ;
  assign n5529 = n957 & n5528 ;
  assign n5530 = n4569 & n5529 ;
  assign n5531 = n5530 ^ x55 ^ 1'b0 ;
  assign n5535 = n3514 ^ n1102 ^ 1'b0 ;
  assign n5536 = n5311 & n5535 ;
  assign n5532 = n2472 ^ n2070 ^ n1708 ;
  assign n5533 = ( n1683 & ~n1928 ) | ( n1683 & n5532 ) | ( ~n1928 & n5532 ) ;
  assign n5534 = n3355 & ~n5533 ;
  assign n5537 = n5536 ^ n5534 ^ 1'b0 ;
  assign n5542 = ( n1646 & ~n2944 ) | ( n1646 & n4074 ) | ( ~n2944 & n4074 ) ;
  assign n5543 = ( n707 & n1850 ) | ( n707 & n4128 ) | ( n1850 & n4128 ) ;
  assign n5544 = ( n781 & ~n2436 ) | ( n781 & n5543 ) | ( ~n2436 & n5543 ) ;
  assign n5545 = n5544 ^ n1783 ^ 1'b0 ;
  assign n5546 = n5545 ^ n2610 ^ 1'b0 ;
  assign n5547 = ( n2096 & n5542 ) | ( n2096 & n5546 ) | ( n5542 & n5546 ) ;
  assign n5538 = n807 | n4653 ;
  assign n5539 = n5538 ^ n1164 ^ 1'b0 ;
  assign n5540 = n1628 | n5539 ;
  assign n5541 = n5540 ^ n3765 ^ 1'b0 ;
  assign n5548 = n5547 ^ n5541 ^ n3186 ;
  assign n5549 = n3753 ^ n625 ^ n401 ;
  assign n5550 = ~n3559 & n5549 ;
  assign n5551 = n5550 ^ n1146 ^ 1'b0 ;
  assign n5552 = n5012 ^ n2273 ^ 1'b0 ;
  assign n5553 = n5145 | n5552 ;
  assign n5554 = n4478 ^ n1634 ^ x121 ;
  assign n5555 = n5554 ^ n3798 ^ n3458 ;
  assign n5556 = n3176 ^ n2094 ^ n683 ;
  assign n5557 = n550 | n5556 ;
  assign n5558 = ( n4192 & n4999 ) | ( n4192 & ~n5061 ) | ( n4999 & ~n5061 ) ;
  assign n5559 = n2497 | n5558 ;
  assign n5560 = n4622 ^ n2809 ^ n711 ;
  assign n5563 = n5265 ^ n1037 ^ 1'b0 ;
  assign n5564 = ~n3174 & n5563 ;
  assign n5565 = n5564 ^ n911 ^ 1'b0 ;
  assign n5561 = n4087 ^ n2525 ^ n1525 ;
  assign n5562 = ( ~x109 & n1971 ) | ( ~x109 & n5561 ) | ( n1971 & n5561 ) ;
  assign n5566 = n5565 ^ n5562 ^ 1'b0 ;
  assign n5567 = ~x128 & n2551 ;
  assign n5569 = n3503 ^ n745 ^ 1'b0 ;
  assign n5570 = n5569 ^ n4681 ^ 1'b0 ;
  assign n5568 = ( x33 & ~x250 ) | ( x33 & n1551 ) | ( ~x250 & n1551 ) ;
  assign n5571 = n5570 ^ n5568 ^ 1'b0 ;
  assign n5572 = n5567 | n5571 ;
  assign n5573 = n5572 ^ n1077 ^ 1'b0 ;
  assign n5579 = n824 & n2648 ;
  assign n5580 = n1789 & n5579 ;
  assign n5574 = n977 ^ n491 ^ x81 ;
  assign n5575 = n5574 ^ n1311 ^ 1'b0 ;
  assign n5576 = ~n2798 & n5575 ;
  assign n5577 = n5220 ^ n1926 ^ 1'b0 ;
  assign n5578 = n5576 & n5577 ;
  assign n5581 = n5580 ^ n5578 ^ n4770 ;
  assign n5582 = n3056 | n4338 ;
  assign n5583 = n5582 ^ n1606 ^ 1'b0 ;
  assign n5584 = n2720 ^ n1827 ^ n564 ;
  assign n5585 = n5584 ^ n1343 ^ n735 ;
  assign n5586 = n697 ^ n511 ^ 1'b0 ;
  assign n5587 = n2453 & ~n5586 ;
  assign n5588 = ~n4804 & n5587 ;
  assign n5589 = n3925 ^ n1284 ^ n941 ;
  assign n5590 = n5589 ^ n1152 ^ n960 ;
  assign n5591 = n2980 | n5590 ;
  assign n5592 = n5591 ^ n923 ^ 1'b0 ;
  assign n5594 = n577 | n851 ;
  assign n5595 = n1365 | n5594 ;
  assign n5593 = n3325 ^ x112 ^ 1'b0 ;
  assign n5596 = n5595 ^ n5593 ^ n4771 ;
  assign n5597 = n683 | n3615 ;
  assign n5598 = n5597 ^ n4111 ^ 1'b0 ;
  assign n5599 = n5598 ^ n511 ^ 1'b0 ;
  assign n5600 = ( ~n941 & n1543 ) | ( ~n941 & n1980 ) | ( n1543 & n1980 ) ;
  assign n5601 = ( n489 & n1030 ) | ( n489 & n5600 ) | ( n1030 & n5600 ) ;
  assign n5602 = ( n2552 & n2769 ) | ( n2552 & n2845 ) | ( n2769 & n2845 ) ;
  assign n5603 = n470 | n5602 ;
  assign n5604 = n5601 | n5603 ;
  assign n5605 = n2004 | n2143 ;
  assign n5606 = n5605 ^ n2589 ^ 1'b0 ;
  assign n5607 = n1410 | n3051 ;
  assign n5608 = n3126 & ~n5607 ;
  assign n5609 = n617 & ~n5608 ;
  assign n5610 = x252 & ~n4375 ;
  assign n5611 = ~x4 & n5610 ;
  assign n5612 = n708 & ~n3445 ;
  assign n5613 = n5612 ^ n1734 ^ 1'b0 ;
  assign n5614 = ~n5611 & n5613 ;
  assign n5615 = ~n5609 & n5614 ;
  assign n5621 = n339 & ~n772 ;
  assign n5622 = n3550 & n5621 ;
  assign n5620 = ( n926 & n3107 ) | ( n926 & ~n3705 ) | ( n3107 & ~n3705 ) ;
  assign n5618 = n1567 | n3662 ;
  assign n5616 = n746 ^ n591 ^ 1'b0 ;
  assign n5617 = n5616 ^ n5251 ^ n4929 ;
  assign n5619 = n5618 ^ n5617 ^ n1784 ;
  assign n5623 = n5622 ^ n5620 ^ n5619 ;
  assign n5634 = ( n388 & n1410 ) | ( n388 & ~n3211 ) | ( n1410 & ~n3211 ) ;
  assign n5624 = n2126 ^ n632 ^ 1'b0 ;
  assign n5625 = n5624 ^ n2946 ^ 1'b0 ;
  assign n5626 = n374 & n5625 ;
  assign n5627 = n1393 ^ x227 ^ 1'b0 ;
  assign n5628 = n852 | n5627 ;
  assign n5629 = ~n1614 & n4065 ;
  assign n5630 = ~n5628 & n5629 ;
  assign n5631 = ~n2691 & n5630 ;
  assign n5632 = n3301 & ~n5631 ;
  assign n5633 = ~n5626 & n5632 ;
  assign n5635 = n5634 ^ n5633 ^ 1'b0 ;
  assign n5636 = n5623 | n5635 ;
  assign n5639 = n4024 ^ n914 ^ 1'b0 ;
  assign n5640 = ~n523 & n5639 ;
  assign n5638 = ( x37 & ~n560 ) | ( x37 & n3199 ) | ( ~n560 & n3199 ) ;
  assign n5637 = ( n947 & n1558 ) | ( n947 & ~n2552 ) | ( n1558 & ~n2552 ) ;
  assign n5641 = n5640 ^ n5638 ^ n5637 ;
  assign n5642 = n5641 ^ n3579 ^ n758 ;
  assign n5643 = n1793 ^ x183 ^ 1'b0 ;
  assign n5644 = n3821 & n5643 ;
  assign n5645 = n5644 ^ n4798 ^ 1'b0 ;
  assign n5646 = ( n1000 & n2709 ) | ( n1000 & n3713 ) | ( n2709 & n3713 ) ;
  assign n5647 = ( n506 & ~n1518 ) | ( n506 & n5646 ) | ( ~n1518 & n5646 ) ;
  assign n5652 = ~n1926 & n4120 ;
  assign n5653 = n5652 ^ x22 ^ 1'b0 ;
  assign n5648 = n2513 ^ n2265 ^ n544 ;
  assign n5649 = ( n315 & n4752 ) | ( n315 & n5648 ) | ( n4752 & n5648 ) ;
  assign n5650 = n582 | n1730 ;
  assign n5651 = ( x108 & n5649 ) | ( x108 & n5650 ) | ( n5649 & n5650 ) ;
  assign n5654 = n5653 ^ n5651 ^ n3306 ;
  assign n5655 = n2874 & ~n5654 ;
  assign n5656 = n1779 | n1895 ;
  assign n5657 = n5656 ^ x60 ^ 1'b0 ;
  assign n5658 = n1502 | n1955 ;
  assign n5659 = n5658 ^ n559 ^ 1'b0 ;
  assign n5660 = n5659 ^ n2184 ^ n1146 ;
  assign n5661 = n5657 & n5660 ;
  assign n5662 = n5661 ^ n1984 ^ 1'b0 ;
  assign n5663 = n3241 & n4754 ;
  assign n5664 = ( ~n1398 & n1504 ) | ( ~n1398 & n3540 ) | ( n1504 & n3540 ) ;
  assign n5665 = n5664 ^ n322 ^ 1'b0 ;
  assign n5666 = n2375 ^ n1221 ^ x101 ;
  assign n5667 = ( n788 & n1536 ) | ( n788 & n5666 ) | ( n1536 & n5666 ) ;
  assign n5668 = n2594 & ~n5667 ;
  assign n5669 = n3486 & n5668 ;
  assign n5670 = ( ~x57 & n5665 ) | ( ~x57 & n5669 ) | ( n5665 & n5669 ) ;
  assign n5671 = n3497 ^ n3166 ^ n971 ;
  assign n5672 = ( ~x142 & n347 ) | ( ~x142 & n3075 ) | ( n347 & n3075 ) ;
  assign n5673 = n5672 ^ n4409 ^ n2417 ;
  assign n5674 = n5671 & ~n5673 ;
  assign n5675 = n5674 ^ n975 ^ 1'b0 ;
  assign n5676 = ( n4086 & ~n5670 ) | ( n4086 & n5675 ) | ( ~n5670 & n5675 ) ;
  assign n5677 = n4064 ^ n1171 ^ x1 ;
  assign n5683 = n1089 & ~n2567 ;
  assign n5681 = ( n346 & ~n670 ) | ( n346 & n5309 ) | ( ~n670 & n5309 ) ;
  assign n5678 = n1652 & ~n2575 ;
  assign n5679 = ~n1225 & n5678 ;
  assign n5680 = ( n1894 & n4433 ) | ( n1894 & ~n5679 ) | ( n4433 & ~n5679 ) ;
  assign n5682 = n5681 ^ n5680 ^ n525 ;
  assign n5684 = n5683 ^ n5682 ^ n4532 ;
  assign n5685 = ~n877 & n1753 ;
  assign n5686 = n4549 ^ n2672 ^ 1'b0 ;
  assign n5687 = ( ~n4371 & n5685 ) | ( ~n4371 & n5686 ) | ( n5685 & n5686 ) ;
  assign n5688 = n3042 & n4562 ;
  assign n5689 = n5688 ^ n566 ^ 1'b0 ;
  assign n5690 = n5687 & n5689 ;
  assign n5692 = n2192 ^ n1768 ^ n1567 ;
  assign n5691 = x215 & ~n551 ;
  assign n5693 = n5692 ^ n5691 ^ 1'b0 ;
  assign n5694 = n613 | n5693 ;
  assign n5695 = n5694 ^ n1279 ^ 1'b0 ;
  assign n5696 = ( n1592 & n2371 ) | ( n1592 & ~n4942 ) | ( n2371 & ~n4942 ) ;
  assign n5697 = n3018 ^ n713 ^ 1'b0 ;
  assign n5698 = n2112 | n5697 ;
  assign n5699 = n5698 ^ n4393 ^ 1'b0 ;
  assign n5700 = n5696 | n5699 ;
  assign n5703 = ( x3 & n712 ) | ( x3 & n2187 ) | ( n712 & n2187 ) ;
  assign n5701 = n2142 ^ n1621 ^ n591 ;
  assign n5702 = n270 & ~n5701 ;
  assign n5704 = n5703 ^ n5702 ^ 1'b0 ;
  assign n5705 = ~n1524 & n5704 ;
  assign n5706 = n4255 ^ x54 ^ 1'b0 ;
  assign n5707 = n1081 & ~n5706 ;
  assign n5708 = n5707 ^ n805 ^ n656 ;
  assign n5709 = ( n1198 & ~n1216 ) | ( n1198 & n1626 ) | ( ~n1216 & n1626 ) ;
  assign n5710 = ( n2576 & n3815 ) | ( n2576 & ~n4162 ) | ( n3815 & ~n4162 ) ;
  assign n5711 = ( n4104 & n5709 ) | ( n4104 & ~n5710 ) | ( n5709 & ~n5710 ) ;
  assign n5712 = ( n3051 & n5708 ) | ( n3051 & n5711 ) | ( n5708 & n5711 ) ;
  assign n5713 = n1856 ^ n903 ^ n460 ;
  assign n5714 = n3139 ^ n2583 ^ n1990 ;
  assign n5715 = n5714 ^ n3443 ^ n2739 ;
  assign n5716 = n2992 & ~n5715 ;
  assign n5717 = n5716 ^ n3826 ^ 1'b0 ;
  assign n5718 = ( n2118 & n2256 ) | ( n2118 & ~n3283 ) | ( n2256 & ~n3283 ) ;
  assign n5719 = n5718 ^ n5351 ^ n1639 ;
  assign n5720 = ( n843 & ~n933 ) | ( n843 & n5719 ) | ( ~n933 & n5719 ) ;
  assign n5721 = ( n5713 & ~n5717 ) | ( n5713 & n5720 ) | ( ~n5717 & n5720 ) ;
  assign n5722 = n3900 ^ n3787 ^ n2605 ;
  assign n5723 = n5341 ^ n2028 ^ 1'b0 ;
  assign n5724 = n5723 ^ n4401 ^ n462 ;
  assign n5725 = ( n789 & ~n5465 ) | ( n789 & n5724 ) | ( ~n5465 & n5724 ) ;
  assign n5726 = ( n1637 & n2359 ) | ( n1637 & n2530 ) | ( n2359 & n2530 ) ;
  assign n5727 = ( x126 & n2899 ) | ( x126 & n5726 ) | ( n2899 & n5726 ) ;
  assign n5728 = n5727 ^ n2174 ^ 1'b0 ;
  assign n5729 = n5728 ^ n3455 ^ n1815 ;
  assign n5730 = ( x108 & n2347 ) | ( x108 & ~n5729 ) | ( n2347 & ~n5729 ) ;
  assign n5731 = ~n1620 & n2501 ;
  assign n5732 = n796 & ~n1771 ;
  assign n5733 = ( n914 & n4499 ) | ( n914 & ~n5732 ) | ( n4499 & ~n5732 ) ;
  assign n5734 = ~n5112 & n5733 ;
  assign n5735 = n5386 ^ n4027 ^ n2635 ;
  assign n5736 = n917 | n3268 ;
  assign n5737 = n5736 ^ n2979 ^ 1'b0 ;
  assign n5738 = n1163 | n5737 ;
  assign n5739 = ( ~n2639 & n4645 ) | ( ~n2639 & n4775 ) | ( n4645 & n4775 ) ;
  assign n5744 = n2424 | n3087 ;
  assign n5740 = ( ~n526 & n671 ) | ( ~n526 & n795 ) | ( n671 & n795 ) ;
  assign n5741 = n2775 ^ n2130 ^ 1'b0 ;
  assign n5742 = ( n3240 & n3540 ) | ( n3240 & ~n5741 ) | ( n3540 & ~n5741 ) ;
  assign n5743 = n5740 & ~n5742 ;
  assign n5745 = n5744 ^ n5743 ^ 1'b0 ;
  assign n5746 = ( x172 & n5739 ) | ( x172 & ~n5745 ) | ( n5739 & ~n5745 ) ;
  assign n5748 = n3204 | n4293 ;
  assign n5747 = n4408 ^ n2828 ^ n422 ;
  assign n5749 = n5748 ^ n5747 ^ n4011 ;
  assign n5750 = ( n884 & ~n5746 ) | ( n884 & n5749 ) | ( ~n5746 & n5749 ) ;
  assign n5751 = n5738 & ~n5750 ;
  assign n5752 = n5751 ^ n1923 ^ 1'b0 ;
  assign n5753 = ( n1393 & n1776 ) | ( n1393 & ~n2191 ) | ( n1776 & ~n2191 ) ;
  assign n5754 = n3747 ^ n3664 ^ 1'b0 ;
  assign n5755 = n5754 ^ n2635 ^ n1460 ;
  assign n5756 = n5027 ^ n4007 ^ n1022 ;
  assign n5757 = ( n580 & ~n3200 ) | ( n580 & n5221 ) | ( ~n3200 & n5221 ) ;
  assign n5758 = n5757 ^ n3877 ^ n1690 ;
  assign n5759 = ( n296 & n1064 ) | ( n296 & n2111 ) | ( n1064 & n2111 ) ;
  assign n5760 = n5759 ^ n1639 ^ 1'b0 ;
  assign n5761 = ~n2679 & n5760 ;
  assign n5762 = n2819 ^ n654 ^ x104 ;
  assign n5763 = n3771 ^ x35 ^ 1'b0 ;
  assign n5764 = n1670 & ~n5763 ;
  assign n5765 = n5764 ^ n4136 ^ n3051 ;
  assign n5766 = n5765 ^ n2448 ^ 1'b0 ;
  assign n5767 = n2853 & n5766 ;
  assign n5768 = ~n1670 & n2552 ;
  assign n5769 = ( ~n2768 & n3466 ) | ( ~n2768 & n5768 ) | ( n3466 & n5768 ) ;
  assign n5770 = n713 | n3375 ;
  assign n5771 = n5770 ^ n5372 ^ 1'b0 ;
  assign n5772 = n2172 ^ n666 ^ 1'b0 ;
  assign n5775 = n3502 ^ n363 ^ x11 ;
  assign n5773 = ( ~n488 & n1581 ) | ( ~n488 & n2393 ) | ( n1581 & n2393 ) ;
  assign n5774 = n5329 & ~n5773 ;
  assign n5776 = n5775 ^ n5774 ^ 1'b0 ;
  assign n5777 = n665 | n5776 ;
  assign n5778 = n5772 & ~n5777 ;
  assign n5779 = n5544 ^ n5074 ^ n707 ;
  assign n5780 = ~n5588 & n5779 ;
  assign n5782 = ( x86 & n981 ) | ( x86 & n1328 ) | ( n981 & n1328 ) ;
  assign n5781 = ( n981 & n2402 ) | ( n981 & ~n5584 ) | ( n2402 & ~n5584 ) ;
  assign n5783 = n5782 ^ n5781 ^ n1691 ;
  assign n5784 = n5176 ^ n2077 ^ 1'b0 ;
  assign n5785 = n5783 | n5784 ;
  assign n5786 = n5785 ^ n2422 ^ x38 ;
  assign n5787 = x5 & ~n2967 ;
  assign n5788 = n5787 ^ n3026 ^ x41 ;
  assign n5789 = ( n1440 & n2506 ) | ( n1440 & n3731 ) | ( n2506 & n3731 ) ;
  assign n5790 = n3567 | n4653 ;
  assign n5791 = n5790 ^ n1516 ^ 1'b0 ;
  assign n5792 = n2664 & n3497 ;
  assign n5793 = n5791 & n5792 ;
  assign n5794 = n3261 & n4517 ;
  assign n5795 = n2148 & n5794 ;
  assign n5796 = n3339 ^ n1797 ^ 1'b0 ;
  assign n5797 = ~n2009 & n5796 ;
  assign n5798 = n3309 ^ n1887 ^ n1061 ;
  assign n5799 = n465 & n5798 ;
  assign n5800 = ( n1918 & ~n4554 ) | ( n1918 & n5799 ) | ( ~n4554 & n5799 ) ;
  assign n5801 = n5797 & ~n5800 ;
  assign n5802 = n5801 ^ n393 ^ 1'b0 ;
  assign n5803 = ~n337 & n5802 ;
  assign n5804 = n3340 ^ n2400 ^ x40 ;
  assign n5805 = n1476 | n1843 ;
  assign n5806 = x218 | n5805 ;
  assign n5807 = x205 & ~n4551 ;
  assign n5808 = ~n1625 & n5807 ;
  assign n5809 = ( n3566 & n5176 ) | ( n3566 & n5808 ) | ( n5176 & n5808 ) ;
  assign n5810 = ( n557 & n5806 ) | ( n557 & n5809 ) | ( n5806 & n5809 ) ;
  assign n5811 = n5804 | n5810 ;
  assign n5812 = n5803 | n5811 ;
  assign n5813 = ~n5795 & n5812 ;
  assign n5814 = n5813 ^ n1310 ^ 1'b0 ;
  assign n5815 = ( n690 & n2183 ) | ( n690 & n3718 ) | ( n2183 & n3718 ) ;
  assign n5816 = n4197 ^ n4084 ^ 1'b0 ;
  assign n5817 = ( n997 & n5815 ) | ( n997 & n5816 ) | ( n5815 & n5816 ) ;
  assign n5818 = ~n3056 & n3818 ;
  assign n5819 = n843 & ~n5818 ;
  assign n5820 = ~n5817 & n5819 ;
  assign n5825 = ( ~x29 & n545 ) | ( ~x29 & n1841 ) | ( n545 & n1841 ) ;
  assign n5821 = n1768 ^ n893 ^ 1'b0 ;
  assign n5822 = n1450 & n2356 ;
  assign n5823 = n5822 ^ n1749 ^ 1'b0 ;
  assign n5824 = ( ~x58 & n5821 ) | ( ~x58 & n5823 ) | ( n5821 & n5823 ) ;
  assign n5826 = n5825 ^ n5824 ^ 1'b0 ;
  assign n5827 = n5826 ^ n5609 ^ 1'b0 ;
  assign n5828 = ( n1188 & n3229 ) | ( n1188 & n4784 ) | ( n3229 & n4784 ) ;
  assign n5830 = n5671 ^ n3113 ^ n2497 ;
  assign n5831 = n5830 ^ n5420 ^ n1179 ;
  assign n5832 = n787 & ~n5831 ;
  assign n5829 = n2782 | n3983 ;
  assign n5833 = n5832 ^ n5829 ^ 1'b0 ;
  assign n5834 = n4359 ^ n1364 ^ 1'b0 ;
  assign n5835 = n4065 ^ n3025 ^ n1387 ;
  assign n5836 = ( n5215 & n5834 ) | ( n5215 & ~n5835 ) | ( n5834 & ~n5835 ) ;
  assign n5837 = n3897 ^ n3209 ^ x137 ;
  assign n5838 = n5837 ^ n4333 ^ 1'b0 ;
  assign n5839 = n5454 ^ n602 ^ 1'b0 ;
  assign n5840 = n3942 ^ n3369 ^ n331 ;
  assign n5841 = n1275 & ~n5840 ;
  assign n5842 = n5841 ^ n5244 ^ 1'b0 ;
  assign n5843 = n1235 & ~n5782 ;
  assign n5844 = n3364 & n5843 ;
  assign n5845 = n5844 ^ n3114 ^ n1792 ;
  assign n5846 = ( n1188 & n2996 ) | ( n1188 & n5845 ) | ( n2996 & n5845 ) ;
  assign n5847 = ~n546 & n2052 ;
  assign n5848 = n916 | n5847 ;
  assign n5849 = n4307 ^ n3431 ^ 1'b0 ;
  assign n5850 = n5848 & ~n5849 ;
  assign n5851 = n3144 & ~n5755 ;
  assign n5852 = n2076 ^ n381 ^ 1'b0 ;
  assign n5853 = ~n727 & n5852 ;
  assign n5854 = ( x220 & n2508 ) | ( x220 & ~n5853 ) | ( n2508 & ~n5853 ) ;
  assign n5855 = ( n3069 & n4470 ) | ( n3069 & n4670 ) | ( n4470 & n4670 ) ;
  assign n5856 = ( ~n4066 & n5854 ) | ( ~n4066 & n5855 ) | ( n5854 & n5855 ) ;
  assign n5859 = n2374 ^ n639 ^ 1'b0 ;
  assign n5860 = n3056 | n5859 ;
  assign n5861 = x217 & ~n3732 ;
  assign n5862 = n5860 & n5861 ;
  assign n5857 = ( n525 & ~n1669 ) | ( n525 & n3515 ) | ( ~n1669 & n3515 ) ;
  assign n5858 = ~n1839 & n5857 ;
  assign n5863 = n5862 ^ n5858 ^ 1'b0 ;
  assign n5864 = n5670 ^ n5252 ^ n1312 ;
  assign n5865 = ( ~n1056 & n5620 ) | ( ~n1056 & n5864 ) | ( n5620 & n5864 ) ;
  assign n5866 = n5670 ^ n1531 ^ 1'b0 ;
  assign n5867 = n5866 ^ n3681 ^ n2071 ;
  assign n5868 = n2701 ^ n671 ^ 1'b0 ;
  assign n5869 = n4649 ^ n707 ^ 1'b0 ;
  assign n5870 = n4085 ^ n1599 ^ 1'b0 ;
  assign n5871 = n5869 & n5870 ;
  assign n5872 = n868 & ~n2824 ;
  assign n5873 = ~n3147 & n5872 ;
  assign n5874 = n5873 ^ n3398 ^ n2080 ;
  assign n5875 = ~n1061 & n5874 ;
  assign n5876 = n5875 ^ n4257 ^ n650 ;
  assign n5877 = ~n1561 & n4093 ;
  assign n5878 = ~n2673 & n5877 ;
  assign n5879 = n995 & ~n2070 ;
  assign n5880 = n5879 ^ n3997 ^ 1'b0 ;
  assign n5881 = n4071 ^ n1438 ^ n639 ;
  assign n5882 = n1574 ^ n767 ^ n433 ;
  assign n5883 = ( n3818 & n4420 ) | ( n3818 & ~n5882 ) | ( n4420 & ~n5882 ) ;
  assign n5884 = ( n2084 & ~n5881 ) | ( n2084 & n5883 ) | ( ~n5881 & n5883 ) ;
  assign n5887 = n3365 & ~n5385 ;
  assign n5888 = n5887 ^ n2114 ^ 1'b0 ;
  assign n5885 = n3213 ^ n1400 ^ n657 ;
  assign n5886 = ( ~n1121 & n2410 ) | ( ~n1121 & n5885 ) | ( n2410 & n5885 ) ;
  assign n5889 = n5888 ^ n5886 ^ n3258 ;
  assign n5890 = n5889 ^ n1261 ^ n854 ;
  assign n5893 = n1156 ^ n748 ^ 1'b0 ;
  assign n5894 = x219 & n5893 ;
  assign n5895 = n5894 ^ n345 ^ x165 ;
  assign n5891 = n393 & n1196 ;
  assign n5892 = n3059 & n5891 ;
  assign n5896 = n5895 ^ n5892 ^ 1'b0 ;
  assign n5897 = ( n4142 & n5890 ) | ( n4142 & ~n5896 ) | ( n5890 & ~n5896 ) ;
  assign n5910 = n5329 ^ n4945 ^ 1'b0 ;
  assign n5911 = ( n4099 & ~n5205 ) | ( n4099 & n5910 ) | ( ~n5205 & n5910 ) ;
  assign n5898 = ~n642 & n3044 ;
  assign n5899 = n5898 ^ n1109 ^ 1'b0 ;
  assign n5900 = n4103 ^ n3753 ^ n2503 ;
  assign n5901 = n2655 | n4138 ;
  assign n5902 = ( x50 & n5900 ) | ( x50 & n5901 ) | ( n5900 & n5901 ) ;
  assign n5904 = n458 | n3397 ;
  assign n5905 = ( x236 & n733 ) | ( x236 & n2943 ) | ( n733 & n2943 ) ;
  assign n5906 = ( n1722 & ~n5904 ) | ( n1722 & n5905 ) | ( ~n5904 & n5905 ) ;
  assign n5907 = n5906 ^ n1861 ^ 1'b0 ;
  assign n5903 = ~n1210 & n3679 ;
  assign n5908 = n5907 ^ n5903 ^ n4012 ;
  assign n5909 = ( ~n5899 & n5902 ) | ( ~n5899 & n5908 ) | ( n5902 & n5908 ) ;
  assign n5912 = n5911 ^ n5909 ^ n2951 ;
  assign n5913 = ( n308 & n671 ) | ( n308 & n1030 ) | ( n671 & n1030 ) ;
  assign n5914 = ~n1388 & n5913 ;
  assign n5915 = n2814 ^ n2150 ^ 1'b0 ;
  assign n5916 = n1770 & ~n5915 ;
  assign n5917 = n1152 ^ x69 ^ 1'b0 ;
  assign n5918 = n5917 ^ n2840 ^ n799 ;
  assign n5919 = n5918 ^ n3067 ^ n476 ;
  assign n5920 = n5919 ^ n4705 ^ 1'b0 ;
  assign n5921 = n5916 & n5920 ;
  assign n5922 = n5914 & n5921 ;
  assign n5923 = n815 & n5922 ;
  assign n5924 = ( n1670 & n2844 ) | ( n1670 & n5386 ) | ( n2844 & n5386 ) ;
  assign n5925 = n1702 ^ n640 ^ 1'b0 ;
  assign n5926 = n5924 & ~n5925 ;
  assign n5927 = n2831 ^ n2436 ^ n1197 ;
  assign n5928 = n4023 ^ n606 ^ 1'b0 ;
  assign n5929 = ( x67 & n2455 ) | ( x67 & ~n2755 ) | ( n2455 & ~n2755 ) ;
  assign n5930 = n5929 ^ n5798 ^ n955 ;
  assign n5931 = n1771 | n5930 ;
  assign n5932 = x59 & n1625 ;
  assign n5933 = n5932 ^ n1673 ^ 1'b0 ;
  assign n5934 = n5933 ^ n5499 ^ n5363 ;
  assign n5935 = ~n2711 & n5934 ;
  assign n5937 = n3293 ^ n2237 ^ 1'b0 ;
  assign n5936 = n1786 & n2105 ;
  assign n5938 = n5937 ^ n5936 ^ 1'b0 ;
  assign n5939 = n5938 ^ n5126 ^ n3078 ;
  assign n5940 = n3696 | n5939 ;
  assign n5941 = n5940 ^ n2286 ^ 1'b0 ;
  assign n5942 = n2360 | n5116 ;
  assign n5943 = n4305 | n5942 ;
  assign n5944 = ( n2609 & n5941 ) | ( n2609 & ~n5943 ) | ( n5941 & ~n5943 ) ;
  assign n5945 = n5935 & n5944 ;
  assign n5946 = n2071 ^ n642 ^ 1'b0 ;
  assign n5947 = ( ~n1588 & n5667 ) | ( ~n1588 & n5946 ) | ( n5667 & n5946 ) ;
  assign n5948 = n4555 ^ n2945 ^ 1'b0 ;
  assign n5949 = n701 ^ x127 ^ x47 ;
  assign n5950 = n5949 ^ n4371 ^ n3229 ;
  assign n5951 = n5914 & n5950 ;
  assign n5952 = n5951 ^ n5091 ^ 1'b0 ;
  assign n5953 = ( n1172 & n1692 ) | ( n1172 & n4598 ) | ( n1692 & n4598 ) ;
  assign n5954 = n5953 ^ n3856 ^ n1854 ;
  assign n5955 = ( n3279 & n3645 ) | ( n3279 & ~n4950 ) | ( n3645 & ~n4950 ) ;
  assign n5959 = n310 & n1264 ;
  assign n5960 = n5527 & n5959 ;
  assign n5961 = n1012 & n5960 ;
  assign n5962 = ( ~n2165 & n5180 ) | ( ~n2165 & n5961 ) | ( n5180 & n5961 ) ;
  assign n5956 = ( x71 & n1883 ) | ( x71 & ~n5708 ) | ( n1883 & ~n5708 ) ;
  assign n5957 = ( n2615 & ~n3910 ) | ( n2615 & n5956 ) | ( ~n3910 & n5956 ) ;
  assign n5958 = n5957 ^ n3838 ^ 1'b0 ;
  assign n5963 = n5962 ^ n5958 ^ n2110 ;
  assign n5964 = x210 & n440 ;
  assign n5965 = ~n741 & n5964 ;
  assign n5966 = n5965 ^ n2896 ^ n1146 ;
  assign n5969 = n2024 | n3046 ;
  assign n5970 = n3005 | n5969 ;
  assign n5967 = ( n2506 & ~n3237 ) | ( n2506 & n5701 ) | ( ~n3237 & n5701 ) ;
  assign n5968 = ( ~n1190 & n2998 ) | ( ~n1190 & n5967 ) | ( n2998 & n5967 ) ;
  assign n5971 = n5970 ^ n5968 ^ 1'b0 ;
  assign n5972 = n4316 ^ n1863 ^ x30 ;
  assign n5973 = n5392 ^ n1738 ^ 1'b0 ;
  assign n5974 = n5973 ^ n5881 ^ 1'b0 ;
  assign n5975 = n5974 ^ n440 ^ 1'b0 ;
  assign n5976 = n5972 & ~n5975 ;
  assign n5977 = n3052 & ~n4626 ;
  assign n5978 = n5977 ^ n986 ^ 1'b0 ;
  assign n5979 = n5978 ^ n3726 ^ 1'b0 ;
  assign n5980 = n5208 ^ n4652 ^ 1'b0 ;
  assign n5982 = ~n257 & n1908 ;
  assign n5983 = n3762 & n5982 ;
  assign n5981 = ( ~n2562 & n2593 ) | ( ~n2562 & n3383 ) | ( n2593 & n3383 ) ;
  assign n5984 = n5983 ^ n5981 ^ 1'b0 ;
  assign n5988 = n1985 ^ n534 ^ 1'b0 ;
  assign n5989 = ~n2928 & n5988 ;
  assign n5990 = n5989 ^ n4038 ^ n2276 ;
  assign n5985 = n763 ^ n618 ^ 1'b0 ;
  assign n5986 = n895 & ~n5985 ;
  assign n5987 = ~x97 & n5986 ;
  assign n5991 = n5990 ^ n5987 ^ n4061 ;
  assign n5992 = ~x186 & n5991 ;
  assign n5993 = n4465 & ~n5992 ;
  assign n5994 = n5993 ^ n3444 ^ 1'b0 ;
  assign n5995 = n2777 ^ n929 ^ 1'b0 ;
  assign n5996 = n5102 ^ n2883 ^ n1419 ;
  assign n5997 = ( n3219 & n5995 ) | ( n3219 & n5996 ) | ( n5995 & n5996 ) ;
  assign n5998 = n5160 ^ n2134 ^ n394 ;
  assign n5999 = n3847 ^ n1225 ^ n311 ;
  assign n6000 = n2224 & ~n5999 ;
  assign n6001 = ( n3494 & ~n3629 ) | ( n3494 & n4240 ) | ( ~n3629 & n4240 ) ;
  assign n6002 = n5818 | n6001 ;
  assign n6003 = ( n1669 & n2634 ) | ( n1669 & n5276 ) | ( n2634 & n5276 ) ;
  assign n6004 = ( ~n1683 & n2228 ) | ( ~n1683 & n3545 ) | ( n2228 & n3545 ) ;
  assign n6005 = n6004 ^ n2335 ^ n559 ;
  assign n6006 = n3445 ^ n2824 ^ n816 ;
  assign n6007 = n6006 ^ n934 ^ n901 ;
  assign n6008 = n6005 & n6007 ;
  assign n6009 = n6008 ^ n1540 ^ 1'b0 ;
  assign n6010 = ( n1145 & n3840 ) | ( n1145 & n4840 ) | ( n3840 & n4840 ) ;
  assign n6011 = n6010 ^ n4874 ^ 1'b0 ;
  assign n6012 = n2456 | n6011 ;
  assign n6015 = ( n1485 & ~n1675 ) | ( n1485 & n2154 ) | ( ~n1675 & n2154 ) ;
  assign n6013 = ~n784 & n2737 ;
  assign n6014 = ~n3616 & n6013 ;
  assign n6016 = n6015 ^ n6014 ^ 1'b0 ;
  assign n6017 = n425 & n6016 ;
  assign n6018 = n6017 ^ n4774 ^ n443 ;
  assign n6019 = n4525 | n6018 ;
  assign n6020 = n6019 ^ n664 ^ 1'b0 ;
  assign n6021 = n3705 ^ n2445 ^ 1'b0 ;
  assign n6026 = ( n795 & ~n1914 ) | ( n795 & n3081 ) | ( ~n1914 & n3081 ) ;
  assign n6027 = n6026 ^ n4189 ^ n1041 ;
  assign n6023 = ( ~n2283 & n2732 ) | ( ~n2283 & n3684 ) | ( n2732 & n3684 ) ;
  assign n6024 = ( n1058 & n3385 ) | ( n1058 & ~n6023 ) | ( n3385 & ~n6023 ) ;
  assign n6025 = n895 & n6024 ;
  assign n6022 = n897 | n2736 ;
  assign n6028 = n6027 ^ n6025 ^ n6022 ;
  assign n6029 = ( n3058 & n6021 ) | ( n3058 & n6028 ) | ( n6021 & n6028 ) ;
  assign n6030 = n370 ^ n273 ^ 1'b0 ;
  assign n6032 = ( n974 & n1894 ) | ( n974 & ~n2069 ) | ( n1894 & ~n2069 ) ;
  assign n6033 = n6032 ^ n3677 ^ n3126 ;
  assign n6031 = n356 | n2172 ;
  assign n6034 = n6033 ^ n6031 ^ 1'b0 ;
  assign n6035 = n6030 & ~n6034 ;
  assign n6037 = n843 & n990 ;
  assign n6036 = n3737 ^ n1846 ^ 1'b0 ;
  assign n6038 = n6037 ^ n6036 ^ n1775 ;
  assign n6039 = n3840 | n6038 ;
  assign n6040 = n4688 ^ n4231 ^ n3774 ;
  assign n6041 = ( x25 & n633 ) | ( x25 & n6040 ) | ( n633 & n6040 ) ;
  assign n6042 = ~n2898 & n6041 ;
  assign n6043 = n400 & ~n877 ;
  assign n6044 = n6043 ^ n2490 ^ 1'b0 ;
  assign n6045 = n3804 ^ n1684 ^ n1067 ;
  assign n6046 = n6045 ^ n555 ^ 1'b0 ;
  assign n6047 = n6044 & n6046 ;
  assign n6048 = n6047 ^ n959 ^ 1'b0 ;
  assign n6049 = n748 & ~n2167 ;
  assign n6050 = x251 | n6049 ;
  assign n6051 = n6050 ^ n3681 ^ n1419 ;
  assign n6052 = n432 & n6051 ;
  assign n6053 = ( x155 & ~n3637 ) | ( x155 & n6052 ) | ( ~n3637 & n6052 ) ;
  assign n6054 = n5305 ^ n2192 ^ 1'b0 ;
  assign n6055 = n528 & n6054 ;
  assign n6056 = ( n4422 & n5200 ) | ( n4422 & n6055 ) | ( n5200 & n6055 ) ;
  assign n6057 = n5314 ^ n2798 ^ n1311 ;
  assign n6058 = ( ~n1380 & n3006 ) | ( ~n1380 & n3060 ) | ( n3006 & n3060 ) ;
  assign n6059 = ~n4495 & n6058 ;
  assign n6060 = n5419 & ~n6059 ;
  assign n6061 = ~n6057 & n6060 ;
  assign n6062 = ~n928 & n5005 ;
  assign n6063 = n711 & ~n6062 ;
  assign n6064 = n6063 ^ n3182 ^ 1'b0 ;
  assign n6065 = n2371 & n4522 ;
  assign n6066 = n6065 ^ n1662 ^ 1'b0 ;
  assign n6067 = ( n3122 & n6064 ) | ( n3122 & ~n6066 ) | ( n6064 & ~n6066 ) ;
  assign n6068 = n4371 ^ n2443 ^ x28 ;
  assign n6069 = n3234 & ~n6068 ;
  assign n6070 = ( n2347 & n2980 ) | ( n2347 & ~n6069 ) | ( n2980 & ~n6069 ) ;
  assign n6071 = ~n2143 & n4570 ;
  assign n6072 = n3081 & ~n5428 ;
  assign n6073 = n6071 & n6072 ;
  assign n6074 = n1645 & ~n3059 ;
  assign n6075 = n6074 ^ n3633 ^ n2464 ;
  assign n6076 = ( n564 & ~n3350 ) | ( n564 & n3736 ) | ( ~n3350 & n3736 ) ;
  assign n6077 = n6076 ^ n2025 ^ 1'b0 ;
  assign n6078 = ( x202 & n6075 ) | ( x202 & n6077 ) | ( n6075 & n6077 ) ;
  assign n6079 = n1699 & n2433 ;
  assign n6080 = n6079 ^ x130 ^ 1'b0 ;
  assign n6082 = ~n885 & n4519 ;
  assign n6083 = n6082 ^ x26 ^ 1'b0 ;
  assign n6081 = n1419 & ~n4960 ;
  assign n6084 = n6083 ^ n6081 ^ 1'b0 ;
  assign n6085 = ~n6080 & n6084 ;
  assign n6086 = n6085 ^ x29 ^ 1'b0 ;
  assign n6087 = n6086 ^ x199 ^ 1'b0 ;
  assign n6088 = n4840 & ~n6087 ;
  assign n6089 = n2367 | n4285 ;
  assign n6090 = n301 | n6089 ;
  assign n6091 = n1358 | n1864 ;
  assign n6092 = ( n2482 & n5933 ) | ( n2482 & n6091 ) | ( n5933 & n6091 ) ;
  assign n6093 = ~n1410 & n2254 ;
  assign n6094 = n6093 ^ n1892 ^ 1'b0 ;
  assign n6099 = ( n1972 & ~n2764 ) | ( n1972 & n3224 ) | ( ~n2764 & n3224 ) ;
  assign n6100 = ( ~n3826 & n4757 ) | ( ~n3826 & n6099 ) | ( n4757 & n6099 ) ;
  assign n6101 = n6100 ^ n5464 ^ n3847 ;
  assign n6095 = n5340 ^ n2863 ^ 1'b0 ;
  assign n6096 = n6095 ^ n313 ^ 1'b0 ;
  assign n6097 = n4634 ^ n2131 ^ 1'b0 ;
  assign n6098 = n6096 & ~n6097 ;
  assign n6102 = n6101 ^ n6098 ^ 1'b0 ;
  assign n6103 = ~n6094 & n6102 ;
  assign n6104 = ~x110 & x181 ;
  assign n6105 = ( x94 & n1863 ) | ( x94 & ~n6104 ) | ( n1863 & ~n6104 ) ;
  assign n6106 = n1438 ^ x208 ^ 1'b0 ;
  assign n6107 = ( n730 & n2676 ) | ( n730 & n6106 ) | ( n2676 & n6106 ) ;
  assign n6108 = n6105 & n6107 ;
  assign n6109 = n1671 & n6108 ;
  assign n6110 = ( n2562 & n3348 ) | ( n2562 & ~n6109 ) | ( n3348 & ~n6109 ) ;
  assign n6111 = ( n4138 & n5003 ) | ( n4138 & ~n5267 ) | ( n5003 & ~n5267 ) ;
  assign n6112 = n4759 ^ n4521 ^ 1'b0 ;
  assign n6113 = n6111 & ~n6112 ;
  assign n6114 = n6113 ^ n5346 ^ n5112 ;
  assign n6115 = ( ~n669 & n4766 ) | ( ~n669 & n6114 ) | ( n4766 & n6114 ) ;
  assign n6116 = ( n1354 & ~n2887 ) | ( n1354 & n4720 ) | ( ~n2887 & n4720 ) ;
  assign n6117 = n6116 ^ n4933 ^ n3319 ;
  assign n6118 = ~n3497 & n6117 ;
  assign n6119 = n5666 ^ n2417 ^ 1'b0 ;
  assign n6120 = ( n2939 & n5715 ) | ( n2939 & n6119 ) | ( n5715 & n6119 ) ;
  assign n6121 = ( ~n332 & n3645 ) | ( ~n332 & n6120 ) | ( n3645 & n6120 ) ;
  assign n6126 = n3103 ^ n370 ^ 1'b0 ;
  assign n6127 = n3216 & ~n6126 ;
  assign n6128 = n6127 ^ n3826 ^ 1'b0 ;
  assign n6129 = ~n2490 & n6128 ;
  assign n6122 = ( n1985 & n3287 ) | ( n1985 & ~n4960 ) | ( n3287 & ~n4960 ) ;
  assign n6123 = ~n5809 & n6122 ;
  assign n6124 = n3360 | n6123 ;
  assign n6125 = n1199 & ~n6124 ;
  assign n6130 = n6129 ^ n6125 ^ 1'b0 ;
  assign n6131 = ( n360 & n704 ) | ( n360 & n1856 ) | ( n704 & n1856 ) ;
  assign n6132 = n1622 ^ n899 ^ 1'b0 ;
  assign n6133 = n1236 & ~n6132 ;
  assign n6134 = n533 & n6133 ;
  assign n6135 = ~n1420 & n5321 ;
  assign n6136 = n3283 ^ n1518 ^ 1'b0 ;
  assign n6137 = n6136 ^ n1336 ^ 1'b0 ;
  assign n6138 = n1150 | n6137 ;
  assign n6139 = n6138 ^ n3741 ^ n1224 ;
  assign n6140 = ~n2353 & n6139 ;
  assign n6141 = ~n3432 & n6140 ;
  assign n6142 = x204 & ~n4086 ;
  assign n6143 = ~n3504 & n6142 ;
  assign n6151 = ( n803 & n1130 ) | ( n803 & n4367 ) | ( n1130 & n4367 ) ;
  assign n6144 = n2814 & n3323 ;
  assign n6145 = n2418 & n6144 ;
  assign n6146 = n2127 ^ n1851 ^ 1'b0 ;
  assign n6147 = n2168 ^ n682 ^ 1'b0 ;
  assign n6148 = n4046 ^ n1893 ^ x200 ;
  assign n6149 = ( n3171 & n6147 ) | ( n3171 & n6148 ) | ( n6147 & n6148 ) ;
  assign n6150 = ( n6145 & n6146 ) | ( n6145 & n6149 ) | ( n6146 & n6149 ) ;
  assign n6152 = n6151 ^ n6150 ^ 1'b0 ;
  assign n6153 = n2853 & n6152 ;
  assign n6154 = ~n1604 & n6153 ;
  assign n6155 = n6143 & n6154 ;
  assign n6156 = ( n6135 & n6141 ) | ( n6135 & ~n6155 ) | ( n6141 & ~n6155 ) ;
  assign n6157 = ( n563 & n1430 ) | ( n563 & ~n6015 ) | ( n1430 & ~n6015 ) ;
  assign n6158 = n4042 ^ n1886 ^ 1'b0 ;
  assign n6161 = n426 & n3190 ;
  assign n6159 = n5034 ^ n335 ^ 1'b0 ;
  assign n6160 = ( x74 & n2060 ) | ( x74 & ~n6159 ) | ( n2060 & ~n6159 ) ;
  assign n6162 = n6161 ^ n6160 ^ n1650 ;
  assign n6163 = n1592 & n3155 ;
  assign n6164 = ( n3214 & n6162 ) | ( n3214 & ~n6163 ) | ( n6162 & ~n6163 ) ;
  assign n6165 = n6158 & n6164 ;
  assign n6166 = n6165 ^ n6141 ^ 1'b0 ;
  assign n6167 = ( n1408 & n6157 ) | ( n1408 & ~n6166 ) | ( n6157 & ~n6166 ) ;
  assign n6168 = n3016 | n5186 ;
  assign n6169 = n5975 ^ n5125 ^ n4249 ;
  assign n6170 = n2174 ^ n1366 ^ x116 ;
  assign n6171 = n5778 & n6170 ;
  assign n6172 = ~n2881 & n4662 ;
  assign n6173 = n6172 ^ n1841 ^ 1'b0 ;
  assign n6174 = n1431 & n4328 ;
  assign n6175 = n1783 | n6174 ;
  assign n6176 = n6175 ^ n5094 ^ 1'b0 ;
  assign n6177 = ( x74 & x198 ) | ( x74 & n2340 ) | ( x198 & n2340 ) ;
  assign n6178 = n6177 ^ n2200 ^ n301 ;
  assign n6179 = ( n1163 & n1749 ) | ( n1163 & n6178 ) | ( n1749 & n6178 ) ;
  assign n6180 = ~n2482 & n3273 ;
  assign n6181 = ( n1627 & n5197 ) | ( n1627 & ~n6180 ) | ( n5197 & ~n6180 ) ;
  assign n6182 = n3956 & n6181 ;
  assign n6183 = ( n293 & n565 ) | ( n293 & n1703 ) | ( n565 & n1703 ) ;
  assign n6184 = ( x219 & ~n6136 ) | ( x219 & n6183 ) | ( ~n6136 & n6183 ) ;
  assign n6185 = n4428 ^ n2635 ^ n604 ;
  assign n6186 = ( ~n1792 & n6184 ) | ( ~n1792 & n6185 ) | ( n6184 & n6185 ) ;
  assign n6188 = n2824 ^ n1714 ^ 1'b0 ;
  assign n6187 = ( ~x62 & n3409 ) | ( ~x62 & n3415 ) | ( n3409 & n3415 ) ;
  assign n6189 = n6188 ^ n6187 ^ n5099 ;
  assign n6190 = ~n1072 & n2045 ;
  assign n6191 = n6037 ^ n2104 ^ 1'b0 ;
  assign n6192 = n6190 & ~n6191 ;
  assign n6193 = n6049 ^ n5373 ^ x130 ;
  assign n6197 = ( n1325 & n2192 ) | ( n1325 & ~n3847 ) | ( n2192 & ~n3847 ) ;
  assign n6196 = n1506 ^ n940 ^ n759 ;
  assign n6194 = n2319 & n3018 ;
  assign n6195 = n6194 ^ n1862 ^ 1'b0 ;
  assign n6198 = n6197 ^ n6196 ^ n6195 ;
  assign n6199 = ~n6193 & n6198 ;
  assign n6200 = n1208 & n6199 ;
  assign n6201 = n3322 ^ n380 ^ 1'b0 ;
  assign n6202 = ( n1671 & ~n4217 ) | ( n1671 & n5824 ) | ( ~n4217 & n5824 ) ;
  assign n6212 = x179 & n3201 ;
  assign n6213 = n6212 ^ n286 ^ 1'b0 ;
  assign n6209 = n3094 ^ n2330 ^ x171 ;
  assign n6210 = n6209 ^ n271 ^ 1'b0 ;
  assign n6211 = n3134 & n6210 ;
  assign n6214 = n6213 ^ n6211 ^ n2293 ;
  assign n6208 = n4530 ^ n2244 ^ 1'b0 ;
  assign n6215 = n6214 ^ n6208 ^ 1'b0 ;
  assign n6207 = ( n1320 & n1724 ) | ( n1320 & ~n5093 ) | ( n1724 & ~n5093 ) ;
  assign n6203 = n1362 | n2859 ;
  assign n6204 = n6203 ^ n6044 ^ n1970 ;
  assign n6205 = n2052 & n6204 ;
  assign n6206 = n6205 ^ n663 ^ 1'b0 ;
  assign n6216 = n6215 ^ n6207 ^ n6206 ;
  assign n6217 = n6216 ^ n2558 ^ 1'b0 ;
  assign n6218 = ~n4150 & n6217 ;
  assign n6219 = n5553 ^ n5316 ^ n3502 ;
  assign n6220 = n1040 & ~n3203 ;
  assign n6221 = n1806 & n5071 ;
  assign n6222 = n4786 & n6221 ;
  assign n6223 = n2250 ^ n1753 ^ n595 ;
  assign n6224 = n2970 & n6223 ;
  assign n6225 = ~n3908 & n6004 ;
  assign n6226 = n6225 ^ n3844 ^ 1'b0 ;
  assign n6227 = ( n1790 & ~n2104 ) | ( n1790 & n4462 ) | ( ~n2104 & n4462 ) ;
  assign n6228 = n822 | n6227 ;
  assign n6229 = n6228 ^ n5212 ^ 1'b0 ;
  assign n6230 = n4700 ^ n2240 ^ x217 ;
  assign n6231 = ~n596 & n2260 ;
  assign n6232 = ~n755 & n6231 ;
  assign n6233 = n6149 & ~n6232 ;
  assign n6234 = ( n3394 & n5686 ) | ( n3394 & n5976 ) | ( n5686 & n5976 ) ;
  assign n6237 = ~x129 & n1331 ;
  assign n6235 = n2706 ^ n2302 ^ n1891 ;
  assign n6236 = ~n1659 & n6235 ;
  assign n6238 = n6237 ^ n6236 ^ n3972 ;
  assign n6239 = n2672 ^ x143 ^ 1'b0 ;
  assign n6240 = ( ~n3768 & n4680 ) | ( ~n3768 & n6239 ) | ( n4680 & n6239 ) ;
  assign n6241 = ( n4237 & n5106 ) | ( n4237 & ~n6240 ) | ( n5106 & ~n6240 ) ;
  assign n6242 = ~n618 & n785 ;
  assign n6243 = n1323 & ~n6242 ;
  assign n6244 = ~n2296 & n6243 ;
  assign n6245 = ( n1461 & ~n3762 ) | ( n1461 & n6244 ) | ( ~n3762 & n6244 ) ;
  assign n6246 = ~n4291 & n6245 ;
  assign n6247 = ( ~x60 & n5363 ) | ( ~x60 & n6246 ) | ( n5363 & n6246 ) ;
  assign n6248 = n1725 ^ x34 ^ 1'b0 ;
  assign n6249 = n1545 | n6248 ;
  assign n6250 = n6006 ^ n4439 ^ n2020 ;
  assign n6251 = n6250 ^ n3561 ^ n2311 ;
  assign n6252 = n3255 & n6251 ;
  assign n6253 = n6249 & n6252 ;
  assign n6254 = n1186 & ~n4542 ;
  assign n6255 = n6254 ^ n4638 ^ 1'b0 ;
  assign n6256 = ( n3927 & ~n6118 ) | ( n3927 & n6255 ) | ( ~n6118 & n6255 ) ;
  assign n6257 = ( ~n286 & n917 ) | ( ~n286 & n2213 ) | ( n917 & n2213 ) ;
  assign n6258 = n6251 ^ n1709 ^ 1'b0 ;
  assign n6259 = ~n6257 & n6258 ;
  assign n6260 = n6259 ^ n4576 ^ n1623 ;
  assign n6261 = n3348 | n4885 ;
  assign n6262 = n5183 ^ n3051 ^ 1'b0 ;
  assign n6263 = n2887 | n6262 ;
  assign n6264 = n2354 ^ n2315 ^ 1'b0 ;
  assign n6265 = n4618 | n6264 ;
  assign n6266 = n6265 ^ n2265 ^ 1'b0 ;
  assign n6267 = n6263 & ~n6266 ;
  assign n6268 = n1404 ^ n279 ^ 1'b0 ;
  assign n6269 = n6268 ^ n4606 ^ 1'b0 ;
  assign n6270 = ( n3580 & n4905 ) | ( n3580 & n6269 ) | ( n4905 & n6269 ) ;
  assign n6271 = x192 & ~n6270 ;
  assign n6272 = n6267 & n6271 ;
  assign n6273 = ~n4070 & n6032 ;
  assign n6274 = ( n542 & n3147 ) | ( n542 & ~n6273 ) | ( n3147 & ~n6273 ) ;
  assign n6275 = ( x9 & n2064 ) | ( x9 & n2265 ) | ( n2064 & n2265 ) ;
  assign n6276 = n6275 ^ x186 ^ 1'b0 ;
  assign n6277 = x2 & n6276 ;
  assign n6278 = n1942 ^ n870 ^ 1'b0 ;
  assign n6279 = n6277 & n6278 ;
  assign n6280 = n599 & n6279 ;
  assign n6281 = ~n6274 & n6280 ;
  assign n6282 = n5933 ^ n4989 ^ n3349 ;
  assign n6283 = n4068 | n4706 ;
  assign n6284 = n2853 ^ n2327 ^ 1'b0 ;
  assign n6285 = n2104 & ~n6284 ;
  assign n6287 = n1592 ^ n505 ^ n480 ;
  assign n6286 = ( x202 & n745 ) | ( x202 & n1155 ) | ( n745 & n1155 ) ;
  assign n6288 = n6287 ^ n6286 ^ 1'b0 ;
  assign n6289 = n868 & ~n6288 ;
  assign n6290 = n6289 ^ n3267 ^ 1'b0 ;
  assign n6291 = n4844 & ~n6290 ;
  assign n6292 = ( n751 & n3029 ) | ( n751 & ~n6291 ) | ( n3029 & ~n6291 ) ;
  assign n6293 = n5539 ^ n572 ^ x156 ;
  assign n6296 = n1331 & n5049 ;
  assign n6297 = n6296 ^ n2800 ^ 1'b0 ;
  assign n6294 = n4650 ^ n3701 ^ 1'b0 ;
  assign n6295 = x234 & ~n6294 ;
  assign n6298 = n6297 ^ n6295 ^ 1'b0 ;
  assign n6299 = ( x145 & n6293 ) | ( x145 & n6298 ) | ( n6293 & n6298 ) ;
  assign n6302 = n4892 ^ n2567 ^ n1587 ;
  assign n6303 = n6302 ^ x14 ^ 1'b0 ;
  assign n6304 = n498 & ~n6303 ;
  assign n6300 = n1718 | n4498 ;
  assign n6301 = n6300 ^ n5288 ^ n3113 ;
  assign n6305 = n6304 ^ n6301 ^ n4139 ;
  assign n6307 = n4350 & ~n4640 ;
  assign n6306 = n474 & ~n2396 ;
  assign n6308 = n6307 ^ n6306 ^ 1'b0 ;
  assign n6309 = x152 & ~n5088 ;
  assign n6310 = n6309 ^ n4687 ^ 1'b0 ;
  assign n6311 = n5133 ^ n4691 ^ n3779 ;
  assign n6312 = n3008 ^ n2042 ^ 1'b0 ;
  assign n6313 = n1966 & n2557 ;
  assign n6314 = n1943 & ~n3241 ;
  assign n6315 = n1722 & ~n6314 ;
  assign n6316 = n3801 ^ n462 ^ 1'b0 ;
  assign n6317 = n362 | n6316 ;
  assign n6318 = ( n1315 & n1755 ) | ( n1315 & n6317 ) | ( n1755 & n6317 ) ;
  assign n6319 = n1139 ^ n831 ^ n506 ;
  assign n6320 = ( n1725 & n2635 ) | ( n1725 & ~n6319 ) | ( n2635 & ~n6319 ) ;
  assign n6321 = ~n516 & n5775 ;
  assign n6322 = ~n6320 & n6321 ;
  assign n6323 = n1916 ^ n1816 ^ 1'b0 ;
  assign n6324 = n1716 ^ n1249 ^ n959 ;
  assign n6325 = ( ~n5499 & n6323 ) | ( ~n5499 & n6324 ) | ( n6323 & n6324 ) ;
  assign n6326 = n3480 ^ n3363 ^ x108 ;
  assign n6327 = n2406 & ~n5727 ;
  assign n6328 = ( n4084 & n6326 ) | ( n4084 & ~n6327 ) | ( n6326 & ~n6327 ) ;
  assign n6329 = ( n775 & n883 ) | ( n775 & n2608 ) | ( n883 & n2608 ) ;
  assign n6330 = n1131 & ~n1145 ;
  assign n6331 = n885 & n6330 ;
  assign n6332 = ~n6329 & n6331 ;
  assign n6333 = ( n1614 & n2217 ) | ( n1614 & ~n2642 ) | ( n2217 & ~n2642 ) ;
  assign n6334 = ( x41 & n1184 ) | ( x41 & n6333 ) | ( n1184 & n6333 ) ;
  assign n6335 = n1542 & ~n6334 ;
  assign n6336 = n5490 & n6335 ;
  assign n6338 = x150 & n1516 ;
  assign n6337 = ( n1489 & n1794 ) | ( n1489 & ~n2373 ) | ( n1794 & ~n2373 ) ;
  assign n6339 = n6338 ^ n6337 ^ n4987 ;
  assign n6340 = n1592 | n3503 ;
  assign n6341 = n6340 ^ n1373 ^ 1'b0 ;
  assign n6342 = n4937 ^ n2502 ^ n1054 ;
  assign n6343 = n2256 | n6342 ;
  assign n6344 = n6341 & ~n6343 ;
  assign n6345 = n5913 ^ n2850 ^ 1'b0 ;
  assign n6346 = n3718 | n5701 ;
  assign n6347 = n6346 ^ n2750 ^ 1'b0 ;
  assign n6348 = n615 | n6347 ;
  assign n6349 = n6348 ^ n4079 ^ n1779 ;
  assign n6350 = ( ~n4876 & n6345 ) | ( ~n4876 & n6349 ) | ( n6345 & n6349 ) ;
  assign n6351 = ( x5 & n431 ) | ( x5 & ~n633 ) | ( n431 & ~n633 ) ;
  assign n6352 = n6351 ^ x193 ^ 1'b0 ;
  assign n6353 = n2926 & ~n6352 ;
  assign n6354 = ( n3078 & ~n4569 ) | ( n3078 & n6353 ) | ( ~n4569 & n6353 ) ;
  assign n6355 = n3952 ^ n849 ^ 1'b0 ;
  assign n6356 = ( n2266 & n6354 ) | ( n2266 & n6355 ) | ( n6354 & n6355 ) ;
  assign n6357 = n4582 ^ n2777 ^ n341 ;
  assign n6358 = n1169 | n6357 ;
  assign n6359 = n6358 ^ n3185 ^ 1'b0 ;
  assign n6360 = ( x44 & ~n634 ) | ( x44 & n981 ) | ( ~n634 & n981 ) ;
  assign n6361 = ~n957 & n6360 ;
  assign n6362 = n6361 ^ n5549 ^ 1'b0 ;
  assign n6364 = n2905 ^ n2090 ^ n349 ;
  assign n6365 = n6364 ^ n5050 ^ n706 ;
  assign n6363 = n540 & ~n1916 ;
  assign n6366 = n6365 ^ n6363 ^ 1'b0 ;
  assign n6367 = n1162 | n3285 ;
  assign n6368 = ( n6362 & n6366 ) | ( n6362 & ~n6367 ) | ( n6366 & ~n6367 ) ;
  assign n6369 = ( n351 & n2271 ) | ( n351 & ~n3878 ) | ( n2271 & ~n3878 ) ;
  assign n6370 = n3796 & n6369 ;
  assign n6371 = x60 & ~n6370 ;
  assign n6372 = ~n6319 & n6371 ;
  assign n6373 = n1904 ^ x113 ^ 1'b0 ;
  assign n6374 = n1515 & n6373 ;
  assign n6375 = n6374 ^ n4389 ^ 1'b0 ;
  assign n6376 = n3095 & ~n6375 ;
  assign n6377 = ~n2886 & n6376 ;
  assign n6378 = ~n946 & n6377 ;
  assign n6379 = ~n986 & n2749 ;
  assign n6380 = ~n2259 & n6379 ;
  assign n6381 = ~n1262 & n6380 ;
  assign n6382 = ( n2552 & n4118 ) | ( n2552 & n5281 ) | ( n4118 & n5281 ) ;
  assign n6383 = n932 & ~n2524 ;
  assign n6384 = n6383 ^ n1561 ^ 1'b0 ;
  assign n6385 = n3707 & ~n6384 ;
  assign n6386 = x186 & ~n2053 ;
  assign n6387 = ( ~n6382 & n6385 ) | ( ~n6382 & n6386 ) | ( n6385 & n6386 ) ;
  assign n6388 = n3209 ^ n2324 ^ n1037 ;
  assign n6389 = n6388 ^ n5836 ^ 1'b0 ;
  assign n6390 = n3398 ^ n483 ^ x48 ;
  assign n6391 = n6390 ^ n3184 ^ n3111 ;
  assign n6392 = n6391 ^ n4224 ^ n1643 ;
  assign n6394 = ~n2791 & n4144 ;
  assign n6395 = ~n2697 & n6394 ;
  assign n6393 = n3330 ^ n3166 ^ n304 ;
  assign n6396 = n6395 ^ n6393 ^ x91 ;
  assign n6403 = n5351 ^ n4086 ^ n3148 ;
  assign n6399 = ( ~n1133 & n1995 ) | ( ~n1133 & n3555 ) | ( n1995 & n3555 ) ;
  assign n6400 = n6399 ^ x213 ^ x104 ;
  assign n6397 = ~n315 & n2587 ;
  assign n6398 = ~x21 & n6397 ;
  assign n6401 = n6400 ^ n6398 ^ n5948 ;
  assign n6402 = n403 & n6401 ;
  assign n6404 = n6403 ^ n6402 ^ 1'b0 ;
  assign n6405 = ~n910 & n4488 ;
  assign n6406 = n4904 & n6405 ;
  assign n6407 = n1831 ^ x206 ^ 1'b0 ;
  assign n6408 = ( n675 & ~n1761 ) | ( n675 & n6407 ) | ( ~n1761 & n6407 ) ;
  assign n6411 = n4191 ^ n2705 ^ n2034 ;
  assign n6409 = n974 | n4974 ;
  assign n6410 = n4797 | n6409 ;
  assign n6412 = n6411 ^ n6410 ^ n587 ;
  assign n6413 = n6408 | n6412 ;
  assign n6416 = n5195 ^ n4272 ^ n2859 ;
  assign n6414 = ( x203 & n1478 ) | ( x203 & n3902 ) | ( n1478 & n3902 ) ;
  assign n6415 = ~n1924 & n6414 ;
  assign n6417 = n6416 ^ n6415 ^ 1'b0 ;
  assign n6418 = n5613 ^ n4580 ^ 1'b0 ;
  assign n6419 = ~n2949 & n4510 ;
  assign n6420 = n6419 ^ n6000 ^ 1'b0 ;
  assign n6423 = ( ~n1664 & n4071 ) | ( ~n1664 & n4473 ) | ( n4071 & n4473 ) ;
  assign n6421 = n394 & ~n6074 ;
  assign n6422 = n6421 ^ n4530 ^ n4209 ;
  assign n6424 = n6423 ^ n6422 ^ n2039 ;
  assign n6425 = ( ~n2298 & n2397 ) | ( ~n2298 & n4875 ) | ( n2397 & n4875 ) ;
  assign n6426 = n1036 & ~n2348 ;
  assign n6427 = n6425 & n6426 ;
  assign n6428 = n3374 & ~n6214 ;
  assign n6431 = ( n1794 & ~n1826 ) | ( n1794 & n2649 ) | ( ~n1826 & n2649 ) ;
  assign n6429 = n2528 & ~n4216 ;
  assign n6430 = n6429 ^ n2729 ^ 1'b0 ;
  assign n6432 = n6431 ^ n6430 ^ n1818 ;
  assign n6433 = n6432 ^ n3138 ^ 1'b0 ;
  assign n6434 = n1108 ^ x171 ^ 1'b0 ;
  assign n6435 = ( x217 & n2215 ) | ( x217 & ~n6434 ) | ( n2215 & ~n6434 ) ;
  assign n6436 = n2467 ^ n1884 ^ 1'b0 ;
  assign n6437 = n458 | n6436 ;
  assign n6438 = n6435 & ~n6437 ;
  assign n6439 = n6438 ^ n4582 ^ 1'b0 ;
  assign n6440 = n3152 & n4814 ;
  assign n6441 = n2114 | n2794 ;
  assign n6442 = n3569 & ~n6441 ;
  assign n6443 = ~n5401 & n6442 ;
  assign n6444 = n6235 ^ n1010 ^ 1'b0 ;
  assign n6445 = ( n929 & n3087 ) | ( n929 & ~n6444 ) | ( n3087 & ~n6444 ) ;
  assign n6454 = n360 ^ x157 ^ 1'b0 ;
  assign n6455 = ~n456 & n6454 ;
  assign n6446 = n3094 ^ n2248 ^ 1'b0 ;
  assign n6447 = ~n2020 & n6446 ;
  assign n6448 = n6447 ^ n693 ^ 1'b0 ;
  assign n6449 = n6448 ^ n5991 ^ n3705 ;
  assign n6450 = n6449 ^ n4892 ^ n4087 ;
  assign n6451 = ( n4769 & ~n5072 ) | ( n4769 & n6450 ) | ( ~n5072 & n6450 ) ;
  assign n6452 = ( n3310 & n3538 ) | ( n3310 & ~n6451 ) | ( n3538 & ~n6451 ) ;
  assign n6453 = n1582 & ~n6452 ;
  assign n6456 = n6455 ^ n6453 ^ 1'b0 ;
  assign n6457 = ( n1617 & ~n2816 ) | ( n1617 & n5093 ) | ( ~n2816 & n5093 ) ;
  assign n6458 = n6457 ^ n1034 ^ 1'b0 ;
  assign n6459 = n6458 ^ n5392 ^ n1251 ;
  assign n6460 = ( n1309 & n1545 ) | ( n1309 & n6459 ) | ( n1545 & n6459 ) ;
  assign n6461 = n3798 & n6460 ;
  assign n6462 = n6461 ^ n2054 ^ 1'b0 ;
  assign n6475 = n260 & ~n1524 ;
  assign n6476 = n6475 ^ n1306 ^ 1'b0 ;
  assign n6477 = ( ~n1786 & n1995 ) | ( ~n1786 & n6476 ) | ( n1995 & n6476 ) ;
  assign n6473 = n358 | n3310 ;
  assign n6474 = n6473 ^ n1367 ^ 1'b0 ;
  assign n6478 = n6477 ^ n6474 ^ n2077 ;
  assign n6471 = ( n499 & n712 ) | ( n499 & ~n4129 ) | ( n712 & ~n4129 ) ;
  assign n6463 = ~n1005 & n2425 ;
  assign n6464 = n4807 ^ n3285 ^ n933 ;
  assign n6465 = n6464 ^ n2422 ^ 1'b0 ;
  assign n6466 = n6463 & ~n6465 ;
  assign n6467 = n4812 ^ n363 ^ 1'b0 ;
  assign n6468 = n6466 & ~n6467 ;
  assign n6469 = n6468 ^ n5617 ^ n2620 ;
  assign n6470 = n6289 & ~n6469 ;
  assign n6472 = n6471 ^ n6470 ^ 1'b0 ;
  assign n6479 = n6478 ^ n6472 ^ n529 ;
  assign n6480 = n2856 & n6479 ;
  assign n6481 = n5248 ^ n4788 ^ 1'b0 ;
  assign n6482 = n2733 & ~n6310 ;
  assign n6483 = ( x137 & n1266 ) | ( x137 & ~n2261 ) | ( n1266 & ~n2261 ) ;
  assign n6484 = ( ~n995 & n3654 ) | ( ~n995 & n6483 ) | ( n3654 & n6483 ) ;
  assign n6485 = ( n1225 & n3963 ) | ( n1225 & ~n6484 ) | ( n3963 & ~n6484 ) ;
  assign n6486 = n6485 ^ n3833 ^ n2155 ;
  assign n6488 = n2828 ^ n2273 ^ n1510 ;
  assign n6489 = ( ~n1998 & n2903 ) | ( ~n1998 & n6488 ) | ( n2903 & n6488 ) ;
  assign n6487 = n2217 & n2283 ;
  assign n6490 = n6489 ^ n6487 ^ 1'b0 ;
  assign n6491 = n6042 ^ n1776 ^ n1068 ;
  assign n6494 = n6423 ^ n3330 ^ n1320 ;
  assign n6495 = n2501 ^ n1275 ^ x158 ;
  assign n6496 = ~n6450 & n6495 ;
  assign n6497 = ( n658 & n6494 ) | ( n658 & ~n6496 ) | ( n6494 & ~n6496 ) ;
  assign n6492 = ( x78 & n1412 ) | ( x78 & ~n5146 ) | ( n1412 & ~n5146 ) ;
  assign n6493 = ( n4471 & ~n5799 ) | ( n4471 & n6492 ) | ( ~n5799 & n6492 ) ;
  assign n6498 = n6497 ^ n6493 ^ n4960 ;
  assign n6499 = ( x169 & n3475 ) | ( x169 & ~n6279 ) | ( n3475 & ~n6279 ) ;
  assign n6500 = n5397 ^ n933 ^ n554 ;
  assign n6501 = ( n2831 & n3213 ) | ( n2831 & n6500 ) | ( n3213 & n6500 ) ;
  assign n6502 = n6501 ^ n5330 ^ 1'b0 ;
  assign n6503 = ~n570 & n4522 ;
  assign n6504 = n6503 ^ n5278 ^ 1'b0 ;
  assign n6515 = ( n1160 & n3839 ) | ( n1160 & n5294 ) | ( n3839 & n5294 ) ;
  assign n6510 = ~n2681 & n2874 ;
  assign n6508 = ~n1634 & n4065 ;
  assign n6509 = n6508 ^ n819 ^ 1'b0 ;
  assign n6511 = n6510 ^ n6509 ^ n4373 ;
  assign n6512 = n6511 ^ n1401 ^ x61 ;
  assign n6505 = n2167 ^ n1138 ^ n508 ;
  assign n6506 = n4204 & n6505 ;
  assign n6507 = n4516 & n6506 ;
  assign n6513 = n6512 ^ n6507 ^ 1'b0 ;
  assign n6514 = ~n870 & n6513 ;
  assign n6516 = n6515 ^ n6514 ^ n5458 ;
  assign n6517 = n5906 ^ n2770 ^ n744 ;
  assign n6518 = n3484 ^ n698 ^ 1'b0 ;
  assign n6519 = ~n2346 & n6518 ;
  assign n6520 = ~n598 & n6519 ;
  assign n6521 = ( x128 & n6434 ) | ( x128 & ~n6520 ) | ( n6434 & ~n6520 ) ;
  assign n6522 = n2292 ^ n2160 ^ 1'b0 ;
  assign n6523 = n6145 ^ n569 ^ 1'b0 ;
  assign n6524 = n6523 ^ n5557 ^ 1'b0 ;
  assign n6525 = ~n3972 & n6524 ;
  assign n6528 = n1646 & n2182 ;
  assign n6526 = x185 & n4375 ;
  assign n6527 = ( n3760 & n3864 ) | ( n3760 & ~n6526 ) | ( n3864 & ~n6526 ) ;
  assign n6529 = n6528 ^ n6527 ^ n1945 ;
  assign n6530 = n922 ^ x100 ^ 1'b0 ;
  assign n6531 = n4333 | n6530 ;
  assign n6532 = ( n1363 & n3813 ) | ( n1363 & n6531 ) | ( n3813 & n6531 ) ;
  assign n6533 = ~n1180 & n3394 ;
  assign n6534 = ~n6532 & n6533 ;
  assign n6535 = n6534 ^ n4471 ^ 1'b0 ;
  assign n6536 = n6529 | n6535 ;
  assign n6537 = n4807 ^ n1945 ^ 1'b0 ;
  assign n6538 = n6537 ^ n3721 ^ 1'b0 ;
  assign n6539 = ~n6536 & n6538 ;
  assign n6540 = n4767 ^ n3059 ^ n1428 ;
  assign n6541 = n6540 ^ n5701 ^ n2230 ;
  assign n6542 = n6541 ^ n3767 ^ 1'b0 ;
  assign n6543 = n2206 & n6542 ;
  assign n6545 = n3181 ^ n1150 ^ 1'b0 ;
  assign n6546 = x208 & ~n6545 ;
  assign n6547 = n610 | n3076 ;
  assign n6548 = n6547 ^ n2912 ^ 1'b0 ;
  assign n6549 = ( x161 & n6546 ) | ( x161 & n6548 ) | ( n6546 & n6548 ) ;
  assign n6544 = n5086 ^ n4516 ^ n643 ;
  assign n6550 = n6549 ^ n6544 ^ n3271 ;
  assign n6551 = ~n753 & n1599 ;
  assign n6552 = n6550 | n6551 ;
  assign n6553 = n5183 | n6552 ;
  assign n6554 = ~n4298 & n5757 ;
  assign n6555 = n6485 ^ n5718 ^ n5042 ;
  assign n6556 = n6555 ^ n3279 ^ 1'b0 ;
  assign n6557 = n6554 | n6556 ;
  assign n6559 = n2419 ^ n2367 ^ 1'b0 ;
  assign n6560 = n6559 ^ n2676 ^ 1'b0 ;
  assign n6558 = n4043 ^ x143 ^ 1'b0 ;
  assign n6561 = n6560 ^ n6558 ^ n3567 ;
  assign n6562 = n2943 ^ n2417 ^ n1468 ;
  assign n6563 = ( n1072 & n3264 ) | ( n1072 & ~n6562 ) | ( n3264 & ~n6562 ) ;
  assign n6564 = n3090 & n3813 ;
  assign n6565 = ( ~n4518 & n5713 ) | ( ~n4518 & n6564 ) | ( n5713 & n6564 ) ;
  assign n6566 = ( n3057 & n6563 ) | ( n3057 & ~n6565 ) | ( n6563 & ~n6565 ) ;
  assign n6567 = n5808 ^ n3878 ^ n874 ;
  assign n6568 = ~n557 & n6567 ;
  assign n6569 = ~n4761 & n6568 ;
  assign n6575 = ~x220 & n4888 ;
  assign n6576 = n6468 ^ n1743 ^ 1'b0 ;
  assign n6577 = n6575 & n6576 ;
  assign n6572 = ~n1387 & n1840 ;
  assign n6573 = n6572 ^ n458 ^ 1'b0 ;
  assign n6571 = x68 & ~n3034 ;
  assign n6574 = n6573 ^ n6571 ^ 1'b0 ;
  assign n6570 = ~n698 & n1831 ;
  assign n6578 = n6577 ^ n6574 ^ n6570 ;
  assign n6579 = ( n2891 & ~n4636 ) | ( n2891 & n4776 ) | ( ~n4636 & n4776 ) ;
  assign n6581 = n890 | n3122 ;
  assign n6582 = ( n2210 & ~n5542 ) | ( n2210 & n6581 ) | ( ~n5542 & n6581 ) ;
  assign n6583 = n2822 ^ x189 ^ 1'b0 ;
  assign n6584 = n6583 ^ n2633 ^ 1'b0 ;
  assign n6585 = n6582 & ~n6584 ;
  assign n6580 = n3706 | n6208 ;
  assign n6586 = n6585 ^ n6580 ^ 1'b0 ;
  assign n6587 = n3273 & ~n6586 ;
  assign n6588 = n387 & ~n2091 ;
  assign n6589 = n6588 ^ n4761 ^ 1'b0 ;
  assign n6599 = ~n326 & n4312 ;
  assign n6600 = ( n401 & ~n1301 ) | ( n401 & n6599 ) | ( ~n1301 & n6599 ) ;
  assign n6590 = ( ~n1139 & n1858 ) | ( ~n1139 & n2595 ) | ( n1858 & n2595 ) ;
  assign n6591 = n4489 ^ n3586 ^ x103 ;
  assign n6592 = ( ~n3226 & n6590 ) | ( ~n3226 & n6591 ) | ( n6590 & n6591 ) ;
  assign n6593 = n1014 & ~n6177 ;
  assign n6594 = n6593 ^ n5500 ^ n4161 ;
  assign n6595 = n2182 & n6594 ;
  assign n6596 = ~n6592 & n6595 ;
  assign n6597 = n1798 & ~n6596 ;
  assign n6598 = n6597 ^ n4599 ^ 1'b0 ;
  assign n6601 = n6600 ^ n6598 ^ 1'b0 ;
  assign n6602 = n6589 & ~n6601 ;
  assign n6603 = n3803 ^ n2562 ^ 1'b0 ;
  assign n6604 = n3476 & n6603 ;
  assign n6605 = n6604 ^ n1864 ^ 1'b0 ;
  assign n6606 = n2251 & n6605 ;
  assign n6607 = ( n920 & ~n6566 ) | ( n920 & n6606 ) | ( ~n6566 & n6606 ) ;
  assign n6608 = ( n700 & n799 ) | ( n700 & ~n1010 ) | ( n799 & ~n1010 ) ;
  assign n6609 = n6608 ^ n5700 ^ 1'b0 ;
  assign n6610 = n6021 ^ n3718 ^ x55 ;
  assign n6611 = n2942 ^ n1549 ^ n499 ;
  assign n6612 = n6611 ^ n5881 ^ n4155 ;
  assign n6613 = ( ~n634 & n1229 ) | ( ~n634 & n6612 ) | ( n1229 & n6612 ) ;
  assign n6614 = n2278 ^ n1512 ^ 1'b0 ;
  assign n6615 = n1124 | n6614 ;
  assign n6616 = n6615 ^ n4138 ^ n1216 ;
  assign n6617 = ( ~n1803 & n3945 ) | ( ~n1803 & n6616 ) | ( n3945 & n6616 ) ;
  assign n6618 = n6617 ^ n723 ^ 1'b0 ;
  assign n6627 = n3857 | n6469 ;
  assign n6628 = n1114 & ~n6627 ;
  assign n6629 = n343 & n4136 ;
  assign n6630 = n6629 ^ n1623 ^ 1'b0 ;
  assign n6631 = n6630 ^ n3709 ^ 1'b0 ;
  assign n6632 = ( ~n565 & n6628 ) | ( ~n565 & n6631 ) | ( n6628 & n6631 ) ;
  assign n6624 = n978 | n6095 ;
  assign n6625 = n6624 ^ n5017 ^ 1'b0 ;
  assign n6626 = n6625 ^ n5097 ^ n645 ;
  assign n6633 = n6632 ^ n6626 ^ n638 ;
  assign n6619 = ~n2510 & n5224 ;
  assign n6620 = n6619 ^ n734 ^ 1'b0 ;
  assign n6621 = ( x227 & n1550 ) | ( x227 & ~n6620 ) | ( n1550 & ~n6620 ) ;
  assign n6622 = n6621 ^ n5119 ^ n2733 ;
  assign n6623 = x219 & ~n6622 ;
  assign n6634 = n6633 ^ n6623 ^ 1'b0 ;
  assign n6635 = n5767 ^ n2975 ^ n2417 ;
  assign n6636 = n3776 ^ n2881 ^ 1'b0 ;
  assign n6637 = n4980 & n6636 ;
  assign n6638 = n6635 | n6637 ;
  assign n6639 = n6293 ^ n6242 ^ n1748 ;
  assign n6640 = n6639 ^ n6091 ^ n5650 ;
  assign n6641 = n1837 | n2266 ;
  assign n6642 = n6641 ^ n2980 ^ 1'b0 ;
  assign n6643 = n6642 ^ n4449 ^ n322 ;
  assign n6644 = n435 & ~n3003 ;
  assign n6645 = n1951 & n6644 ;
  assign n6646 = ( x249 & n3439 ) | ( x249 & n6645 ) | ( n3439 & n6645 ) ;
  assign n6647 = n6187 | n6646 ;
  assign n6648 = x236 & n557 ;
  assign n6649 = n1792 ^ n666 ^ x187 ;
  assign n6650 = ( ~n3655 & n6648 ) | ( ~n3655 & n6649 ) | ( n6648 & n6649 ) ;
  assign n6651 = n4209 ^ n1891 ^ 1'b0 ;
  assign n6652 = n6650 | n6651 ;
  assign n6653 = n2589 ^ n1410 ^ 1'b0 ;
  assign n6654 = n2416 & n5536 ;
  assign n6655 = ( n454 & ~n6653 ) | ( n454 & n6654 ) | ( ~n6653 & n6654 ) ;
  assign n6657 = ( ~n933 & n1282 ) | ( ~n933 & n4414 ) | ( n1282 & n4414 ) ;
  assign n6656 = n5412 ^ n4965 ^ x233 ;
  assign n6658 = n6657 ^ n6656 ^ n1276 ;
  assign n6659 = n5034 ^ n1816 ^ n1543 ;
  assign n6660 = n2726 ^ n353 ^ 1'b0 ;
  assign n6661 = n6660 ^ n6474 ^ n674 ;
  assign n6662 = n6661 ^ n6549 ^ n1228 ;
  assign n6663 = ~n6659 & n6662 ;
  assign n6664 = ~n3130 & n6663 ;
  assign n6665 = ( n1928 & n5077 ) | ( n1928 & n6119 ) | ( n5077 & n6119 ) ;
  assign n6666 = n6665 ^ n443 ^ 1'b0 ;
  assign n6667 = n3638 ^ n3425 ^ n1179 ;
  assign n6668 = ( n337 & n6450 ) | ( n337 & n6667 ) | ( n6450 & n6667 ) ;
  assign n6669 = ~n3028 & n4999 ;
  assign n6670 = n6669 ^ x172 ^ 1'b0 ;
  assign n6671 = n1130 ^ n897 ^ n752 ;
  assign n6672 = n5823 & n6671 ;
  assign n6673 = n6672 ^ n5128 ^ 1'b0 ;
  assign n6674 = ( n5619 & n6670 ) | ( n5619 & ~n6673 ) | ( n6670 & ~n6673 ) ;
  assign n6675 = n1638 & ~n5798 ;
  assign n6676 = ( n736 & ~n4346 ) | ( n736 & n6675 ) | ( ~n4346 & n6675 ) ;
  assign n6677 = n2013 ^ n1566 ^ 1'b0 ;
  assign n6678 = n2804 ^ n2051 ^ n1095 ;
  assign n6679 = n4774 & n6678 ;
  assign n6680 = n5382 & ~n6679 ;
  assign n6681 = ~n6677 & n6680 ;
  assign n6682 = n5918 ^ n296 ^ n260 ;
  assign n6683 = n6682 ^ n4476 ^ n2232 ;
  assign n6684 = ~n2160 & n6484 ;
  assign n6685 = n6684 ^ n1258 ^ 1'b0 ;
  assign n6686 = ( n638 & n1071 ) | ( n638 & n3051 ) | ( n1071 & n3051 ) ;
  assign n6690 = n5601 ^ n323 ^ 1'b0 ;
  assign n6691 = ~n5590 & n6690 ;
  assign n6687 = n5904 ^ x223 ^ 1'b0 ;
  assign n6688 = n4950 | n6687 ;
  assign n6689 = n6688 ^ n4090 ^ n1005 ;
  assign n6692 = n6691 ^ n6689 ^ n1351 ;
  assign n6693 = ( ~n5675 & n5808 ) | ( ~n5675 & n6692 ) | ( n5808 & n6692 ) ;
  assign n6694 = n6686 | n6693 ;
  assign n6695 = n6685 | n6694 ;
  assign n6696 = n3624 ^ n1922 ^ x135 ;
  assign n6697 = x13 & n271 ;
  assign n6698 = n6697 ^ n3820 ^ n1288 ;
  assign n6699 = ~n6696 & n6698 ;
  assign n6700 = ~n1595 & n6699 ;
  assign n6701 = ( n2896 & ~n3022 ) | ( n2896 & n6700 ) | ( ~n3022 & n6700 ) ;
  assign n6703 = ~n920 & n3654 ;
  assign n6704 = n3869 & n6703 ;
  assign n6702 = ( n2988 & ~n5036 ) | ( n2988 & n5795 ) | ( ~n5036 & n5795 ) ;
  assign n6705 = n6704 ^ n6702 ^ n1910 ;
  assign n6706 = n724 & ~n4118 ;
  assign n6707 = n6706 ^ n6261 ^ 1'b0 ;
  assign n6708 = n3717 & ~n6707 ;
  assign n6719 = n303 | n1418 ;
  assign n6720 = n1832 | n6719 ;
  assign n6715 = ~n257 & n2085 ;
  assign n6716 = n685 & n6715 ;
  assign n6711 = ( n1705 & n2349 ) | ( n1705 & ~n4782 ) | ( n2349 & ~n4782 ) ;
  assign n6712 = n3381 ^ n2145 ^ x254 ;
  assign n6713 = ( n318 & n6711 ) | ( n318 & n6712 ) | ( n6711 & n6712 ) ;
  assign n6709 = n1032 & ~n1340 ;
  assign n6710 = n1405 | n6709 ;
  assign n6714 = n6713 ^ n6710 ^ 1'b0 ;
  assign n6717 = n6716 ^ n6714 ^ n5008 ;
  assign n6718 = n6717 ^ n3552 ^ n3319 ;
  assign n6721 = n6720 ^ n6718 ^ x196 ;
  assign n6722 = n5034 ^ n1056 ^ 1'b0 ;
  assign n6723 = n562 | n6722 ;
  assign n6724 = n6723 ^ n2388 ^ 1'b0 ;
  assign n6725 = n883 & ~n6724 ;
  assign n6726 = n6725 ^ n1668 ^ 1'b0 ;
  assign n6727 = n4378 ^ n1055 ^ 1'b0 ;
  assign n6728 = n6726 | n6727 ;
  assign n6729 = ( x167 & n2433 ) | ( x167 & n6018 ) | ( n2433 & n6018 ) ;
  assign n6730 = n2691 ^ n1550 ^ n1122 ;
  assign n6733 = n3280 & n5347 ;
  assign n6734 = n4431 & n6733 ;
  assign n6731 = n4738 ^ n2021 ^ x13 ;
  assign n6732 = ~n2751 & n6731 ;
  assign n6735 = n6734 ^ n6732 ^ 1'b0 ;
  assign n6736 = ( n961 & n1428 ) | ( n961 & ~n3494 ) | ( n1428 & ~n3494 ) ;
  assign n6737 = n6736 ^ n5248 ^ n2553 ;
  assign n6738 = x73 & n6737 ;
  assign n6739 = n6738 ^ n3219 ^ 1'b0 ;
  assign n6740 = ( n1728 & ~n3924 ) | ( n1728 & n6739 ) | ( ~n3924 & n6739 ) ;
  assign n6741 = n550 | n1755 ;
  assign n6744 = n902 ^ n572 ^ x103 ;
  assign n6742 = n5278 ^ n854 ^ 1'b0 ;
  assign n6743 = ~n4277 & n6742 ;
  assign n6745 = n6744 ^ n6743 ^ n1227 ;
  assign n6746 = n6745 ^ n1786 ^ 1'b0 ;
  assign n6747 = n4014 & ~n6746 ;
  assign n6748 = x80 ^ x43 ^ x42 ;
  assign n6749 = n6748 ^ x173 ^ 1'b0 ;
  assign n6750 = n6749 ^ n2510 ^ 1'b0 ;
  assign n6751 = n475 & ~n1190 ;
  assign n6752 = n604 & n6751 ;
  assign n6753 = n6752 ^ n4936 ^ n3214 ;
  assign n6754 = n643 | n3679 ;
  assign n6755 = n6753 & ~n6754 ;
  assign n6756 = ( n1549 & ~n2043 ) | ( n1549 & n5234 ) | ( ~n2043 & n5234 ) ;
  assign n6757 = n718 | n1418 ;
  assign n6758 = n4816 | n6757 ;
  assign n6759 = n2557 ^ n1758 ^ 1'b0 ;
  assign n6760 = n6758 & n6759 ;
  assign n6763 = n1691 | n2146 ;
  assign n6761 = n6319 ^ n2550 ^ 1'b0 ;
  assign n6762 = n6761 ^ n3939 ^ n1508 ;
  assign n6764 = n6763 ^ n6762 ^ 1'b0 ;
  assign n6765 = n6760 & n6764 ;
  assign n6766 = n1988 & n2954 ;
  assign n6767 = n6766 ^ n3218 ^ 1'b0 ;
  assign n6768 = ( n427 & n3255 ) | ( n427 & ~n6767 ) | ( n3255 & ~n6767 ) ;
  assign n6769 = ~n1766 & n4290 ;
  assign n6770 = n1050 | n4401 ;
  assign n6771 = n4791 & ~n6770 ;
  assign n6772 = ( n329 & ~n975 ) | ( n329 & n4217 ) | ( ~n975 & n4217 ) ;
  assign n6773 = n6772 ^ n4224 ^ n4138 ;
  assign n6774 = ( n712 & n4300 ) | ( n712 & ~n6773 ) | ( n4300 & ~n6773 ) ;
  assign n6775 = ( n1848 & n4231 ) | ( n1848 & n6774 ) | ( n4231 & n6774 ) ;
  assign n6776 = n4789 & n5883 ;
  assign n6777 = x75 & n266 ;
  assign n6778 = n6777 ^ n5589 ^ 1'b0 ;
  assign n6779 = n2325 | n6778 ;
  assign n6780 = n6779 ^ n521 ^ 1'b0 ;
  assign n6781 = n3367 ^ n2397 ^ n1829 ;
  assign n6782 = n2623 & n6781 ;
  assign n6783 = n6782 ^ n789 ^ 1'b0 ;
  assign n6784 = n6783 ^ n3313 ^ n2292 ;
  assign n6785 = n6784 ^ n4192 ^ 1'b0 ;
  assign n6786 = ( n1767 & n3231 ) | ( n1767 & n6785 ) | ( n3231 & n6785 ) ;
  assign n6787 = n3254 & n6786 ;
  assign n6788 = n1887 & ~n6787 ;
  assign n6789 = ~n6780 & n6788 ;
  assign n6790 = n1188 & ~n1853 ;
  assign n6791 = n6269 & n6790 ;
  assign n6792 = ~n2592 & n6711 ;
  assign n6793 = n6792 ^ n4230 ^ 1'b0 ;
  assign n6794 = n4279 & n6793 ;
  assign n6795 = n5193 & n6794 ;
  assign n6796 = n2393 ^ n1690 ^ n1122 ;
  assign n6797 = n6796 ^ n2960 ^ 1'b0 ;
  assign n6798 = n2631 & n6311 ;
  assign n6799 = ~n6797 & n6798 ;
  assign n6800 = n1487 ^ n426 ^ n353 ;
  assign n6801 = n2565 | n6800 ;
  assign n6802 = n6801 ^ n3253 ^ 1'b0 ;
  assign n6803 = ( n2537 & n5329 ) | ( n2537 & ~n5420 ) | ( n5329 & ~n5420 ) ;
  assign n6804 = ~n2031 & n6803 ;
  assign n6805 = n1474 & n6804 ;
  assign n6806 = n3507 ^ n1104 ^ 1'b0 ;
  assign n6807 = n6806 ^ x15 ^ 1'b0 ;
  assign n6808 = n6807 ^ n6652 ^ n310 ;
  assign n6809 = n4505 & n4599 ;
  assign n6810 = n6809 ^ n2978 ^ 1'b0 ;
  assign n6811 = ( ~x162 & n6214 ) | ( ~x162 & n6810 ) | ( n6214 & n6810 ) ;
  assign n6812 = n3612 ^ n1098 ^ 1'b0 ;
  assign n6813 = n1511 & ~n6812 ;
  assign n6823 = n2649 ^ n1200 ^ 1'b0 ;
  assign n6824 = n3167 & ~n6823 ;
  assign n6814 = n1629 ^ n1504 ^ 1'b0 ;
  assign n6815 = n2178 | n6814 ;
  assign n6816 = n5996 ^ n3075 ^ 1'b0 ;
  assign n6817 = x193 & ~n6816 ;
  assign n6818 = n6365 ^ n4384 ^ 1'b0 ;
  assign n6819 = n2880 & n6818 ;
  assign n6820 = ( n4697 & n6817 ) | ( n4697 & ~n6819 ) | ( n6817 & ~n6819 ) ;
  assign n6821 = n6815 | n6820 ;
  assign n6822 = n3650 & ~n6821 ;
  assign n6825 = n6824 ^ n6822 ^ n3003 ;
  assign n6826 = n4128 ^ n1693 ^ n654 ;
  assign n6827 = n6826 ^ n5135 ^ n1113 ;
  assign n6828 = n3933 ^ x213 ^ 1'b0 ;
  assign n6829 = n6268 ^ n4141 ^ n2234 ;
  assign n6830 = n6829 ^ x254 ^ x130 ;
  assign n6831 = ( n1900 & n2273 ) | ( n1900 & n6390 ) | ( n2273 & n6390 ) ;
  assign n6832 = n6831 ^ x32 ^ 1'b0 ;
  assign n6833 = ~n1961 & n3209 ;
  assign n6834 = n6832 & n6833 ;
  assign n6835 = n4828 & n6834 ;
  assign n6836 = n2145 & ~n6835 ;
  assign n6837 = n2418 & n6836 ;
  assign n6838 = n5020 ^ n3564 ^ n3187 ;
  assign n6839 = ( n1620 & ~n1887 ) | ( n1620 & n2073 ) | ( ~n1887 & n2073 ) ;
  assign n6840 = ( x197 & n4420 ) | ( x197 & ~n6839 ) | ( n4420 & ~n6839 ) ;
  assign n6841 = n6840 ^ n4908 ^ 1'b0 ;
  assign n6842 = n5412 & ~n6841 ;
  assign n6843 = ( n702 & n796 ) | ( n702 & ~n4848 ) | ( n796 & ~n4848 ) ;
  assign n6844 = n6843 ^ n2657 ^ 1'b0 ;
  assign n6845 = n1755 | n6483 ;
  assign n6846 = ~n1763 & n4439 ;
  assign n6847 = ( n525 & n1436 ) | ( n525 & ~n6463 ) | ( n1436 & ~n6463 ) ;
  assign n6848 = ( ~n1322 & n2669 ) | ( ~n1322 & n6847 ) | ( n2669 & n6847 ) ;
  assign n6849 = ( n2723 & ~n6846 ) | ( n2723 & n6848 ) | ( ~n6846 & n6848 ) ;
  assign n6850 = ( ~n991 & n1935 ) | ( ~n991 & n6849 ) | ( n1935 & n6849 ) ;
  assign n6851 = ( n799 & n3353 ) | ( n799 & n4738 ) | ( n3353 & n4738 ) ;
  assign n6854 = n2652 ^ n1949 ^ 1'b0 ;
  assign n6855 = n326 & n6854 ;
  assign n6852 = n5991 ^ n3391 ^ 1'b0 ;
  assign n6853 = n2157 & ~n6852 ;
  assign n6856 = n6855 ^ n6853 ^ n4164 ;
  assign n6857 = ( ~n2784 & n2861 ) | ( ~n2784 & n6856 ) | ( n2861 & n6856 ) ;
  assign n6858 = n5526 ^ n5204 ^ n1355 ;
  assign n6862 = x126 & ~n2224 ;
  assign n6863 = ~n4822 & n6862 ;
  assign n6859 = n542 & ~n4089 ;
  assign n6860 = n5748 & n6859 ;
  assign n6861 = n6860 ^ n4844 ^ n3499 ;
  assign n6864 = n6863 ^ n6861 ^ 1'b0 ;
  assign n6865 = n1104 | n2000 ;
  assign n6866 = ~n5713 & n6544 ;
  assign n6867 = n6866 ^ n1485 ^ 1'b0 ;
  assign n6868 = n6865 & ~n6867 ;
  assign n6869 = ( n793 & n2006 ) | ( n793 & n2709 ) | ( n2006 & n2709 ) ;
  assign n6870 = n6869 ^ n2207 ^ n2009 ;
  assign n6871 = n6870 ^ n3245 ^ n500 ;
  assign n6872 = n6726 ^ n4608 ^ n2350 ;
  assign n6873 = n1249 ^ n1186 ^ n550 ;
  assign n6874 = ( n1158 & ~n2800 ) | ( n1158 & n6873 ) | ( ~n2800 & n6873 ) ;
  assign n6875 = ~n865 & n6874 ;
  assign n6876 = ~n6873 & n6875 ;
  assign n6877 = n6872 & ~n6876 ;
  assign n6878 = ( x177 & n2598 ) | ( x177 & n4553 ) | ( n2598 & n4553 ) ;
  assign n6879 = n5168 ^ n2917 ^ 1'b0 ;
  assign n6880 = ( n502 & n1697 ) | ( n502 & ~n3306 ) | ( n1697 & ~n3306 ) ;
  assign n6881 = ( n6203 & n6879 ) | ( n6203 & n6880 ) | ( n6879 & n6880 ) ;
  assign n6882 = ( n5370 & n6878 ) | ( n5370 & ~n6881 ) | ( n6878 & ~n6881 ) ;
  assign n6883 = n3013 ^ n735 ^ 1'b0 ;
  assign n6884 = n2551 ^ n1214 ^ 1'b0 ;
  assign n6885 = n6883 & n6884 ;
  assign n6886 = n1042 & ~n5949 ;
  assign n6887 = n6886 ^ n3593 ^ 1'b0 ;
  assign n6888 = ( n2755 & n5110 ) | ( n2755 & n6887 ) | ( n5110 & n6887 ) ;
  assign n6889 = ( ~n1887 & n3660 ) | ( ~n1887 & n4160 ) | ( n3660 & n4160 ) ;
  assign n6890 = n4529 | n5480 ;
  assign n6891 = n887 | n6890 ;
  assign n6892 = n6891 ^ n5121 ^ n3151 ;
  assign n6893 = n6892 ^ n2756 ^ 1'b0 ;
  assign n6894 = ~n6889 & n6893 ;
  assign n6895 = n6894 ^ n1336 ^ 1'b0 ;
  assign n6896 = ( n4228 & n6888 ) | ( n4228 & ~n6895 ) | ( n6888 & ~n6895 ) ;
  assign n6897 = ( n567 & n965 ) | ( n567 & n1260 ) | ( n965 & n1260 ) ;
  assign n6898 = ( n3401 & ~n4301 ) | ( n3401 & n6897 ) | ( ~n4301 & n6897 ) ;
  assign n6899 = n3554 ^ n1387 ^ x28 ;
  assign n6900 = n1329 | n6899 ;
  assign n6901 = n287 | n6900 ;
  assign n6902 = n6901 ^ n4989 ^ 1'b0 ;
  assign n6903 = ( n1055 & n4524 ) | ( n1055 & ~n6902 ) | ( n4524 & ~n6902 ) ;
  assign n6904 = n1086 & ~n6317 ;
  assign n6905 = ( n1989 & n2700 ) | ( n1989 & ~n4681 ) | ( n2700 & ~n4681 ) ;
  assign n6906 = n6905 ^ n874 ^ 1'b0 ;
  assign n6907 = n628 & n6906 ;
  assign n6908 = ( n2063 & ~n2193 ) | ( n2063 & n6907 ) | ( ~n2193 & n6907 ) ;
  assign n6910 = n2453 & ~n3203 ;
  assign n6911 = n6910 ^ n2071 ^ 1'b0 ;
  assign n6912 = ( x129 & n1833 ) | ( x129 & n6911 ) | ( n1833 & n6911 ) ;
  assign n6913 = n2372 ^ n2355 ^ x129 ;
  assign n6914 = n6912 & ~n6913 ;
  assign n6915 = n6914 ^ n842 ^ 1'b0 ;
  assign n6909 = n6642 ^ n4274 ^ n2655 ;
  assign n6916 = n6915 ^ n6909 ^ n3690 ;
  assign n6917 = n1107 ^ n407 ^ 1'b0 ;
  assign n6918 = ( ~n2712 & n2845 ) | ( ~n2712 & n6917 ) | ( n2845 & n6917 ) ;
  assign n6919 = n6918 ^ n2190 ^ n1457 ;
  assign n6920 = n6919 ^ n5907 ^ n5388 ;
  assign n6921 = ( n1505 & n2237 ) | ( n1505 & ~n4460 ) | ( n2237 & ~n4460 ) ;
  assign n6922 = n6921 ^ n1628 ^ 1'b0 ;
  assign n6923 = n2749 & ~n6922 ;
  assign n6925 = n2810 ^ n1396 ^ 1'b0 ;
  assign n6926 = n6925 ^ n765 ^ 1'b0 ;
  assign n6924 = n1511 & ~n3037 ;
  assign n6927 = n6926 ^ n6924 ^ 1'b0 ;
  assign n6928 = ( n636 & n3954 ) | ( n636 & ~n5176 ) | ( n3954 & ~n5176 ) ;
  assign n6929 = ( n2875 & n6918 ) | ( n2875 & n6928 ) | ( n6918 & n6928 ) ;
  assign n6930 = ( n358 & n1676 ) | ( n358 & ~n5176 ) | ( n1676 & ~n5176 ) ;
  assign n6931 = n6930 ^ n2144 ^ 1'b0 ;
  assign n6932 = ~n6929 & n6931 ;
  assign n6933 = n6932 ^ n6796 ^ n1362 ;
  assign n6935 = n2681 ^ n2263 ^ n308 ;
  assign n6936 = n5146 & n6935 ;
  assign n6937 = ~n2645 & n6936 ;
  assign n6934 = ( ~n592 & n3280 ) | ( ~n592 & n3775 ) | ( n3280 & n3775 ) ;
  assign n6938 = n6937 ^ n6934 ^ n2690 ;
  assign n6939 = n6938 ^ n4771 ^ 1'b0 ;
  assign n6940 = n5031 & n6939 ;
  assign n6941 = ( ~n5272 & n5517 ) | ( ~n5272 & n6940 ) | ( n5517 & n6940 ) ;
  assign n6943 = n416 & ~n3080 ;
  assign n6944 = ~n2645 & n6943 ;
  assign n6945 = n6944 ^ n4131 ^ n1010 ;
  assign n6942 = ~n1561 & n5789 ;
  assign n6946 = n6945 ^ n6942 ^ 1'b0 ;
  assign n6947 = ( n1148 & n1432 ) | ( n1148 & n3720 ) | ( n1432 & n3720 ) ;
  assign n6948 = x208 & ~n4763 ;
  assign n6949 = n6948 ^ n3547 ^ n2598 ;
  assign n6954 = n2796 ^ n1691 ^ x137 ;
  assign n6951 = n4150 ^ n3446 ^ 1'b0 ;
  assign n6952 = n1879 & ~n6951 ;
  assign n6953 = n6952 ^ n2918 ^ 1'b0 ;
  assign n6950 = ( n464 & n1401 ) | ( n464 & ~n4723 ) | ( n1401 & ~n4723 ) ;
  assign n6955 = n6954 ^ n6953 ^ n6950 ;
  assign n6956 = n4922 ^ n3672 ^ n2634 ;
  assign n6957 = ( n1880 & n2545 ) | ( n1880 & ~n6956 ) | ( n2545 & ~n6956 ) ;
  assign n6958 = n2510 | n6957 ;
  assign n6959 = n6955 & ~n6958 ;
  assign n6971 = n4185 ^ n462 ^ 1'b0 ;
  assign n6972 = n6971 ^ n2936 ^ n1320 ;
  assign n6960 = x251 | n3075 ;
  assign n6965 = n4609 ^ n1550 ^ 1'b0 ;
  assign n6966 = n2680 & ~n6965 ;
  assign n6964 = n3166 | n4325 ;
  assign n6967 = n6966 ^ n6964 ^ 1'b0 ;
  assign n6962 = n4171 | n5385 ;
  assign n6961 = n5268 ^ n2708 ^ 1'b0 ;
  assign n6963 = n6962 ^ n6961 ^ 1'b0 ;
  assign n6968 = n6967 ^ n6963 ^ n4653 ;
  assign n6969 = ( ~n1318 & n6083 ) | ( ~n1318 & n6968 ) | ( n6083 & n6968 ) ;
  assign n6970 = n6960 & n6969 ;
  assign n6973 = n6972 ^ n6970 ^ 1'b0 ;
  assign n6974 = n3992 ^ x211 ^ 1'b0 ;
  assign n6975 = ( n1131 & n3037 ) | ( n1131 & ~n3445 ) | ( n3037 & ~n3445 ) ;
  assign n6976 = ( n2079 & n4701 ) | ( n2079 & ~n6975 ) | ( n4701 & ~n6975 ) ;
  assign n6977 = n6348 ^ n3122 ^ n2417 ;
  assign n6978 = ~n6976 & n6977 ;
  assign n6979 = n6978 ^ n2459 ^ 1'b0 ;
  assign n6980 = n2183 & n3399 ;
  assign n6981 = n4155 ^ n3243 ^ n638 ;
  assign n6982 = ( n3415 & n4761 ) | ( n3415 & ~n6981 ) | ( n4761 & ~n6981 ) ;
  assign n6983 = n6032 ^ n5328 ^ n3715 ;
  assign n6984 = n6727 & ~n6983 ;
  assign n6985 = n6984 ^ n4385 ^ 1'b0 ;
  assign n6986 = n2128 | n6985 ;
  assign n6996 = n1428 ^ n599 ^ 1'b0 ;
  assign n6997 = n5972 & ~n6996 ;
  assign n6987 = n3783 ^ n1540 ^ 1'b0 ;
  assign n6988 = ~n1803 & n6987 ;
  assign n6989 = n1592 & n6988 ;
  assign n6990 = ( ~n1763 & n3567 ) | ( ~n1763 & n6989 ) | ( n3567 & n6989 ) ;
  assign n6991 = n1086 ^ n520 ^ 1'b0 ;
  assign n6992 = n5245 | n6991 ;
  assign n6993 = n4294 & ~n6992 ;
  assign n6994 = n6993 ^ n4279 ^ n1587 ;
  assign n6995 = ( n4271 & n6990 ) | ( n4271 & n6994 ) | ( n6990 & n6994 ) ;
  assign n6998 = n6997 ^ n6995 ^ 1'b0 ;
  assign n6999 = n5715 ^ x186 ^ 1'b0 ;
  assign n7000 = n720 & ~n6999 ;
  assign n7001 = n6998 & n7000 ;
  assign n7002 = n1307 & n4756 ;
  assign n7003 = ~x50 & n7002 ;
  assign n7004 = n4018 & ~n7003 ;
  assign n7005 = n4421 ^ n2436 ^ n706 ;
  assign n7006 = ( n902 & n7004 ) | ( n902 & n7005 ) | ( n7004 & n7005 ) ;
  assign n7007 = n811 ^ x182 ^ 1'b0 ;
  assign n7008 = n7007 ^ n5380 ^ n707 ;
  assign n7009 = ( ~n304 & n2811 ) | ( ~n304 & n3167 ) | ( n2811 & n3167 ) ;
  assign n7010 = ( n5945 & ~n7008 ) | ( n5945 & n7009 ) | ( ~n7008 & n7009 ) ;
  assign n7012 = n4111 | n4775 ;
  assign n7013 = n7012 ^ n4529 ^ 1'b0 ;
  assign n7011 = n3666 ^ n2232 ^ n1736 ;
  assign n7014 = n7013 ^ n7011 ^ n268 ;
  assign n7015 = n7014 ^ n4756 ^ 1'b0 ;
  assign n7016 = ~n7010 & n7015 ;
  assign n7023 = ( ~n741 & n1617 ) | ( ~n741 & n1679 ) | ( n1617 & n1679 ) ;
  assign n7024 = n7023 ^ n4342 ^ n2342 ;
  assign n7020 = n1672 | n4998 ;
  assign n7021 = n470 & ~n7020 ;
  assign n7018 = ( n518 & n2105 ) | ( n518 & n6950 ) | ( n2105 & n6950 ) ;
  assign n7017 = x245 & n667 ;
  assign n7019 = n7018 ^ n7017 ^ 1'b0 ;
  assign n7022 = n7021 ^ n7019 ^ n6255 ;
  assign n7025 = n7024 ^ n7022 ^ n1145 ;
  assign n7028 = n2724 & n4595 ;
  assign n7029 = n2813 & n7028 ;
  assign n7030 = n7029 ^ x28 ^ 1'b0 ;
  assign n7026 = n4817 ^ n2162 ^ 1'b0 ;
  assign n7027 = n3151 | n7026 ;
  assign n7031 = n7030 ^ n7027 ^ n3934 ;
  assign n7032 = ~n408 & n1572 ;
  assign n7033 = n916 & n7032 ;
  assign n7034 = n2043 & ~n6998 ;
  assign n7035 = ~x100 & n7034 ;
  assign n7036 = n5957 ^ n5082 ^ n3725 ;
  assign n7037 = n5584 ^ n4222 ^ n1777 ;
  assign n7038 = ( ~n4025 & n6859 ) | ( ~n4025 & n7037 ) | ( n6859 & n7037 ) ;
  assign n7039 = n1367 & n7038 ;
  assign n7040 = ~n7036 & n7039 ;
  assign n7041 = n3159 ^ n1384 ^ 1'b0 ;
  assign n7042 = n4169 & n7041 ;
  assign n7043 = n3662 ^ n300 ^ 1'b0 ;
  assign n7044 = n2577 & n7043 ;
  assign n7045 = ( n2600 & ~n7042 ) | ( n2600 & n7044 ) | ( ~n7042 & n7044 ) ;
  assign n7046 = n7045 ^ x151 ^ 1'b0 ;
  assign n7047 = ~n1570 & n7046 ;
  assign n7048 = n1952 & ~n2782 ;
  assign n7049 = ~n3897 & n7048 ;
  assign n7050 = n638 & ~n7049 ;
  assign n7051 = n3786 & n7050 ;
  assign n7052 = ( n594 & n2267 ) | ( n594 & n2376 ) | ( n2267 & n2376 ) ;
  assign n7053 = n1924 ^ x73 ^ 1'b0 ;
  assign n7054 = n7053 ^ n2348 ^ 1'b0 ;
  assign n7055 = x109 & n7054 ;
  assign n7056 = ( x6 & n7052 ) | ( x6 & ~n7055 ) | ( n7052 & ~n7055 ) ;
  assign n7057 = n6119 ^ n2615 ^ n438 ;
  assign n7058 = n3379 | n7057 ;
  assign n7059 = n1167 | n3306 ;
  assign n7060 = n3790 | n7059 ;
  assign n7061 = n3058 ^ n542 ^ 1'b0 ;
  assign n7062 = n7061 ^ n436 ^ 1'b0 ;
  assign n7063 = n7062 ^ n5259 ^ n1883 ;
  assign n7064 = ~n2791 & n5523 ;
  assign n7065 = n7064 ^ x163 ^ 1'b0 ;
  assign n7066 = n2112 | n7065 ;
  assign n7067 = n7063 & ~n7066 ;
  assign n7074 = ~n1776 & n2648 ;
  assign n7075 = ~n4046 & n7074 ;
  assign n7072 = n4596 ^ n3804 ^ x71 ;
  assign n7073 = n4985 | n7072 ;
  assign n7076 = n7075 ^ n7073 ^ n3167 ;
  assign n7068 = n829 & n1508 ;
  assign n7069 = ~n512 & n7068 ;
  assign n7070 = n5568 ^ n2109 ^ n2090 ;
  assign n7071 = n7069 | n7070 ;
  assign n7077 = n7076 ^ n7071 ^ 1'b0 ;
  assign n7078 = ( n1562 & n3673 ) | ( n1562 & ~n7077 ) | ( n3673 & ~n7077 ) ;
  assign n7079 = n4634 ^ n3397 ^ n1789 ;
  assign n7080 = n7079 ^ n6819 ^ n3879 ;
  assign n7081 = n6113 ^ n3105 ^ x54 ;
  assign n7082 = n5392 ^ n1381 ^ x198 ;
  assign n7083 = ( ~x56 & n1486 ) | ( ~x56 & n7082 ) | ( n1486 & n7082 ) ;
  assign n7084 = n7083 ^ n632 ^ 1'b0 ;
  assign n7085 = n441 & n1087 ;
  assign n7086 = n1114 & n7085 ;
  assign n7087 = n262 | n7086 ;
  assign n7088 = ( n3226 & ~n7084 ) | ( n3226 & n7087 ) | ( ~n7084 & n7087 ) ;
  assign n7089 = n729 ^ n418 ^ 1'b0 ;
  assign n7090 = n2960 & n7089 ;
  assign n7091 = n7090 ^ n6642 ^ 1'b0 ;
  assign n7092 = n7091 ^ n6433 ^ n5340 ;
  assign n7093 = n618 & ~n3133 ;
  assign n7094 = ( ~n740 & n3723 ) | ( ~n740 & n7093 ) | ( n3723 & n7093 ) ;
  assign n7097 = ~x132 & n2301 ;
  assign n7095 = x86 & x115 ;
  assign n7096 = ~n4022 & n7095 ;
  assign n7098 = n7097 ^ n7096 ^ x22 ;
  assign n7099 = n7098 ^ n3010 ^ 1'b0 ;
  assign n7100 = n7099 ^ n5175 ^ n565 ;
  assign n7101 = n1743 ^ n1255 ^ x234 ;
  assign n7102 = n6563 ^ n1470 ^ 1'b0 ;
  assign n7103 = n5634 ^ n2918 ^ n2546 ;
  assign n7104 = ( n751 & n4782 ) | ( n751 & ~n7103 ) | ( n4782 & ~n7103 ) ;
  assign n7105 = n1714 ^ x213 ^ 1'b0 ;
  assign n7106 = n5099 | n7105 ;
  assign n7107 = n4640 | n7106 ;
  assign n7108 = n2050 & ~n7107 ;
  assign n7109 = n5640 ^ n2904 ^ 1'b0 ;
  assign n7110 = ~n7108 & n7109 ;
  assign n7111 = n7110 ^ n3634 ^ n2987 ;
  assign n7112 = n7111 ^ n1239 ^ n661 ;
  assign n7113 = n7112 ^ n2094 ^ n500 ;
  assign n7115 = ~n1534 & n2124 ;
  assign n7116 = n7115 ^ n2174 ^ 1'b0 ;
  assign n7114 = n3126 ^ n1156 ^ x68 ;
  assign n7117 = n7116 ^ n7114 ^ n2731 ;
  assign n7118 = n1745 & ~n7117 ;
  assign n7119 = ( n1077 & n2682 ) | ( n1077 & n4783 ) | ( n2682 & n4783 ) ;
  assign n7120 = n7119 ^ n3317 ^ n1139 ;
  assign n7121 = n7120 ^ n4706 ^ 1'b0 ;
  assign n7122 = ~n7118 & n7121 ;
  assign n7125 = n3364 ^ n2269 ^ n600 ;
  assign n7123 = n683 | n3869 ;
  assign n7124 = n7123 ^ n1546 ^ 1'b0 ;
  assign n7126 = n7125 ^ n7124 ^ n759 ;
  assign n7127 = n7126 ^ n2470 ^ 1'b0 ;
  assign n7128 = ( n399 & ~n2592 ) | ( n399 & n7127 ) | ( ~n2592 & n7127 ) ;
  assign n7129 = n5017 ^ n2500 ^ 1'b0 ;
  assign n7130 = ( n1781 & n7128 ) | ( n1781 & n7129 ) | ( n7128 & n7129 ) ;
  assign n7131 = n3190 ^ n1723 ^ n1585 ;
  assign n7132 = ~n1032 & n7131 ;
  assign n7133 = ~n1073 & n7132 ;
  assign n7134 = ( n2240 & n4510 ) | ( n2240 & ~n7133 ) | ( n4510 & ~n7133 ) ;
  assign n7135 = ~n1180 & n3672 ;
  assign n7136 = n7135 ^ n7007 ^ 1'b0 ;
  assign n7137 = ( n2450 & ~n6304 ) | ( n2450 & n7136 ) | ( ~n6304 & n7136 ) ;
  assign n7138 = ( n1003 & n1673 ) | ( n1003 & ~n1988 ) | ( n1673 & ~n1988 ) ;
  assign n7139 = ( n6277 & n6494 ) | ( n6277 & n7138 ) | ( n6494 & n7138 ) ;
  assign n7140 = n6741 | n6913 ;
  assign n7141 = x157 | n7140 ;
  assign n7142 = n1328 ^ x23 ^ 1'b0 ;
  assign n7143 = n5460 ^ n4680 ^ 1'b0 ;
  assign n7144 = n1311 & ~n7143 ;
  assign n7145 = n7144 ^ n4694 ^ 1'b0 ;
  assign n7146 = n7142 | n7145 ;
  assign n7147 = n7146 ^ n4331 ^ 1'b0 ;
  assign n7148 = n7147 ^ n2602 ^ 1'b0 ;
  assign n7149 = n2546 ^ n945 ^ 1'b0 ;
  assign n7150 = n6235 & n7149 ;
  assign n7151 = n2571 ^ n1395 ^ 1'b0 ;
  assign n7152 = n981 | n7151 ;
  assign n7153 = ( n5867 & n7150 ) | ( n5867 & ~n7152 ) | ( n7150 & ~n7152 ) ;
  assign n7154 = n4465 ^ n1747 ^ 1'b0 ;
  assign n7155 = n3503 | n7154 ;
  assign n7156 = n6915 ^ n3732 ^ 1'b0 ;
  assign n7157 = ~n7155 & n7156 ;
  assign n7158 = n1438 | n3325 ;
  assign n7159 = n7158 ^ n3502 ^ 1'b0 ;
  assign n7160 = n7159 ^ n4078 ^ n3144 ;
  assign n7167 = ~n1260 & n2012 ;
  assign n7161 = n478 & ~n4892 ;
  assign n7162 = ~n2107 & n7161 ;
  assign n7163 = n1367 ^ n1319 ^ n750 ;
  assign n7164 = n4078 & n7163 ;
  assign n7165 = ( ~n4006 & n5709 ) | ( ~n4006 & n7164 ) | ( n5709 & n7164 ) ;
  assign n7166 = n7162 | n7165 ;
  assign n7168 = n7167 ^ n7166 ^ 1'b0 ;
  assign n7174 = ( x185 & n866 ) | ( x185 & ~n1214 ) | ( n866 & ~n1214 ) ;
  assign n7175 = ( n2828 & n5373 ) | ( n2828 & n7174 ) | ( n5373 & n7174 ) ;
  assign n7176 = n7175 ^ n4638 ^ 1'b0 ;
  assign n7177 = n4782 & ~n7176 ;
  assign n7178 = n7177 ^ n6598 ^ n3744 ;
  assign n7169 = n5570 ^ n4068 ^ n2443 ;
  assign n7170 = n7169 ^ n4035 ^ 1'b0 ;
  assign n7171 = ~n3867 & n7170 ;
  assign n7172 = n2434 | n7171 ;
  assign n7173 = n7172 ^ n5696 ^ n3358 ;
  assign n7179 = n7178 ^ n7173 ^ n1826 ;
  assign n7180 = ( n2448 & n3391 ) | ( n2448 & n4608 ) | ( n3391 & n4608 ) ;
  assign n7181 = ( n2333 & ~n5688 ) | ( n2333 & n7180 ) | ( ~n5688 & n7180 ) ;
  assign n7185 = ( n1372 & ~n1481 ) | ( n1372 & n3585 ) | ( ~n1481 & n3585 ) ;
  assign n7186 = x231 & ~n7185 ;
  assign n7187 = n7186 ^ n1304 ^ n672 ;
  assign n7182 = ~n1230 & n2476 ;
  assign n7183 = n7182 ^ n4826 ^ 1'b0 ;
  assign n7184 = n3921 | n7183 ;
  assign n7188 = n7187 ^ n7184 ^ n5919 ;
  assign n7189 = ( n1685 & n2178 ) | ( n1685 & ~n2315 ) | ( n2178 & ~n2315 ) ;
  assign n7190 = n7189 ^ n2910 ^ 1'b0 ;
  assign n7191 = ~n2878 & n7190 ;
  assign n7192 = n1331 ^ x109 ^ 1'b0 ;
  assign n7193 = ~n3771 & n7192 ;
  assign n7194 = n2810 | n5480 ;
  assign n7195 = n6483 | n7194 ;
  assign n7196 = ( n798 & ~n7193 ) | ( n798 & n7195 ) | ( ~n7193 & n7195 ) ;
  assign n7197 = ( n1743 & ~n1948 ) | ( n1743 & n2165 ) | ( ~n1948 & n2165 ) ;
  assign n7198 = ( n1189 & ~n6850 ) | ( n1189 & n7197 ) | ( ~n6850 & n7197 ) ;
  assign n7207 = ( ~x155 & x171 ) | ( ~x155 & n623 ) | ( x171 & n623 ) ;
  assign n7208 = n2765 & n3276 ;
  assign n7209 = n7208 ^ x39 ^ 1'b0 ;
  assign n7210 = n7209 ^ n5806 ^ n1037 ;
  assign n7211 = ( n4071 & n7207 ) | ( n4071 & n7210 ) | ( n7207 & n7210 ) ;
  assign n7205 = n1697 | n2878 ;
  assign n7206 = n1114 & ~n7205 ;
  assign n7202 = n679 | n2272 ;
  assign n7203 = n986 & ~n7202 ;
  assign n7199 = n1821 ^ n1309 ^ x253 ;
  assign n7200 = ( n2077 & n5405 ) | ( n2077 & ~n7199 ) | ( n5405 & ~n7199 ) ;
  assign n7201 = n7200 ^ n4132 ^ n1557 ;
  assign n7204 = n7203 ^ n7201 ^ 1'b0 ;
  assign n7212 = n7211 ^ n7206 ^ n7204 ;
  assign n7213 = ( ~n1185 & n1803 ) | ( ~n1185 & n2681 ) | ( n1803 & n2681 ) ;
  assign n7218 = n2819 ^ n2209 ^ n1358 ;
  assign n7214 = n1315 ^ n831 ^ n772 ;
  assign n7215 = n7214 ^ n2600 ^ n276 ;
  assign n7216 = n3507 ^ n2535 ^ 1'b0 ;
  assign n7217 = ( n6050 & n7215 ) | ( n6050 & n7216 ) | ( n7215 & n7216 ) ;
  assign n7219 = n7218 ^ n7217 ^ 1'b0 ;
  assign n7220 = ( n5412 & n7213 ) | ( n5412 & n7219 ) | ( n7213 & n7219 ) ;
  assign n7221 = n5278 ^ n4902 ^ n2425 ;
  assign n7222 = n7221 ^ n3094 ^ n626 ;
  assign n7223 = n5343 ^ n4421 ^ n2482 ;
  assign n7224 = ~n7222 & n7223 ;
  assign n7225 = n2572 ^ x147 ^ 1'b0 ;
  assign n7226 = n4640 | n7225 ;
  assign n7227 = ( n3075 & n5784 ) | ( n3075 & ~n7226 ) | ( n5784 & ~n7226 ) ;
  assign n7228 = n7227 ^ n1669 ^ 1'b0 ;
  assign n7229 = n7228 ^ n6661 ^ 1'b0 ;
  assign n7230 = n5119 & n5801 ;
  assign n7231 = n3761 ^ n1121 ^ 1'b0 ;
  assign n7232 = n4021 | n7231 ;
  assign n7233 = ( ~n3942 & n5886 ) | ( ~n3942 & n7232 ) | ( n5886 & n7232 ) ;
  assign n7234 = n6036 ^ n5609 ^ 1'b0 ;
  assign n7235 = ( n558 & n1233 ) | ( n558 & ~n3245 ) | ( n1233 & ~n3245 ) ;
  assign n7236 = ( n3400 & n3493 ) | ( n3400 & ~n7235 ) | ( n3493 & ~n7235 ) ;
  assign n7240 = n4771 & n6594 ;
  assign n7241 = ~n5419 & n7240 ;
  assign n7237 = n2300 | n2997 ;
  assign n7238 = n4065 | n7237 ;
  assign n7239 = n7238 ^ n2943 ^ n2803 ;
  assign n7242 = n7241 ^ n7239 ^ 1'b0 ;
  assign n7243 = n7236 & n7242 ;
  assign n7244 = n5065 ^ n4525 ^ n2832 ;
  assign n7245 = n4412 & n7244 ;
  assign n7246 = ~n7243 & n7245 ;
  assign n7247 = n4745 ^ n1676 ^ n856 ;
  assign n7248 = n673 & n4078 ;
  assign n7249 = ( n4464 & n7247 ) | ( n4464 & n7248 ) | ( n7247 & n7248 ) ;
  assign n7253 = ( x240 & n1058 ) | ( x240 & ~n1767 ) | ( n1058 & ~n1767 ) ;
  assign n7254 = n7253 ^ n5710 ^ n2933 ;
  assign n7250 = n2274 | n2337 ;
  assign n7251 = n7250 ^ n5066 ^ n2195 ;
  assign n7252 = ~n2141 & n7251 ;
  assign n7255 = n7254 ^ n7252 ^ 1'b0 ;
  assign n7256 = ~n2187 & n4488 ;
  assign n7257 = ( n3335 & ~n4662 ) | ( n3335 & n7256 ) | ( ~n4662 & n7256 ) ;
  assign n7258 = n3956 ^ n1118 ^ x98 ;
  assign n7259 = ( n5367 & n7253 ) | ( n5367 & n7258 ) | ( n7253 & n7258 ) ;
  assign n7260 = ( x26 & n1821 ) | ( x26 & n6829 ) | ( n1821 & n6829 ) ;
  assign n7261 = ( n658 & n3273 ) | ( n658 & ~n5542 ) | ( n3273 & ~n5542 ) ;
  assign n7262 = n6863 ^ n4085 ^ n2877 ;
  assign n7263 = n4897 & ~n6963 ;
  assign n7264 = n4828 ^ x94 ^ x51 ;
  assign n7265 = n7264 ^ n3129 ^ n3115 ;
  assign n7266 = n7263 & ~n7265 ;
  assign n7267 = n2436 ^ n1037 ^ 1'b0 ;
  assign n7268 = n333 & n7267 ;
  assign n7269 = n7268 ^ n546 ^ 1'b0 ;
  assign n7270 = n7269 ^ n4090 ^ n2222 ;
  assign n7271 = ~n1804 & n7270 ;
  assign n7272 = ~n4044 & n4931 ;
  assign n7273 = n5208 & ~n7272 ;
  assign n7274 = n5560 & n7273 ;
  assign n7275 = n7271 & ~n7274 ;
  assign n7276 = n5332 & n7275 ;
  assign n7277 = n5415 ^ n1930 ^ 1'b0 ;
  assign n7278 = n7277 ^ n2416 ^ x209 ;
  assign n7279 = ( n698 & n910 ) | ( n698 & n3145 ) | ( n910 & n3145 ) ;
  assign n7280 = ( ~n3235 & n4156 ) | ( ~n3235 & n7279 ) | ( n4156 & n7279 ) ;
  assign n7281 = x88 | n7280 ;
  assign n7282 = ( x130 & ~x139 ) | ( x130 & n7281 ) | ( ~x139 & n7281 ) ;
  assign n7283 = n6100 ^ n4853 ^ n613 ;
  assign n7284 = ( n2391 & ~n6178 ) | ( n2391 & n7283 ) | ( ~n6178 & n7283 ) ;
  assign n7285 = ( x208 & n3977 ) | ( x208 & ~n4480 ) | ( n3977 & ~n4480 ) ;
  assign n7286 = ( n642 & ~n6056 ) | ( n642 & n7285 ) | ( ~n6056 & n7285 ) ;
  assign n7287 = n7286 ^ n627 ^ 1'b0 ;
  assign n7288 = n2405 & ~n7287 ;
  assign n7289 = ( x89 & n3971 ) | ( x89 & n6650 ) | ( n3971 & n6650 ) ;
  assign n7290 = n7289 ^ n5300 ^ 1'b0 ;
  assign n7291 = n2927 ^ n750 ^ 1'b0 ;
  assign n7292 = ( n3210 & n4463 ) | ( n3210 & ~n7291 ) | ( n4463 & ~n7291 ) ;
  assign n7294 = n3319 & n5152 ;
  assign n7293 = n545 & ~n1998 ;
  assign n7295 = n7294 ^ n7293 ^ 1'b0 ;
  assign n7296 = ( n2384 & ~n2712 ) | ( n2384 & n7295 ) | ( ~n2712 & n7295 ) ;
  assign n7297 = ( n997 & ~n1192 ) | ( n997 & n2896 ) | ( ~n1192 & n2896 ) ;
  assign n7298 = ~n5353 & n7297 ;
  assign n7299 = n6193 ^ n550 ^ 1'b0 ;
  assign n7300 = n7298 & n7299 ;
  assign n7301 = n7300 ^ n4975 ^ n4298 ;
  assign n7302 = n4426 ^ n1563 ^ 1'b0 ;
  assign n7303 = n485 & ~n7302 ;
  assign n7304 = n7303 ^ n5992 ^ 1'b0 ;
  assign n7305 = n3458 & ~n7304 ;
  assign n7306 = n7227 ^ n6059 ^ n683 ;
  assign n7309 = ~n787 & n2094 ;
  assign n7307 = ~n1863 & n1974 ;
  assign n7308 = ~n6434 & n7307 ;
  assign n7310 = n7309 ^ n7308 ^ 1'b0 ;
  assign n7311 = n7310 ^ n1544 ^ 1'b0 ;
  assign n7312 = ( n5271 & n7306 ) | ( n5271 & ~n7311 ) | ( n7306 & ~n7311 ) ;
  assign n7313 = ~n6459 & n6665 ;
  assign n7314 = n4249 ^ n3838 ^ n2080 ;
  assign n7315 = n7314 ^ n6643 ^ 1'b0 ;
  assign n7316 = x170 & ~n7315 ;
  assign n7317 = ~n1364 & n1942 ;
  assign n7318 = n4603 ^ n3747 ^ n1044 ;
  assign n7319 = n7318 ^ n4450 ^ 1'b0 ;
  assign n7320 = n7317 | n7319 ;
  assign n7321 = n3703 | n7320 ;
  assign n7322 = n2594 | n7321 ;
  assign n7323 = ~n2831 & n7322 ;
  assign n7324 = n925 & ~n6883 ;
  assign n7325 = n1180 & n7324 ;
  assign n7326 = n7325 ^ n2200 ^ 1'b0 ;
  assign n7329 = n3164 ^ n1870 ^ 1'b0 ;
  assign n7327 = n2171 ^ n1823 ^ 1'b0 ;
  assign n7328 = n5996 & n7327 ;
  assign n7330 = n7329 ^ n7328 ^ 1'b0 ;
  assign n7331 = n7330 ^ n983 ^ 1'b0 ;
  assign n7332 = n7326 & n7331 ;
  assign n7333 = ( ~x70 & n1909 ) | ( ~x70 & n2337 ) | ( n1909 & n2337 ) ;
  assign n7334 = n3615 | n7133 ;
  assign n7335 = ( ~n6193 & n7065 ) | ( ~n6193 & n7334 ) | ( n7065 & n7334 ) ;
  assign n7336 = n7335 ^ n3220 ^ 1'b0 ;
  assign n7337 = n2346 | n7336 ;
  assign n7338 = n2892 & n4558 ;
  assign n7339 = n7337 & n7338 ;
  assign n7340 = x142 & n1276 ;
  assign n7341 = n7340 ^ n3905 ^ 1'b0 ;
  assign n7342 = n3561 ^ n1926 ^ 1'b0 ;
  assign n7343 = n3489 & n7325 ;
  assign n7344 = n7343 ^ n4723 ^ n3740 ;
  assign n7345 = n1167 ^ n298 ^ x21 ;
  assign n7346 = n5991 & ~n7345 ;
  assign n7347 = n7346 ^ n4797 ^ n3160 ;
  assign n7348 = n1645 & n4348 ;
  assign n7349 = ~n7347 & n7348 ;
  assign n7350 = n7349 ^ n3828 ^ n2644 ;
  assign n7351 = ( ~n720 & n3154 ) | ( ~n720 & n3516 ) | ( n3154 & n3516 ) ;
  assign n7352 = ( n7344 & n7350 ) | ( n7344 & n7351 ) | ( n7350 & n7351 ) ;
  assign n7353 = n7342 | n7352 ;
  assign n7354 = n7341 | n7353 ;
  assign n7355 = n327 & n7354 ;
  assign n7356 = n7355 ^ n5888 ^ 1'b0 ;
  assign n7357 = ~n1833 & n3439 ;
  assign n7358 = ~n2226 & n7357 ;
  assign n7359 = n7358 ^ n488 ^ x7 ;
  assign n7360 = n4659 & ~n6294 ;
  assign n7361 = ~n1597 & n6211 ;
  assign n7362 = n7361 ^ n1890 ^ 1'b0 ;
  assign n7363 = ( ~n2912 & n7360 ) | ( ~n2912 & n7362 ) | ( n7360 & n7362 ) ;
  assign n7364 = n7346 ^ n2682 ^ n587 ;
  assign n7365 = ( n530 & n6322 ) | ( n530 & ~n7364 ) | ( n6322 & ~n7364 ) ;
  assign n7368 = n2655 ^ n1524 ^ 1'b0 ;
  assign n7369 = n1394 & n7368 ;
  assign n7366 = n2996 ^ n2148 ^ 1'b0 ;
  assign n7367 = n7366 ^ n5278 ^ n3159 ;
  assign n7370 = n7369 ^ n7367 ^ n2212 ;
  assign n7371 = n7370 ^ n1205 ^ 1'b0 ;
  assign n7372 = n3493 & n7371 ;
  assign n7373 = n6760 & n7372 ;
  assign n7374 = ~n3604 & n7373 ;
  assign n7375 = n352 & ~n5061 ;
  assign n7376 = ~n7279 & n7375 ;
  assign n7377 = n7376 ^ n6442 ^ n410 ;
  assign n7378 = n569 | n7377 ;
  assign n7384 = n3834 ^ n3445 ^ n2990 ;
  assign n7379 = ( n433 & ~n1550 ) | ( n433 & n6209 ) | ( ~n1550 & n6209 ) ;
  assign n7380 = x208 & n7379 ;
  assign n7381 = ~n5576 & n7380 ;
  assign n7382 = ( n4046 & n4327 ) | ( n4046 & ~n6640 ) | ( n4327 & ~n6640 ) ;
  assign n7383 = ~n7381 & n7382 ;
  assign n7385 = n7384 ^ n7383 ^ 1'b0 ;
  assign n7387 = n5325 ^ n3620 ^ 1'b0 ;
  assign n7386 = ( ~n1787 & n2177 ) | ( ~n1787 & n2727 ) | ( n2177 & n2727 ) ;
  assign n7388 = n7387 ^ n7386 ^ n1625 ;
  assign n7389 = ( ~x122 & x128 ) | ( ~x122 & n2053 ) | ( x128 & n2053 ) ;
  assign n7390 = n3355 | n7389 ;
  assign n7391 = ( n3371 & n5613 ) | ( n3371 & n7390 ) | ( n5613 & n7390 ) ;
  assign n7392 = ~n2711 & n7391 ;
  assign n7393 = ~n2060 & n5669 ;
  assign n7394 = n1156 ^ x189 ^ 1'b0 ;
  assign n7395 = n6483 & n7394 ;
  assign n7396 = ( n4908 & ~n7393 ) | ( n4908 & n7395 ) | ( ~n7393 & n7395 ) ;
  assign n7397 = n6542 ^ n4556 ^ 1'b0 ;
  assign n7398 = n3117 ^ n2085 ^ 1'b0 ;
  assign n7399 = n1880 ^ x109 ^ x23 ;
  assign n7400 = n5460 & n7399 ;
  assign n7401 = ( n3106 & n3220 ) | ( n3106 & ~n5051 ) | ( n3220 & ~n5051 ) ;
  assign n7402 = ( n3339 & ~n5452 ) | ( n3339 & n6131 ) | ( ~n5452 & n6131 ) ;
  assign n7403 = ( n2666 & ~n5146 ) | ( n2666 & n6177 ) | ( ~n5146 & n6177 ) ;
  assign n7404 = n7403 ^ n2373 ^ n2364 ;
  assign n7405 = n7404 ^ n5769 ^ n2003 ;
  assign n7406 = n1692 & ~n5840 ;
  assign n7407 = ( n646 & n6478 ) | ( n646 & ~n7406 ) | ( n6478 & ~n7406 ) ;
  assign n7408 = n1888 & n7407 ;
  assign n7409 = n7408 ^ n1310 ^ 1'b0 ;
  assign n7410 = ~n1068 & n5230 ;
  assign n7411 = n7410 ^ n4293 ^ n1727 ;
  assign n7412 = ( n317 & n6658 ) | ( n317 & ~n7411 ) | ( n6658 & ~n7411 ) ;
  assign n7413 = n5864 & n7288 ;
  assign n7414 = n5800 ^ x69 ^ 1'b0 ;
  assign n7415 = n4223 | n7414 ;
  assign n7416 = n4239 ^ n1861 ^ 1'b0 ;
  assign n7417 = ~n7415 & n7416 ;
  assign n7418 = n7417 ^ n7082 ^ n5686 ;
  assign n7419 = ( n1739 & ~n5788 ) | ( n1739 & n7055 ) | ( ~n5788 & n7055 ) ;
  assign n7424 = n1693 ^ n1003 ^ 1'b0 ;
  assign n7420 = n1183 & ~n3517 ;
  assign n7421 = n7420 ^ n2367 ^ 1'b0 ;
  assign n7422 = ~n1683 & n7421 ;
  assign n7423 = ~n6720 & n7422 ;
  assign n7425 = n7424 ^ n7423 ^ n5344 ;
  assign n7426 = n7197 ^ n6478 ^ n4772 ;
  assign n7427 = n6987 ^ n2246 ^ n1050 ;
  assign n7428 = n2486 & n7427 ;
  assign n7429 = n7428 ^ n1412 ^ 1'b0 ;
  assign n7430 = n4745 | n7429 ;
  assign n7431 = n6420 ^ n5166 ^ n761 ;
  assign n7432 = n4044 ^ n3955 ^ n3774 ;
  assign n7433 = n7432 ^ n3934 ^ n3648 ;
  assign n7434 = ~n1219 & n5509 ;
  assign n7435 = ( ~n1794 & n4028 ) | ( ~n1794 & n5163 ) | ( n4028 & n5163 ) ;
  assign n7436 = n7435 ^ n2874 ^ x182 ;
  assign n7437 = ~n3550 & n7436 ;
  assign n7438 = n7437 ^ n3465 ^ 1'b0 ;
  assign n7439 = n7434 & n7438 ;
  assign n7444 = ~n562 & n3660 ;
  assign n7445 = n7444 ^ n910 ^ 1'b0 ;
  assign n7440 = n679 & ~n1856 ;
  assign n7441 = n2391 | n7440 ;
  assign n7442 = n7441 ^ n4672 ^ 1'b0 ;
  assign n7443 = n1773 | n7442 ;
  assign n7446 = n7445 ^ n7443 ^ n3629 ;
  assign n7447 = ( n2201 & n6652 ) | ( n2201 & ~n7446 ) | ( n6652 & ~n7446 ) ;
  assign n7461 = ~x203 & n4674 ;
  assign n7453 = ( n826 & ~n3624 ) | ( n826 & n5267 ) | ( ~n3624 & n5267 ) ;
  assign n7448 = n3311 ^ n2163 ^ 1'b0 ;
  assign n7449 = ( n521 & ~n1699 ) | ( n521 & n5249 ) | ( ~n1699 & n5249 ) ;
  assign n7450 = n7449 ^ n5198 ^ n1382 ;
  assign n7451 = n7450 ^ n1190 ^ 1'b0 ;
  assign n7452 = n7448 & ~n7451 ;
  assign n7454 = n7453 ^ n7452 ^ n1145 ;
  assign n7456 = n5317 | n6407 ;
  assign n7457 = n7456 ^ n7203 ^ n6448 ;
  assign n7455 = n3844 & n6731 ;
  assign n7458 = n7457 ^ n7455 ^ 1'b0 ;
  assign n7459 = n7458 ^ n7452 ^ n1884 ;
  assign n7460 = n7454 | n7459 ;
  assign n7462 = n7461 ^ n7460 ^ 1'b0 ;
  assign n7466 = ( n784 & n1570 ) | ( n784 & ~n4294 ) | ( n1570 & ~n4294 ) ;
  assign n7463 = n2986 ^ n1198 ^ 1'b0 ;
  assign n7464 = ( n2172 & n2526 ) | ( n2172 & ~n7463 ) | ( n2526 & ~n7463 ) ;
  assign n7465 = n2100 & n7464 ;
  assign n7467 = n7466 ^ n7465 ^ 1'b0 ;
  assign n7468 = n6797 & n7467 ;
  assign n7469 = n4386 ^ n3130 ^ n2490 ;
  assign n7470 = n1628 ^ n1551 ^ n497 ;
  assign n7471 = n2207 | n5515 ;
  assign n7472 = ( n5901 & ~n7470 ) | ( n5901 & n7471 ) | ( ~n7470 & n7471 ) ;
  assign n7473 = n2539 ^ n1468 ^ x251 ;
  assign n7475 = n6268 ^ n3504 ^ 1'b0 ;
  assign n7476 = n7131 ^ n5873 ^ 1'b0 ;
  assign n7477 = x188 & ~n7476 ;
  assign n7478 = n3154 ^ n1073 ^ 1'b0 ;
  assign n7479 = ( n7475 & n7477 ) | ( n7475 & n7478 ) | ( n7477 & n7478 ) ;
  assign n7474 = ( ~n2671 & n6046 ) | ( ~n2671 & n6472 ) | ( n6046 & n6472 ) ;
  assign n7480 = n7479 ^ n7474 ^ n6917 ;
  assign n7481 = n3210 ^ n2311 ^ 1'b0 ;
  assign n7482 = n3503 | n7481 ;
  assign n7483 = n2042 ^ n1476 ^ n327 ;
  assign n7484 = ~n7482 & n7483 ;
  assign n7485 = ~x204 & n7484 ;
  assign n7486 = n1595 & ~n5697 ;
  assign n7487 = ( ~x151 & n1298 ) | ( ~x151 & n5812 ) | ( n1298 & n5812 ) ;
  assign n7488 = n672 | n7487 ;
  assign n7489 = n7486 | n7488 ;
  assign n7490 = ( ~n325 & n1457 ) | ( ~n325 & n1953 ) | ( n1457 & n1953 ) ;
  assign n7491 = ( x127 & n1580 ) | ( x127 & n2588 ) | ( n1580 & n2588 ) ;
  assign n7492 = n4137 ^ n647 ^ 1'b0 ;
  assign n7493 = n7492 ^ n4744 ^ n2701 ;
  assign n7494 = ( n7490 & n7491 ) | ( n7490 & n7493 ) | ( n7491 & n7493 ) ;
  assign n7495 = n550 | n2681 ;
  assign n7496 = n7495 ^ n2257 ^ 1'b0 ;
  assign n7497 = ( n538 & ~n1355 ) | ( n538 & n4705 ) | ( ~n1355 & n4705 ) ;
  assign n7498 = n7497 ^ n1253 ^ 1'b0 ;
  assign n7499 = n7498 ^ n3198 ^ 1'b0 ;
  assign n7500 = n7496 & ~n7499 ;
  assign n7501 = ~n3028 & n6073 ;
  assign n7502 = n7501 ^ n6135 ^ 1'b0 ;
  assign n7503 = n7106 ^ n977 ^ 1'b0 ;
  assign n7504 = n1845 & ~n7503 ;
  assign n7505 = n2451 & n2936 ;
  assign n7506 = n920 & n7505 ;
  assign n7507 = n4735 ^ n4710 ^ n4122 ;
  assign n7509 = n6213 ^ x145 ^ 1'b0 ;
  assign n7508 = ~n2816 & n7448 ;
  assign n7510 = n7509 ^ n7508 ^ 1'b0 ;
  assign n7511 = ( ~n3535 & n7507 ) | ( ~n3535 & n7510 ) | ( n7507 & n7510 ) ;
  assign n7512 = n7511 ^ n2722 ^ 1'b0 ;
  assign n7513 = n2927 & n7512 ;
  assign n7514 = ( n2450 & n7506 ) | ( n2450 & n7513 ) | ( n7506 & n7513 ) ;
  assign n7515 = n327 | n7108 ;
  assign n7516 = n1516 | n7515 ;
  assign n7517 = n7516 ^ n6443 ^ 1'b0 ;
  assign n7518 = n763 & n4660 ;
  assign n7519 = n6607 & n7518 ;
  assign n7520 = n7519 ^ n4467 ^ 1'b0 ;
  assign n7521 = n3069 & ~n6435 ;
  assign n7522 = n7521 ^ n6424 ^ 1'b0 ;
  assign n7523 = n5739 | n7522 ;
  assign n7524 = n3616 ^ n1313 ^ 1'b0 ;
  assign n7525 = n4897 & n7524 ;
  assign n7526 = n7525 ^ n257 ^ 1'b0 ;
  assign n7527 = n6291 & n7526 ;
  assign n7528 = n3838 & n7527 ;
  assign n7529 = n5657 | n7403 ;
  assign n7530 = n4153 ^ n1912 ^ 1'b0 ;
  assign n7531 = ~n3956 & n7530 ;
  assign n7532 = n7531 ^ n5214 ^ 1'b0 ;
  assign n7533 = n4926 & ~n7532 ;
  assign n7534 = n3323 ^ n2208 ^ n2190 ;
  assign n7535 = n7534 ^ n7463 ^ n2386 ;
  assign n7539 = n6248 ^ n5707 ^ n3154 ;
  assign n7536 = ( n2290 & ~n3547 ) | ( n2290 & n5568 ) | ( ~n3547 & n5568 ) ;
  assign n7537 = n257 | n7536 ;
  assign n7538 = n7211 | n7537 ;
  assign n7540 = n7539 ^ n7538 ^ 1'b0 ;
  assign n7541 = ( n1279 & ~n1367 ) | ( n1279 & n2673 ) | ( ~n1367 & n2673 ) ;
  assign n7542 = ( n541 & ~n4268 ) | ( n541 & n6270 ) | ( ~n4268 & n6270 ) ;
  assign n7543 = n1331 | n7542 ;
  assign n7544 = ( n3939 & ~n7541 ) | ( n3939 & n7543 ) | ( ~n7541 & n7543 ) ;
  assign n7546 = n5545 ^ n436 ^ 1'b0 ;
  assign n7545 = ~n2967 & n4625 ;
  assign n7547 = n7546 ^ n7545 ^ 1'b0 ;
  assign n7548 = ( n3099 & ~n3342 ) | ( n3099 & n5039 ) | ( ~n3342 & n5039 ) ;
  assign n7549 = ( n640 & ~n7314 ) | ( n640 & n7548 ) | ( ~n7314 & n7548 ) ;
  assign n7550 = n3790 ^ n329 ^ x57 ;
  assign n7552 = x188 & ~n5041 ;
  assign n7553 = n7552 ^ n436 ^ 1'b0 ;
  assign n7554 = n7553 ^ n2981 ^ n2267 ;
  assign n7555 = x53 & n7554 ;
  assign n7556 = n7555 ^ n317 ^ 1'b0 ;
  assign n7551 = n5733 ^ n2723 ^ n1900 ;
  assign n7557 = n7556 ^ n7551 ^ 1'b0 ;
  assign n7558 = ( n6348 & ~n7550 ) | ( n6348 & n7557 ) | ( ~n7550 & n7557 ) ;
  assign n7559 = n7558 ^ n4420 ^ n962 ;
  assign n7560 = n3794 & ~n4315 ;
  assign n7561 = ( ~x107 & n2149 ) | ( ~x107 & n7560 ) | ( n2149 & n7560 ) ;
  assign n7562 = n7561 ^ n6802 ^ 1'b0 ;
  assign n7563 = n2467 ^ n901 ^ n483 ;
  assign n7564 = n3198 & ~n7563 ;
  assign n7565 = ~n3324 & n7564 ;
  assign n7566 = n7565 ^ n3218 ^ n1673 ;
  assign n7567 = ( ~n1111 & n3254 ) | ( ~n1111 & n5484 ) | ( n3254 & n5484 ) ;
  assign n7570 = n7013 ^ n3490 ^ 1'b0 ;
  assign n7571 = n3779 | n7570 ;
  assign n7568 = n5672 ^ n1451 ^ 1'b0 ;
  assign n7569 = ( ~x82 & n1052 ) | ( ~x82 & n7568 ) | ( n1052 & n7568 ) ;
  assign n7572 = n7571 ^ n7569 ^ n5508 ;
  assign n7573 = ( n2627 & ~n3179 ) | ( n2627 & n4395 ) | ( ~n3179 & n4395 ) ;
  assign n7574 = ( ~n5897 & n7572 ) | ( ~n5897 & n7573 ) | ( n7572 & n7573 ) ;
  assign n7575 = n7567 | n7574 ;
  assign n7576 = n3267 & ~n7575 ;
  assign n7577 = n6678 ^ n5224 ^ 1'b0 ;
  assign n7578 = n2346 ^ n1771 ^ 1'b0 ;
  assign n7579 = ( n967 & n3879 ) | ( n967 & n6714 ) | ( n3879 & n6714 ) ;
  assign n7580 = ( n3659 & n7578 ) | ( n3659 & ~n7579 ) | ( n7578 & ~n7579 ) ;
  assign n7581 = ( n2107 & ~n5040 ) | ( n2107 & n6596 ) | ( ~n5040 & n6596 ) ;
  assign n7584 = n7097 ^ n3458 ^ 1'b0 ;
  assign n7585 = n5454 & n7584 ;
  assign n7582 = n2229 ^ n1743 ^ n311 ;
  assign n7583 = ~n4581 & n7582 ;
  assign n7586 = n7585 ^ n7583 ^ n2970 ;
  assign n7587 = n3491 | n7376 ;
  assign n7591 = n3905 & n5412 ;
  assign n7588 = n3317 & ~n3355 ;
  assign n7589 = n6287 | n7588 ;
  assign n7590 = n4445 | n7589 ;
  assign n7592 = n7591 ^ n7590 ^ n3747 ;
  assign n7593 = n7592 ^ n4349 ^ n3783 ;
  assign n7596 = x3 & n3567 ;
  assign n7594 = n4421 ^ n1550 ^ 1'b0 ;
  assign n7595 = n5554 & ~n7594 ;
  assign n7597 = n7596 ^ n7595 ^ n3801 ;
  assign n7598 = n1340 | n5128 ;
  assign n7599 = n7598 ^ n3759 ^ 1'b0 ;
  assign n7600 = ~n7597 & n7599 ;
  assign n7601 = n690 & n4272 ;
  assign n7602 = ( ~n1043 & n3515 ) | ( ~n1043 & n6036 ) | ( n3515 & n6036 ) ;
  assign n7603 = n7602 ^ n4593 ^ 1'b0 ;
  assign n7604 = n7603 ^ n4615 ^ 1'b0 ;
  assign n7605 = n4722 ^ n1310 ^ n1239 ;
  assign n7606 = ~n2695 & n7605 ;
  assign n7607 = n7606 ^ n5809 ^ n2734 ;
  assign n7608 = n7607 ^ n5361 ^ n708 ;
  assign n7621 = ( n864 & ~n4885 ) | ( n864 & n5508 ) | ( ~n4885 & n5508 ) ;
  assign n7609 = ( n3075 & n3257 ) | ( n3075 & n3744 ) | ( n3257 & n3744 ) ;
  assign n7610 = n2182 ^ n386 ^ 1'b0 ;
  assign n7611 = n3258 & n7610 ;
  assign n7612 = ( x198 & x230 ) | ( x198 & ~n755 ) | ( x230 & ~n755 ) ;
  assign n7613 = ~n3517 & n7612 ;
  assign n7614 = n7613 ^ n3066 ^ 1'b0 ;
  assign n7615 = n5111 | n7614 ;
  assign n7616 = n7611 & ~n7615 ;
  assign n7617 = n2228 | n7616 ;
  assign n7618 = n7609 & ~n7617 ;
  assign n7619 = n948 & ~n7618 ;
  assign n7620 = ~n6828 & n7619 ;
  assign n7622 = n7621 ^ n7620 ^ n3579 ;
  assign n7623 = ( n393 & n1005 ) | ( n393 & n1382 ) | ( n1005 & n1382 ) ;
  assign n7625 = n3494 ^ n840 ^ n393 ;
  assign n7624 = ~n7185 & n7593 ;
  assign n7626 = n7625 ^ n7624 ^ 1'b0 ;
  assign n7627 = n7114 ^ n4873 ^ n4346 ;
  assign n7628 = ( n4216 & n5549 ) | ( n4216 & n5662 ) | ( n5549 & n5662 ) ;
  assign n7629 = ~n7627 & n7628 ;
  assign n7630 = ( n1768 & n2691 ) | ( n1768 & n2922 ) | ( n2691 & n2922 ) ;
  assign n7631 = n6097 ^ n1502 ^ 1'b0 ;
  assign n7632 = ~n7630 & n7631 ;
  assign n7636 = ( x40 & ~x218 ) | ( x40 & n1474 ) | ( ~x218 & n1474 ) ;
  assign n7635 = n1478 & n5284 ;
  assign n7637 = n7636 ^ n7635 ^ 1'b0 ;
  assign n7638 = n7637 ^ n5125 ^ 1'b0 ;
  assign n7633 = n4014 & n4351 ;
  assign n7634 = n797 | n7633 ;
  assign n7639 = n7638 ^ n7634 ^ n509 ;
  assign n7646 = n3775 & ~n4703 ;
  assign n7640 = ~n3382 & n7111 ;
  assign n7641 = n7640 ^ n6559 ^ n4015 ;
  assign n7642 = ( x174 & n2926 ) | ( x174 & ~n4710 ) | ( n2926 & ~n4710 ) ;
  assign n7643 = n4507 & ~n7642 ;
  assign n7644 = n7643 ^ n4950 ^ 1'b0 ;
  assign n7645 = ( n788 & ~n7641 ) | ( n788 & n7644 ) | ( ~n7641 & n7644 ) ;
  assign n7647 = n7646 ^ n7645 ^ 1'b0 ;
  assign n7648 = x161 & ~n7647 ;
  assign n7649 = n4366 ^ n2100 ^ 1'b0 ;
  assign n7650 = n5643 & ~n7649 ;
  assign n7651 = ~n2635 & n7650 ;
  assign n7652 = n1862 & ~n5772 ;
  assign n7653 = n981 & ~n4327 ;
  assign n7654 = ( n462 & n2121 ) | ( n462 & n7653 ) | ( n2121 & n7653 ) ;
  assign n7655 = ( x110 & ~n739 ) | ( x110 & n2438 ) | ( ~n739 & n2438 ) ;
  assign n7660 = n4989 ^ n3636 ^ 1'b0 ;
  assign n7656 = n2210 & ~n2984 ;
  assign n7657 = ~x182 & n7656 ;
  assign n7658 = ( n897 & ~n1129 ) | ( n897 & n7657 ) | ( ~n1129 & n7657 ) ;
  assign n7659 = n1308 | n7658 ;
  assign n7661 = n7660 ^ n7659 ^ n362 ;
  assign n7662 = ( ~n7295 & n7655 ) | ( ~n7295 & n7661 ) | ( n7655 & n7661 ) ;
  assign n7663 = ~n733 & n5624 ;
  assign n7664 = ( n1424 & ~n5515 ) | ( n1424 & n7663 ) | ( ~n5515 & n7663 ) ;
  assign n7665 = n4948 ^ n1758 ^ x190 ;
  assign n7666 = ~n308 & n7665 ;
  assign n7667 = n7664 & n7666 ;
  assign n7668 = n905 & ~n6237 ;
  assign n7669 = n2990 ^ n2392 ^ n696 ;
  assign n7670 = n7669 ^ n1173 ^ n596 ;
  assign n7671 = ( x72 & ~n3070 ) | ( x72 & n3128 ) | ( ~n3070 & n3128 ) ;
  assign n7672 = n7671 ^ n3219 ^ n1874 ;
  assign n7673 = n2360 ^ n492 ^ 1'b0 ;
  assign n7674 = ~n872 & n7673 ;
  assign n7675 = n7674 ^ n5307 ^ n824 ;
  assign n7676 = ( n7670 & n7672 ) | ( n7670 & ~n7675 ) | ( n7672 & ~n7675 ) ;
  assign n7677 = n2571 & ~n7676 ;
  assign n7678 = ( n1407 & n7668 ) | ( n1407 & ~n7677 ) | ( n7668 & ~n7677 ) ;
  assign n7679 = n1494 & ~n4387 ;
  assign n7680 = ( n410 & ~n3535 ) | ( n410 & n7679 ) | ( ~n3535 & n7679 ) ;
  assign n7681 = ( n2936 & ~n4815 ) | ( n2936 & n7680 ) | ( ~n4815 & n7680 ) ;
  assign n7682 = n7681 ^ n2286 ^ 1'b0 ;
  assign n7683 = n353 & ~n1396 ;
  assign n7684 = n7683 ^ x186 ^ 1'b0 ;
  assign n7685 = n1451 & n3377 ;
  assign n7686 = n7685 ^ n4613 ^ n510 ;
  assign n7687 = ~n1800 & n3078 ;
  assign n7688 = ~n282 & n7687 ;
  assign n7689 = x85 | n7688 ;
  assign n7690 = ~n3640 & n7689 ;
  assign n7691 = n6590 ^ n808 ^ 1'b0 ;
  assign n7692 = n903 | n7691 ;
  assign n7693 = n3122 | n7692 ;
  assign n7694 = n7693 ^ n1007 ^ n712 ;
  assign n7702 = n4222 & n6078 ;
  assign n7695 = n3152 ^ n1776 ^ n1652 ;
  assign n7696 = n5545 ^ n3604 ^ 1'b0 ;
  assign n7697 = ( n1400 & n7695 ) | ( n1400 & n7696 ) | ( n7695 & n7696 ) ;
  assign n7698 = n2059 ^ n1644 ^ n1156 ;
  assign n7699 = n7698 ^ n5823 ^ n4265 ;
  assign n7700 = n7699 ^ n3965 ^ n1270 ;
  assign n7701 = n7697 & ~n7700 ;
  assign n7703 = n7702 ^ n7701 ^ 1'b0 ;
  assign n7707 = n1821 ^ n459 ^ 1'b0 ;
  assign n7706 = n5168 ^ n331 ^ 1'b0 ;
  assign n7704 = ~n520 & n2780 ;
  assign n7705 = ( n4625 & ~n6987 ) | ( n4625 & n7704 ) | ( ~n6987 & n7704 ) ;
  assign n7708 = n7707 ^ n7706 ^ n7705 ;
  assign n7709 = n4802 ^ n3530 ^ n2545 ;
  assign n7710 = ( n723 & n1040 ) | ( n723 & ~n7709 ) | ( n1040 & ~n7709 ) ;
  assign n7711 = n7710 ^ n753 ^ 1'b0 ;
  assign n7712 = n7708 & ~n7711 ;
  assign n7713 = ~n5386 & n6649 ;
  assign n7714 = n7713 ^ n6498 ^ 1'b0 ;
  assign n7715 = n7714 ^ n2885 ^ 1'b0 ;
  assign n7716 = n2187 ^ x2 ^ 1'b0 ;
  assign n7717 = n5536 ^ n3674 ^ 1'b0 ;
  assign n7718 = n655 | n7717 ;
  assign n7719 = n3116 ^ n407 ^ x236 ;
  assign n7720 = n7719 ^ n4070 ^ 1'b0 ;
  assign n7721 = n7718 | n7720 ;
  assign n7722 = ( n3499 & n3853 ) | ( n3499 & n6648 ) | ( n3853 & n6648 ) ;
  assign n7723 = ( n1935 & n4208 ) | ( n1935 & ~n6630 ) | ( n4208 & ~n6630 ) ;
  assign n7724 = n630 | n7723 ;
  assign n7725 = n7724 ^ n3114 ^ 1'b0 ;
  assign n7726 = n1684 ^ n1199 ^ 1'b0 ;
  assign n7727 = ( ~n640 & n6459 ) | ( ~n640 & n7061 ) | ( n6459 & n7061 ) ;
  assign n7728 = n7727 ^ n3560 ^ 1'b0 ;
  assign n7729 = n3627 & ~n7728 ;
  assign n7730 = n7729 ^ n4671 ^ 1'b0 ;
  assign n7731 = ~n5242 & n7730 ;
  assign n7732 = n7726 | n7731 ;
  assign n7733 = n7725 & ~n7732 ;
  assign n7734 = n7733 ^ n6520 ^ 1'b0 ;
  assign n7735 = ( ~n7721 & n7722 ) | ( ~n7721 & n7734 ) | ( n7722 & n7734 ) ;
  assign n7736 = x233 | n2086 ;
  assign n7737 = ( ~x242 & n2371 ) | ( ~x242 & n7736 ) | ( n2371 & n7736 ) ;
  assign n7738 = n7737 ^ n5424 ^ 1'b0 ;
  assign n7739 = n3991 ^ n3279 ^ n536 ;
  assign n7740 = n3128 | n7739 ;
  assign n7741 = n866 | n7740 ;
  assign n7742 = n3891 ^ n268 ^ 1'b0 ;
  assign n7743 = n1810 & n7742 ;
  assign n7744 = ~n7741 & n7743 ;
  assign n7761 = ~n394 & n5392 ;
  assign n7762 = n7761 ^ n4359 ^ 1'b0 ;
  assign n7763 = n4547 & n7762 ;
  assign n7745 = n1361 ^ n345 ^ 1'b0 ;
  assign n7746 = n5929 & ~n7745 ;
  assign n7747 = n5268 ^ n2250 ^ 1'b0 ;
  assign n7748 = n2273 | n7747 ;
  assign n7755 = x43 & n6338 ;
  assign n7756 = ~n1649 & n7755 ;
  assign n7757 = n7756 ^ n3202 ^ 1'b0 ;
  assign n7749 = x170 & ~n966 ;
  assign n7750 = n7749 ^ n491 ^ 1'b0 ;
  assign n7751 = n4360 ^ n2640 ^ 1'b0 ;
  assign n7752 = ~n807 & n7751 ;
  assign n7753 = n7752 ^ n7003 ^ n4038 ;
  assign n7754 = ( ~n4582 & n7750 ) | ( ~n4582 & n7753 ) | ( n7750 & n7753 ) ;
  assign n7758 = n7757 ^ n7754 ^ n1651 ;
  assign n7759 = ( n7746 & n7748 ) | ( n7746 & n7758 ) | ( n7748 & n7758 ) ;
  assign n7760 = ~n7266 & n7759 ;
  assign n7764 = n7763 ^ n7760 ^ 1'b0 ;
  assign n7765 = n439 & ~n7466 ;
  assign n7766 = n5115 & n7765 ;
  assign n7767 = n2533 & ~n7766 ;
  assign n7768 = n7767 ^ n4998 ^ 1'b0 ;
  assign n7769 = n3353 | n7768 ;
  assign n7770 = ~n293 & n933 ;
  assign n7771 = n7770 ^ n3701 ^ 1'b0 ;
  assign n7772 = n4863 ^ n1036 ^ 1'b0 ;
  assign n7773 = n4943 | n7772 ;
  assign n7774 = n7773 ^ n3335 ^ 1'b0 ;
  assign n7775 = n7774 ^ n4782 ^ 1'b0 ;
  assign n7776 = n7771 & ~n7775 ;
  assign n7777 = n1140 & n2285 ;
  assign n7778 = n7777 ^ x206 ^ 1'b0 ;
  assign n7779 = n7778 ^ n401 ^ 1'b0 ;
  assign n7780 = n4363 & ~n7779 ;
  assign n7781 = ~n2217 & n2401 ;
  assign n7782 = n4176 & n7781 ;
  assign n7783 = ( n1617 & ~n4173 ) | ( n1617 & n7782 ) | ( ~n4173 & n7782 ) ;
  assign n7784 = ( n2500 & n4556 ) | ( n2500 & ~n7783 ) | ( n4556 & ~n7783 ) ;
  assign n7785 = n7784 ^ n2633 ^ 1'b0 ;
  assign n7786 = n7780 | n7785 ;
  assign n7787 = n1087 & n4813 ;
  assign n7788 = n4137 & n7787 ;
  assign n7789 = ( ~n1373 & n3087 ) | ( ~n1373 & n5683 ) | ( n3087 & n5683 ) ;
  assign n7790 = n7789 ^ n6753 ^ n3190 ;
  assign n7791 = ( ~n1526 & n5314 ) | ( ~n1526 & n7790 ) | ( n5314 & n7790 ) ;
  assign n7792 = ( n7080 & ~n7788 ) | ( n7080 & n7791 ) | ( ~n7788 & n7791 ) ;
  assign n7793 = ( n418 & n2594 ) | ( n418 & n3309 ) | ( n2594 & n3309 ) ;
  assign n7796 = n3367 ^ n1314 ^ n689 ;
  assign n7797 = n5114 & ~n7796 ;
  assign n7794 = ~x148 & n6720 ;
  assign n7795 = ( n5097 & ~n5557 ) | ( n5097 & n7794 ) | ( ~n5557 & n7794 ) ;
  assign n7798 = n7797 ^ n7795 ^ n3655 ;
  assign n7799 = ( n3730 & n4802 ) | ( n3730 & n5536 ) | ( n4802 & n5536 ) ;
  assign n7800 = n2668 ^ n2527 ^ x238 ;
  assign n7801 = n6307 ^ n5357 ^ n1610 ;
  assign n7802 = ~n765 & n4405 ;
  assign n7803 = ~n7243 & n7802 ;
  assign n7807 = ~n681 & n3775 ;
  assign n7808 = n7807 ^ n4359 ^ 1'b0 ;
  assign n7809 = n7808 ^ n6918 ^ n4563 ;
  assign n7804 = n2714 ^ n2494 ^ 1'b0 ;
  assign n7805 = ~n2923 & n7804 ;
  assign n7806 = ( n1330 & ~n4816 ) | ( n1330 & n7805 ) | ( ~n4816 & n7805 ) ;
  assign n7810 = n7809 ^ n7806 ^ n1760 ;
  assign n7811 = n7810 ^ n5133 ^ n4664 ;
  assign n7815 = n7595 ^ n7096 ^ n3188 ;
  assign n7812 = n5643 ^ n3620 ^ n903 ;
  assign n7813 = n4777 & ~n7812 ;
  assign n7814 = ~n1652 & n7813 ;
  assign n7816 = n7815 ^ n7814 ^ 1'b0 ;
  assign n7817 = n6977 & n7816 ;
  assign n7818 = n3922 ^ n1943 ^ x176 ;
  assign n7819 = ( n5236 & n6420 ) | ( n5236 & ~n7818 ) | ( n6420 & ~n7818 ) ;
  assign n7828 = ( n434 & n1894 ) | ( n434 & n4230 ) | ( n1894 & n4230 ) ;
  assign n7829 = ( ~n4999 & n5234 ) | ( ~n4999 & n7828 ) | ( n5234 & n7828 ) ;
  assign n7820 = ~n2354 & n2701 ;
  assign n7821 = ( ~n2401 & n4692 ) | ( ~n2401 & n7820 ) | ( n4692 & n7820 ) ;
  assign n7822 = ~n2049 & n2373 ;
  assign n7823 = n4694 ^ n1985 ^ 1'b0 ;
  assign n7824 = ~n3706 & n7823 ;
  assign n7825 = n7824 ^ n6294 ^ 1'b0 ;
  assign n7826 = n7822 | n7825 ;
  assign n7827 = n7821 & ~n7826 ;
  assign n7830 = n7829 ^ n7827 ^ 1'b0 ;
  assign n7831 = n5385 ^ n3169 ^ 1'b0 ;
  assign n7832 = n7042 & n7831 ;
  assign n7833 = n7832 ^ n4724 ^ n3229 ;
  assign n7834 = n6370 ^ n6301 ^ n5283 ;
  assign n7835 = ( n1970 & n6483 ) | ( n1970 & n7834 ) | ( n6483 & n7834 ) ;
  assign n7836 = ( n896 & ~n2814 ) | ( n896 & n4020 ) | ( ~n2814 & n4020 ) ;
  assign n7837 = n7836 ^ n7152 ^ n6589 ;
  assign n7838 = n7470 ^ n4230 ^ n1816 ;
  assign n7839 = n1872 & ~n4075 ;
  assign n7840 = ( ~n6723 & n7838 ) | ( ~n6723 & n7839 ) | ( n7838 & n7839 ) ;
  assign n7845 = ( x225 & n1880 ) | ( x225 & ~n3489 ) | ( n1880 & ~n3489 ) ;
  assign n7846 = n7539 & n7845 ;
  assign n7842 = n3339 ^ n2513 ^ n1975 ;
  assign n7843 = ( n905 & n7317 ) | ( n905 & ~n7842 ) | ( n7317 & ~n7842 ) ;
  assign n7841 = ~n556 & n3269 ;
  assign n7844 = n7843 ^ n7841 ^ 1'b0 ;
  assign n7847 = n7846 ^ n7844 ^ n6945 ;
  assign n7848 = n4251 & n6882 ;
  assign n7849 = ~n7442 & n7848 ;
  assign n7850 = n2918 ^ n2097 ^ 1'b0 ;
  assign n7851 = n1892 ^ n1103 ^ x81 ;
  assign n7852 = n3829 ^ n1152 ^ 1'b0 ;
  assign n7853 = n7851 | n7852 ;
  assign n7854 = ( n3342 & n4438 ) | ( n3342 & n6585 ) | ( n4438 & n6585 ) ;
  assign n7855 = n7854 ^ n5013 ^ n438 ;
  assign n7856 = ( ~n690 & n7853 ) | ( ~n690 & n7855 ) | ( n7853 & n7855 ) ;
  assign n7857 = n3445 ^ n3200 ^ n410 ;
  assign n7858 = n5524 ^ n2603 ^ n300 ;
  assign n7859 = n6631 ^ n6540 ^ n3437 ;
  assign n7860 = n5380 ^ n2064 ^ n679 ;
  assign n7861 = n2322 & n7860 ;
  assign n7862 = ~n7859 & n7861 ;
  assign n7863 = n4161 & n7862 ;
  assign n7864 = ( n523 & n6755 ) | ( n523 & n7144 ) | ( n6755 & n7144 ) ;
  assign n7865 = n1998 & ~n3320 ;
  assign n7873 = n3013 ^ n1928 ^ n843 ;
  assign n7866 = x46 & ~n7772 ;
  assign n7867 = n7866 ^ n4747 ^ 1'b0 ;
  assign n7868 = n1655 ^ n896 ^ 1'b0 ;
  assign n7869 = n7659 & ~n7836 ;
  assign n7870 = n7868 & n7869 ;
  assign n7871 = n7870 ^ n3394 ^ 1'b0 ;
  assign n7872 = n7867 & n7871 ;
  assign n7874 = n7873 ^ n7872 ^ 1'b0 ;
  assign n7875 = n4884 | n5557 ;
  assign n7876 = n7746 & ~n7875 ;
  assign n7878 = n4735 ^ n4486 ^ x226 ;
  assign n7877 = n2837 ^ n1538 ^ n685 ;
  assign n7879 = n7878 ^ n7877 ^ 1'b0 ;
  assign n7880 = ( n684 & ~n4989 ) | ( n684 & n6548 ) | ( ~n4989 & n6548 ) ;
  assign n7881 = ( x101 & n3550 ) | ( x101 & ~n7880 ) | ( n3550 & ~n7880 ) ;
  assign n7882 = n7881 ^ n5163 ^ 1'b0 ;
  assign n7883 = n961 & ~n4119 ;
  assign n7884 = n7883 ^ n2469 ^ 1'b0 ;
  assign n7885 = ( n687 & n7602 ) | ( n687 & ~n7884 ) | ( n7602 & ~n7884 ) ;
  assign n7886 = n746 & ~n1355 ;
  assign n7887 = n3707 & n6437 ;
  assign n7888 = n5443 | n7887 ;
  assign n7889 = n6338 ^ x56 ^ 1'b0 ;
  assign n7890 = n3206 & n7889 ;
  assign n7892 = n6817 ^ n5854 ^ n1189 ;
  assign n7893 = n7892 ^ n4788 ^ 1'b0 ;
  assign n7894 = n4956 | n7893 ;
  assign n7895 = ( n4453 & n5868 ) | ( n4453 & n7894 ) | ( n5868 & n7894 ) ;
  assign n7896 = n7895 ^ n7584 ^ 1'b0 ;
  assign n7891 = n5929 ^ n3947 ^ 1'b0 ;
  assign n7897 = n7896 ^ n7891 ^ n4500 ;
  assign n7899 = n898 ^ n896 ^ 1'b0 ;
  assign n7900 = n7899 ^ n3466 ^ n1765 ;
  assign n7901 = ( ~n322 & n3484 ) | ( ~n322 & n7900 ) | ( n3484 & n7900 ) ;
  assign n7898 = x14 & ~n2464 ;
  assign n7902 = n7901 ^ n7898 ^ 1'b0 ;
  assign n7903 = n1918 | n7902 ;
  assign n7904 = ( ~x51 & n5787 ) | ( ~x51 & n7903 ) | ( n5787 & n7903 ) ;
  assign n7905 = n6246 ^ n854 ^ 1'b0 ;
  assign n7906 = n7905 ^ n7159 ^ 1'b0 ;
  assign n7907 = n7906 ^ n7447 ^ n4344 ;
  assign n7908 = n6355 ^ n3666 ^ 1'b0 ;
  assign n7912 = n5608 ^ n2565 ^ x126 ;
  assign n7909 = n4745 ^ n1732 ^ 1'b0 ;
  assign n7910 = n2503 | n7909 ;
  assign n7911 = n3236 | n7910 ;
  assign n7913 = n7912 ^ n7911 ^ n6562 ;
  assign n7914 = ( ~n6602 & n7908 ) | ( ~n6602 & n7913 ) | ( n7908 & n7913 ) ;
  assign n7915 = ( ~n1255 & n2142 ) | ( ~n1255 & n5145 ) | ( n2142 & n5145 ) ;
  assign n7916 = n2338 ^ n2035 ^ 1'b0 ;
  assign n7917 = n6127 & ~n7916 ;
  assign n7918 = n7917 ^ n7685 ^ 1'b0 ;
  assign n7919 = ~n7915 & n7918 ;
  assign n7920 = ~n351 & n2979 ;
  assign n7921 = n7920 ^ n6374 ^ 1'b0 ;
  assign n7922 = x29 & ~n7921 ;
  assign n7923 = ~n7342 & n7922 ;
  assign n7935 = ( n1720 & n2497 ) | ( n1720 & n2657 ) | ( n2497 & n2657 ) ;
  assign n7931 = ( ~n595 & n7085 ) | ( ~n595 & n7098 ) | ( n7085 & n7098 ) ;
  assign n7926 = ( n1162 & n3199 ) | ( n1162 & ~n5576 ) | ( n3199 & ~n5576 ) ;
  assign n7927 = n7926 ^ n7185 ^ n1404 ;
  assign n7924 = n991 ^ n660 ^ n295 ;
  assign n7925 = n471 & n7924 ;
  assign n7928 = n7927 ^ n7925 ^ 1'b0 ;
  assign n7929 = n5082 ^ n2585 ^ 1'b0 ;
  assign n7930 = n7928 & ~n7929 ;
  assign n7932 = n7931 ^ n7930 ^ 1'b0 ;
  assign n7933 = n7932 ^ n5164 ^ 1'b0 ;
  assign n7934 = n1078 & ~n7933 ;
  assign n7936 = n7935 ^ n7934 ^ 1'b0 ;
  assign n7937 = n914 & ~n3208 ;
  assign n7938 = n7937 ^ n1221 ^ 1'b0 ;
  assign n7939 = n7938 ^ n5740 ^ 1'b0 ;
  assign n7940 = ~n6709 & n7939 ;
  assign n7941 = ~n6870 & n7940 ;
  assign n7942 = n7941 ^ n2869 ^ 1'b0 ;
  assign n7943 = n7942 ^ n2029 ^ 1'b0 ;
  assign n7944 = n1629 & n7943 ;
  assign n7945 = n4382 & n7098 ;
  assign n7946 = n7945 ^ n2763 ^ 1'b0 ;
  assign n7947 = ( x11 & n6529 ) | ( x11 & n7946 ) | ( n6529 & n7946 ) ;
  assign n7948 = n1753 & n6504 ;
  assign n7949 = n525 | n7948 ;
  assign n7950 = n7949 ^ n601 ^ 1'b0 ;
  assign n7951 = ~n5115 & n5569 ;
  assign n7952 = ( ~n5071 & n6683 ) | ( ~n5071 & n7951 ) | ( n6683 & n7951 ) ;
  assign n7953 = n1967 & n2480 ;
  assign n7955 = n4917 ^ n2964 ^ 1'b0 ;
  assign n7954 = ( n4421 & n6864 ) | ( n4421 & ~n7698 ) | ( n6864 & ~n7698 ) ;
  assign n7956 = n7955 ^ n7954 ^ n2912 ;
  assign n7958 = n2764 ^ n1122 ^ n701 ;
  assign n7959 = n7958 ^ n2448 ^ 1'b0 ;
  assign n7960 = x194 & n7959 ;
  assign n7961 = ( n1028 & n3515 ) | ( n1028 & ~n7960 ) | ( n3515 & ~n7960 ) ;
  assign n7957 = ( ~n4313 & n5065 ) | ( ~n4313 & n5310 ) | ( n5065 & n5310 ) ;
  assign n7962 = n7961 ^ n7957 ^ 1'b0 ;
  assign n7963 = n342 | n1893 ;
  assign n7964 = n7963 ^ n4010 ^ 1'b0 ;
  assign n7965 = n740 & ~n7964 ;
  assign n7966 = x169 & n7965 ;
  assign n7967 = n5401 ^ n4060 ^ 1'b0 ;
  assign n7968 = ~n7966 & n7967 ;
  assign n7969 = ~n5541 & n7968 ;
  assign n7970 = n7969 ^ x154 ^ 1'b0 ;
  assign n7971 = n6540 ^ n5732 ^ n2306 ;
  assign n7972 = ~n3620 & n7971 ;
  assign n7973 = ( n2266 & n4969 ) | ( n2266 & n5205 ) | ( n4969 & n5205 ) ;
  assign n7974 = n2631 | n7973 ;
  assign n7975 = n688 & ~n2000 ;
  assign n7976 = n7975 ^ n3486 ^ 1'b0 ;
  assign n7977 = ( ~n1914 & n5155 ) | ( ~n1914 & n7976 ) | ( n5155 & n7976 ) ;
  assign n7978 = n7179 ^ n5919 ^ x71 ;
  assign n7983 = n4972 ^ n2034 ^ 1'b0 ;
  assign n7984 = ~n1258 & n7983 ;
  assign n7981 = n2796 ^ x37 ^ 1'b0 ;
  assign n7982 = n6314 & n7981 ;
  assign n7979 = n4065 ^ n287 ^ 1'b0 ;
  assign n7980 = n7979 ^ n1598 ^ 1'b0 ;
  assign n7985 = n7984 ^ n7982 ^ n7980 ;
  assign n7986 = n2695 | n5762 ;
  assign n7987 = n7986 ^ n6527 ^ 1'b0 ;
  assign n7991 = n2544 ^ n1628 ^ n286 ;
  assign n7990 = ( n3449 & n3887 ) | ( n3449 & n4137 ) | ( n3887 & n4137 ) ;
  assign n7988 = n2539 & n2988 ;
  assign n7989 = ( n4300 & n7851 ) | ( n4300 & ~n7988 ) | ( n7851 & ~n7988 ) ;
  assign n7992 = n7991 ^ n7990 ^ n7989 ;
  assign n7993 = n7072 ^ n2205 ^ 1'b0 ;
  assign n7994 = n7218 ^ n5061 ^ 1'b0 ;
  assign n7995 = n6058 | n7994 ;
  assign n8002 = n6752 ^ n5500 ^ n5484 ;
  assign n7996 = n323 & n593 ;
  assign n7997 = n7996 ^ n887 ^ 1'b0 ;
  assign n7998 = ~n563 & n882 ;
  assign n7999 = n7605 & n7998 ;
  assign n8000 = n7999 ^ n3838 ^ 1'b0 ;
  assign n8001 = ~n7997 & n8000 ;
  assign n8003 = n8002 ^ n8001 ^ 1'b0 ;
  assign n8004 = n3863 & n8003 ;
  assign n8005 = n3603 & ~n4473 ;
  assign n8006 = ~n8004 & n8005 ;
  assign n8007 = ( n487 & n751 ) | ( n487 & ~n1772 ) | ( n751 & ~n1772 ) ;
  assign n8008 = n8007 ^ n3942 ^ n536 ;
  assign n8015 = n2718 ^ n2278 ^ n2139 ;
  assign n8016 = n4598 & ~n5539 ;
  assign n8017 = ~n8015 & n8016 ;
  assign n8010 = n4225 ^ n1949 ^ n588 ;
  assign n8009 = n5134 & n5173 ;
  assign n8011 = n8010 ^ n8009 ^ 1'b0 ;
  assign n8012 = n7591 ^ n3294 ^ 1'b0 ;
  assign n8013 = n4481 | n8012 ;
  assign n8014 = n8011 | n8013 ;
  assign n8018 = n8017 ^ n8014 ^ 1'b0 ;
  assign n8019 = x0 | n8018 ;
  assign n8020 = n3886 ^ n622 ^ 1'b0 ;
  assign n8021 = n6096 & n8020 ;
  assign n8022 = n1543 & n8021 ;
  assign n8023 = n6548 & n8022 ;
  assign n8024 = ~n3128 & n5499 ;
  assign n8025 = n8024 ^ n2033 ^ 1'b0 ;
  assign n8031 = n4376 | n6362 ;
  assign n8032 = n8031 ^ n2604 ^ 1'b0 ;
  assign n8027 = n6907 ^ n2131 ^ n834 ;
  assign n8026 = n7726 ^ n4285 ^ 1'b0 ;
  assign n8028 = n8027 ^ n8026 ^ n1436 ;
  assign n8029 = ~n1816 & n8028 ;
  assign n8030 = n8029 ^ n2553 ^ 1'b0 ;
  assign n8033 = n8032 ^ n8030 ^ 1'b0 ;
  assign n8034 = ( ~n297 & n4868 ) | ( ~n297 & n6462 ) | ( n4868 & n6462 ) ;
  assign n8035 = n7609 ^ n7591 ^ n3673 ;
  assign n8036 = n7114 ^ n5685 ^ n1098 ;
  assign n8037 = n683 & n1831 ;
  assign n8038 = ( n536 & ~n1326 ) | ( n536 & n8037 ) | ( ~n1326 & n8037 ) ;
  assign n8039 = n6410 ^ n4685 ^ n844 ;
  assign n8041 = n290 | n6749 ;
  assign n8042 = n8041 ^ n841 ^ 1'b0 ;
  assign n8040 = ( x135 & n565 ) | ( x135 & n3021 ) | ( n565 & n3021 ) ;
  assign n8043 = n8042 ^ n8040 ^ n4518 ;
  assign n8044 = n8043 ^ n5032 ^ 1'b0 ;
  assign n8045 = n7500 & ~n8044 ;
  assign n8047 = ( ~n1761 & n2070 ) | ( ~n1761 & n6017 ) | ( n2070 & n6017 ) ;
  assign n8048 = n8047 ^ n266 ^ 1'b0 ;
  assign n8046 = n2712 & n3348 ;
  assign n8049 = n8048 ^ n8046 ^ 1'b0 ;
  assign n8053 = ( n957 & ~n4575 ) | ( n957 & n6360 ) | ( ~n4575 & n6360 ) ;
  assign n8054 = n5851 & n8053 ;
  assign n8055 = n8054 ^ n1196 ^ 1'b0 ;
  assign n8050 = n2367 ^ n683 ^ 1'b0 ;
  assign n8051 = ~n5535 & n8050 ;
  assign n8052 = n8051 ^ n3305 ^ 1'b0 ;
  assign n8056 = n8055 ^ n8052 ^ n2991 ;
  assign n8057 = n3632 ^ x227 ^ 1'b0 ;
  assign n8058 = x54 & ~n2015 ;
  assign n8059 = n8058 ^ n1309 ^ 1'b0 ;
  assign n8060 = ( n1760 & ~n2875 ) | ( n1760 & n8059 ) | ( ~n2875 & n8059 ) ;
  assign n8061 = ~n1915 & n4430 ;
  assign n8062 = n8061 ^ n1491 ^ 1'b0 ;
  assign n8063 = n2309 | n7189 ;
  assign n8064 = n8063 ^ n3013 ^ x70 ;
  assign n8065 = n8064 ^ n3765 ^ 1'b0 ;
  assign n8066 = ~n2315 & n8065 ;
  assign n8067 = n7049 & n8066 ;
  assign n8068 = n8062 & n8067 ;
  assign n8069 = n8068 ^ n4987 ^ 1'b0 ;
  assign n8070 = ( n3058 & n3929 ) | ( n3058 & ~n8069 ) | ( n3929 & ~n8069 ) ;
  assign n8071 = ( ~n277 & n4338 ) | ( ~n277 & n7217 ) | ( n4338 & n7217 ) ;
  assign n8072 = n2098 ^ n661 ^ x250 ;
  assign n8073 = n8071 | n8072 ;
  assign n8074 = ( n8060 & ~n8070 ) | ( n8060 & n8073 ) | ( ~n8070 & n8073 ) ;
  assign n8077 = ( n816 & ~n5415 ) | ( n816 & n5559 ) | ( ~n5415 & n5559 ) ;
  assign n8075 = n909 & ~n3951 ;
  assign n8076 = ~n2296 & n8075 ;
  assign n8078 = n8077 ^ n8076 ^ 1'b0 ;
  assign n8079 = n2195 ^ n1279 ^ n446 ;
  assign n8080 = n8079 ^ n3188 ^ 1'b0 ;
  assign n8081 = n788 | n4542 ;
  assign n8082 = n1067 & ~n8081 ;
  assign n8083 = n8082 ^ n5350 ^ n3992 ;
  assign n8084 = n5990 ^ n3084 ^ 1'b0 ;
  assign n8085 = ( x36 & ~x240 ) | ( x36 & n4938 ) | ( ~x240 & n4938 ) ;
  assign n8086 = ( n485 & n7999 ) | ( n485 & ~n8085 ) | ( n7999 & ~n8085 ) ;
  assign n8087 = n928 & n8086 ;
  assign n8088 = n5581 ^ n1396 ^ 1'b0 ;
  assign n8089 = n8087 & n8088 ;
  assign n8090 = ~n8084 & n8089 ;
  assign n8092 = n4740 ^ n4182 ^ n1367 ;
  assign n8093 = ( n432 & ~n1432 ) | ( n432 & n8092 ) | ( ~n1432 & n8092 ) ;
  assign n8094 = n1892 | n4040 ;
  assign n8095 = ( n690 & ~n8093 ) | ( n690 & n8094 ) | ( ~n8093 & n8094 ) ;
  assign n8091 = n5899 ^ n2530 ^ 1'b0 ;
  assign n8096 = n8095 ^ n8091 ^ 1'b0 ;
  assign n8097 = n6078 & n8096 ;
  assign n8098 = n946 & ~n981 ;
  assign n8099 = n8098 ^ n6796 ^ 1'b0 ;
  assign n8100 = n1978 & ~n2810 ;
  assign n8101 = ( n2693 & n6190 ) | ( n2693 & ~n8100 ) | ( n6190 & ~n8100 ) ;
  assign n8102 = ( ~n803 & n1171 ) | ( ~n803 & n1597 ) | ( n1171 & n1597 ) ;
  assign n8103 = n8102 ^ n2134 ^ 1'b0 ;
  assign n8104 = ( n883 & n1388 ) | ( n883 & n8103 ) | ( n1388 & n8103 ) ;
  assign n8105 = ( ~n1527 & n5617 ) | ( ~n1527 & n6575 ) | ( n5617 & n6575 ) ;
  assign n8106 = n8105 ^ n6099 ^ n3218 ;
  assign n8107 = n5660 ^ n4824 ^ n4651 ;
  assign n8108 = n4153 ^ n3900 ^ 1'b0 ;
  assign n8109 = n2100 & ~n8108 ;
  assign n8110 = n6412 | n8109 ;
  assign n8111 = ( ~n2498 & n2787 ) | ( ~n2498 & n2979 ) | ( n2787 & n2979 ) ;
  assign n8112 = ~n952 & n8111 ;
  assign n8113 = n8112 ^ n6389 ^ n4521 ;
  assign n8114 = n8113 ^ n3512 ^ n3339 ;
  assign n8116 = x187 & n5651 ;
  assign n8117 = n8116 ^ n1734 ^ 1'b0 ;
  assign n8115 = n2375 & ~n2776 ;
  assign n8118 = n8117 ^ n8115 ^ 1'b0 ;
  assign n8119 = n2331 ^ n2272 ^ 1'b0 ;
  assign n8120 = x34 & n8119 ;
  assign n8121 = n8120 ^ n2671 ^ 1'b0 ;
  assign n8122 = ( n1910 & ~n7871 ) | ( n1910 & n8121 ) | ( ~n7871 & n8121 ) ;
  assign n8123 = ~n4157 & n8122 ;
  assign n8124 = n5241 ^ n631 ^ 1'b0 ;
  assign n8125 = n8124 ^ n6560 ^ 1'b0 ;
  assign n8126 = x171 & n8125 ;
  assign n8127 = n5780 | n8126 ;
  assign n8128 = n2598 | n3481 ;
  assign n8129 = x101 & ~n4272 ;
  assign n8130 = ~n3069 & n8129 ;
  assign n8131 = n8128 & ~n8130 ;
  assign n8132 = n940 & n8131 ;
  assign n8133 = n879 & ~n8132 ;
  assign n8134 = ( n1885 & n6170 ) | ( n1885 & ~n7583 ) | ( n6170 & ~n7583 ) ;
  assign n8135 = n7516 ^ n6195 ^ n5114 ;
  assign n8139 = n2196 & n4825 ;
  assign n8138 = n3910 & n7009 ;
  assign n8136 = n8028 ^ n2624 ^ n335 ;
  assign n8137 = ~n6702 & n8136 ;
  assign n8140 = n8139 ^ n8138 ^ n8137 ;
  assign n8141 = n7381 ^ n5769 ^ n4893 ;
  assign n8144 = n1415 & ~n1573 ;
  assign n8145 = n8144 ^ n798 ^ 1'b0 ;
  assign n8146 = n6311 & ~n7013 ;
  assign n8147 = n8145 & n8146 ;
  assign n8148 = n8147 ^ n6585 ^ 1'b0 ;
  assign n8142 = n2744 & n6424 ;
  assign n8143 = n8142 ^ n2574 ^ 1'b0 ;
  assign n8149 = n8148 ^ n8143 ^ n2315 ;
  assign n8150 = ( n3721 & n5693 ) | ( n3721 & ~n8149 ) | ( n5693 & ~n8149 ) ;
  assign n8151 = n4740 | n5628 ;
  assign n8152 = n8151 ^ n1376 ^ 1'b0 ;
  assign n8153 = n5914 & ~n6868 ;
  assign n8154 = ~n8152 & n8153 ;
  assign n8156 = n5459 ^ n2724 ^ n1148 ;
  assign n8157 = n3493 ^ n1617 ^ n1032 ;
  assign n8158 = n8157 ^ n3627 ^ n2384 ;
  assign n8159 = ( n2144 & n8156 ) | ( n2144 & ~n8158 ) | ( n8156 & ~n8158 ) ;
  assign n8155 = n3408 ^ n1049 ^ 1'b0 ;
  assign n8160 = n8159 ^ n8155 ^ x178 ;
  assign n8161 = n2169 ^ n1222 ^ 1'b0 ;
  assign n8162 = n3036 & ~n8161 ;
  assign n8167 = n2553 ^ x226 ^ 1'b0 ;
  assign n8168 = n7314 & n8167 ;
  assign n8163 = n2576 ^ n1791 ^ n511 ;
  assign n8164 = n2355 | n8163 ;
  assign n8165 = ~n2720 & n8164 ;
  assign n8166 = ~n506 & n8165 ;
  assign n8169 = n8168 ^ n8166 ^ n3927 ;
  assign n8170 = n1644 & ~n8169 ;
  assign n8171 = ( ~n1044 & n8162 ) | ( ~n1044 & n8170 ) | ( n8162 & n8170 ) ;
  assign n8172 = n3840 ^ n3159 ^ 1'b0 ;
  assign n8173 = n5411 & ~n8172 ;
  assign n8176 = ~n490 & n1061 ;
  assign n8177 = n8176 ^ n3759 ^ 1'b0 ;
  assign n8175 = n3779 & ~n5242 ;
  assign n8178 = n8177 ^ n8175 ^ 1'b0 ;
  assign n8179 = ( n4234 & n7195 ) | ( n4234 & n8178 ) | ( n7195 & n8178 ) ;
  assign n8174 = n3843 ^ n577 ^ 1'b0 ;
  assign n8180 = n8179 ^ n8174 ^ n3427 ;
  assign n8181 = n6029 | n8180 ;
  assign n8182 = n8181 ^ n6211 ^ 1'b0 ;
  assign n8183 = ( n3949 & n8173 ) | ( n3949 & ~n8182 ) | ( n8173 & ~n8182 ) ;
  assign n8184 = n2529 ^ n1642 ^ 1'b0 ;
  assign n8185 = ( n5266 & n6468 ) | ( n5266 & n6550 ) | ( n6468 & n6550 ) ;
  assign n8186 = n5713 ^ n587 ^ 1'b0 ;
  assign n8187 = n381 | n8186 ;
  assign n8188 = ( n1508 & n5622 ) | ( n1508 & n8187 ) | ( n5622 & n8187 ) ;
  assign n8189 = ( x203 & n2139 ) | ( x203 & n8188 ) | ( n2139 & n8188 ) ;
  assign n8190 = n7475 ^ n7113 ^ n5935 ;
  assign n8192 = n2102 ^ n1836 ^ 1'b0 ;
  assign n8193 = n2980 | n8192 ;
  assign n8191 = n7554 ^ n5110 ^ 1'b0 ;
  assign n8194 = n8193 ^ n8191 ^ 1'b0 ;
  assign n8195 = n8190 | n8194 ;
  assign n8196 = n8195 ^ n6685 ^ 1'b0 ;
  assign n8200 = n2352 & n2712 ;
  assign n8198 = n1536 | n3121 ;
  assign n8199 = n6162 & ~n8198 ;
  assign n8197 = ( ~n2662 & n3278 ) | ( ~n2662 & n3961 ) | ( n3278 & n3961 ) ;
  assign n8201 = n8200 ^ n8199 ^ n8197 ;
  assign n8202 = n1307 ^ n633 ^ 1'b0 ;
  assign n8203 = n6323 & n8202 ;
  assign n8204 = n483 & ~n1921 ;
  assign n8205 = ~x113 & n8204 ;
  assign n8206 = n2132 ^ n2003 ^ n1197 ;
  assign n8209 = n6884 ^ n2442 ^ 1'b0 ;
  assign n8207 = n6211 ^ x133 ^ 1'b0 ;
  assign n8208 = n1255 & n8207 ;
  assign n8210 = n8209 ^ n8208 ^ x57 ;
  assign n8211 = ( n6244 & n8206 ) | ( n6244 & ~n8210 ) | ( n8206 & ~n8210 ) ;
  assign n8212 = ( ~n425 & n652 ) | ( ~n425 & n6591 ) | ( n652 & n6591 ) ;
  assign n8213 = ( ~x205 & n2692 ) | ( ~x205 & n8212 ) | ( n2692 & n8212 ) ;
  assign n8214 = ( n2651 & n6090 ) | ( n2651 & n8213 ) | ( n6090 & n8213 ) ;
  assign n8215 = n3241 & n3791 ;
  assign n8216 = n8215 ^ n6963 ^ n4132 ;
  assign n8217 = n5997 | n8216 ;
  assign n8218 = ( n3380 & n3763 ) | ( n3380 & n4147 ) | ( n3763 & n4147 ) ;
  assign n8219 = ( n2743 & n2954 ) | ( n2743 & ~n8218 ) | ( n2954 & ~n8218 ) ;
  assign n8221 = n4582 ^ n3225 ^ n1693 ;
  assign n8222 = ( n3637 & ~n6148 ) | ( n3637 & n8221 ) | ( ~n6148 & n8221 ) ;
  assign n8220 = n6873 ^ n6273 ^ n1826 ;
  assign n8223 = n8222 ^ n8220 ^ 1'b0 ;
  assign n8224 = n8219 & ~n8223 ;
  assign n8225 = n8217 & n8224 ;
  assign n8226 = ~n3813 & n8225 ;
  assign n8230 = n7971 ^ n1825 ^ 1'b0 ;
  assign n8231 = n4255 | n8230 ;
  assign n8232 = n8231 ^ n4142 ^ n296 ;
  assign n8227 = n774 & ~n1118 ;
  assign n8228 = n8227 ^ x232 ^ 1'b0 ;
  assign n8229 = ( n5958 & n7088 ) | ( n5958 & n8228 ) | ( n7088 & n8228 ) ;
  assign n8233 = n8232 ^ n8229 ^ 1'b0 ;
  assign n8234 = n1519 ^ n1068 ^ 1'b0 ;
  assign n8235 = n5882 ^ n4693 ^ n3138 ;
  assign n8236 = ( n6488 & n6565 ) | ( n6488 & n8235 ) | ( n6565 & n8235 ) ;
  assign n8237 = n8236 ^ n1172 ^ 1'b0 ;
  assign n8238 = n989 ^ n933 ^ 1'b0 ;
  assign n8239 = n1806 & n8238 ;
  assign n8240 = n4189 & n8239 ;
  assign n8241 = n6773 & n8240 ;
  assign n8242 = n8241 ^ n6458 ^ 1'b0 ;
  assign n8243 = n7091 & ~n8242 ;
  assign n8244 = n6004 & ~n6018 ;
  assign n8245 = n8244 ^ n5654 ^ 1'b0 ;
  assign n8246 = n1540 & ~n4611 ;
  assign n8247 = n1272 & n8246 ;
  assign n8248 = n8245 & n8247 ;
  assign n8249 = n4853 ^ n4753 ^ n3383 ;
  assign n8250 = ~n5458 & n8249 ;
  assign n8251 = ( n2411 & n8248 ) | ( n2411 & ~n8250 ) | ( n8248 & ~n8250 ) ;
  assign n8256 = n4384 ^ n2979 ^ x106 ;
  assign n8257 = ( x77 & ~n806 ) | ( x77 & n5900 ) | ( ~n806 & n5900 ) ;
  assign n8258 = n8257 ^ n2369 ^ 1'b0 ;
  assign n8259 = n8256 | n8258 ;
  assign n8253 = n1908 & n2652 ;
  assign n8252 = x179 & ~n8216 ;
  assign n8254 = n8253 ^ n8252 ^ 1'b0 ;
  assign n8255 = ~n7265 & n8254 ;
  assign n8260 = n8259 ^ n8255 ^ 1'b0 ;
  assign n8261 = n8198 ^ n1208 ^ 1'b0 ;
  assign n8262 = n4445 & n8261 ;
  assign n8263 = ~n986 & n5523 ;
  assign n8264 = n8263 ^ n6673 ^ 1'b0 ;
  assign n8265 = n4344 ^ n599 ^ 1'b0 ;
  assign n8266 = n8264 & n8265 ;
  assign n8267 = ( n8164 & ~n8262 ) | ( n8164 & n8266 ) | ( ~n8262 & n8266 ) ;
  assign n8268 = x234 | n658 ;
  assign n8269 = ~n1412 & n3406 ;
  assign n8270 = ~n403 & n8269 ;
  assign n8271 = n1779 | n3322 ;
  assign n8272 = n261 | n8271 ;
  assign n8273 = ~n7325 & n8272 ;
  assign n8274 = n8270 & n8273 ;
  assign n8275 = n1294 | n8274 ;
  assign n8276 = n8268 | n8275 ;
  assign n8277 = n8276 ^ n606 ^ 1'b0 ;
  assign n8278 = n8267 & ~n8277 ;
  assign n8279 = n318 & n7366 ;
  assign n8280 = n8279 ^ n4906 ^ 1'b0 ;
  assign n8281 = n8280 ^ n6251 ^ n2276 ;
  assign n8282 = ( n862 & n986 ) | ( n862 & n8281 ) | ( n986 & n8281 ) ;
  assign n8283 = n1693 ^ n1012 ^ 1'b0 ;
  assign n8284 = n2701 & ~n8283 ;
  assign n8285 = ~n7706 & n8284 ;
  assign n8286 = n3368 & n8285 ;
  assign n8287 = n8286 ^ n6090 ^ 1'b0 ;
  assign n8288 = n6667 & n7536 ;
  assign n8289 = x74 & ~n495 ;
  assign n8290 = n8289 ^ n6484 ^ 1'b0 ;
  assign n8291 = n4195 & n8290 ;
  assign n8292 = n8288 & ~n8291 ;
  assign n8293 = n2899 & n8292 ;
  assign n8294 = n1846 ^ n566 ^ 1'b0 ;
  assign n8295 = n1984 | n6642 ;
  assign n8296 = n8295 ^ n3959 ^ 1'b0 ;
  assign n8297 = n5022 ^ n4692 ^ 1'b0 ;
  assign n8298 = x4 & ~n8297 ;
  assign n8299 = ~n8296 & n8298 ;
  assign n8300 = n8294 | n8299 ;
  assign n8301 = n7612 | n8300 ;
  assign n8302 = n8083 | n8188 ;
  assign n8305 = n1927 & ~n4068 ;
  assign n8303 = n4603 ^ n1289 ^ n656 ;
  assign n8304 = ( n7612 & ~n8000 ) | ( n7612 & n8303 ) | ( ~n8000 & n8303 ) ;
  assign n8306 = n8305 ^ n8304 ^ n3320 ;
  assign n8307 = ( n668 & n796 ) | ( n668 & n5268 ) | ( n796 & n5268 ) ;
  assign n8308 = ( ~n2963 & n7044 ) | ( ~n2963 & n8307 ) | ( n7044 & n8307 ) ;
  assign n8312 = n3550 ^ n2878 ^ 1'b0 ;
  assign n8313 = n1772 & n8312 ;
  assign n8309 = n7490 ^ n2671 ^ n1317 ;
  assign n8310 = n8309 ^ n6983 ^ 1'b0 ;
  assign n8311 = ~n1304 & n8310 ;
  assign n8314 = n8313 ^ n8311 ^ 1'b0 ;
  assign n8315 = n1937 & n8314 ;
  assign n8316 = n8315 ^ n6048 ^ n5477 ;
  assign n8317 = n7301 | n8316 ;
  assign n8318 = n8317 ^ n500 ^ 1'b0 ;
  assign n8319 = n1478 ^ n1227 ^ 1'b0 ;
  assign n8320 = n8319 ^ n2398 ^ n1760 ;
  assign n8321 = n6878 ^ n2812 ^ n1760 ;
  assign n8322 = n7116 ^ n3556 ^ 1'b0 ;
  assign n8323 = n1945 & ~n8322 ;
  assign n8324 = ( ~n2796 & n2882 ) | ( ~n2796 & n8323 ) | ( n2882 & n8323 ) ;
  assign n8325 = ( ~n8320 & n8321 ) | ( ~n8320 & n8324 ) | ( n8321 & n8324 ) ;
  assign n8326 = n8325 ^ n7602 ^ n1759 ;
  assign n8327 = n5114 ^ n3899 ^ n3256 ;
  assign n8328 = ( n2040 & ~n8326 ) | ( n2040 & n8327 ) | ( ~n8326 & n8327 ) ;
  assign n8329 = n696 & n1185 ;
  assign n8330 = ( ~x1 & n877 ) | ( ~x1 & n1432 ) | ( n877 & n1432 ) ;
  assign n8331 = n1627 & ~n8330 ;
  assign n8332 = n8331 ^ n4784 ^ x39 ;
  assign n8333 = ~n2948 & n6122 ;
  assign n8334 = n8333 ^ n5278 ^ n2178 ;
  assign n8335 = x37 & ~n8334 ;
  assign n8336 = n8335 ^ n5063 ^ 1'b0 ;
  assign n8337 = n7741 ^ n1007 ^ x102 ;
  assign n8338 = ( n2246 & ~n4863 ) | ( n2246 & n8337 ) | ( ~n4863 & n8337 ) ;
  assign n8339 = n1381 ^ n1083 ^ 1'b0 ;
  assign n8340 = ~n704 & n8339 ;
  assign n8341 = ( n3110 & n5527 ) | ( n3110 & ~n8340 ) | ( n5527 & ~n8340 ) ;
  assign n8342 = n8341 ^ n5350 ^ 1'b0 ;
  assign n8343 = n8342 ^ x201 ^ 1'b0 ;
  assign n8344 = n8338 & ~n8343 ;
  assign n8345 = ( ~n6411 & n8336 ) | ( ~n6411 & n8344 ) | ( n8336 & n8344 ) ;
  assign n8346 = n2669 ^ x126 ^ 1'b0 ;
  assign n8347 = ~n4386 & n5237 ;
  assign n8348 = n2021 | n3662 ;
  assign n8349 = n8348 ^ n2607 ^ 1'b0 ;
  assign n8350 = ( n1859 & n3061 ) | ( n1859 & ~n8349 ) | ( n3061 & ~n8349 ) ;
  assign n8351 = n8350 ^ n7150 ^ n331 ;
  assign n8352 = n6289 ^ n2229 ^ 1'b0 ;
  assign n8353 = ( ~n5385 & n6369 ) | ( ~n5385 & n8352 ) | ( n6369 & n8352 ) ;
  assign n8360 = n2936 ^ n1158 ^ 1'b0 ;
  assign n8355 = ( ~n3157 & n5036 ) | ( ~n3157 & n5640 ) | ( n5036 & n5640 ) ;
  assign n8356 = n8355 ^ x30 ^ 1'b0 ;
  assign n8357 = n6459 ^ n2212 ^ n1432 ;
  assign n8358 = n5018 & n8357 ;
  assign n8359 = ~n8356 & n8358 ;
  assign n8354 = n7322 ^ n5927 ^ 1'b0 ;
  assign n8361 = n8360 ^ n8359 ^ n8354 ;
  assign n8362 = n1982 & n8361 ;
  assign n8363 = ~n8353 & n8362 ;
  assign n8364 = n2248 ^ n1447 ^ 1'b0 ;
  assign n8365 = n7113 | n8364 ;
  assign n8366 = n2132 & ~n8365 ;
  assign n8367 = n8366 ^ n5149 ^ 1'b0 ;
  assign n8368 = n1487 | n8367 ;
  assign n8369 = n1506 | n2168 ;
  assign n8370 = ( n1672 & n2743 ) | ( n1672 & ~n8369 ) | ( n2743 & ~n8369 ) ;
  assign n8371 = n3726 | n8370 ;
  assign n8372 = n8371 ^ n3476 ^ 1'b0 ;
  assign n8373 = n3202 ^ n2666 ^ 1'b0 ;
  assign n8374 = n8373 ^ n4462 ^ n2444 ;
  assign n8375 = n8374 ^ n3294 ^ 1'b0 ;
  assign n8376 = n8011 ^ n5121 ^ n4858 ;
  assign n8377 = n798 & ~n5543 ;
  assign n8378 = n811 & n8377 ;
  assign n8379 = n8378 ^ n7946 ^ n1642 ;
  assign n8380 = ( n5477 & n8376 ) | ( n5477 & ~n8379 ) | ( n8376 & ~n8379 ) ;
  assign n8381 = n7463 & n8272 ;
  assign n8382 = n8381 ^ n2844 ^ 1'b0 ;
  assign n8383 = n8382 ^ n4032 ^ 1'b0 ;
  assign n8384 = n8380 | n8383 ;
  assign n8385 = ~n1010 & n1374 ;
  assign n8386 = n8385 ^ n822 ^ 1'b0 ;
  assign n8387 = n2489 ^ n1084 ^ 1'b0 ;
  assign n8388 = n6349 & ~n8387 ;
  assign n8389 = ~n5079 & n8388 ;
  assign n8390 = n8389 ^ x240 ^ 1'b0 ;
  assign n8391 = ~n4474 & n8390 ;
  assign n8392 = ~n2412 & n8391 ;
  assign n8393 = ~n8386 & n8392 ;
  assign n8394 = n8393 ^ n4328 ^ 1'b0 ;
  assign n8396 = n2633 & n4622 ;
  assign n8395 = n1296 & ~n3810 ;
  assign n8397 = n8396 ^ n8395 ^ 1'b0 ;
  assign n8398 = n1883 & ~n5744 ;
  assign n8399 = ~n5225 & n6589 ;
  assign n8400 = n8399 ^ n1118 ^ 1'b0 ;
  assign n8401 = n8400 ^ n7089 ^ n5471 ;
  assign n8402 = ( n3188 & ~n8398 ) | ( n3188 & n8401 ) | ( ~n8398 & n8401 ) ;
  assign n8403 = ( n741 & n2192 ) | ( n741 & n7236 ) | ( n2192 & n7236 ) ;
  assign n8404 = n3600 & n4902 ;
  assign n8405 = n8403 & n8404 ;
  assign n8406 = n8405 ^ n2855 ^ 1'b0 ;
  assign n8407 = n4073 ^ n2191 ^ n984 ;
  assign n8408 = n8407 ^ n2382 ^ n1755 ;
  assign n8409 = ( ~n4156 & n6088 ) | ( ~n4156 & n8408 ) | ( n6088 & n8408 ) ;
  assign n8410 = n2855 & ~n3753 ;
  assign n8411 = ~n8409 & n8410 ;
  assign n8412 = n1122 ^ n1014 ^ 1'b0 ;
  assign n8413 = x158 & n8412 ;
  assign n8414 = n8413 ^ n5159 ^ n3633 ;
  assign n8415 = n4844 ^ n1416 ^ n640 ;
  assign n8416 = n8415 ^ n1628 ^ 1'b0 ;
  assign n8417 = ~n2819 & n8416 ;
  assign n8418 = ( n3529 & n6995 ) | ( n3529 & n8417 ) | ( n6995 & n8417 ) ;
  assign n8419 = ( x36 & n320 ) | ( x36 & ~n1308 ) | ( n320 & ~n1308 ) ;
  assign n8420 = ( n4831 & n8272 ) | ( n4831 & n8419 ) | ( n8272 & n8419 ) ;
  assign n8421 = n4933 & ~n7406 ;
  assign n8422 = ~n8420 & n8421 ;
  assign n8423 = n4301 ^ n1580 ^ 1'b0 ;
  assign n8424 = n1599 & ~n8423 ;
  assign n8425 = n2688 ^ n1921 ^ 1'b0 ;
  assign n8426 = ( ~n2642 & n3732 ) | ( ~n2642 & n8425 ) | ( n3732 & n8425 ) ;
  assign n8427 = ( x112 & ~n5792 ) | ( x112 & n8426 ) | ( ~n5792 & n8426 ) ;
  assign n8428 = ( n1714 & ~n5685 ) | ( n1714 & n7372 ) | ( ~n5685 & n7372 ) ;
  assign n8430 = x42 & ~n781 ;
  assign n8431 = n8430 ^ n4752 ^ 1'b0 ;
  assign n8429 = n7596 ^ n2553 ^ n2229 ;
  assign n8432 = n8431 ^ n8429 ^ n2146 ;
  assign n8433 = x79 & ~n2042 ;
  assign n8434 = n8433 ^ n419 ^ 1'b0 ;
  assign n8435 = n4407 ^ n3736 ^ n2765 ;
  assign n8436 = ( x173 & n8434 ) | ( x173 & n8435 ) | ( n8434 & n8435 ) ;
  assign n8437 = n7598 ^ n4099 ^ 1'b0 ;
  assign n8438 = n1633 ^ n715 ^ 1'b0 ;
  assign n8439 = n8438 ^ n6837 ^ 1'b0 ;
  assign n8440 = n8437 & n8439 ;
  assign n8441 = x7 & n2167 ;
  assign n8442 = ~n2701 & n8441 ;
  assign n8443 = n8442 ^ n2139 ^ 1'b0 ;
  assign n8447 = ~n1781 & n4354 ;
  assign n8444 = n2672 & ~n4363 ;
  assign n8445 = n8444 ^ n4611 ^ 1'b0 ;
  assign n8446 = ( n1343 & n1921 ) | ( n1343 & ~n8445 ) | ( n1921 & ~n8445 ) ;
  assign n8448 = n8447 ^ n8446 ^ 1'b0 ;
  assign n8449 = ~n2999 & n8448 ;
  assign n8450 = n461 | n1126 ;
  assign n8451 = n1797 | n8450 ;
  assign n8452 = ( x88 & n5587 ) | ( x88 & n8451 ) | ( n5587 & n8451 ) ;
  assign n8453 = n487 ^ n469 ^ 1'b0 ;
  assign n8454 = n2111 | n3335 ;
  assign n8455 = n8453 | n8454 ;
  assign n8456 = ( n2320 & n7433 ) | ( n2320 & ~n8455 ) | ( n7433 & ~n8455 ) ;
  assign n8457 = n7259 ^ n6659 ^ n2372 ;
  assign n8459 = n414 & n5258 ;
  assign n8458 = ~n2391 & n3983 ;
  assign n8460 = n8459 ^ n8458 ^ n6549 ;
  assign n8461 = n4659 ^ n2907 ^ n2843 ;
  assign n8462 = ( ~n4035 & n4939 ) | ( ~n4035 & n8461 ) | ( n4939 & n8461 ) ;
  assign n8463 = ~n2113 & n2978 ;
  assign n8464 = n4136 ^ n1527 ^ 1'b0 ;
  assign n8465 = x130 & n8464 ;
  assign n8466 = n5604 & ~n8465 ;
  assign n8467 = ( n4929 & n8463 ) | ( n4929 & ~n8466 ) | ( n8463 & ~n8466 ) ;
  assign n8468 = n3422 & n7646 ;
  assign n8469 = n8468 ^ n7879 ^ 1'b0 ;
  assign n8470 = n8467 & ~n8469 ;
  assign n8473 = ( n864 & n2169 ) | ( n864 & n3865 ) | ( n2169 & n3865 ) ;
  assign n8474 = n3146 ^ x147 ^ 1'b0 ;
  assign n8475 = ~n8473 & n8474 ;
  assign n8471 = n2620 & ~n5285 ;
  assign n8472 = n8471 ^ n4945 ^ 1'b0 ;
  assign n8476 = n8475 ^ n8472 ^ n6218 ;
  assign n8477 = n4001 & ~n6706 ;
  assign n8478 = ( ~n335 & n416 ) | ( ~n335 & n3185 ) | ( n416 & n3185 ) ;
  assign n8479 = ( ~n5701 & n6146 ) | ( ~n5701 & n6645 ) | ( n6146 & n6645 ) ;
  assign n8480 = ~n6657 & n8479 ;
  assign n8481 = ( ~n8124 & n8478 ) | ( ~n8124 & n8480 ) | ( n8478 & n8480 ) ;
  assign n8485 = n2732 & ~n3353 ;
  assign n8486 = n8485 ^ n1245 ^ 1'b0 ;
  assign n8487 = n6523 ^ n5958 ^ 1'b0 ;
  assign n8488 = n3352 | n8487 ;
  assign n8489 = n8486 | n8488 ;
  assign n8482 = n2873 ^ x65 ^ 1'b0 ;
  assign n8483 = n7406 ^ n966 ^ 1'b0 ;
  assign n8484 = n8482 | n8483 ;
  assign n8490 = n8489 ^ n8484 ^ 1'b0 ;
  assign n8491 = n8481 & ~n8490 ;
  assign n8492 = ( n1346 & n2220 ) | ( n1346 & n3933 ) | ( n2220 & n3933 ) ;
  assign n8493 = n8492 ^ n8076 ^ x110 ;
  assign n8494 = ( x82 & n559 ) | ( x82 & ~n3747 ) | ( n559 & ~n3747 ) ;
  assign n8495 = n6417 ^ n6075 ^ n2865 ;
  assign n8496 = ( n1188 & n4210 ) | ( n1188 & ~n6203 ) | ( n4210 & ~n6203 ) ;
  assign n8497 = n5264 & ~n7894 ;
  assign n8498 = n1201 & n8497 ;
  assign n8499 = ( n2553 & n8496 ) | ( n2553 & ~n8498 ) | ( n8496 & ~n8498 ) ;
  assign n8500 = ( x222 & n1766 ) | ( x222 & n3252 ) | ( n1766 & n3252 ) ;
  assign n8501 = n4237 ^ n1298 ^ 1'b0 ;
  assign n8502 = n8501 ^ n4837 ^ 1'b0 ;
  assign n8503 = ~n8500 & n8502 ;
  assign n8504 = n6839 ^ n3835 ^ 1'b0 ;
  assign n8505 = n8503 & n8504 ;
  assign n8506 = ~n2670 & n8505 ;
  assign n8507 = ~x59 & n1096 ;
  assign n8509 = n1968 | n7294 ;
  assign n8508 = n1581 ^ n1373 ^ 1'b0 ;
  assign n8510 = n8509 ^ n8508 ^ n7390 ;
  assign n8511 = ~n8507 & n8510 ;
  assign n8512 = ( n1625 & n2639 ) | ( n1625 & n2885 ) | ( n2639 & n2885 ) ;
  assign n8513 = ~n7266 & n8512 ;
  assign n8514 = n5314 ^ n4526 ^ n3962 ;
  assign n8515 = ( n2501 & n4848 ) | ( n2501 & ~n8514 ) | ( n4848 & ~n8514 ) ;
  assign n8516 = n8515 ^ x110 ^ 1'b0 ;
  assign n8517 = n3431 ^ n2711 ^ 1'b0 ;
  assign n8518 = n8350 & ~n8517 ;
  assign n8519 = n8516 & n8518 ;
  assign n8521 = ~n1393 & n5703 ;
  assign n8522 = ~n4066 & n8521 ;
  assign n8520 = ~n1274 & n4322 ;
  assign n8523 = n8522 ^ n8520 ^ 1'b0 ;
  assign n8524 = n8523 ^ n7631 ^ n2367 ;
  assign n8525 = n2451 & ~n8524 ;
  assign n8526 = n3686 & n5248 ;
  assign n8527 = n1028 & ~n8526 ;
  assign n8528 = ( ~n7445 & n7604 ) | ( ~n7445 & n8527 ) | ( n7604 & n8527 ) ;
  assign n8529 = n8528 ^ n7680 ^ n2292 ;
  assign n8530 = n7116 ^ n3313 ^ x200 ;
  assign n8531 = n6274 & ~n8530 ;
  assign n8532 = n3591 ^ n1978 ^ 1'b0 ;
  assign n8533 = n6839 & ~n8532 ;
  assign n8534 = n3391 | n8533 ;
  assign n8535 = n5808 ^ n4033 ^ 1'b0 ;
  assign n8536 = x49 & ~n8535 ;
  assign n8537 = n6510 ^ n4153 ^ 1'b0 ;
  assign n8538 = ( x191 & ~n2098 ) | ( x191 & n6242 ) | ( ~n2098 & n6242 ) ;
  assign n8539 = ( x151 & n8537 ) | ( x151 & ~n8538 ) | ( n8537 & ~n8538 ) ;
  assign n8540 = n8539 ^ n3660 ^ n2444 ;
  assign n8541 = n8536 & ~n8540 ;
  assign n8542 = n8541 ^ n2569 ^ 1'b0 ;
  assign n8543 = ( ~n2046 & n2928 ) | ( ~n2046 & n4445 ) | ( n2928 & n4445 ) ;
  assign n8544 = ~n2419 & n8128 ;
  assign n8545 = n6950 & n8544 ;
  assign n8546 = ( n1228 & n6611 ) | ( n1228 & ~n8545 ) | ( n6611 & ~n8545 ) ;
  assign n8547 = ~n8543 & n8546 ;
  assign n8548 = n8542 & n8547 ;
  assign n8550 = n1243 & ~n4972 ;
  assign n8551 = ( n1366 & ~n2327 ) | ( n1366 & n8550 ) | ( ~n2327 & n8550 ) ;
  assign n8549 = n5686 ^ n618 ^ x12 ;
  assign n8552 = n8551 ^ n8549 ^ n7364 ;
  assign n8553 = ~n4441 & n7984 ;
  assign n8554 = n5001 ^ n2331 ^ 1'b0 ;
  assign n8555 = n4569 & n8554 ;
  assign n8565 = x152 ^ x2 ^ 1'b0 ;
  assign n8562 = ( ~n1578 & n1600 ) | ( ~n1578 & n2098 ) | ( n1600 & n2098 ) ;
  assign n8563 = ( n713 & n1364 ) | ( n713 & ~n8562 ) | ( n1364 & ~n8562 ) ;
  assign n8564 = ~n1856 & n8563 ;
  assign n8566 = n8565 ^ n8564 ^ 1'b0 ;
  assign n8567 = n8566 ^ n8257 ^ n5646 ;
  assign n8556 = n1800 ^ n1466 ^ 1'b0 ;
  assign n8557 = n3326 | n8556 ;
  assign n8558 = ~n595 & n4505 ;
  assign n8559 = n1004 & n8558 ;
  assign n8560 = ~x130 & n8559 ;
  assign n8561 = ( n3232 & n8557 ) | ( n3232 & ~n8560 ) | ( n8557 & ~n8560 ) ;
  assign n8568 = n8567 ^ n8561 ^ n6989 ;
  assign n8569 = n8555 & ~n8568 ;
  assign n8570 = n8569 ^ n3310 ^ 1'b0 ;
  assign n8571 = n643 | n5722 ;
  assign n8572 = n7577 | n8571 ;
  assign n8573 = n3193 & n6820 ;
  assign n8574 = n7171 ^ n2576 ^ n1819 ;
  assign n8575 = n8574 ^ n2998 ^ 1'b0 ;
  assign n8576 = n6505 ^ n3847 ^ n2688 ;
  assign n8577 = ( n2759 & n7706 ) | ( n2759 & ~n8576 ) | ( n7706 & ~n8576 ) ;
  assign n8580 = n861 & ~n1691 ;
  assign n8578 = x78 & n3073 ;
  assign n8579 = n1245 & n8578 ;
  assign n8581 = n8580 ^ n8579 ^ n7845 ;
  assign n8582 = n8581 ^ n1439 ^ 1'b0 ;
  assign n8583 = ( ~n1328 & n2517 ) | ( ~n1328 & n4261 ) | ( n2517 & n4261 ) ;
  assign n8584 = ( ~x111 & n5007 ) | ( ~x111 & n8583 ) | ( n5007 & n8583 ) ;
  assign n8585 = n8584 ^ n5198 ^ 1'b0 ;
  assign n8586 = n6901 & ~n8585 ;
  assign n8587 = n1592 ^ n1465 ^ 1'b0 ;
  assign n8588 = n8587 ^ n3728 ^ n1841 ;
  assign n8589 = n8588 ^ n3460 ^ n2131 ;
  assign n8590 = n8589 ^ n5388 ^ 1'b0 ;
  assign n8591 = n8586 & ~n8590 ;
  assign n8592 = n485 & ~n1172 ;
  assign n8593 = ( n8373 & n8561 ) | ( n8373 & ~n8592 ) | ( n8561 & ~n8592 ) ;
  assign n8594 = n3918 ^ n2530 ^ 1'b0 ;
  assign n8595 = ( ~n1010 & n5687 ) | ( ~n1010 & n8594 ) | ( n5687 & n8594 ) ;
  assign n8596 = ( ~n2114 & n2266 ) | ( ~n2114 & n8595 ) | ( n2266 & n8595 ) ;
  assign n8597 = ( n1796 & n5256 ) | ( n1796 & ~n8596 ) | ( n5256 & ~n8596 ) ;
  assign n8598 = n1189 & n4138 ;
  assign n8599 = n8597 & n8598 ;
  assign n8600 = n6752 ^ n384 ^ 1'b0 ;
  assign n8601 = n8600 ^ n6897 ^ n502 ;
  assign n8602 = ( ~n4529 & n6284 ) | ( ~n4529 & n8601 ) | ( n6284 & n8601 ) ;
  assign n8603 = ( n5490 & n7987 ) | ( n5490 & ~n8602 ) | ( n7987 & ~n8602 ) ;
  assign n8604 = n5421 ^ n3667 ^ n1980 ;
  assign n8605 = n8604 ^ n8288 ^ 1'b0 ;
  assign n8606 = n3504 ^ n3049 ^ n563 ;
  assign n8607 = ( n600 & ~n2271 ) | ( n600 & n4778 ) | ( ~n2271 & n4778 ) ;
  assign n8608 = n8607 ^ n5426 ^ n1642 ;
  assign n8609 = n8608 ^ n4613 ^ n1940 ;
  assign n8610 = n8609 ^ n4735 ^ 1'b0 ;
  assign n8611 = n8606 & ~n8610 ;
  assign n8612 = ( n1675 & n2672 ) | ( n1675 & ~n4492 ) | ( n2672 & ~n4492 ) ;
  assign n8613 = n8612 ^ n6413 ^ 1'b0 ;
  assign n8614 = n8611 & ~n8613 ;
  assign n8615 = n1598 & n2963 ;
  assign n8616 = n773 ^ x192 ^ 1'b0 ;
  assign n8617 = n2527 & ~n8616 ;
  assign n8618 = ~n433 & n4300 ;
  assign n8619 = n8618 ^ n2733 ^ 1'b0 ;
  assign n8620 = n8619 ^ n1838 ^ 1'b0 ;
  assign n8621 = n3948 & ~n8620 ;
  assign n8622 = ~n8617 & n8621 ;
  assign n8623 = n8622 ^ n8371 ^ 1'b0 ;
  assign n8624 = n8015 & ~n8623 ;
  assign n8625 = ~n2142 & n8624 ;
  assign n8626 = n3775 & n7550 ;
  assign n8627 = n8626 ^ n3408 ^ 1'b0 ;
  assign n8628 = n8627 ^ n3707 ^ n870 ;
  assign n8630 = n1689 & ~n4071 ;
  assign n8631 = n8630 ^ n3044 ^ 1'b0 ;
  assign n8629 = n1403 & ~n4196 ;
  assign n8632 = n8631 ^ n8629 ^ 1'b0 ;
  assign n8633 = ( n2085 & ~n3945 ) | ( n2085 & n5245 ) | ( ~n3945 & n5245 ) ;
  assign n8635 = n4249 ^ n2288 ^ 1'b0 ;
  assign n8636 = ~n2040 & n8635 ;
  assign n8634 = n7924 & ~n8059 ;
  assign n8637 = n8636 ^ n8634 ^ 1'b0 ;
  assign n8638 = ( ~n1061 & n7541 ) | ( ~n1061 & n8637 ) | ( n7541 & n8637 ) ;
  assign n8639 = n335 | n1352 ;
  assign n8640 = ( n4981 & ~n8638 ) | ( n4981 & n8639 ) | ( ~n8638 & n8639 ) ;
  assign n8641 = n8633 & ~n8640 ;
  assign n8642 = n8641 ^ n6204 ^ 1'b0 ;
  assign n8643 = x24 & ~n4674 ;
  assign n8644 = n8643 ^ n7749 ^ n500 ;
  assign n8645 = n8644 ^ n4601 ^ n910 ;
  assign n8646 = n6574 ^ n2394 ^ 1'b0 ;
  assign n8647 = n7065 | n8646 ;
  assign n8648 = ( n1353 & n7411 ) | ( n1353 & n8647 ) | ( n7411 & n8647 ) ;
  assign n8649 = n3261 ^ n1603 ^ n1097 ;
  assign n8650 = n930 & ~n2020 ;
  assign n8651 = ~n6667 & n8650 ;
  assign n8652 = ( n546 & n8649 ) | ( n546 & ~n8651 ) | ( n8649 & ~n8651 ) ;
  assign n8653 = ( ~n4067 & n5188 ) | ( ~n4067 & n8652 ) | ( n5188 & n8652 ) ;
  assign n8654 = n1052 & ~n2076 ;
  assign n8655 = n363 | n7003 ;
  assign n8656 = ( n2655 & n4922 ) | ( n2655 & n8655 ) | ( n4922 & n8655 ) ;
  assign n8658 = n3963 ^ n491 ^ n363 ;
  assign n8657 = n2184 & ~n4085 ;
  assign n8659 = n8658 ^ n8657 ^ n4471 ;
  assign n8660 = n5947 ^ n4801 ^ 1'b0 ;
  assign n8661 = n6039 & ~n8660 ;
  assign n8662 = n8659 & n8661 ;
  assign n8663 = ~n7369 & n8662 ;
  assign n8664 = n7468 ^ n3148 ^ 1'b0 ;
  assign n8665 = n2318 ^ n946 ^ 1'b0 ;
  assign n8666 = n995 & n8665 ;
  assign n8667 = n6919 ^ n2779 ^ 1'b0 ;
  assign n8668 = n450 | n5449 ;
  assign n8669 = n8668 ^ n3531 ^ 1'b0 ;
  assign n8670 = n8669 ^ n1063 ^ 1'b0 ;
  assign n8671 = ~n8667 & n8670 ;
  assign n8672 = ( ~n1446 & n2705 ) | ( ~n1446 & n3546 ) | ( n2705 & n3546 ) ;
  assign n8673 = n8672 ^ n5787 ^ n481 ;
  assign n8674 = n4271 & n8673 ;
  assign n8675 = n8674 ^ n3983 ^ n2889 ;
  assign n8676 = n2250 ^ n2196 ^ n1325 ;
  assign n8677 = ( ~n4746 & n8536 ) | ( ~n4746 & n8676 ) | ( n8536 & n8676 ) ;
  assign n8678 = n8010 | n8677 ;
  assign n8679 = n696 & ~n3529 ;
  assign n8680 = n3777 ^ n2589 ^ 1'b0 ;
  assign n8681 = n8680 ^ n2620 ^ 1'b0 ;
  assign n8683 = n1137 ^ x203 ^ 1'b0 ;
  assign n8682 = n6298 ^ n5507 ^ 1'b0 ;
  assign n8684 = n8683 ^ n8682 ^ n7650 ;
  assign n8685 = n1030 ^ n930 ^ 1'b0 ;
  assign n8686 = n682 & n8685 ;
  assign n8687 = ~n2769 & n8686 ;
  assign n8688 = n8687 ^ n4156 ^ 1'b0 ;
  assign n8690 = x66 & ~n2412 ;
  assign n8691 = n8690 ^ n949 ^ 1'b0 ;
  assign n8689 = ( n3783 & ~n4966 ) | ( n3783 & n6390 ) | ( ~n4966 & n6390 ) ;
  assign n8692 = n8691 ^ n8689 ^ x228 ;
  assign n8693 = n4674 ^ n1245 ^ x127 ;
  assign n8694 = n8693 ^ n5298 ^ n2631 ;
  assign n8695 = n1772 & n8694 ;
  assign n8696 = n8695 ^ n6329 ^ n2348 ;
  assign n8697 = n7407 ^ n615 ^ 1'b0 ;
  assign n8698 = n8696 & ~n8697 ;
  assign n8700 = n2720 ^ n1236 ^ n807 ;
  assign n8701 = ( n560 & ~n1881 ) | ( n560 & n8700 ) | ( ~n1881 & n8700 ) ;
  assign n8699 = ( n1401 & ~n4680 ) | ( n1401 & n5792 ) | ( ~n4680 & n5792 ) ;
  assign n8702 = n8701 ^ n8699 ^ 1'b0 ;
  assign n8704 = ( ~n385 & n1061 ) | ( ~n385 & n2176 ) | ( n1061 & n2176 ) ;
  assign n8703 = n4255 ^ n3314 ^ 1'b0 ;
  assign n8705 = n8704 ^ n8703 ^ n1231 ;
  assign n8706 = n6701 & ~n7997 ;
  assign n8707 = n6784 ^ n2248 ^ n1351 ;
  assign n8708 = n5659 | n6705 ;
  assign n8709 = n1367 & n3380 ;
  assign n8710 = n8709 ^ n7218 ^ 1'b0 ;
  assign n8711 = n8710 ^ n5460 ^ n860 ;
  assign n8712 = n6525 ^ n3140 ^ 1'b0 ;
  assign n8713 = x22 & ~n8712 ;
  assign n8714 = n3487 & n4779 ;
  assign n8715 = n1243 | n8714 ;
  assign n8716 = n1716 & ~n4889 ;
  assign n8718 = ( ~n2962 & n3923 ) | ( ~n2962 & n6015 ) | ( n3923 & n6015 ) ;
  assign n8719 = n8718 ^ n5899 ^ n3359 ;
  assign n8717 = ~n1362 & n6602 ;
  assign n8720 = n8719 ^ n8717 ^ 1'b0 ;
  assign n8722 = n2167 & ~n4696 ;
  assign n8723 = n8722 ^ n4346 ^ n1866 ;
  assign n8721 = n4504 ^ n3899 ^ n1863 ;
  assign n8724 = n8723 ^ n8721 ^ n2419 ;
  assign n8725 = n8724 ^ n7531 ^ n3590 ;
  assign n8726 = ( n640 & n1655 ) | ( n640 & n2160 ) | ( n1655 & n2160 ) ;
  assign n8727 = ( n2832 & n5407 ) | ( n2832 & n8726 ) | ( n5407 & n8726 ) ;
  assign n8728 = n5839 | n8727 ;
  assign n8729 = n8728 ^ n1137 ^ 1'b0 ;
  assign n8739 = ( n870 & n1073 ) | ( n870 & ~n3261 ) | ( n1073 & ~n3261 ) ;
  assign n8740 = ( x202 & n1469 ) | ( x202 & n8739 ) | ( n1469 & n8739 ) ;
  assign n8730 = n718 ^ x180 ^ 1'b0 ;
  assign n8731 = ( ~n883 & n7330 ) | ( ~n883 & n8730 ) | ( n7330 & n8730 ) ;
  assign n8732 = n1975 ^ x145 ^ 1'b0 ;
  assign n8733 = n8732 ^ n5899 ^ n4078 ;
  assign n8734 = n3136 | n8733 ;
  assign n8735 = ~n4990 & n8734 ;
  assign n8736 = n8735 ^ n3066 ^ 1'b0 ;
  assign n8737 = n8736 ^ n969 ^ 1'b0 ;
  assign n8738 = ~n8731 & n8737 ;
  assign n8741 = n8740 ^ n8738 ^ n432 ;
  assign n8742 = ( ~x146 & x176 ) | ( ~x146 & n3942 ) | ( x176 & n3942 ) ;
  assign n8743 = ( n5252 & ~n7747 ) | ( n5252 & n8742 ) | ( ~n7747 & n8742 ) ;
  assign n8744 = n6963 & ~n8743 ;
  assign n8745 = n5548 ^ n4378 ^ 1'b0 ;
  assign n8746 = ~n4786 & n8745 ;
  assign n8747 = n8744 & n8746 ;
  assign n8749 = n2644 ^ n1034 ^ 1'b0 ;
  assign n8750 = n3762 | n8749 ;
  assign n8751 = ( ~n4100 & n5956 ) | ( ~n4100 & n8750 ) | ( n5956 & n8750 ) ;
  assign n8752 = n8751 ^ n4486 ^ n2924 ;
  assign n8748 = n6106 ^ n3818 ^ n1970 ;
  assign n8753 = n8752 ^ n8748 ^ n1346 ;
  assign n8754 = n5972 ^ n3448 ^ n1305 ;
  assign n8755 = n8754 ^ n7182 ^ n3779 ;
  assign n8756 = n8755 ^ n5285 ^ n3476 ;
  assign n8757 = ( ~n1028 & n1585 ) | ( ~n1028 & n8756 ) | ( n1585 & n8756 ) ;
  assign n8758 = n523 | n7007 ;
  assign n8759 = n1796 & ~n8758 ;
  assign n8760 = n8759 ^ n4562 ^ 1'b0 ;
  assign n8761 = ~n6892 & n8760 ;
  assign n8762 = ( ~n2727 & n8757 ) | ( ~n2727 & n8761 ) | ( n8757 & n8761 ) ;
  assign n8769 = n1550 | n2536 ;
  assign n8770 = n2471 | n8769 ;
  assign n8771 = n8770 ^ n5724 ^ 1'b0 ;
  assign n8765 = n2138 & ~n8608 ;
  assign n8766 = n8765 ^ n3947 ^ 1'b0 ;
  assign n8767 = n8766 ^ n3645 ^ 1'b0 ;
  assign n8768 = n5643 & n8767 ;
  assign n8763 = n1295 ^ n932 ^ 1'b0 ;
  assign n8764 = n8763 ^ n3801 ^ n2152 ;
  assign n8772 = n8771 ^ n8768 ^ n8764 ;
  assign n8773 = n1603 | n6111 ;
  assign n8774 = ~n4851 & n8773 ;
  assign n8775 = n1888 & n5293 ;
  assign n8776 = n8216 ^ n5279 ^ 1'b0 ;
  assign n8777 = ~n8775 & n8776 ;
  assign n8778 = n4533 ^ n768 ^ 1'b0 ;
  assign n8779 = ( n579 & ~n883 ) | ( n579 & n1076 ) | ( ~n883 & n1076 ) ;
  assign n8780 = n7200 ^ n4599 ^ n3546 ;
  assign n8781 = ( n2617 & ~n8779 ) | ( n2617 & n8780 ) | ( ~n8779 & n8780 ) ;
  assign n8782 = ( n1518 & ~n8778 ) | ( n1518 & n8781 ) | ( ~n8778 & n8781 ) ;
  assign n8783 = n8782 ^ n3093 ^ 1'b0 ;
  assign n8784 = ~n2611 & n7648 ;
  assign n8785 = n946 | n1359 ;
  assign n8786 = ~n3141 & n4326 ;
  assign n8787 = ~n8785 & n8786 ;
  assign n8791 = ( n370 & ~n4831 ) | ( n370 & n6630 ) | ( ~n4831 & n6630 ) ;
  assign n8792 = n8791 ^ n6780 ^ n572 ;
  assign n8788 = n3145 ^ x57 ^ 1'b0 ;
  assign n8789 = n4018 & ~n8788 ;
  assign n8790 = ( ~n2434 & n3763 ) | ( ~n2434 & n8789 ) | ( n3763 & n8789 ) ;
  assign n8793 = n8792 ^ n8790 ^ n5741 ;
  assign n8794 = n8793 ^ n7346 ^ 1'b0 ;
  assign n8795 = ( n2176 & ~n6302 ) | ( n2176 & n8484 ) | ( ~n6302 & n8484 ) ;
  assign n8796 = n2288 ^ n1910 ^ n885 ;
  assign n8797 = n6575 ^ n4171 ^ n3498 ;
  assign n8798 = ( n2135 & ~n5737 ) | ( n2135 & n8797 ) | ( ~n5737 & n8797 ) ;
  assign n8799 = n8798 ^ n4378 ^ n1597 ;
  assign n8800 = n5060 | n5895 ;
  assign n8801 = n737 | n8800 ;
  assign n8802 = ( ~n1427 & n1599 ) | ( ~n1427 & n8801 ) | ( n1599 & n8801 ) ;
  assign n8803 = ( n3856 & n4312 ) | ( n3856 & ~n8802 ) | ( n4312 & ~n8802 ) ;
  assign n8805 = ( ~n326 & n4441 ) | ( ~n326 & n7393 ) | ( n4441 & n7393 ) ;
  assign n8804 = ( n1526 & n3560 ) | ( n1526 & n6139 ) | ( n3560 & n6139 ) ;
  assign n8806 = n8805 ^ n8804 ^ n4185 ;
  assign n8807 = ( n1846 & n5989 ) | ( n1846 & n7173 ) | ( n5989 & n7173 ) ;
  assign n8808 = n8806 | n8807 ;
  assign n8809 = ~n5930 & n8808 ;
  assign n8810 = n8803 & n8809 ;
  assign n8811 = ( n8796 & n8799 ) | ( n8796 & n8810 ) | ( n8799 & n8810 ) ;
  assign n8812 = n5376 ^ n3408 ^ 1'b0 ;
  assign n8813 = n7491 ^ n2553 ^ n2337 ;
  assign n8814 = n8812 & ~n8813 ;
  assign n8816 = n541 | n5697 ;
  assign n8815 = x169 & n2688 ;
  assign n8817 = n8816 ^ n8815 ^ 1'b0 ;
  assign n8818 = n4175 & n8284 ;
  assign n8819 = n8818 ^ n1865 ^ 1'b0 ;
  assign n8820 = n8819 ^ n2757 ^ n1478 ;
  assign n8821 = n8820 ^ n8805 ^ n6431 ;
  assign n8825 = ~n1101 & n1710 ;
  assign n8826 = n949 & n8825 ;
  assign n8823 = n3809 & ~n5567 ;
  assign n8824 = n8823 ^ n6532 ^ 1'b0 ;
  assign n8827 = n8826 ^ n8824 ^ n6305 ;
  assign n8828 = n8827 ^ n5192 ^ 1'b0 ;
  assign n8822 = ( ~n2148 & n4659 ) | ( ~n2148 & n6458 ) | ( n4659 & n6458 ) ;
  assign n8829 = n8828 ^ n8822 ^ 1'b0 ;
  assign n8830 = n8821 & n8829 ;
  assign n8834 = ( n3899 & n5223 ) | ( n3899 & n8701 ) | ( n5223 & n8701 ) ;
  assign n8831 = n1438 ^ n1096 ^ 1'b0 ;
  assign n8832 = n2735 | n8831 ;
  assign n8833 = n2954 & ~n8832 ;
  assign n8835 = n8834 ^ n8833 ^ 1'b0 ;
  assign n8836 = n1515 | n4785 ;
  assign n8837 = n914 & ~n2475 ;
  assign n8838 = n8837 ^ n3136 ^ 1'b0 ;
  assign n8839 = n5913 & n8838 ;
  assign n8840 = ~n1953 & n8839 ;
  assign n8841 = n8840 ^ n2625 ^ n1918 ;
  assign n8842 = ( x126 & n8836 ) | ( x126 & n8841 ) | ( n8836 & n8841 ) ;
  assign n8851 = n1138 | n1890 ;
  assign n8852 = n8851 ^ n7322 ^ n5133 ;
  assign n8850 = ~n3402 & n6532 ;
  assign n8853 = n8852 ^ n8850 ^ 1'b0 ;
  assign n8845 = n4020 ^ n3848 ^ 1'b0 ;
  assign n8846 = n5486 & n8845 ;
  assign n8847 = ( n786 & ~n2084 ) | ( n786 & n8846 ) | ( ~n2084 & n8846 ) ;
  assign n8843 = n2950 ^ n1184 ^ 1'b0 ;
  assign n8844 = n2428 & n8843 ;
  assign n8848 = n8847 ^ n8844 ^ 1'b0 ;
  assign n8849 = n1984 & ~n8848 ;
  assign n8854 = n8853 ^ n8849 ^ n3323 ;
  assign n8855 = ( ~n8835 & n8842 ) | ( ~n8835 & n8854 ) | ( n8842 & n8854 ) ;
  assign n8856 = ( n5288 & ~n5295 ) | ( n5288 & n7700 ) | ( ~n5295 & n7700 ) ;
  assign n8857 = ( n1156 & n3261 ) | ( n1156 & ~n6649 ) | ( n3261 & ~n6649 ) ;
  assign n8858 = ~n1361 & n4054 ;
  assign n8859 = n3484 ^ n1069 ^ n1014 ;
  assign n8860 = n7739 | n8859 ;
  assign n8861 = n8860 ^ n8627 ^ 1'b0 ;
  assign n8862 = ( n868 & n6120 ) | ( n868 & n8861 ) | ( n6120 & n8861 ) ;
  assign n8863 = ( ~n8857 & n8858 ) | ( ~n8857 & n8862 ) | ( n8858 & n8862 ) ;
  assign n8867 = n7642 ^ n1403 ^ 1'b0 ;
  assign n8868 = n5269 & n5890 ;
  assign n8869 = n8867 & n8868 ;
  assign n8870 = n7280 & ~n8869 ;
  assign n8864 = n4405 & ~n5666 ;
  assign n8865 = n3143 ^ n2549 ^ n289 ;
  assign n8866 = n8864 | n8865 ;
  assign n8871 = n8870 ^ n8866 ^ 1'b0 ;
  assign n8880 = n1773 & n3475 ;
  assign n8881 = n8843 ^ n795 ^ n329 ;
  assign n8882 = ( n2983 & n8880 ) | ( n2983 & ~n8881 ) | ( n8880 & ~n8881 ) ;
  assign n8883 = n8882 ^ n6596 ^ n4613 ;
  assign n8884 = n8883 ^ n3798 ^ 1'b0 ;
  assign n8877 = n3007 ^ n1504 ^ x107 ;
  assign n8872 = n2806 & ~n7616 ;
  assign n8873 = n8872 ^ n7270 ^ 1'b0 ;
  assign n8874 = ~n2240 & n5460 ;
  assign n8875 = n8874 ^ n5783 ^ 1'b0 ;
  assign n8876 = ~n8873 & n8875 ;
  assign n8878 = n8877 ^ n8876 ^ n7393 ;
  assign n8879 = n1653 & ~n8878 ;
  assign n8885 = n8884 ^ n8879 ^ 1'b0 ;
  assign n8886 = n1156 ^ n327 ^ 1'b0 ;
  assign n8887 = n8886 ^ n672 ^ 1'b0 ;
  assign n8888 = n8887 ^ n5880 ^ n4049 ;
  assign n8889 = n446 & ~n5947 ;
  assign n8890 = n8889 ^ n7212 ^ 1'b0 ;
  assign n8891 = n3971 & n8179 ;
  assign n8892 = n8891 ^ n7743 ^ n1387 ;
  assign n8893 = n8592 ^ n6562 ^ 1'b0 ;
  assign n8894 = ( ~n3796 & n8007 ) | ( ~n3796 & n8893 ) | ( n8007 & n8893 ) ;
  assign n8895 = n4027 ^ n2362 ^ n1814 ;
  assign n8896 = n6416 & n8895 ;
  assign n8897 = n962 & ~n2141 ;
  assign n8898 = ( n7903 & n8896 ) | ( n7903 & ~n8897 ) | ( n8896 & ~n8897 ) ;
  assign n8899 = ( n4094 & n8101 ) | ( n4094 & n8898 ) | ( n8101 & n8898 ) ;
  assign n8901 = n7629 ^ n2154 ^ 1'b0 ;
  assign n8900 = ( n3991 & n6334 ) | ( n3991 & n8338 ) | ( n6334 & n8338 ) ;
  assign n8902 = n8901 ^ n8900 ^ n4071 ;
  assign n8903 = n6503 ^ n2042 ^ n1314 ;
  assign n8904 = ( n1610 & n1802 ) | ( n1610 & ~n2799 ) | ( n1802 & ~n2799 ) ;
  assign n8905 = n4428 & n8904 ;
  assign n8906 = n3016 & n8905 ;
  assign n8907 = n6031 & n8580 ;
  assign n8908 = n830 & ~n888 ;
  assign n8909 = n911 & n8908 ;
  assign n8910 = n8909 ^ n1979 ^ 1'b0 ;
  assign n8911 = n1203 | n8910 ;
  assign n8912 = n3381 & ~n8911 ;
  assign n8913 = ~n8907 & n8912 ;
  assign n8914 = ( n713 & n8906 ) | ( n713 & ~n8913 ) | ( n8906 & ~n8913 ) ;
  assign n8916 = ~n647 & n6319 ;
  assign n8917 = n8916 ^ n2404 ^ 1'b0 ;
  assign n8915 = ( ~n551 & n3069 ) | ( ~n551 & n6158 ) | ( n3069 & n6158 ) ;
  assign n8918 = n8917 ^ n8915 ^ 1'b0 ;
  assign n8919 = ~n4390 & n8918 ;
  assign n8920 = n1685 & n8919 ;
  assign n8921 = ( ~n2453 & n3643 ) | ( ~n2453 & n8920 ) | ( n3643 & n8920 ) ;
  assign n8922 = ( n8903 & n8914 ) | ( n8903 & ~n8921 ) | ( n8914 & ~n8921 ) ;
  assign n8923 = n8922 ^ n4006 ^ n1260 ;
  assign n8924 = n570 & ~n3536 ;
  assign n8925 = n7520 ^ n639 ^ 1'b0 ;
  assign n8926 = ( n1739 & n1775 ) | ( n1739 & n2422 ) | ( n1775 & n2422 ) ;
  assign n8927 = ( n4390 & n5821 ) | ( n4390 & ~n8926 ) | ( n5821 & ~n8926 ) ;
  assign n8928 = n8927 ^ n7590 ^ 1'b0 ;
  assign n8929 = n3094 ^ n2866 ^ n1040 ;
  assign n8930 = n6049 | n8929 ;
  assign n8931 = n8930 ^ n7490 ^ 1'b0 ;
  assign n8932 = n1969 ^ n1354 ^ n1200 ;
  assign n8933 = n3252 & n3515 ;
  assign n8934 = n3172 | n7325 ;
  assign n8935 = n1296 & ~n8934 ;
  assign n8936 = n5609 ^ n1381 ^ 1'b0 ;
  assign n8937 = n8935 | n8936 ;
  assign n8938 = n2123 & ~n8937 ;
  assign n8939 = n8597 & n8938 ;
  assign n8940 = ( n1393 & n2433 ) | ( n1393 & n3785 ) | ( n2433 & n3785 ) ;
  assign n8941 = n8940 ^ n3604 ^ 1'b0 ;
  assign n8942 = n2824 ^ n536 ^ x81 ;
  assign n8943 = n8942 ^ n1105 ^ 1'b0 ;
  assign n8944 = ( n1935 & n3112 ) | ( n1935 & n8943 ) | ( n3112 & n8943 ) ;
  assign n8945 = n8944 ^ n8043 ^ n1791 ;
  assign n8946 = n1772 & ~n8945 ;
  assign n8947 = ( n3076 & n5227 ) | ( n3076 & n8508 ) | ( n5227 & n8508 ) ;
  assign n8948 = n2520 ^ n683 ^ 1'b0 ;
  assign n8949 = ~n2705 & n8948 ;
  assign n8950 = n4816 & n8949 ;
  assign n8951 = ~n8947 & n8950 ;
  assign n8952 = n7659 ^ n6737 ^ n4113 ;
  assign n8953 = n3811 | n5426 ;
  assign n8954 = n8952 & ~n8953 ;
  assign n8955 = n8954 ^ n1628 ^ n1266 ;
  assign n8956 = n7456 ^ n5129 ^ 1'b0 ;
  assign n8957 = ( ~n454 & n3728 ) | ( ~n454 & n8331 ) | ( n3728 & n8331 ) ;
  assign n8958 = n8957 ^ n7892 ^ n1609 ;
  assign n8959 = n4045 & ~n8958 ;
  assign n8973 = ( n1872 & n2797 ) | ( n1872 & n2869 ) | ( n2797 & n2869 ) ;
  assign n8960 = n5218 ^ n5101 ^ 1'b0 ;
  assign n8967 = x163 & ~n3899 ;
  assign n8968 = n8967 ^ n1258 ^ 1'b0 ;
  assign n8966 = ( ~n1018 & n3181 ) | ( ~n1018 & n7269 ) | ( n3181 & n7269 ) ;
  assign n8964 = ~n4180 & n4370 ;
  assign n8963 = n337 | n2866 ;
  assign n8965 = n8964 ^ n8963 ^ 1'b0 ;
  assign n8969 = n8968 ^ n8966 ^ n8965 ;
  assign n8961 = x182 & n1497 ;
  assign n8962 = n4572 & n8961 ;
  assign n8970 = n8969 ^ n8962 ^ n2593 ;
  assign n8971 = n8960 & n8970 ;
  assign n8972 = ~n4206 & n8971 ;
  assign n8974 = n8973 ^ n8972 ^ 1'b0 ;
  assign n8975 = n8959 & n8974 ;
  assign n8977 = n2466 ^ n630 ^ 1'b0 ;
  assign n8978 = n1803 | n8977 ;
  assign n8979 = n8978 ^ n3891 ^ n1375 ;
  assign n8980 = ( x12 & ~n3352 ) | ( x12 & n8979 ) | ( ~n3352 & n8979 ) ;
  assign n8981 = n2523 ^ n2131 ^ 1'b0 ;
  assign n8982 = n8980 & n8981 ;
  assign n8976 = n2750 & ~n5430 ;
  assign n8983 = n8982 ^ n8976 ^ 1'b0 ;
  assign n8987 = n4173 ^ n3474 ^ n1922 ;
  assign n8984 = n1089 ^ n678 ^ 1'b0 ;
  assign n8985 = n8984 ^ n570 ^ 1'b0 ;
  assign n8986 = ( n3764 & ~n6025 ) | ( n3764 & n8985 ) | ( ~n6025 & n8985 ) ;
  assign n8988 = n8987 ^ n8986 ^ n2335 ;
  assign n8989 = x59 & ~n8988 ;
  assign n8990 = n8989 ^ n5667 ^ 1'b0 ;
  assign n8991 = ( ~n4591 & n8983 ) | ( ~n4591 & n8990 ) | ( n8983 & n8990 ) ;
  assign n8996 = ~n401 & n2448 ;
  assign n8993 = n6667 ^ n3753 ^ 1'b0 ;
  assign n8994 = n1288 & ~n8993 ;
  assign n8995 = ( ~n1163 & n6716 ) | ( ~n1163 & n8994 ) | ( n6716 & n8994 ) ;
  assign n8992 = ( x82 & ~n2191 ) | ( x82 & n5731 ) | ( ~n2191 & n5731 ) ;
  assign n8997 = n8996 ^ n8995 ^ n8992 ;
  assign n8998 = ( n4495 & ~n4893 ) | ( n4495 & n5333 ) | ( ~n4893 & n5333 ) ;
  assign n8999 = n2577 & n6242 ;
  assign n9000 = ( n1472 & ~n5099 ) | ( n1472 & n8480 ) | ( ~n5099 & n8480 ) ;
  assign n9001 = n933 & ~n5881 ;
  assign n9002 = n3670 ^ n1651 ^ 1'b0 ;
  assign n9003 = n6963 ^ n2525 ^ 1'b0 ;
  assign n9006 = n3663 ^ n1183 ^ 1'b0 ;
  assign n9007 = ~n8649 & n9006 ;
  assign n9004 = n5913 & ~n8909 ;
  assign n9005 = n9004 ^ n4598 ^ 1'b0 ;
  assign n9008 = n9007 ^ n9005 ^ 1'b0 ;
  assign n9009 = n1861 | n9008 ;
  assign n9010 = n8085 ^ n1955 ^ 1'b0 ;
  assign n9011 = n9010 ^ n4448 ^ n1073 ;
  assign n9020 = n2850 ^ n1100 ^ 1'b0 ;
  assign n9021 = n750 | n9020 ;
  assign n9022 = ( x100 & ~n6472 ) | ( x100 & n9021 ) | ( ~n6472 & n9021 ) ;
  assign n9023 = ( n2085 & ~n5415 ) | ( n2085 & n7961 ) | ( ~n5415 & n7961 ) ;
  assign n9024 = n9023 ^ n3815 ^ 1'b0 ;
  assign n9025 = x187 & n9024 ;
  assign n9026 = ( n6151 & n9022 ) | ( n6151 & n9025 ) | ( n9022 & n9025 ) ;
  assign n9027 = ( ~n3817 & n5753 ) | ( ~n3817 & n7195 ) | ( n5753 & n7195 ) ;
  assign n9028 = n9026 & ~n9027 ;
  assign n9012 = ( n2070 & ~n2498 ) | ( n2070 & n3611 ) | ( ~n2498 & n3611 ) ;
  assign n9013 = ( n5299 & n5970 ) | ( n5299 & n9012 ) | ( n5970 & n9012 ) ;
  assign n9014 = ( n807 & n7443 ) | ( n807 & ~n9013 ) | ( n7443 & ~n9013 ) ;
  assign n9015 = n737 & ~n3281 ;
  assign n9016 = ~n2402 & n9015 ;
  assign n9017 = n9016 ^ n3234 ^ 1'b0 ;
  assign n9018 = n9017 ^ n4032 ^ n3981 ;
  assign n9019 = ( n8616 & n9014 ) | ( n8616 & n9018 ) | ( n9014 & n9018 ) ;
  assign n9029 = n9028 ^ n9019 ^ n2820 ;
  assign n9030 = n3322 ^ n1659 ^ 1'b0 ;
  assign n9031 = n5520 | n9030 ;
  assign n9032 = n4053 & ~n9031 ;
  assign n9033 = ~n6428 & n9032 ;
  assign n9034 = n6519 ^ n5299 ^ 1'b0 ;
  assign n9035 = ~n6257 & n9034 ;
  assign n9036 = n9035 ^ n2638 ^ n707 ;
  assign n9041 = n1511 ^ n1195 ^ 1'b0 ;
  assign n9042 = n9041 ^ n5275 ^ 1'b0 ;
  assign n9037 = n8778 ^ n1000 ^ n490 ;
  assign n9038 = n2539 & n9037 ;
  assign n9039 = n9038 ^ n8177 ^ 1'b0 ;
  assign n9040 = ( ~x116 & n3186 ) | ( ~x116 & n9039 ) | ( n3186 & n9039 ) ;
  assign n9043 = n9042 ^ n9040 ^ n5279 ;
  assign n9044 = n9043 ^ n1202 ^ 1'b0 ;
  assign n9045 = ( n1747 & ~n5426 ) | ( n1747 & n8722 ) | ( ~n5426 & n8722 ) ;
  assign n9046 = n5782 ^ n5346 ^ n2735 ;
  assign n9047 = ( n3512 & ~n4661 ) | ( n3512 & n9046 ) | ( ~n4661 & n9046 ) ;
  assign n9048 = n4962 ^ x103 ^ 1'b0 ;
  assign n9049 = ( n6451 & n9047 ) | ( n6451 & ~n9048 ) | ( n9047 & ~n9048 ) ;
  assign n9050 = n7423 ^ n1900 ^ 1'b0 ;
  assign n9051 = n4793 ^ n3113 ^ 1'b0 ;
  assign n9052 = ( n1793 & n8449 ) | ( n1793 & n8562 ) | ( n8449 & n8562 ) ;
  assign n9053 = n662 | n967 ;
  assign n9054 = ~n448 & n9053 ;
  assign n9055 = n9054 ^ n1891 ^ 1'b0 ;
  assign n9057 = ~n630 & n2194 ;
  assign n9058 = ~n5005 & n9057 ;
  assign n9056 = n2346 ^ x115 ^ 1'b0 ;
  assign n9059 = n9058 ^ n9056 ^ 1'b0 ;
  assign n9060 = n9059 ^ n541 ^ 1'b0 ;
  assign n9061 = n1870 & ~n9060 ;
  assign n9062 = ( n7500 & n9055 ) | ( n7500 & ~n9061 ) | ( n9055 & ~n9061 ) ;
  assign n9068 = ~n624 & n1851 ;
  assign n9069 = n9068 ^ n642 ^ 1'b0 ;
  assign n9067 = ( ~n1370 & n1553 ) | ( ~n1370 & n6357 ) | ( n1553 & n6357 ) ;
  assign n9063 = n6183 ^ n3397 ^ n1272 ;
  assign n9064 = n1974 & n9063 ;
  assign n9065 = n2635 & ~n9064 ;
  assign n9066 = n9065 ^ n4862 ^ 1'b0 ;
  assign n9070 = n9069 ^ n9067 ^ n9066 ;
  assign n9071 = n1076 & ~n1812 ;
  assign n9072 = n7317 ^ n4075 ^ 1'b0 ;
  assign n9073 = n3470 ^ n2471 ^ 1'b0 ;
  assign n9074 = ( ~n2874 & n9072 ) | ( ~n2874 & n9073 ) | ( n9072 & n9073 ) ;
  assign n9075 = ( n1419 & n1683 ) | ( n1419 & n6006 ) | ( n1683 & n6006 ) ;
  assign n9076 = n9075 ^ n2664 ^ n1991 ;
  assign n9077 = n1668 & ~n6437 ;
  assign n9078 = n9077 ^ n1832 ^ n488 ;
  assign n9079 = n2529 & n9078 ;
  assign n9080 = ~n2425 & n9079 ;
  assign n9081 = n7376 ^ n6785 ^ 1'b0 ;
  assign n9082 = ( n824 & n6253 ) | ( n824 & n9081 ) | ( n6253 & n9081 ) ;
  assign n9089 = ~n784 & n793 ;
  assign n9090 = n9089 ^ n7697 ^ n5245 ;
  assign n9085 = ( ~x190 & n2614 ) | ( ~x190 & n4709 ) | ( n2614 & n4709 ) ;
  assign n9083 = n6748 ^ n3193 ^ n2720 ;
  assign n9084 = n9083 ^ n7344 ^ n309 ;
  assign n9086 = n9085 ^ n9084 ^ n1941 ;
  assign n9087 = n4441 ^ n4014 ^ n1416 ;
  assign n9088 = n9086 & n9087 ;
  assign n9091 = n9090 ^ n9088 ^ 1'b0 ;
  assign n9092 = n1643 ^ n1010 ^ n774 ;
  assign n9093 = ~n2907 & n9092 ;
  assign n9094 = n9093 ^ n3198 ^ 1'b0 ;
  assign n9095 = n926 | n1534 ;
  assign n9096 = n9095 ^ n1787 ^ 1'b0 ;
  assign n9097 = n4908 | n9096 ;
  assign n9098 = n6912 | n9097 ;
  assign n9099 = ~n3444 & n9098 ;
  assign n9100 = n9094 & n9099 ;
  assign n9101 = n9100 ^ n4983 ^ n2404 ;
  assign n9102 = n3798 ^ n2126 ^ n1222 ;
  assign n9103 = n9102 ^ n4298 ^ 1'b0 ;
  assign n9104 = n1217 & ~n6940 ;
  assign n9110 = n974 | n3253 ;
  assign n9111 = n3253 & ~n9110 ;
  assign n9112 = n317 & ~n9111 ;
  assign n9105 = ~n279 & n841 ;
  assign n9106 = ~n841 & n9105 ;
  assign n9107 = n1105 | n5845 ;
  assign n9108 = n9107 ^ n2569 ^ 1'b0 ;
  assign n9109 = n9106 | n9108 ;
  assign n9113 = n9112 ^ n9109 ^ n1686 ;
  assign n9114 = n4204 ^ n2453 ^ n551 ;
  assign n9115 = n857 | n9114 ;
  assign n9116 = n2602 ^ n1560 ^ n1382 ;
  assign n9117 = ( x130 & x144 ) | ( x130 & ~n3807 ) | ( x144 & ~n3807 ) ;
  assign n9118 = ( ~n3272 & n8978 ) | ( ~n3272 & n9117 ) | ( n8978 & n9117 ) ;
  assign n9119 = n7926 ^ n4522 ^ 1'b0 ;
  assign n9120 = n9119 ^ n7193 ^ n4800 ;
  assign n9121 = n2945 ^ n2924 ^ n1337 ;
  assign n9122 = ( x180 & n8036 ) | ( x180 & ~n9121 ) | ( n8036 & ~n9121 ) ;
  assign n9123 = n2600 & ~n6219 ;
  assign n9124 = n7178 & n9123 ;
  assign n9130 = ( x125 & n1888 ) | ( x125 & ~n3844 ) | ( n1888 & ~n3844 ) ;
  assign n9129 = ~n1984 & n2349 ;
  assign n9131 = n9130 ^ n9129 ^ 1'b0 ;
  assign n9125 = ( n634 & n1079 ) | ( n634 & ~n2733 ) | ( n1079 & ~n2733 ) ;
  assign n9126 = n3561 ^ n2557 ^ n1790 ;
  assign n9127 = n9125 | n9126 ;
  assign n9128 = n5853 | n9127 ;
  assign n9132 = n9131 ^ n9128 ^ n1095 ;
  assign n9133 = ~n2847 & n9132 ;
  assign n9134 = ~n1086 & n9133 ;
  assign n9135 = n3157 ^ x156 ^ x88 ;
  assign n9136 = ( n905 & ~n962 ) | ( n905 & n7612 ) | ( ~n962 & n7612 ) ;
  assign n9137 = n3374 & n9136 ;
  assign n9138 = n9135 & n9137 ;
  assign n9139 = ( x165 & ~n3525 ) | ( x165 & n9138 ) | ( ~n3525 & n9138 ) ;
  assign n9140 = n6279 ^ n3807 ^ n890 ;
  assign n9141 = n9139 & n9140 ;
  assign n9142 = n9141 ^ n1086 ^ 1'b0 ;
  assign n9143 = n9134 | n9142 ;
  assign n9144 = x51 & n5084 ;
  assign n9145 = n9144 ^ n5038 ^ 1'b0 ;
  assign n9146 = ( n1061 & ~n3798 ) | ( n1061 & n9145 ) | ( ~n3798 & n9145 ) ;
  assign n9147 = ( ~n4696 & n7705 ) | ( ~n4696 & n8130 ) | ( n7705 & n8130 ) ;
  assign n9148 = n9147 ^ n5646 ^ n3391 ;
  assign n9149 = ~n3410 & n3512 ;
  assign n9150 = n7150 ^ n6686 ^ n5622 ;
  assign n9152 = n1077 & ~n3520 ;
  assign n9153 = n9152 ^ n1309 ^ 1'b0 ;
  assign n9154 = ( n3273 & n4053 ) | ( n3273 & n9153 ) | ( n4053 & n9153 ) ;
  assign n9151 = n4522 ^ n2012 ^ 1'b0 ;
  assign n9155 = n9154 ^ n9151 ^ n1587 ;
  assign n9156 = n9155 ^ n4471 ^ x103 ;
  assign n9157 = n8740 ^ x34 ^ 1'b0 ;
  assign n9158 = x105 & ~n9157 ;
  assign n9159 = ~n3458 & n9158 ;
  assign n9160 = ( n1677 & n2008 ) | ( n1677 & ~n9159 ) | ( n2008 & ~n9159 ) ;
  assign n9161 = n6904 ^ n4225 ^ x169 ;
  assign n9162 = n957 & n9161 ;
  assign n9163 = n9160 & ~n9162 ;
  assign n9164 = ~n5629 & n9163 ;
  assign n9165 = n2700 | n8874 ;
  assign n9166 = n1508 | n9165 ;
  assign n9169 = n946 & ~n2901 ;
  assign n9170 = n1803 & n9169 ;
  assign n9171 = n9170 ^ n8213 ^ 1'b0 ;
  assign n9167 = n4709 ^ n4053 ^ x137 ;
  assign n9168 = ~n8895 & n9167 ;
  assign n9172 = n9171 ^ n9168 ^ 1'b0 ;
  assign n9173 = n7786 ^ n4930 ^ n2415 ;
  assign n9174 = n6163 ^ n3105 ^ n520 ;
  assign n9175 = x198 | n9174 ;
  assign n9176 = ( n1475 & ~n5623 ) | ( n1475 & n9175 ) | ( ~n5623 & n9175 ) ;
  assign n9177 = ( n2998 & n3544 ) | ( n2998 & ~n4606 ) | ( n3544 & ~n4606 ) ;
  assign n9178 = ( n2347 & ~n7270 ) | ( n2347 & n9177 ) | ( ~n7270 & n9177 ) ;
  assign n9179 = n9178 ^ n3090 ^ n2117 ;
  assign n9180 = n6691 ^ n4696 ^ n672 ;
  assign n9181 = x73 & n1794 ;
  assign n9182 = n9181 ^ n2233 ^ 1'b0 ;
  assign n9183 = n3821 & n6399 ;
  assign n9184 = ~x8 & n9183 ;
  assign n9185 = ( n2864 & n8341 ) | ( n2864 & ~n9184 ) | ( n8341 & ~n9184 ) ;
  assign n9192 = ( n2706 & n3565 ) | ( n2706 & ~n8732 ) | ( n3565 & ~n8732 ) ;
  assign n9186 = n525 | n2079 ;
  assign n9187 = n2942 & ~n9186 ;
  assign n9188 = n1709 & n9187 ;
  assign n9189 = ( x95 & n8580 ) | ( x95 & n9188 ) | ( n8580 & n9188 ) ;
  assign n9190 = n9189 ^ n2064 ^ 1'b0 ;
  assign n9191 = ~n4524 & n9190 ;
  assign n9193 = n9192 ^ n9191 ^ n8768 ;
  assign n9194 = ( n9182 & ~n9185 ) | ( n9182 & n9193 ) | ( ~n9185 & n9193 ) ;
  assign n9195 = n5086 ^ n1475 ^ 1'b0 ;
  assign n9201 = n7708 ^ n5863 ^ n1145 ;
  assign n9196 = ~n686 & n4443 ;
  assign n9197 = n7900 & n9196 ;
  assign n9198 = n1733 & ~n4950 ;
  assign n9199 = n9198 ^ n9014 ^ 1'b0 ;
  assign n9200 = ( ~n9130 & n9197 ) | ( ~n9130 & n9199 ) | ( n9197 & n9199 ) ;
  assign n9202 = n9201 ^ n9200 ^ 1'b0 ;
  assign n9203 = n9195 & n9202 ;
  assign n9204 = n2714 ^ n2595 ^ n2476 ;
  assign n9205 = ( n1968 & ~n7588 ) | ( n1968 & n9204 ) | ( ~n7588 & n9204 ) ;
  assign n9206 = n9205 ^ n8778 ^ 1'b0 ;
  assign n9207 = x87 & x158 ;
  assign n9208 = n9207 ^ x81 ^ 1'b0 ;
  assign n9209 = n4734 ^ n2273 ^ 1'b0 ;
  assign n9210 = n3026 & n9209 ;
  assign n9211 = n1391 ^ n1102 ^ 1'b0 ;
  assign n9212 = n9211 ^ n8995 ^ n3906 ;
  assign n9213 = ( n9208 & ~n9210 ) | ( n9208 & n9212 ) | ( ~n9210 & n9212 ) ;
  assign n9214 = n2520 ^ n2455 ^ n271 ;
  assign n9215 = n6523 | n9214 ;
  assign n9216 = n9213 & ~n9215 ;
  assign n9217 = n6007 & ~n9216 ;
  assign n9218 = n7928 ^ n2753 ^ 1'b0 ;
  assign n9219 = n9218 ^ n5458 ^ 1'b0 ;
  assign n9220 = n2769 ^ n851 ^ x208 ;
  assign n9221 = ( n6236 & n9148 ) | ( n6236 & ~n9220 ) | ( n9148 & ~n9220 ) ;
  assign n9222 = n290 | n1979 ;
  assign n9223 = ( n1280 & n3897 ) | ( n1280 & n9222 ) | ( n3897 & n9222 ) ;
  assign n9224 = n9223 ^ n2895 ^ 1'b0 ;
  assign n9225 = n2817 & ~n9224 ;
  assign n9226 = n6662 ^ n6557 ^ 1'b0 ;
  assign n9227 = n5713 & ~n6002 ;
  assign n9228 = n1722 ^ n1703 ^ 1'b0 ;
  assign n9229 = n2169 | n9228 ;
  assign n9230 = n4844 ^ n930 ^ 1'b0 ;
  assign n9231 = n5373 ^ n3609 ^ n3484 ;
  assign n9232 = ( n2814 & ~n9230 ) | ( n2814 & n9231 ) | ( ~n9230 & n9231 ) ;
  assign n9233 = ( n8196 & n9229 ) | ( n8196 & ~n9232 ) | ( n9229 & ~n9232 ) ;
  assign n9234 = n9233 ^ n8528 ^ n1732 ;
  assign n9235 = ( n1077 & n1343 ) | ( n1077 & n2319 ) | ( n1343 & n2319 ) ;
  assign n9236 = n6074 ^ n3992 ^ 1'b0 ;
  assign n9237 = n1200 & n9236 ;
  assign n9238 = ( n2180 & n5542 ) | ( n2180 & n9237 ) | ( n5542 & n9237 ) ;
  assign n9239 = n9235 & n9238 ;
  assign n9240 = n1141 & n9239 ;
  assign n9241 = n4619 ^ n2817 ^ 1'b0 ;
  assign n9242 = n9240 | n9241 ;
  assign n9243 = ~n4762 & n9212 ;
  assign n9244 = n9242 & n9243 ;
  assign n9245 = n544 | n6406 ;
  assign n9246 = n6353 | n9245 ;
  assign n9247 = n5055 ^ n3198 ^ n3162 ;
  assign n9248 = n2932 ^ n950 ^ 1'b0 ;
  assign n9249 = ~n615 & n9248 ;
  assign n9250 = n9249 ^ n6785 ^ 1'b0 ;
  assign n9251 = n7657 | n9250 ;
  assign n9252 = n9247 | n9251 ;
  assign n9253 = ~n1138 & n4650 ;
  assign n9254 = n3353 ^ n872 ^ 1'b0 ;
  assign n9255 = n6183 ^ n5799 ^ 1'b0 ;
  assign n9256 = n4975 & n9255 ;
  assign n9257 = ( n356 & ~n4109 ) | ( n356 & n5598 ) | ( ~n4109 & n5598 ) ;
  assign n9258 = ( n1961 & n2638 ) | ( n1961 & ~n9257 ) | ( n2638 & ~n9257 ) ;
  assign n9259 = ( n434 & ~n5069 ) | ( n434 & n9258 ) | ( ~n5069 & n9258 ) ;
  assign n9260 = n7424 & n9259 ;
  assign n9261 = ( n3504 & ~n4502 ) | ( n3504 & n6209 ) | ( ~n4502 & n6209 ) ;
  assign n9262 = ( ~n3313 & n8579 ) | ( ~n3313 & n9261 ) | ( n8579 & n9261 ) ;
  assign n9263 = n5890 & ~n9262 ;
  assign n9266 = n6639 ^ n5799 ^ n893 ;
  assign n9265 = n1419 & n6083 ;
  assign n9267 = n9266 ^ n9265 ^ 1'b0 ;
  assign n9268 = ( n1208 & n1677 ) | ( n1208 & n9267 ) | ( n1677 & n9267 ) ;
  assign n9264 = n2817 & ~n3214 ;
  assign n9269 = n9268 ^ n9264 ^ n8779 ;
  assign n9270 = ( n518 & n2229 ) | ( n518 & ~n6248 ) | ( n2229 & ~n6248 ) ;
  assign n9271 = ( n690 & ~n3609 ) | ( n690 & n7828 ) | ( ~n3609 & n7828 ) ;
  assign n9272 = ( n4375 & ~n7911 ) | ( n4375 & n9271 ) | ( ~n7911 & n9271 ) ;
  assign n9273 = ( n421 & n1248 ) | ( n421 & n3326 ) | ( n1248 & n3326 ) ;
  assign n9274 = n6878 & ~n9273 ;
  assign n9275 = n9274 ^ n5050 ^ 1'b0 ;
  assign n9276 = ( n1980 & ~n3867 ) | ( n1980 & n9275 ) | ( ~n3867 & n9275 ) ;
  assign n9277 = n754 & ~n791 ;
  assign n9278 = ( ~n5446 & n6355 ) | ( ~n5446 & n9277 ) | ( n6355 & n9277 ) ;
  assign n9279 = n3122 | n6532 ;
  assign n9280 = ( n2515 & n5278 ) | ( n2515 & n6448 ) | ( n5278 & n6448 ) ;
  assign n9281 = x192 | n9280 ;
  assign n9282 = ~n9279 & n9281 ;
  assign n9283 = n3540 ^ n898 ^ 1'b0 ;
  assign n9284 = n9283 ^ n4362 ^ 1'b0 ;
  assign n9285 = n9282 & ~n9284 ;
  assign n9286 = ~n1526 & n9285 ;
  assign n9287 = n9278 & ~n9286 ;
  assign n9289 = n1648 | n8750 ;
  assign n9290 = n9289 ^ n1573 ^ 1'b0 ;
  assign n9291 = n9290 ^ n3190 ^ 1'b0 ;
  assign n9288 = n6298 ^ n5913 ^ 1'b0 ;
  assign n9292 = n9291 ^ n9288 ^ 1'b0 ;
  assign n9293 = x177 & ~n5226 ;
  assign n9294 = n2365 & n9293 ;
  assign n9295 = n9294 ^ n7743 ^ n6888 ;
  assign n9296 = n1708 | n9295 ;
  assign n9297 = n1867 & ~n2895 ;
  assign n9298 = n5779 | n9297 ;
  assign n9299 = ~n1713 & n2010 ;
  assign n9300 = n1277 & ~n6448 ;
  assign n9301 = ~n9299 & n9300 ;
  assign n9302 = n7276 ^ n2627 ^ 1'b0 ;
  assign n9303 = n9301 | n9302 ;
  assign n9304 = n7073 ^ n962 ^ 1'b0 ;
  assign n9305 = ( n303 & ~n6116 ) | ( n303 & n9304 ) | ( ~n6116 & n9304 ) ;
  assign n9306 = n4713 & ~n9305 ;
  assign n9310 = ( n307 & n2908 ) | ( n307 & n4410 ) | ( n2908 & n4410 ) ;
  assign n9311 = n2726 & n9310 ;
  assign n9312 = n9311 ^ n3514 ^ x126 ;
  assign n9307 = n5269 & n7536 ;
  assign n9308 = n9307 ^ n7966 ^ 1'b0 ;
  assign n9309 = ~n8774 & n9308 ;
  assign n9313 = n9312 ^ n9309 ^ 1'b0 ;
  assign n9314 = n2418 ^ x221 ^ 1'b0 ;
  assign n9315 = n8749 ^ n4179 ^ 1'b0 ;
  assign n9316 = ~n9314 & n9315 ;
  assign n9317 = n9316 ^ n333 ^ 1'b0 ;
  assign n9318 = ( n1307 & n6472 ) | ( n1307 & ~n6774 ) | ( n6472 & ~n6774 ) ;
  assign n9319 = n4566 | n5350 ;
  assign n9320 = n9319 ^ n1454 ^ 1'b0 ;
  assign n9321 = n7277 ^ n5183 ^ n436 ;
  assign n9322 = n9320 | n9321 ;
  assign n9323 = ~n2990 & n5783 ;
  assign n9327 = n750 | n4623 ;
  assign n9328 = n1478 | n9327 ;
  assign n9324 = n6159 ^ n750 ^ 1'b0 ;
  assign n9325 = ( x88 & ~n3351 ) | ( x88 & n9324 ) | ( ~n3351 & n9324 ) ;
  assign n9326 = n8599 | n9325 ;
  assign n9329 = n9328 ^ n9326 ^ 1'b0 ;
  assign n9331 = n1449 & ~n1957 ;
  assign n9330 = ~n1336 & n6760 ;
  assign n9332 = n9331 ^ n9330 ^ 1'b0 ;
  assign n9333 = n2108 & n9332 ;
  assign n9334 = ( n2666 & n5592 ) | ( n2666 & n9333 ) | ( n5592 & n9333 ) ;
  assign n9335 = n4483 & ~n9334 ;
  assign n9336 = n9335 ^ n6577 ^ 1'b0 ;
  assign n9337 = n9336 ^ n5142 ^ n2755 ;
  assign n9344 = ( n1616 & ~n3049 ) | ( n1616 & n6102 ) | ( ~n3049 & n6102 ) ;
  assign n9345 = n2764 | n9344 ;
  assign n9346 = n3259 | n9345 ;
  assign n9338 = n1676 | n5392 ;
  assign n9339 = ~n325 & n9338 ;
  assign n9340 = n9339 ^ n3776 ^ 1'b0 ;
  assign n9341 = n729 ^ n565 ^ n560 ;
  assign n9342 = n9341 ^ n2171 ^ 1'b0 ;
  assign n9343 = n9340 & ~n9342 ;
  assign n9347 = n9346 ^ n9343 ^ 1'b0 ;
  assign n9351 = n6058 ^ n5821 ^ 1'b0 ;
  assign n9352 = n7042 & n9351 ;
  assign n9353 = n9352 ^ n2280 ^ 1'b0 ;
  assign n9348 = n1457 ^ n555 ^ 1'b0 ;
  assign n9349 = n362 & n9348 ;
  assign n9350 = n9349 ^ n8309 ^ 1'b0 ;
  assign n9354 = n9353 ^ n9350 ^ 1'b0 ;
  assign n9355 = x191 & n3955 ;
  assign n9356 = n685 & n9355 ;
  assign n9357 = n9356 ^ n4686 ^ n1271 ;
  assign n9358 = x176 | n9357 ;
  assign n9359 = n2669 & n4859 ;
  assign n9360 = n1184 & n9359 ;
  assign n9361 = n9360 ^ n8288 ^ n7710 ;
  assign n9362 = ( n613 & n3994 ) | ( n613 & ~n9361 ) | ( n3994 & ~n9361 ) ;
  assign n9364 = n4351 ^ n3246 ^ 1'b0 ;
  assign n9365 = n2780 & n9364 ;
  assign n9366 = ( n1635 & n8693 ) | ( n1635 & ~n9365 ) | ( n8693 & ~n9365 ) ;
  assign n9367 = n1255 & ~n9366 ;
  assign n9368 = n9367 ^ n4478 ^ 1'b0 ;
  assign n9369 = n9368 ^ n1854 ^ 1'b0 ;
  assign n9363 = ~n1289 & n2448 ;
  assign n9370 = n9369 ^ n9363 ^ 1'b0 ;
  assign n9371 = n9185 ^ n572 ^ 1'b0 ;
  assign n9372 = n4783 ^ n1346 ^ 1'b0 ;
  assign n9373 = n4586 & n9372 ;
  assign n9374 = n9373 ^ n3813 ^ 1'b0 ;
  assign n9375 = n8686 ^ n1457 ^ n1347 ;
  assign n9376 = n9375 ^ n7880 ^ n6791 ;
  assign n9377 = n7098 & n9376 ;
  assign n9378 = n7277 & n9377 ;
  assign n9380 = n2020 ^ n339 ^ 1'b0 ;
  assign n9379 = ~n2999 & n3471 ;
  assign n9381 = n9380 ^ n9379 ^ 1'b0 ;
  assign n9382 = n9381 ^ n2889 ^ 1'b0 ;
  assign n9383 = ~n8515 & n9382 ;
  assign n9384 = ~n4814 & n6291 ;
  assign n9385 = n9384 ^ n1609 ^ 1'b0 ;
  assign n9386 = ( n5056 & ~n5633 ) | ( n5056 & n6159 ) | ( ~n5633 & n6159 ) ;
  assign n9387 = x58 & ~n2400 ;
  assign n9388 = n9386 & ~n9387 ;
  assign n9389 = ~n5208 & n9388 ;
  assign n9390 = ( ~n5494 & n9385 ) | ( ~n5494 & n9389 ) | ( n9385 & n9389 ) ;
  assign n9391 = ( ~n2967 & n4878 ) | ( ~n2967 & n9390 ) | ( n4878 & n9390 ) ;
  assign n9392 = n761 & n7494 ;
  assign n9393 = n366 | n422 ;
  assign n9394 = n9393 ^ x39 ^ 1'b0 ;
  assign n9395 = n9394 ^ n2797 ^ 1'b0 ;
  assign n9396 = ~n4265 & n9395 ;
  assign n9397 = n594 | n9396 ;
  assign n9398 = n5495 ^ n5214 ^ 1'b0 ;
  assign n9399 = n830 & ~n9398 ;
  assign n9400 = n9399 ^ n8418 ^ 1'b0 ;
  assign n9401 = n9072 & ~n9400 ;
  assign n9402 = n1322 & ~n5017 ;
  assign n9412 = n8777 ^ n7990 ^ n7262 ;
  assign n9403 = ( n4055 & n5424 ) | ( n4055 & ~n8750 ) | ( n5424 & ~n8750 ) ;
  assign n9404 = ( n1007 & n7289 ) | ( n1007 & n9403 ) | ( n7289 & n9403 ) ;
  assign n9408 = x154 & n4428 ;
  assign n9409 = n3870 & n9408 ;
  assign n9405 = n7899 ^ n5532 ^ n3156 ;
  assign n9406 = n7779 & n9405 ;
  assign n9407 = ~n4846 & n9406 ;
  assign n9410 = n9409 ^ n9407 ^ 1'b0 ;
  assign n9411 = ~n9404 & n9410 ;
  assign n9413 = n9412 ^ n9411 ^ 1'b0 ;
  assign n9414 = n4842 ^ n2863 ^ n1084 ;
  assign n9415 = ( n840 & n2490 ) | ( n840 & n6404 ) | ( n2490 & n6404 ) ;
  assign n9416 = ~n2728 & n5955 ;
  assign n9417 = n9416 ^ n5419 ^ n2735 ;
  assign n9418 = n9415 & n9417 ;
  assign n9419 = n744 | n8757 ;
  assign n9420 = n1235 & ~n9419 ;
  assign n9421 = n7254 & ~n8663 ;
  assign n9422 = n9421 ^ n4814 ^ 1'b0 ;
  assign n9423 = ~n609 & n9422 ;
  assign n9424 = n2558 & n9423 ;
  assign n9425 = n1400 & n5683 ;
  assign n9426 = n5050 | n9344 ;
  assign n9427 = n8174 ^ n6411 ^ 1'b0 ;
  assign n9428 = n2609 | n4546 ;
  assign n9429 = n9428 ^ n2829 ^ n2497 ;
  assign n9431 = n6246 ^ n1563 ^ n1213 ;
  assign n9430 = n1572 & ~n4571 ;
  assign n9432 = n9431 ^ n9430 ^ 1'b0 ;
  assign n9446 = n879 & n4672 ;
  assign n9447 = n9446 ^ n1164 ^ 1'b0 ;
  assign n9448 = ( n576 & ~n2370 ) | ( n576 & n9447 ) | ( ~n2370 & n9447 ) ;
  assign n9433 = n3982 ^ n3806 ^ x74 ;
  assign n9434 = n9433 ^ n5378 ^ 1'b0 ;
  assign n9435 = n9434 ^ n7961 ^ n5946 ;
  assign n9438 = n4791 ^ n2128 ^ 1'b0 ;
  assign n9439 = n8447 ^ n4285 ^ n2127 ;
  assign n9440 = n9439 ^ n4812 ^ 1'b0 ;
  assign n9441 = n9438 & ~n9440 ;
  assign n9436 = n4467 & n6542 ;
  assign n9437 = ( n824 & n3269 ) | ( n824 & ~n9436 ) | ( n3269 & ~n9436 ) ;
  assign n9442 = n9441 ^ n9437 ^ 1'b0 ;
  assign n9443 = n1440 & n9442 ;
  assign n9444 = ~n9435 & n9443 ;
  assign n9445 = n8215 | n9444 ;
  assign n9449 = n9448 ^ n9445 ^ 1'b0 ;
  assign n9450 = n4080 & ~n6615 ;
  assign n9453 = n2214 ^ n2050 ^ 1'b0 ;
  assign n9454 = ~n1000 & n9453 ;
  assign n9451 = ( n640 & n5564 ) | ( n640 & n5613 ) | ( n5564 & n5613 ) ;
  assign n9452 = n6379 & ~n9451 ;
  assign n9455 = n9454 ^ n9452 ^ 1'b0 ;
  assign n9456 = n9455 ^ n2112 ^ 1'b0 ;
  assign n9457 = n5354 ^ n3523 ^ n1293 ;
  assign n9458 = n1916 | n9457 ;
  assign n9459 = n6065 | n9458 ;
  assign n9460 = x231 & n2625 ;
  assign n9461 = ( n1226 & n5772 ) | ( n1226 & n9460 ) | ( n5772 & n9460 ) ;
  assign n9462 = ~n4281 & n6153 ;
  assign n9463 = ( n2843 & n9461 ) | ( n2843 & n9462 ) | ( n9461 & n9462 ) ;
  assign n9464 = n7087 ^ n6294 ^ n2707 ;
  assign n9465 = n8858 & ~n8894 ;
  assign n9466 = n9465 ^ n5567 ^ 1'b0 ;
  assign n9472 = n3005 & n3573 ;
  assign n9473 = ~n6993 & n9472 ;
  assign n9467 = n2643 ^ n2160 ^ 1'b0 ;
  assign n9468 = ( n4106 & ~n4866 ) | ( n4106 & n8985 ) | ( ~n4866 & n8985 ) ;
  assign n9469 = ( ~n3420 & n6033 ) | ( ~n3420 & n7318 ) | ( n6033 & n7318 ) ;
  assign n9470 = n9468 & ~n9469 ;
  assign n9471 = ~n9467 & n9470 ;
  assign n9474 = n9473 ^ n9471 ^ n5085 ;
  assign n9475 = n8444 ^ n1691 ^ 1'b0 ;
  assign n9476 = n3010 ^ n1143 ^ 1'b0 ;
  assign n9477 = ( n2648 & n8015 ) | ( n2648 & ~n9476 ) | ( n8015 & ~n9476 ) ;
  assign n9478 = n9477 ^ n6328 ^ 1'b0 ;
  assign n9479 = x89 & ~n683 ;
  assign n9480 = n9479 ^ n6526 ^ 1'b0 ;
  assign n9481 = n9478 | n9480 ;
  assign n9495 = n8526 ^ n2562 ^ 1'b0 ;
  assign n9496 = n3608 | n9495 ;
  assign n9497 = n9496 ^ n8836 ^ 1'b0 ;
  assign n9482 = n4211 ^ n2150 ^ n1626 ;
  assign n9483 = n345 | n9482 ;
  assign n9484 = ( n1649 & n3627 ) | ( n1649 & ~n5277 ) | ( n3627 & ~n5277 ) ;
  assign n9490 = ( ~x30 & n2611 ) | ( ~x30 & n3103 ) | ( n2611 & n3103 ) ;
  assign n9487 = n2278 & ~n4435 ;
  assign n9488 = n2301 & ~n9487 ;
  assign n9489 = n9488 ^ n1982 ^ 1'b0 ;
  assign n9491 = n9490 ^ n9489 ^ n2987 ;
  assign n9485 = n3965 ^ n3369 ^ x227 ;
  assign n9486 = ( n1133 & n4390 ) | ( n1133 & ~n9485 ) | ( n4390 & ~n9485 ) ;
  assign n9492 = n9491 ^ n9486 ^ 1'b0 ;
  assign n9493 = ( n1401 & n9484 ) | ( n1401 & ~n9492 ) | ( n9484 & ~n9492 ) ;
  assign n9494 = n9483 & ~n9493 ;
  assign n9498 = n9497 ^ n9494 ^ 1'b0 ;
  assign n9499 = ( ~n1625 & n2918 ) | ( ~n1625 & n5034 ) | ( n2918 & n5034 ) ;
  assign n9500 = n5745 ^ n1394 ^ 1'b0 ;
  assign n9501 = n603 | n2196 ;
  assign n9502 = n9501 ^ n5629 ^ 1'b0 ;
  assign n9503 = n9222 ^ n4120 ^ n3905 ;
  assign n9504 = n9502 & n9503 ;
  assign n9505 = n9504 ^ n450 ^ 1'b0 ;
  assign n9506 = n598 | n1081 ;
  assign n9507 = n9506 ^ n2466 ^ n2114 ;
  assign n9508 = n9507 ^ n7899 ^ 1'b0 ;
  assign n9509 = n6534 ^ n4199 ^ n2715 ;
  assign n9510 = n7563 ^ n5179 ^ 1'b0 ;
  assign n9511 = n2095 & n9510 ;
  assign n9512 = ( n1093 & ~n9509 ) | ( n1093 & n9511 ) | ( ~n9509 & n9511 ) ;
  assign n9513 = n4672 ^ n1139 ^ n851 ;
  assign n9514 = ~n3459 & n8415 ;
  assign n9515 = n9513 & n9514 ;
  assign n9516 = n3348 & n3522 ;
  assign n9517 = n2105 & n3996 ;
  assign n9518 = ( n435 & n9516 ) | ( n435 & ~n9517 ) | ( n9516 & ~n9517 ) ;
  assign n9519 = ( ~n688 & n2072 ) | ( ~n688 & n4085 ) | ( n2072 & n4085 ) ;
  assign n9520 = ( ~n2917 & n3651 ) | ( ~n2917 & n9519 ) | ( n3651 & n9519 ) ;
  assign n9521 = n5180 & ~n9520 ;
  assign n9522 = n8466 & n9521 ;
  assign n9523 = n882 | n8527 ;
  assign n9524 = n285 & n9523 ;
  assign n9525 = n2834 & n9085 ;
  assign n9526 = ~n4486 & n6075 ;
  assign n9527 = ( n2892 & ~n7521 ) | ( n2892 & n9526 ) | ( ~n7521 & n9526 ) ;
  assign n9528 = n9527 ^ n6797 ^ 1'b0 ;
  assign n9529 = n2283 & ~n5275 ;
  assign n9530 = ~n1637 & n9529 ;
  assign n9531 = ( n7376 & ~n8040 ) | ( n7376 & n8051 ) | ( ~n8040 & n8051 ) ;
  assign n9532 = n9413 & n9531 ;
  assign n9533 = n9532 ^ n1632 ^ 1'b0 ;
  assign n9534 = ( ~n3401 & n4286 ) | ( ~n3401 & n8102 ) | ( n4286 & n8102 ) ;
  assign n9535 = n435 | n1874 ;
  assign n9536 = n1864 & n9535 ;
  assign n9537 = ~n9534 & n9536 ;
  assign n9538 = n9537 ^ n8565 ^ n4208 ;
  assign n9539 = n7096 ^ n4727 ^ n1837 ;
  assign n9548 = n4422 ^ n4409 ^ n4398 ;
  assign n9543 = n8444 ^ n7679 ^ n7636 ;
  assign n9540 = n2386 & ~n3810 ;
  assign n9541 = n4974 & n9540 ;
  assign n9542 = n9541 ^ n7490 ^ n3787 ;
  assign n9544 = n9543 ^ n9542 ^ n936 ;
  assign n9545 = n2528 & n9544 ;
  assign n9546 = n6244 & n9545 ;
  assign n9547 = n9546 ^ n6102 ^ n4826 ;
  assign n9549 = n9548 ^ n9547 ^ n4851 ;
  assign n9550 = n3561 ^ n432 ^ 1'b0 ;
  assign n9551 = n6190 & n9550 ;
  assign n9553 = n2829 ^ n967 ^ 1'b0 ;
  assign n9554 = n2670 & n9553 ;
  assign n9552 = ~n4490 & n6362 ;
  assign n9555 = n9554 ^ n9552 ^ n1246 ;
  assign n9556 = ( n2671 & ~n9266 ) | ( n2671 & n9555 ) | ( ~n9266 & n9555 ) ;
  assign n9557 = ( x32 & n291 ) | ( x32 & ~n489 ) | ( n291 & ~n489 ) ;
  assign n9558 = ( ~n550 & n6937 ) | ( ~n550 & n9557 ) | ( n6937 & n9557 ) ;
  assign n9559 = n2388 & n9558 ;
  assign n9560 = ~n9556 & n9559 ;
  assign n9561 = n9551 & ~n9560 ;
  assign n9562 = n7737 & n9561 ;
  assign n9563 = n8294 & ~n9562 ;
  assign n9564 = ( n3046 & ~n5043 ) | ( n3046 & n6171 ) | ( ~n5043 & n6171 ) ;
  assign n9565 = n5549 ^ n4393 ^ 1'b0 ;
  assign n9566 = n4551 ^ n3271 ^ n2450 ;
  assign n9567 = n3828 & n9566 ;
  assign n9568 = ( n1951 & ~n9565 ) | ( n1951 & n9567 ) | ( ~n9565 & n9567 ) ;
  assign n9569 = n7928 ^ n4492 ^ n727 ;
  assign n9570 = n546 & ~n559 ;
  assign n9571 = ~x244 & n9570 ;
  assign n9572 = n9569 & ~n9571 ;
  assign n9573 = n9572 ^ n4827 ^ n2905 ;
  assign n9574 = n9573 ^ n3803 ^ n453 ;
  assign n9575 = x252 & n1129 ;
  assign n9576 = n9575 ^ n4878 ^ n3485 ;
  assign n9577 = n6744 ^ n3430 ^ n2978 ;
  assign n9578 = n8903 ^ n5618 ^ 1'b0 ;
  assign n9579 = n9577 | n9578 ;
  assign n9580 = ( n3090 & ~n4158 ) | ( n3090 & n5608 ) | ( ~n4158 & n5608 ) ;
  assign n9581 = n9580 ^ n9247 ^ n6761 ;
  assign n9584 = n1505 | n2731 ;
  assign n9582 = n3629 ^ n688 ^ 1'b0 ;
  assign n9583 = n9582 ^ n7391 ^ n1889 ;
  assign n9585 = n9584 ^ n9583 ^ 1'b0 ;
  assign n9586 = n9581 & n9585 ;
  assign n9587 = ( n3187 & ~n7960 ) | ( n3187 & n9586 ) | ( ~n7960 & n9586 ) ;
  assign n9588 = n3112 & ~n4475 ;
  assign n9589 = n9588 ^ n3651 ^ 1'b0 ;
  assign n9590 = n9589 ^ n8742 ^ 1'b0 ;
  assign n9591 = ~n4324 & n9590 ;
  assign n9592 = n4365 ^ n3315 ^ 1'b0 ;
  assign n9593 = ~n7493 & n9592 ;
  assign n9594 = n9591 & n9593 ;
  assign n9595 = n9594 ^ n1920 ^ 1'b0 ;
  assign n9596 = n9595 ^ n1830 ^ 1'b0 ;
  assign n9597 = ( n707 & n3196 ) | ( n707 & ~n3906 ) | ( n3196 & ~n3906 ) ;
  assign n9598 = n2583 | n9597 ;
  assign n9599 = n8796 & ~n9598 ;
  assign n9600 = n9599 ^ n6544 ^ 1'b0 ;
  assign n9601 = n2103 & ~n9600 ;
  assign n9602 = n9601 ^ n8607 ^ n8171 ;
  assign n9606 = ( ~n1780 & n2338 ) | ( ~n1780 & n7203 ) | ( n2338 & n7203 ) ;
  assign n9603 = n1211 ^ n745 ^ 1'b0 ;
  assign n9604 = n5616 & n9603 ;
  assign n9605 = ( n3441 & n4497 ) | ( n3441 & ~n9604 ) | ( n4497 & ~n9604 ) ;
  assign n9607 = n9606 ^ n9605 ^ 1'b0 ;
  assign n9608 = n4892 & ~n8333 ;
  assign n9609 = ~n8356 & n9261 ;
  assign n9610 = ( n3269 & n4245 ) | ( n3269 & ~n4569 ) | ( n4245 & ~n4569 ) ;
  assign n9611 = n8686 & n9610 ;
  assign n9612 = n1758 & n3672 ;
  assign n9613 = n9612 ^ n7658 ^ 1'b0 ;
  assign n9614 = n1427 & n7506 ;
  assign n9615 = n6042 ^ n1524 ^ 1'b0 ;
  assign n9616 = n8799 & ~n9615 ;
  assign n9617 = n9614 | n9616 ;
  assign n9618 = n3831 ^ n1700 ^ x189 ;
  assign n9619 = ~n2418 & n4365 ;
  assign n9620 = ~n9618 & n9619 ;
  assign n9621 = n9620 ^ n2187 ^ 1'b0 ;
  assign n9622 = ( x64 & n3049 ) | ( x64 & ~n4630 ) | ( n3049 & ~n4630 ) ;
  assign n9623 = n9622 ^ n8213 ^ n6114 ;
  assign n9624 = ~n7018 & n9623 ;
  assign n9625 = n9175 ^ n4178 ^ n3681 ;
  assign n9626 = n9625 ^ n8107 ^ 1'b0 ;
  assign n9627 = ( ~x95 & n565 ) | ( ~x95 & n6268 ) | ( n565 & n6268 ) ;
  assign n9628 = ( x138 & n5263 ) | ( x138 & ~n9627 ) | ( n5263 & ~n9627 ) ;
  assign n9629 = n9259 ^ n5926 ^ n3703 ;
  assign n9630 = n7248 ^ n3162 ^ n1282 ;
  assign n9631 = x10 & n9630 ;
  assign n9632 = n9631 ^ n3961 ^ 1'b0 ;
  assign n9633 = n6474 ^ n1696 ^ 1'b0 ;
  assign n9634 = n9633 ^ n8294 ^ 1'b0 ;
  assign n9635 = n4555 & n9634 ;
  assign n9636 = n9635 ^ n2271 ^ 1'b0 ;
  assign n9637 = ( ~n2207 & n4277 ) | ( ~n2207 & n6581 ) | ( n4277 & n6581 ) ;
  assign n9638 = n7735 & ~n9637 ;
  assign n9639 = n9638 ^ n7260 ^ 1'b0 ;
  assign n9640 = n4950 ^ n2331 ^ 1'b0 ;
  assign n9641 = ~n1143 & n9640 ;
  assign n9642 = n9641 ^ n394 ^ 1'b0 ;
  assign n9643 = n8978 ^ n2158 ^ n1665 ;
  assign n9644 = n9643 ^ n933 ^ 1'b0 ;
  assign n9645 = n9644 ^ n3214 ^ n834 ;
  assign n9646 = n3016 ^ x97 ^ 1'b0 ;
  assign n9647 = n9645 & ~n9646 ;
  assign n9648 = ( n469 & n2139 ) | ( n469 & n2914 ) | ( n2139 & n2914 ) ;
  assign n9649 = n9648 ^ n2350 ^ 1'b0 ;
  assign n9650 = n2627 & n9649 ;
  assign n9651 = n6145 ^ n3624 ^ n567 ;
  assign n9652 = ( n9647 & ~n9650 ) | ( n9647 & n9651 ) | ( ~n9650 & n9651 ) ;
  assign n9653 = n5299 ^ n2148 ^ 1'b0 ;
  assign n9654 = n277 | n9653 ;
  assign n9655 = n6147 | n8309 ;
  assign n9656 = n9654 | n9655 ;
  assign n9657 = x7 & n5094 ;
  assign n9658 = n9657 ^ n9036 ^ 1'b0 ;
  assign n9659 = n7139 ^ n5212 ^ 1'b0 ;
  assign n9660 = ~n401 & n819 ;
  assign n9661 = n2346 & n9660 ;
  assign n9662 = n9661 ^ n652 ^ 1'b0 ;
  assign n9665 = n608 | n5535 ;
  assign n9663 = n8851 ^ n3140 ^ 1'b0 ;
  assign n9664 = ~n8507 & n9663 ;
  assign n9666 = n9665 ^ n9664 ^ 1'b0 ;
  assign n9667 = n9662 & n9666 ;
  assign n9668 = x56 & n2409 ;
  assign n9669 = n9668 ^ n4764 ^ 1'b0 ;
  assign n9672 = ( n483 & ~n2392 ) | ( n483 & n3921 ) | ( ~n2392 & n3921 ) ;
  assign n9671 = n6772 ^ n6649 ^ n647 ;
  assign n9673 = n9672 ^ n9671 ^ n2804 ;
  assign n9670 = n4596 ^ n2310 ^ n2085 ;
  assign n9674 = n9673 ^ n9670 ^ n7602 ;
  assign n9675 = n2020 ^ n1016 ^ 1'b0 ;
  assign n9676 = ~n642 & n1975 ;
  assign n9677 = n9676 ^ n5886 ^ 1'b0 ;
  assign n9678 = n1104 & ~n9677 ;
  assign n9679 = n9678 ^ n6104 ^ 1'b0 ;
  assign n9680 = n9675 | n9679 ;
  assign n9681 = n9680 ^ n1745 ^ 1'b0 ;
  assign n9682 = n8384 ^ n1676 ^ 1'b0 ;
  assign n9683 = n3412 ^ n1920 ^ 1'b0 ;
  assign n9684 = ~n4475 & n9683 ;
  assign n9685 = ~n2163 & n9684 ;
  assign n9686 = n2793 ^ x16 ^ 1'b0 ;
  assign n9687 = n3233 & ~n9686 ;
  assign n9688 = ~n9685 & n9687 ;
  assign n9689 = n9688 ^ n3567 ^ 1'b0 ;
  assign n9690 = n4633 & n6046 ;
  assign n9691 = n9690 ^ n7297 ^ 1'b0 ;
  assign n9692 = n9691 ^ n2999 ^ 1'b0 ;
  assign n9693 = n9692 ^ n7491 ^ 1'b0 ;
  assign n9694 = ~n1010 & n5815 ;
  assign n9695 = n1903 ^ n1624 ^ 1'b0 ;
  assign n9696 = n902 & ~n9695 ;
  assign n9697 = ( n2371 & ~n9694 ) | ( n2371 & n9696 ) | ( ~n9694 & n9696 ) ;
  assign n9698 = n2638 & ~n7178 ;
  assign n9699 = n1007 | n4776 ;
  assign n9700 = n9699 ^ n858 ^ 1'b0 ;
  assign n9701 = ~n2527 & n9700 ;
  assign n9702 = ~n3130 & n9701 ;
  assign n9703 = n9702 ^ n3743 ^ 1'b0 ;
  assign n9704 = n9698 | n9703 ;
  assign n9705 = n9697 | n9704 ;
  assign n9706 = n9705 ^ n5568 ^ 1'b0 ;
  assign n9707 = n9651 ^ n3076 ^ 1'b0 ;
  assign n9708 = n4596 & ~n9707 ;
  assign n9720 = n2950 ^ n1854 ^ n1162 ;
  assign n9721 = ~n2008 & n9720 ;
  assign n9722 = ~n7108 & n9721 ;
  assign n9723 = ~n2537 & n9722 ;
  assign n9717 = ( ~n647 & n1078 ) | ( ~n647 & n1863 ) | ( n1078 & n1863 ) ;
  assign n9718 = n9717 ^ n2532 ^ 1'b0 ;
  assign n9719 = n5419 & n9718 ;
  assign n9724 = n9723 ^ n9719 ^ 1'b0 ;
  assign n9714 = n5513 ^ n5505 ^ 1'b0 ;
  assign n9715 = n7958 & n9714 ;
  assign n9709 = n4305 ^ n1499 ^ 1'b0 ;
  assign n9710 = n1688 ^ n838 ^ 1'b0 ;
  assign n9711 = n6304 & ~n9710 ;
  assign n9712 = n9711 ^ n1893 ^ 1'b0 ;
  assign n9713 = n9709 & ~n9712 ;
  assign n9716 = n9715 ^ n9713 ^ n8164 ;
  assign n9725 = n9724 ^ n9716 ^ 1'b0 ;
  assign n9727 = n3271 ^ n2537 ^ n1748 ;
  assign n9726 = n868 & n5486 ;
  assign n9728 = n9727 ^ n9726 ^ 1'b0 ;
  assign n9729 = n7155 ^ n1375 ^ 1'b0 ;
  assign n9730 = n2878 | n9729 ;
  assign n9731 = ( n2513 & ~n4313 ) | ( n2513 & n9730 ) | ( ~n4313 & n9730 ) ;
  assign n9732 = ( x108 & n3919 ) | ( x108 & ~n9731 ) | ( n3919 & ~n9731 ) ;
  assign n9733 = n9732 ^ n2229 ^ 1'b0 ;
  assign n9734 = n9728 & ~n9733 ;
  assign n9735 = ~n2561 & n2668 ;
  assign n9736 = n9735 ^ n2329 ^ 1'b0 ;
  assign n9737 = n1989 | n6541 ;
  assign n9738 = n9737 ^ n7155 ^ 1'b0 ;
  assign n9739 = n9738 ^ n2657 ^ 1'b0 ;
  assign n9740 = ( n1331 & n1937 ) | ( n1331 & n3696 ) | ( n1937 & n3696 ) ;
  assign n9741 = ( ~n5720 & n6667 ) | ( ~n5720 & n9740 ) | ( n6667 & n9740 ) ;
  assign n9742 = ( ~n9736 & n9739 ) | ( ~n9736 & n9741 ) | ( n9739 & n9741 ) ;
  assign n9743 = n3917 & ~n3943 ;
  assign n9744 = ~n9742 & n9743 ;
  assign n9745 = n8904 ^ n3426 ^ 1'b0 ;
  assign n9746 = ~n1361 & n9745 ;
  assign n9747 = ( ~n1304 & n4358 ) | ( ~n1304 & n9746 ) | ( n4358 & n9746 ) ;
  assign n9748 = n9747 ^ n4187 ^ 1'b0 ;
  assign n9749 = ~n8657 & n9748 ;
  assign n9750 = n2859 ^ n2543 ^ n2009 ;
  assign n9751 = ( ~n630 & n1011 ) | ( ~n630 & n3705 ) | ( n1011 & n3705 ) ;
  assign n9752 = ( n8644 & n9750 ) | ( n8644 & ~n9751 ) | ( n9750 & ~n9751 ) ;
  assign n9753 = n9752 ^ n1299 ^ 1'b0 ;
  assign n9754 = n2444 & n9753 ;
  assign n9755 = ( x131 & n1626 ) | ( x131 & ~n3274 ) | ( n1626 & ~n3274 ) ;
  assign n9756 = n6423 | n9755 ;
  assign n9757 = n9756 ^ n9378 ^ n1610 ;
  assign n9761 = n6724 ^ n1616 ^ n1473 ;
  assign n9758 = n7595 ^ n6180 ^ n2428 ;
  assign n9759 = n4601 & ~n9758 ;
  assign n9760 = n9759 ^ n4022 ^ 1'b0 ;
  assign n9762 = n9761 ^ n9760 ^ n4220 ;
  assign n9763 = n628 & ~n5516 ;
  assign n9764 = x106 & ~n9763 ;
  assign n9765 = n9577 & n9764 ;
  assign n9766 = n9765 ^ n3432 ^ 1'b0 ;
  assign n9768 = n546 | n789 ;
  assign n9769 = n9768 ^ x159 ^ 1'b0 ;
  assign n9767 = n1150 | n1423 ;
  assign n9770 = n9769 ^ n9767 ^ n2828 ;
  assign n9771 = n4307 & n9770 ;
  assign n9772 = ~x79 & n9771 ;
  assign n9773 = n7091 | n9772 ;
  assign n9774 = n4428 & ~n7506 ;
  assign n9775 = n8601 & n9774 ;
  assign n9776 = ( x35 & n6498 ) | ( x35 & n9775 ) | ( n6498 & n9775 ) ;
  assign n9777 = ( n9766 & n9773 ) | ( n9766 & ~n9776 ) | ( n9773 & ~n9776 ) ;
  assign n9783 = n9717 ^ n1743 ^ 1'b0 ;
  assign n9784 = ~n9672 & n9783 ;
  assign n9780 = n6714 ^ n4542 ^ 1'b0 ;
  assign n9778 = n6092 ^ n2135 ^ n866 ;
  assign n9779 = n9778 ^ n1562 ^ 1'b0 ;
  assign n9781 = n9780 ^ n9779 ^ 1'b0 ;
  assign n9782 = ~n685 & n9781 ;
  assign n9785 = n9784 ^ n9782 ^ 1'b0 ;
  assign n9786 = n8935 | n9785 ;
  assign n9787 = n8937 ^ n1820 ^ x8 ;
  assign n9788 = n963 | n9787 ;
  assign n9789 = n5935 ^ n2835 ^ 1'b0 ;
  assign n9790 = n5918 | n9789 ;
  assign n9791 = ( ~n3375 & n6989 ) | ( ~n3375 & n9790 ) | ( n6989 & n9790 ) ;
  assign n9792 = ~n3322 & n3919 ;
  assign n9793 = ~x32 & n9792 ;
  assign n9794 = n885 & ~n9793 ;
  assign n9795 = ( n2453 & n5601 ) | ( n2453 & n5834 ) | ( n5601 & n5834 ) ;
  assign n9796 = n4317 ^ n1370 ^ n807 ;
  assign n9797 = n3037 | n9796 ;
  assign n9798 = n9797 ^ n5025 ^ 1'b0 ;
  assign n9799 = ( n2103 & n2400 ) | ( n2103 & ~n9798 ) | ( n2400 & ~n9798 ) ;
  assign n9800 = n8995 ^ n8342 ^ 1'b0 ;
  assign n9801 = n8587 & ~n9800 ;
  assign n9802 = n530 & n2611 ;
  assign n9803 = n9802 ^ n7595 ^ 1'b0 ;
  assign n9804 = ~n4410 & n9803 ;
  assign n9805 = ~n6075 & n9804 ;
  assign n9806 = n8567 ^ n7436 ^ 1'b0 ;
  assign n9807 = x64 & ~n9806 ;
  assign n9808 = n7977 ^ n3491 ^ 1'b0 ;
  assign n9809 = ~n9761 & n9808 ;
  assign n9810 = n7709 ^ n1069 ^ 1'b0 ;
  assign n9811 = n6348 & ~n9810 ;
  assign n9812 = n5059 & n9811 ;
  assign n9813 = n4280 | n5903 ;
  assign n9814 = n3554 & ~n9813 ;
  assign n9815 = ( ~n7557 & n9076 ) | ( ~n7557 & n9363 ) | ( n9076 & n9363 ) ;
  assign n9816 = n5477 ^ n5076 ^ n3353 ;
  assign n9817 = ( n2335 & n3255 ) | ( n2335 & n9816 ) | ( n3255 & n9816 ) ;
  assign n9818 = n9461 ^ n3858 ^ 1'b0 ;
  assign n9819 = n1600 & ~n9818 ;
  assign n9820 = n9819 ^ n3870 ^ 1'b0 ;
  assign n9822 = x158 & n1731 ;
  assign n9823 = ~n2426 & n9822 ;
  assign n9821 = n7732 ^ n585 ^ n372 ;
  assign n9824 = n9823 ^ n9821 ^ n8636 ;
  assign n9825 = n463 & ~n1452 ;
  assign n9826 = n1452 & n9825 ;
  assign n9827 = n1243 & n2097 ;
  assign n9828 = n9826 & n9827 ;
  assign n9829 = n9828 ^ n3255 ^ 1'b0 ;
  assign n9830 = ( n1128 & n4182 ) | ( n1128 & ~n9829 ) | ( n4182 & ~n9829 ) ;
  assign n9831 = n5924 & n9650 ;
  assign n9832 = n9831 ^ n6592 ^ 1'b0 ;
  assign n9833 = n9832 ^ n7904 ^ n3979 ;
  assign n9834 = n267 | n667 ;
  assign n9835 = ( n596 & n2257 ) | ( n596 & n5618 ) | ( n2257 & n5618 ) ;
  assign n9836 = n9835 ^ n3941 ^ n2329 ;
  assign n9837 = ( ~n2107 & n7314 ) | ( ~n2107 & n9836 ) | ( n7314 & n9836 ) ;
  assign n9838 = x30 & n3416 ;
  assign n9839 = ~n9837 & n9838 ;
  assign n9840 = n3069 ^ n2244 ^ n999 ;
  assign n9841 = n5949 | n9840 ;
  assign n9842 = n9841 ^ n5242 ^ 1'b0 ;
  assign n9843 = n9842 ^ n3556 ^ 1'b0 ;
  assign n9844 = n7083 | n9843 ;
  assign n9845 = ( n1684 & n3460 ) | ( n1684 & ~n5640 ) | ( n3460 & ~n5640 ) ;
  assign n9846 = n5377 ^ n1262 ^ n633 ;
  assign n9847 = ~n2563 & n9846 ;
  assign n9848 = ~x105 & n9847 ;
  assign n9849 = n9845 | n9848 ;
  assign n9850 = n9844 & ~n9849 ;
  assign n9851 = n9018 & n9850 ;
  assign n9852 = ( n9834 & n9839 ) | ( n9834 & n9851 ) | ( n9839 & n9851 ) ;
  assign n9853 = n7686 ^ n3527 ^ n2957 ;
  assign n9855 = n3984 ^ n1408 ^ 1'b0 ;
  assign n9856 = n1536 | n9855 ;
  assign n9857 = n9856 ^ n5450 ^ n816 ;
  assign n9854 = ( x79 & n3485 ) | ( x79 & n7195 ) | ( n3485 & n7195 ) ;
  assign n9858 = n9857 ^ n9854 ^ n8957 ;
  assign n9859 = n969 ^ n566 ^ 1'b0 ;
  assign n9860 = n3552 | n9859 ;
  assign n9861 = ( ~n1593 & n2417 ) | ( ~n1593 & n7882 ) | ( n2417 & n7882 ) ;
  assign n9862 = n9861 ^ n3934 ^ 1'b0 ;
  assign n9863 = n9862 ^ n1266 ^ 1'b0 ;
  assign n9864 = ~n9860 & n9863 ;
  assign n9866 = n4888 & ~n7281 ;
  assign n9867 = n9866 ^ n8451 ^ 1'b0 ;
  assign n9865 = n6356 & ~n8155 ;
  assign n9868 = n9867 ^ n9865 ^ n1203 ;
  assign n9869 = ( ~n917 & n1836 ) | ( ~n917 & n7688 ) | ( n1836 & n7688 ) ;
  assign n9870 = n8331 ^ n5784 ^ x151 ;
  assign n9871 = n1627 ^ n1044 ^ x78 ;
  assign n9872 = ( x58 & n1445 ) | ( x58 & n9871 ) | ( n1445 & n9871 ) ;
  assign n9873 = n9872 ^ n2551 ^ x13 ;
  assign n9874 = n6173 ^ n4453 ^ 1'b0 ;
  assign n9875 = ~n9873 & n9874 ;
  assign n9876 = ( ~n9869 & n9870 ) | ( ~n9869 & n9875 ) | ( n9870 & n9875 ) ;
  assign n9877 = n644 | n1294 ;
  assign n9878 = n853 & ~n5502 ;
  assign n9879 = n9878 ^ n9860 ^ 1'b0 ;
  assign n9880 = n511 & ~n4681 ;
  assign n9881 = n2312 & n9880 ;
  assign n9882 = ~n1025 & n1036 ;
  assign n9883 = n9881 & n9882 ;
  assign n9884 = n5880 & ~n9883 ;
  assign n9885 = n518 ^ x147 ^ 1'b0 ;
  assign n9886 = n788 | n8017 ;
  assign n9887 = n9885 & ~n9886 ;
  assign n9888 = n5884 & ~n9887 ;
  assign n9889 = n9888 ^ n2571 ^ 1'b0 ;
  assign n9893 = n8084 ^ n4989 ^ n313 ;
  assign n9894 = ~n5502 & n9893 ;
  assign n9895 = n9894 ^ n5179 ^ 1'b0 ;
  assign n9890 = n4886 ^ n4725 ^ n1928 ;
  assign n9891 = x81 & n9890 ;
  assign n9892 = ~n3707 & n9891 ;
  assign n9896 = n9895 ^ n9892 ^ 1'b0 ;
  assign n9897 = ~n9889 & n9896 ;
  assign n9898 = n8425 & n9897 ;
  assign n9899 = n9884 & ~n9898 ;
  assign n9900 = n9899 ^ n5284 ^ 1'b0 ;
  assign n9901 = n9879 & n9900 ;
  assign n9902 = n9237 ^ n8778 ^ 1'b0 ;
  assign n9903 = n5443 ^ n450 ^ 1'b0 ;
  assign n9904 = ~n6497 & n9903 ;
  assign n9905 = n5549 ^ n711 ^ n459 ;
  assign n9906 = n9185 | n9905 ;
  assign n9907 = ( n5031 & n8867 ) | ( n5031 & n8968 ) | ( n8867 & n8968 ) ;
  assign n9908 = n9907 ^ n467 ^ n301 ;
  assign n9909 = n9569 ^ n2808 ^ 1'b0 ;
  assign n9910 = n9909 ^ n7638 ^ 1'b0 ;
  assign n9911 = x39 & n9910 ;
  assign n9912 = n4635 | n4798 ;
  assign n9913 = x136 & n3806 ;
  assign n9914 = n9912 & n9913 ;
  assign n9915 = n5520 ^ n1281 ^ 1'b0 ;
  assign n9916 = n425 & ~n9915 ;
  assign n9917 = ( n1736 & n9914 ) | ( n1736 & n9916 ) | ( n9914 & n9916 ) ;
  assign n9924 = n322 & ~n3087 ;
  assign n9920 = ~x174 & n838 ;
  assign n9921 = n828 & n9920 ;
  assign n9919 = n3848 ^ x28 ^ 1'b0 ;
  assign n9922 = n9921 ^ n9919 ^ 1'b0 ;
  assign n9918 = ( ~n5104 & n5307 ) | ( ~n5104 & n6659 ) | ( n5307 & n6659 ) ;
  assign n9923 = n9922 ^ n9918 ^ n1434 ;
  assign n9925 = n9924 ^ n9923 ^ n5825 ;
  assign n9926 = n9622 ^ n6053 ^ n2337 ;
  assign n9927 = ( n3540 & n9444 ) | ( n3540 & ~n9926 ) | ( n9444 & ~n9926 ) ;
  assign n9928 = ( x203 & n816 ) | ( x203 & n3163 ) | ( n816 & n3163 ) ;
  assign n9929 = n5313 & ~n9928 ;
  assign n9930 = ~n1922 & n9929 ;
  assign n9931 = n9930 ^ n6410 ^ 1'b0 ;
  assign n9932 = n2110 & ~n6373 ;
  assign n9933 = n1889 ^ n331 ^ 1'b0 ;
  assign n9934 = n9932 & n9933 ;
  assign n9935 = n2409 | n5748 ;
  assign n9936 = n5131 & n5234 ;
  assign n9937 = n1815 | n4021 ;
  assign n9938 = n9937 ^ n7763 ^ 1'b0 ;
  assign n9939 = n9938 ^ n6002 ^ 1'b0 ;
  assign n9940 = n9936 & n9939 ;
  assign n9941 = ( n465 & n6127 ) | ( n465 & ~n9940 ) | ( n6127 & ~n9940 ) ;
  assign n9942 = ( n1953 & ~n3713 ) | ( n1953 & n4802 ) | ( ~n3713 & n4802 ) ;
  assign n9943 = n9942 ^ n9467 ^ n8607 ;
  assign n9944 = n9943 ^ n3543 ^ 1'b0 ;
  assign n9945 = n2880 & ~n5222 ;
  assign n9946 = n9945 ^ n8540 ^ n5050 ;
  assign n9947 = ( n8193 & n9944 ) | ( n8193 & ~n9946 ) | ( n9944 & ~n9946 ) ;
  assign n9948 = n5567 ^ x3 ^ 1'b0 ;
  assign n9949 = n9948 ^ n1903 ^ n1468 ;
  assign n9950 = n6559 ^ n3148 ^ 1'b0 ;
  assign n9951 = ~n4078 & n9950 ;
  assign n9952 = ( n6515 & n9949 ) | ( n6515 & ~n9951 ) | ( n9949 & ~n9951 ) ;
  assign n9953 = ( n526 & n9947 ) | ( n526 & n9952 ) | ( n9947 & n9952 ) ;
  assign n9956 = n7487 ^ n4997 ^ n498 ;
  assign n9954 = x247 & n7598 ;
  assign n9955 = n9954 ^ n6414 ^ 1'b0 ;
  assign n9957 = n9956 ^ n9955 ^ n4298 ;
  assign n9958 = n9957 ^ n2469 ^ 1'b0 ;
  assign n9959 = n5043 & n9810 ;
  assign n9960 = n3939 & ~n9959 ;
  assign n9961 = n9960 ^ n8525 ^ 1'b0 ;
  assign n9962 = n9961 ^ n5365 ^ 1'b0 ;
  assign n9963 = ( ~n426 & n2176 ) | ( ~n426 & n3794 ) | ( n2176 & n3794 ) ;
  assign n9964 = n3037 | n6065 ;
  assign n9965 = n9964 ^ n4442 ^ 1'b0 ;
  assign n9966 = n9965 ^ n1848 ^ 1'b0 ;
  assign n9967 = ~n9963 & n9966 ;
  assign n9968 = ~n3169 & n3609 ;
  assign n9969 = n3346 ^ n1867 ^ n471 ;
  assign n9970 = n2194 & ~n3820 ;
  assign n9971 = n9970 ^ n6466 ^ 1'b0 ;
  assign n9972 = n1967 & ~n9971 ;
  assign n9973 = ( n1590 & n1990 ) | ( n1590 & n2487 ) | ( n1990 & n2487 ) ;
  assign n9974 = ( ~x61 & n9153 ) | ( ~x61 & n9973 ) | ( n9153 & n9973 ) ;
  assign n9975 = n2867 | n9974 ;
  assign n9976 = n9972 | n9975 ;
  assign n9977 = n9969 & ~n9976 ;
  assign n9978 = n9977 ^ n7737 ^ 1'b0 ;
  assign n9979 = n3741 | n9978 ;
  assign n9980 = n9979 ^ n4147 ^ 1'b0 ;
  assign n9981 = n4549 | n8784 ;
  assign n9982 = n9980 & ~n9981 ;
  assign n9983 = n6464 ^ n4068 ^ 1'b0 ;
  assign n9984 = n9983 ^ n5916 ^ 1'b0 ;
  assign n9985 = n9963 ^ n1381 ^ 1'b0 ;
  assign n9986 = ~n9984 & n9985 ;
  assign n9990 = ~x137 & n667 ;
  assign n9991 = n4351 & ~n9990 ;
  assign n9988 = n4956 | n7075 ;
  assign n9989 = n3007 | n9988 ;
  assign n9992 = n9991 ^ n9989 ^ n8431 ;
  assign n9987 = n3751 ^ n2782 ^ 1'b0 ;
  assign n9993 = n9992 ^ n9987 ^ n6887 ;
  assign n9994 = n1219 ^ x210 ^ 1'b0 ;
  assign n9995 = n5587 ^ n1636 ^ 1'b0 ;
  assign n9996 = ~n9994 & n9995 ;
  assign n9997 = ~n4139 & n9996 ;
  assign n9998 = n3406 & n9997 ;
  assign n9999 = ~n4319 & n9349 ;
  assign n10000 = n9614 ^ n7912 ^ n4996 ;
  assign n10001 = n887 | n1609 ;
  assign n10002 = ~n2139 & n10001 ;
  assign n10003 = n10002 ^ n4060 ^ 1'b0 ;
  assign n10004 = ~n6458 & n10003 ;
  assign n10005 = n1834 ^ n1573 ^ 1'b0 ;
  assign n10006 = n10005 ^ n5387 ^ 1'b0 ;
  assign n10007 = n261 & ~n10006 ;
  assign n10008 = n10007 ^ n4053 ^ 1'b0 ;
  assign n10009 = n8644 ^ n7630 ^ n4351 ;
  assign n10010 = ( ~n10004 & n10008 ) | ( ~n10004 & n10009 ) | ( n10008 & n10009 ) ;
  assign n10011 = n3988 | n10010 ;
  assign n10013 = ~n1792 & n7211 ;
  assign n10012 = ( ~n670 & n1731 ) | ( ~n670 & n2984 ) | ( n1731 & n2984 ) ;
  assign n10014 = n10013 ^ n10012 ^ n1375 ;
  assign n10015 = n10014 ^ n7840 ^ 1'b0 ;
  assign n10016 = ( n2244 & n4078 ) | ( n2244 & n5821 ) | ( n4078 & n5821 ) ;
  assign n10017 = n10016 ^ n9126 ^ n7631 ;
  assign n10018 = n1886 & n3117 ;
  assign n10019 = ~n5418 & n10018 ;
  assign n10020 = ( ~n1387 & n2120 ) | ( ~n1387 & n2700 ) | ( n2120 & n2700 ) ;
  assign n10021 = ( n4178 & n10019 ) | ( n4178 & n10020 ) | ( n10019 & n10020 ) ;
  assign n10022 = n6496 & ~n10021 ;
  assign n10023 = n2937 ^ n473 ^ n342 ;
  assign n10024 = n6259 & ~n10023 ;
  assign n10025 = n10024 ^ n7763 ^ 1'b0 ;
  assign n10026 = n4312 & ~n10025 ;
  assign n10027 = n10022 & n10026 ;
  assign n10032 = n1737 ^ n286 ^ x185 ;
  assign n10028 = n1227 | n3465 ;
  assign n10029 = n2587 | n10028 ;
  assign n10030 = n3264 ^ n2187 ^ x156 ;
  assign n10031 = n10029 & n10030 ;
  assign n10033 = n10032 ^ n10031 ^ 1'b0 ;
  assign n10034 = n6423 ^ n1915 ^ 1'b0 ;
  assign n10035 = ~n5140 & n10034 ;
  assign n10036 = n10035 ^ n8237 ^ 1'b0 ;
  assign n10037 = n5430 | n5975 ;
  assign n10038 = n2495 | n10037 ;
  assign n10042 = n4103 & n4151 ;
  assign n10041 = n4145 ^ n2367 ^ 1'b0 ;
  assign n10043 = n10042 ^ n10041 ^ n4407 ;
  assign n10044 = ~n5930 & n10043 ;
  assign n10045 = n10044 ^ n4067 ^ 1'b0 ;
  assign n10039 = n9944 ^ n8423 ^ n798 ;
  assign n10040 = ( n7736 & n9526 ) | ( n7736 & ~n10039 ) | ( n9526 & ~n10039 ) ;
  assign n10046 = n10045 ^ n10040 ^ n7665 ;
  assign n10047 = n10038 | n10046 ;
  assign n10058 = n5556 ^ n4754 ^ n1968 ;
  assign n10054 = n7235 ^ n2061 ^ n997 ;
  assign n10055 = n2333 ^ n1427 ^ n1068 ;
  assign n10056 = ( n7726 & ~n10054 ) | ( n7726 & n10055 ) | ( ~n10054 & n10055 ) ;
  assign n10057 = n10056 ^ n8342 ^ n5631 ;
  assign n10051 = n3658 ^ n1634 ^ 1'b0 ;
  assign n10052 = n2614 & n10051 ;
  assign n10048 = n326 ^ x207 ^ 1'b0 ;
  assign n10049 = n6279 & n10048 ;
  assign n10050 = ~n6472 & n10049 ;
  assign n10053 = n10052 ^ n10050 ^ 1'b0 ;
  assign n10059 = n10058 ^ n10057 ^ n10053 ;
  assign n10060 = n8633 ^ n1129 ^ n337 ;
  assign n10061 = n9340 & ~n9680 ;
  assign n10075 = n4376 ^ n1068 ^ 1'b0 ;
  assign n10062 = n523 & ~n1226 ;
  assign n10063 = n10062 ^ n5256 ^ x235 ;
  assign n10064 = n690 & ~n8703 ;
  assign n10065 = n10064 ^ n5529 ^ 1'b0 ;
  assign n10066 = n9031 ^ n5076 ^ 1'b0 ;
  assign n10067 = x181 & n2099 ;
  assign n10068 = ( n1666 & n2796 ) | ( n1666 & ~n3123 ) | ( n2796 & ~n3123 ) ;
  assign n10069 = n3682 ^ n2735 ^ 1'b0 ;
  assign n10070 = n10069 ^ n6279 ^ n6236 ;
  assign n10071 = n10068 & n10070 ;
  assign n10072 = ( n1154 & n10067 ) | ( n1154 & ~n10071 ) | ( n10067 & ~n10071 ) ;
  assign n10073 = ( n10065 & n10066 ) | ( n10065 & n10072 ) | ( n10066 & n10072 ) ;
  assign n10074 = n10063 & n10073 ;
  assign n10076 = n10075 ^ n10074 ^ 1'b0 ;
  assign n10085 = n774 & ~n5095 ;
  assign n10086 = n5069 & n10085 ;
  assign n10080 = ( n2149 & ~n4274 ) | ( n2149 & n5244 ) | ( ~n4274 & n5244 ) ;
  assign n10077 = ~n4516 & n5036 ;
  assign n10078 = n7698 ^ n5153 ^ 1'b0 ;
  assign n10079 = n10077 & n10078 ;
  assign n10081 = n10080 ^ n10079 ^ 1'b0 ;
  assign n10082 = n786 & ~n4441 ;
  assign n10083 = ~n5421 & n10082 ;
  assign n10084 = n10081 | n10083 ;
  assign n10087 = n10086 ^ n10084 ^ 1'b0 ;
  assign n10088 = n8000 ^ n6855 ^ n1326 ;
  assign n10089 = n9124 ^ n8759 ^ 1'b0 ;
  assign n10090 = n4194 & ~n5628 ;
  assign n10091 = x128 & n10090 ;
  assign n10094 = ( n1229 & n2309 ) | ( n1229 & ~n8718 ) | ( n2309 & ~n8718 ) ;
  assign n10092 = ( n894 & n2359 ) | ( n894 & n6021 ) | ( n2359 & n6021 ) ;
  assign n10093 = ( n683 & n4593 ) | ( n683 & ~n10092 ) | ( n4593 & ~n10092 ) ;
  assign n10095 = n10094 ^ n10093 ^ 1'b0 ;
  assign n10096 = ( n3923 & n5458 ) | ( n3923 & n10095 ) | ( n5458 & n10095 ) ;
  assign n10097 = n355 & n5071 ;
  assign n10098 = n7721 & ~n10097 ;
  assign n10099 = n2574 ^ n1699 ^ 1'b0 ;
  assign n10100 = n10099 ^ x239 ^ 1'b0 ;
  assign n10102 = n3404 & ~n4508 ;
  assign n10103 = n10102 ^ n2029 ^ 1'b0 ;
  assign n10104 = n10103 ^ n4268 ^ n3707 ;
  assign n10101 = n7648 ^ n7478 ^ n3145 ;
  assign n10105 = n10104 ^ n10101 ^ 1'b0 ;
  assign n10106 = n10055 ^ n8260 ^ n854 ;
  assign n10107 = n5921 ^ n3531 ^ n1952 ;
  assign n10108 = n10107 ^ n5337 ^ n3772 ;
  assign n10109 = n10108 ^ n8248 ^ n8076 ;
  assign n10110 = n1968 & ~n2373 ;
  assign n10111 = n10110 ^ n6420 ^ 1'b0 ;
  assign n10112 = n7931 ^ n7901 ^ n7303 ;
  assign n10113 = n6450 ^ n4468 ^ n1101 ;
  assign n10114 = ~n10072 & n10113 ;
  assign n10115 = ( n3278 & n3319 ) | ( n3278 & n3762 ) | ( n3319 & n3762 ) ;
  assign n10116 = n673 & ~n10115 ;
  assign n10117 = x43 & n4781 ;
  assign n10118 = n6800 & n10117 ;
  assign n10119 = n10118 ^ n4113 ^ 1'b0 ;
  assign n10120 = n10116 | n10119 ;
  assign n10121 = n7062 | n7815 ;
  assign n10122 = n2360 & ~n6857 ;
  assign n10123 = n1088 & ~n7224 ;
  assign n10124 = n2844 ^ n1192 ^ 1'b0 ;
  assign n10125 = n10124 ^ n7833 ^ x74 ;
  assign n10126 = n1662 ^ n817 ^ 1'b0 ;
  assign n10127 = n1545 | n10126 ;
  assign n10128 = n10127 ^ n5338 ^ 1'b0 ;
  assign n10130 = n1731 & ~n7053 ;
  assign n10131 = n10130 ^ n3787 ^ 1'b0 ;
  assign n10129 = n1561 ^ n518 ^ 1'b0 ;
  assign n10132 = n10131 ^ n10129 ^ 1'b0 ;
  assign n10133 = n464 & n3672 ;
  assign n10134 = n10133 ^ n2712 ^ 1'b0 ;
  assign n10135 = n10134 ^ n2411 ^ 1'b0 ;
  assign n10136 = n2406 & ~n10135 ;
  assign n10137 = ( n5938 & n10132 ) | ( n5938 & n10136 ) | ( n10132 & n10136 ) ;
  assign n10138 = ( n5983 & n10128 ) | ( n5983 & n10137 ) | ( n10128 & n10137 ) ;
  assign n10139 = n6839 ^ n2316 ^ 1'b0 ;
  assign n10140 = ~n911 & n2751 ;
  assign n10141 = ( n1549 & n2976 ) | ( n1549 & ~n10140 ) | ( n2976 & ~n10140 ) ;
  assign n10142 = ~n4441 & n9479 ;
  assign n10143 = ~n10141 & n10142 ;
  assign n10144 = ( n2121 & n10139 ) | ( n2121 & n10143 ) | ( n10139 & n10143 ) ;
  assign n10145 = n2065 & ~n9125 ;
  assign n10146 = n10145 ^ n4876 ^ 1'b0 ;
  assign n10147 = n1297 | n1433 ;
  assign n10148 = n10146 | n10147 ;
  assign n10149 = ( ~n3187 & n7929 ) | ( ~n3187 & n10148 ) | ( n7929 & n10148 ) ;
  assign n10150 = n10149 ^ n8960 ^ 1'b0 ;
  assign n10151 = n840 & ~n1122 ;
  assign n10152 = n2711 ^ n2002 ^ 1'b0 ;
  assign n10153 = n10152 ^ n8710 ^ 1'b0 ;
  assign n10154 = ( x215 & ~n10151 ) | ( x215 & n10153 ) | ( ~n10151 & n10153 ) ;
  assign n10155 = n9793 ^ n829 ^ n421 ;
  assign n10156 = ( n6667 & ~n9518 ) | ( n6667 & n10155 ) | ( ~n9518 & n10155 ) ;
  assign n10158 = x190 & n4180 ;
  assign n10159 = n539 & n10158 ;
  assign n10157 = n4374 | n8043 ;
  assign n10160 = n10159 ^ n10157 ^ 1'b0 ;
  assign n10161 = ~n3010 & n10160 ;
  assign n10162 = n10161 ^ n3746 ^ n2406 ;
  assign n10163 = n5056 ^ n801 ^ 1'b0 ;
  assign n10164 = n1419 & ~n4126 ;
  assign n10165 = ~n10163 & n10164 ;
  assign n10166 = n10165 ^ n6928 ^ 1'b0 ;
  assign n10167 = n10162 | n10166 ;
  assign n10168 = ~n1697 & n2540 ;
  assign n10169 = n10168 ^ n894 ^ 1'b0 ;
  assign n10170 = n10169 ^ n2828 ^ n1676 ;
  assign n10171 = n5065 ^ n940 ^ 1'b0 ;
  assign n10172 = n10170 & ~n10171 ;
  assign n10173 = n4999 ^ n2226 ^ 1'b0 ;
  assign n10174 = x17 & ~n10173 ;
  assign n10177 = ( ~n307 & n2936 ) | ( ~n307 & n7069 ) | ( n2936 & n7069 ) ;
  assign n10178 = ( n5001 & n10021 ) | ( n5001 & ~n10177 ) | ( n10021 & ~n10177 ) ;
  assign n10175 = n268 & ~n1884 ;
  assign n10176 = n10175 ^ n1217 ^ x208 ;
  assign n10179 = n10178 ^ n10176 ^ 1'b0 ;
  assign n10180 = n5814 ^ n2362 ^ n523 ;
  assign n10181 = n2530 & ~n10180 ;
  assign n10182 = n10163 ^ n4839 ^ n1236 ;
  assign n10184 = n1004 & ~n1901 ;
  assign n10185 = n4197 & n10184 ;
  assign n10183 = n256 & ~n4487 ;
  assign n10186 = n10185 ^ n10183 ^ 1'b0 ;
  assign n10187 = n3744 ^ n2657 ^ 1'b0 ;
  assign n10188 = ( n2905 & ~n7829 ) | ( n2905 & n10187 ) | ( ~n7829 & n10187 ) ;
  assign n10189 = n3906 & ~n10188 ;
  assign n10190 = ~n4949 & n10189 ;
  assign n10191 = ( n647 & n2734 ) | ( n647 & n6744 ) | ( n2734 & n6744 ) ;
  assign n10192 = ~n364 & n10191 ;
  assign n10193 = n10192 ^ n7359 ^ n662 ;
  assign n10194 = n1189 & ~n4153 ;
  assign n10195 = n10194 ^ n5601 ^ 1'b0 ;
  assign n10196 = n10195 ^ n6265 ^ n5764 ;
  assign n10197 = n3377 & n5101 ;
  assign n10198 = n10197 ^ n6577 ^ 1'b0 ;
  assign n10199 = n9522 | n10198 ;
  assign n10200 = n10196 & ~n10199 ;
  assign n10201 = n2388 ^ n1372 ^ 1'b0 ;
  assign n10202 = n9865 | n10201 ;
  assign n10203 = n2459 ^ n648 ^ 1'b0 ;
  assign n10204 = n10203 ^ n6915 ^ 1'b0 ;
  assign n10205 = n7779 & ~n10204 ;
  assign n10206 = ( ~n1676 & n7445 ) | ( ~n1676 & n10205 ) | ( n7445 & n10205 ) ;
  assign n10208 = ( ~n4615 & n6458 ) | ( ~n4615 & n8703 ) | ( n6458 & n8703 ) ;
  assign n10207 = n4370 ^ n2594 ^ n295 ;
  assign n10209 = n10208 ^ n10207 ^ 1'b0 ;
  assign n10210 = n10206 & n10209 ;
  assign n10211 = n1492 | n9842 ;
  assign n10212 = n10211 ^ n2822 ^ 1'b0 ;
  assign n10213 = ~n1340 & n4198 ;
  assign n10214 = n598 & n10213 ;
  assign n10215 = n2999 & ~n10214 ;
  assign n10216 = n10215 ^ n6201 ^ 1'b0 ;
  assign n10217 = ~n10212 & n10216 ;
  assign n10218 = n10217 ^ n2641 ^ 1'b0 ;
  assign n10219 = ( ~n5911 & n7229 ) | ( ~n5911 & n10218 ) | ( n7229 & n10218 ) ;
  assign n10220 = n3767 ^ n1286 ^ 1'b0 ;
  assign n10221 = n4463 ^ n2160 ^ 1'b0 ;
  assign n10222 = ( x94 & n2351 ) | ( x94 & n5665 ) | ( n2351 & n5665 ) ;
  assign n10223 = n10222 ^ n9568 ^ n9519 ;
  assign n10224 = n10223 ^ n5928 ^ n2242 ;
  assign n10229 = ~n3322 & n3375 ;
  assign n10225 = n9672 ^ n3398 ^ 1'b0 ;
  assign n10226 = x142 & n10225 ;
  assign n10227 = n4769 ^ n2662 ^ 1'b0 ;
  assign n10228 = n10226 & n10227 ;
  assign n10230 = n10229 ^ n10228 ^ n1455 ;
  assign n10231 = ~n2330 & n5234 ;
  assign n10232 = ~n5421 & n10231 ;
  assign n10233 = n10232 ^ n6948 ^ n3567 ;
  assign n10234 = n7952 ^ n270 ^ 1'b0 ;
  assign n10235 = n6763 | n10234 ;
  assign n10236 = ~n4396 & n5129 ;
  assign n10237 = n10236 ^ n9686 ^ n2834 ;
  assign n10238 = n7209 ^ n1958 ^ n1211 ;
  assign n10239 = n1784 | n10238 ;
  assign n10240 = n10239 ^ n4130 ^ n529 ;
  assign n10241 = ( n1116 & ~n8369 ) | ( n1116 & n10240 ) | ( ~n8369 & n10240 ) ;
  assign n10242 = ( n7257 & n10098 ) | ( n7257 & n10241 ) | ( n10098 & n10241 ) ;
  assign n10243 = ( n504 & n1699 ) | ( n504 & ~n4783 ) | ( n1699 & ~n4783 ) ;
  assign n10244 = n8779 ^ n525 ^ 1'b0 ;
  assign n10245 = ~n610 & n2734 ;
  assign n10246 = n517 & n10245 ;
  assign n10247 = n10246 ^ n2059 ^ n358 ;
  assign n10248 = ~n7022 & n10247 ;
  assign n10249 = ~n10244 & n10248 ;
  assign n10250 = n3896 & ~n10249 ;
  assign n10251 = n10250 ^ n8768 ^ 1'b0 ;
  assign n10252 = ( n2001 & ~n2301 ) | ( n2001 & n7659 ) | ( ~n2301 & n7659 ) ;
  assign n10253 = n9802 ^ n3989 ^ 1'b0 ;
  assign n10254 = n6505 & n10253 ;
  assign n10255 = n10254 ^ n3525 ^ n1461 ;
  assign n10264 = ~n5336 & n6203 ;
  assign n10265 = n10264 ^ n2099 ^ 1'b0 ;
  assign n10261 = n306 & ~n2458 ;
  assign n10262 = n10261 ^ n5093 ^ 1'b0 ;
  assign n10263 = n7805 & ~n10262 ;
  assign n10266 = n10265 ^ n10263 ^ n6418 ;
  assign n10256 = ( ~n1543 & n2814 ) | ( ~n1543 & n3825 ) | ( n2814 & n3825 ) ;
  assign n10257 = n5066 ^ n4932 ^ 1'b0 ;
  assign n10258 = n8239 & ~n10257 ;
  assign n10259 = ( n1010 & ~n4816 ) | ( n1010 & n10258 ) | ( ~n4816 & n10258 ) ;
  assign n10260 = n10256 | n10259 ;
  assign n10267 = n10266 ^ n10260 ^ 1'b0 ;
  assign n10268 = n10255 | n10267 ;
  assign n10269 = ( n840 & n10252 ) | ( n840 & n10268 ) | ( n10252 & n10268 ) ;
  assign n10274 = n1921 | n4465 ;
  assign n10270 = n2624 ^ n1173 ^ n591 ;
  assign n10271 = n5580 ^ n534 ^ 1'b0 ;
  assign n10272 = ~n8455 & n10271 ;
  assign n10273 = n10270 & n10272 ;
  assign n10275 = n10274 ^ n10273 ^ 1'b0 ;
  assign n10276 = n7214 ^ n4623 ^ 1'b0 ;
  assign n10277 = n1217 & n10276 ;
  assign n10278 = n6496 ^ n957 ^ n656 ;
  assign n10279 = n10278 ^ n6634 ^ 1'b0 ;
  assign n10280 = n10277 & ~n10279 ;
  assign n10281 = n1858 ^ n324 ^ 1'b0 ;
  assign n10282 = n7146 | n10281 ;
  assign n10283 = n6712 & ~n10282 ;
  assign n10285 = ( n916 & n4315 ) | ( n916 & n4660 ) | ( n4315 & n4660 ) ;
  assign n10284 = ~n4262 & n7040 ;
  assign n10286 = n10285 ^ n10284 ^ n1768 ;
  assign n10287 = n4209 ^ n684 ^ 1'b0 ;
  assign n10288 = n4902 & n5617 ;
  assign n10289 = ~n4626 & n10288 ;
  assign n10290 = n10287 & n10289 ;
  assign n10291 = n1114 | n6540 ;
  assign n10292 = n10291 ^ n10030 ^ 1'b0 ;
  assign n10298 = ~n557 & n7550 ;
  assign n10299 = n10298 ^ n6369 ^ 1'b0 ;
  assign n10293 = n5168 ^ n2838 ^ 1'b0 ;
  assign n10294 = n10191 ^ n9834 ^ n7347 ;
  assign n10295 = n10294 ^ x205 ^ 1'b0 ;
  assign n10296 = n10293 & n10295 ;
  assign n10297 = n4015 & n10296 ;
  assign n10300 = n10299 ^ n10297 ^ 1'b0 ;
  assign n10301 = ( n4439 & ~n10292 ) | ( n4439 & n10300 ) | ( ~n10292 & n10300 ) ;
  assign n10304 = n2086 | n5115 ;
  assign n10302 = n1213 & ~n1226 ;
  assign n10303 = n2694 | n10302 ;
  assign n10305 = n10304 ^ n10303 ^ n8664 ;
  assign n10306 = ( n6381 & n7390 ) | ( n6381 & n8952 ) | ( n7390 & n8952 ) ;
  assign n10307 = ( n509 & n5617 ) | ( n509 & ~n10306 ) | ( n5617 & ~n10306 ) ;
  assign n10308 = ~n3268 & n4786 ;
  assign n10309 = n10308 ^ n6855 ^ 1'b0 ;
  assign n10310 = n8078 ^ n7253 ^ n3080 ;
  assign n10311 = ( ~n2338 & n5634 ) | ( ~n2338 & n10310 ) | ( n5634 & n10310 ) ;
  assign n10312 = n3699 & ~n3810 ;
  assign n10314 = ( x223 & n2562 ) | ( x223 & ~n7195 ) | ( n2562 & ~n7195 ) ;
  assign n10315 = ( n2817 & ~n5676 ) | ( n2817 & n10314 ) | ( ~n5676 & n10314 ) ;
  assign n10313 = ~n3000 & n6320 ;
  assign n10316 = n10315 ^ n10313 ^ 1'b0 ;
  assign n10317 = ( n1901 & n4166 ) | ( n1901 & n6665 ) | ( n4166 & n6665 ) ;
  assign n10318 = n10317 ^ n6410 ^ n3898 ;
  assign n10319 = n8492 ^ n593 ^ 1'b0 ;
  assign n10320 = ( ~x64 & n1258 ) | ( ~x64 & n3314 ) | ( n1258 & n3314 ) ;
  assign n10321 = ( ~n4866 & n10319 ) | ( ~n4866 & n10320 ) | ( n10319 & n10320 ) ;
  assign n10322 = ( n3139 & ~n9376 ) | ( n3139 & n10321 ) | ( ~n9376 & n10321 ) ;
  assign n10323 = ~n884 & n3828 ;
  assign n10324 = ( n8575 & ~n8955 ) | ( n8575 & n10260 ) | ( ~n8955 & n10260 ) ;
  assign n10325 = n2984 ^ n394 ^ 1'b0 ;
  assign n10326 = ~n2424 & n10325 ;
  assign n10327 = n10201 ^ n710 ^ 1'b0 ;
  assign n10328 = n10327 ^ n2619 ^ n1245 ;
  assign n10329 = n485 & n6410 ;
  assign n10330 = n10329 ^ n6496 ^ 1'b0 ;
  assign n10331 = n10330 ^ n6825 ^ 1'b0 ;
  assign n10332 = ( n1877 & ~n9287 ) | ( n1877 & n9530 ) | ( ~n9287 & n9530 ) ;
  assign n10333 = n10094 ^ n4951 ^ n2428 ;
  assign n10334 = n1129 ^ n422 ^ x227 ;
  assign n10335 = n10334 ^ n9987 ^ n3219 ;
  assign n10337 = n2550 ^ n1526 ^ n1450 ;
  assign n10336 = ( x89 & n3163 ) | ( x89 & n5419 ) | ( n3163 & n5419 ) ;
  assign n10338 = n10337 ^ n10336 ^ 1'b0 ;
  assign n10339 = n10335 & n10338 ;
  assign n10340 = n6412 & n10339 ;
  assign n10341 = ~n3352 & n3439 ;
  assign n10342 = n10341 ^ n6876 ^ 1'b0 ;
  assign n10343 = ( n4546 & ~n4762 ) | ( n4546 & n10342 ) | ( ~n4762 & n10342 ) ;
  assign n10344 = n6181 ^ n5681 ^ 1'b0 ;
  assign n10345 = n6645 ^ n3546 ^ 1'b0 ;
  assign n10346 = ( n3109 & n10344 ) | ( n3109 & n10345 ) | ( n10344 & n10345 ) ;
  assign n10347 = n5093 | n10346 ;
  assign n10348 = n10343 | n10347 ;
  assign n10349 = n8042 ^ n6248 ^ 1'b0 ;
  assign n10351 = n1849 | n3495 ;
  assign n10350 = n7707 ^ n3482 ^ 1'b0 ;
  assign n10352 = n10351 ^ n10350 ^ 1'b0 ;
  assign n10353 = ( ~n4544 & n5615 ) | ( ~n4544 & n10352 ) | ( n5615 & n10352 ) ;
  assign n10354 = n10349 | n10353 ;
  assign n10355 = n6450 | n10354 ;
  assign n10356 = ( n1722 & n4300 ) | ( n1722 & ~n5839 ) | ( n4300 & ~n5839 ) ;
  assign n10357 = n2467 & n10356 ;
  assign n10358 = ~n1157 & n10357 ;
  assign n10359 = ~n3416 & n10358 ;
  assign n10360 = n10355 & ~n10359 ;
  assign n10361 = ~n8514 & n10360 ;
  assign n10362 = n5397 ^ n2460 ^ n1900 ;
  assign n10363 = ( n858 & ~n6476 ) | ( n858 & n10362 ) | ( ~n6476 & n10362 ) ;
  assign n10364 = n10363 ^ n8607 ^ n1054 ;
  assign n10365 = n10364 ^ n9616 ^ 1'b0 ;
  assign n10366 = n8651 | n10365 ;
  assign n10372 = n5007 & ~n6349 ;
  assign n10373 = ( n905 & ~n4752 ) | ( n905 & n10372 ) | ( ~n4752 & n10372 ) ;
  assign n10371 = n6756 ^ n5355 ^ n1624 ;
  assign n10367 = n4328 ^ n2637 ^ 1'b0 ;
  assign n10368 = n4221 & ~n10367 ;
  assign n10369 = n10368 ^ n9765 ^ n5427 ;
  assign n10370 = ( n5935 & ~n7947 ) | ( n5935 & n10369 ) | ( ~n7947 & n10369 ) ;
  assign n10374 = n10373 ^ n10371 ^ n10370 ;
  assign n10375 = ( x138 & ~n1130 ) | ( x138 & n1185 ) | ( ~n1130 & n1185 ) ;
  assign n10376 = ( n1118 & n4881 ) | ( n1118 & n10375 ) | ( n4881 & n10375 ) ;
  assign n10377 = ~n497 & n4924 ;
  assign n10378 = n4938 & ~n9526 ;
  assign n10379 = n10378 ^ n4767 ^ 1'b0 ;
  assign n10380 = n9403 ^ n3081 ^ n1271 ;
  assign n10381 = ( n8736 & n10379 ) | ( n8736 & n10380 ) | ( n10379 & n10380 ) ;
  assign n10382 = ( n2552 & ~n10377 ) | ( n2552 & n10381 ) | ( ~n10377 & n10381 ) ;
  assign n10383 = n5718 ^ n5355 ^ 1'b0 ;
  assign n10384 = n362 ^ n345 ^ 1'b0 ;
  assign n10385 = ( n3643 & ~n8596 ) | ( n3643 & n10384 ) | ( ~n8596 & n10384 ) ;
  assign n10386 = n10385 ^ n8324 ^ 1'b0 ;
  assign n10387 = n10383 | n10386 ;
  assign n10388 = n10387 ^ n3419 ^ 1'b0 ;
  assign n10389 = n6956 | n10388 ;
  assign n10390 = n10389 ^ n4757 ^ 1'b0 ;
  assign n10391 = n1616 | n7828 ;
  assign n10392 = n10391 ^ x183 ^ 1'b0 ;
  assign n10393 = n6499 & ~n10392 ;
  assign n10394 = ~n1226 & n1243 ;
  assign n10395 = n10394 ^ n556 ^ 1'b0 ;
  assign n10396 = ( n2960 & n9443 ) | ( n2960 & ~n10395 ) | ( n9443 & ~n10395 ) ;
  assign n10397 = n8028 & ~n10396 ;
  assign n10398 = n9089 ^ n2461 ^ 1'b0 ;
  assign n10399 = ~n3161 & n10398 ;
  assign n10400 = n975 & n8982 ;
  assign n10401 = n10400 ^ n4672 ^ n1199 ;
  assign n10402 = n1028 & n10401 ;
  assign n10403 = ~n10399 & n10402 ;
  assign n10404 = n10403 ^ n7942 ^ n3248 ;
  assign n10405 = ( n1556 & ~n5565 ) | ( n1556 & n8806 ) | ( ~n5565 & n8806 ) ;
  assign n10406 = n10405 ^ n8492 ^ n5747 ;
  assign n10407 = n5906 ^ n2027 ^ 1'b0 ;
  assign n10408 = n2571 & ~n10407 ;
  assign n10409 = n10408 ^ n9755 ^ n5655 ;
  assign n10410 = ( n1267 & n1346 ) | ( n1267 & ~n6761 ) | ( n1346 & ~n6761 ) ;
  assign n10411 = n3942 & n10410 ;
  assign n10412 = ~n2421 & n8199 ;
  assign n10413 = n3849 ^ n3710 ^ 1'b0 ;
  assign n10414 = n10412 | n10413 ;
  assign n10415 = n10414 ^ n3417 ^ 1'b0 ;
  assign n10416 = n10415 ^ n8219 ^ 1'b0 ;
  assign n10417 = n372 & ~n10416 ;
  assign n10418 = ( n1056 & n1734 ) | ( n1056 & n10417 ) | ( n1734 & n10417 ) ;
  assign n10419 = n10411 & n10418 ;
  assign n10420 = n7611 & n10419 ;
  assign n10421 = n7809 ^ n4131 ^ 1'b0 ;
  assign n10427 = n841 & n8138 ;
  assign n10428 = n2367 & n10427 ;
  assign n10426 = n9222 ^ n4995 ^ n1415 ;
  assign n10424 = n3715 & n8710 ;
  assign n10422 = ~n1528 & n2311 ;
  assign n10423 = n10422 ^ n3883 ^ 1'b0 ;
  assign n10425 = n10424 ^ n10423 ^ n6432 ;
  assign n10429 = n10428 ^ n10426 ^ n10425 ;
  assign n10430 = n9227 ^ n6468 ^ n2652 ;
  assign n10431 = n2416 & ~n10177 ;
  assign n10432 = n2121 & n10431 ;
  assign n10433 = n1078 & n10432 ;
  assign n10434 = n10433 ^ n6768 ^ 1'b0 ;
  assign n10435 = n5041 | n10434 ;
  assign n10436 = ( n765 & ~n2178 ) | ( n765 & n10435 ) | ( ~n2178 & n10435 ) ;
  assign n10437 = n4728 | n6872 ;
  assign n10438 = n9188 & ~n10437 ;
  assign n10439 = n1593 | n10438 ;
  assign n10440 = x5 & x25 ;
  assign n10441 = ( n4011 & n5433 ) | ( n4011 & ~n10440 ) | ( n5433 & ~n10440 ) ;
  assign n10442 = n2470 | n8510 ;
  assign n10443 = n10442 ^ n1724 ^ 1'b0 ;
  assign n10444 = ( n9842 & ~n10441 ) | ( n9842 & n10443 ) | ( ~n10441 & n10443 ) ;
  assign n10448 = ~n1226 & n3490 ;
  assign n10449 = ~n8419 & n10448 ;
  assign n10445 = ( ~n1418 & n2257 ) | ( ~n1418 & n6147 ) | ( n2257 & n6147 ) ;
  assign n10446 = n10445 ^ n5086 ^ n4923 ;
  assign n10447 = ~n6131 & n10446 ;
  assign n10450 = n10449 ^ n10447 ^ 1'b0 ;
  assign n10451 = n10450 ^ n9905 ^ n2061 ;
  assign n10456 = n8773 ^ n4210 ^ n346 ;
  assign n10455 = ~n2455 & n6878 ;
  assign n10457 = n10456 ^ n10455 ^ 1'b0 ;
  assign n10458 = x237 & ~n10457 ;
  assign n10452 = n5071 ^ n1030 ^ n948 ;
  assign n10453 = ( n4122 & n4642 ) | ( n4122 & n10452 ) | ( n4642 & n10452 ) ;
  assign n10454 = ( n491 & n564 ) | ( n491 & ~n10453 ) | ( n564 & ~n10453 ) ;
  assign n10459 = n10458 ^ n10454 ^ n3586 ;
  assign n10460 = n6030 & ~n8180 ;
  assign n10461 = ( ~n946 & n1518 ) | ( ~n946 & n2206 ) | ( n1518 & n2206 ) ;
  assign n10462 = n10461 ^ n9845 ^ n936 ;
  assign n10463 = ( n9238 & n10460 ) | ( n9238 & ~n10462 ) | ( n10460 & ~n10462 ) ;
  assign n10464 = x89 & ~n3796 ;
  assign n10465 = ( ~n1608 & n3273 ) | ( ~n1608 & n10464 ) | ( n3273 & n10464 ) ;
  assign n10466 = n6177 ^ n5068 ^ 1'b0 ;
  assign n10467 = n2045 & ~n10466 ;
  assign n10468 = n10467 ^ n4301 ^ x63 ;
  assign n10469 = n10465 | n10468 ;
  assign n10470 = n4283 ^ n1784 ^ 1'b0 ;
  assign n10471 = n7936 ^ n1304 ^ 1'b0 ;
  assign n10472 = n10470 & n10471 ;
  assign n10473 = ( ~n5213 & n10469 ) | ( ~n5213 & n10472 ) | ( n10469 & n10472 ) ;
  assign n10474 = n10463 & n10473 ;
  assign n10479 = ~n4268 & n9433 ;
  assign n10480 = n7381 & n10479 ;
  assign n10481 = n6399 & n10480 ;
  assign n10482 = ( n3590 & ~n8743 ) | ( n3590 & n10481 ) | ( ~n8743 & n10481 ) ;
  assign n10478 = n6161 | n6432 ;
  assign n10483 = n10482 ^ n10478 ^ 1'b0 ;
  assign n10475 = ~n2286 & n5213 ;
  assign n10476 = n6023 ^ n3655 ^ n481 ;
  assign n10477 = ~n10475 & n10476 ;
  assign n10484 = n10483 ^ n10477 ^ 1'b0 ;
  assign n10485 = ( ~n559 & n1800 ) | ( ~n559 & n5298 ) | ( n1800 & n5298 ) ;
  assign n10486 = n10186 & ~n10485 ;
  assign n10487 = n10486 ^ n8867 ^ 1'b0 ;
  assign n10488 = n4027 ^ n3151 ^ 1'b0 ;
  assign n10489 = n3425 | n4399 ;
  assign n10490 = n4629 | n10489 ;
  assign n10491 = ~n504 & n8357 ;
  assign n10492 = ( n10488 & ~n10490 ) | ( n10488 & n10491 ) | ( ~n10490 & n10491 ) ;
  assign n10493 = n4409 ^ n1331 ^ 1'b0 ;
  assign n10494 = x252 & ~n10493 ;
  assign n10495 = n6474 | n8649 ;
  assign n10496 = n10495 ^ n1914 ^ 1'b0 ;
  assign n10497 = n10494 & n10496 ;
  assign n10498 = n10497 ^ n8109 ^ n7471 ;
  assign n10499 = n2998 & n5601 ;
  assign n10500 = n5717 & n6481 ;
  assign n10501 = ( n2493 & n10499 ) | ( n2493 & n10500 ) | ( n10499 & n10500 ) ;
  assign n10509 = n6297 | n9513 ;
  assign n10510 = n4951 & ~n10509 ;
  assign n10503 = n8601 ^ n2903 ^ 1'b0 ;
  assign n10504 = n8750 | n10503 ;
  assign n10505 = n10504 ^ n7169 ^ n5531 ;
  assign n10502 = n6238 & ~n10197 ;
  assign n10506 = n10505 ^ n10502 ^ 1'b0 ;
  assign n10507 = n10506 ^ n6022 ^ 1'b0 ;
  assign n10508 = ( ~n6649 & n9769 ) | ( ~n6649 & n10507 ) | ( n9769 & n10507 ) ;
  assign n10511 = n10510 ^ n10508 ^ n1210 ;
  assign n10512 = ~n1511 & n2614 ;
  assign n10513 = n2199 & ~n3557 ;
  assign n10514 = n5214 & n10513 ;
  assign n10515 = n10512 & ~n10514 ;
  assign n10516 = n10515 ^ n9599 ^ 1'b0 ;
  assign n10517 = ( ~n3699 & n5799 ) | ( ~n3699 & n10197 ) | ( n5799 & n10197 ) ;
  assign n10518 = ( n9206 & ~n9738 ) | ( n9206 & n10517 ) | ( ~n9738 & n10517 ) ;
  assign n10519 = n7174 & ~n8886 ;
  assign n10520 = ~n6162 & n10519 ;
  assign n10521 = n10520 ^ n4816 ^ n593 ;
  assign n10522 = n6249 ^ n4635 ^ n897 ;
  assign n10523 = ( ~n971 & n10521 ) | ( ~n971 & n10522 ) | ( n10521 & n10522 ) ;
  assign n10524 = n8801 ^ n5726 ^ n3989 ;
  assign n10525 = n10524 ^ n10492 ^ n7671 ;
  assign n10530 = n6245 ^ n3663 ^ n603 ;
  assign n10531 = n10530 ^ n7376 ^ n1326 ;
  assign n10528 = n304 | n793 ;
  assign n10529 = n636 & ~n10528 ;
  assign n10532 = n10531 ^ n10529 ^ n941 ;
  assign n10533 = n10488 ^ n8893 ^ n6246 ;
  assign n10534 = n4580 ^ n2734 ^ 1'b0 ;
  assign n10535 = n10533 & ~n10534 ;
  assign n10536 = ( n454 & n10532 ) | ( n454 & n10535 ) | ( n10532 & n10535 ) ;
  assign n10526 = n7692 ^ n7429 ^ 1'b0 ;
  assign n10527 = ~n7290 & n10526 ;
  assign n10537 = n10536 ^ n10527 ^ 1'b0 ;
  assign n10538 = ~n3090 & n10155 ;
  assign n10539 = ( n5347 & n9688 ) | ( n5347 & ~n10538 ) | ( n9688 & ~n10538 ) ;
  assign n10540 = n10539 ^ n10397 ^ 1'b0 ;
  assign n10541 = n4672 & ~n7079 ;
  assign n10542 = n974 | n10541 ;
  assign n10543 = n5072 | n10542 ;
  assign n10544 = n9623 ^ n1434 ^ 1'b0 ;
  assign n10545 = n10544 ^ n270 ^ 1'b0 ;
  assign n10546 = n4198 ^ n2180 ^ x221 ;
  assign n10547 = n1089 & n7507 ;
  assign n10548 = ( n7835 & n10546 ) | ( n7835 & n10547 ) | ( n10546 & n10547 ) ;
  assign n10549 = n6709 | n8376 ;
  assign n10550 = ( n1310 & n5981 ) | ( n1310 & ~n8027 ) | ( n5981 & ~n8027 ) ;
  assign n10551 = n10134 ^ n5896 ^ 1'b0 ;
  assign n10552 = n10551 ^ n6051 ^ n1543 ;
  assign n10553 = n10552 ^ n9351 ^ n8060 ;
  assign n10554 = n10550 & ~n10553 ;
  assign n10555 = n10549 & n10554 ;
  assign n10556 = n10555 ^ n9167 ^ n4582 ;
  assign n10557 = n10548 & ~n10556 ;
  assign n10558 = n10557 ^ n1587 ^ 1'b0 ;
  assign n10559 = n2083 & ~n6621 ;
  assign n10560 = n4274 ^ n3309 ^ n3204 ;
  assign n10561 = ( n5480 & n8896 ) | ( n5480 & n9144 ) | ( n8896 & n9144 ) ;
  assign n10562 = n7475 ^ n883 ^ 1'b0 ;
  assign n10563 = ~n7527 & n10562 ;
  assign n10564 = ( n10560 & n10561 ) | ( n10560 & ~n10563 ) | ( n10561 & ~n10563 ) ;
  assign n10565 = ( n6501 & ~n10523 ) | ( n6501 & n10564 ) | ( ~n10523 & n10564 ) ;
  assign n10566 = ~n4193 & n5806 ;
  assign n10567 = n7440 & n10566 ;
  assign n10568 = n4744 & ~n10567 ;
  assign n10569 = n10568 ^ n8956 ^ 1'b0 ;
  assign n10570 = n5886 ^ n1109 ^ 1'b0 ;
  assign n10571 = n10570 ^ n5755 ^ n1848 ;
  assign n10572 = ( n3117 & ~n5323 ) | ( n3117 & n10571 ) | ( ~n5323 & n10571 ) ;
  assign n10578 = n6702 ^ n4430 ^ 1'b0 ;
  assign n10579 = n10578 ^ n5848 ^ 1'b0 ;
  assign n10573 = ( n2392 & n3713 ) | ( n2392 & ~n5732 ) | ( n3713 & ~n5732 ) ;
  assign n10574 = n1489 & n10573 ;
  assign n10575 = n4594 | n5310 ;
  assign n10576 = n10575 ^ n7503 ^ 1'b0 ;
  assign n10577 = ( n3527 & n10574 ) | ( n3527 & ~n10576 ) | ( n10574 & ~n10576 ) ;
  assign n10580 = n10579 ^ n10577 ^ 1'b0 ;
  assign n10581 = n4813 ^ n3939 ^ 1'b0 ;
  assign n10582 = n2166 & n10581 ;
  assign n10583 = ~n2770 & n10582 ;
  assign n10584 = n10583 ^ n1430 ^ 1'b0 ;
  assign n10585 = ( n3061 & n4996 ) | ( n3061 & ~n10584 ) | ( n4996 & ~n10584 ) ;
  assign n10586 = x153 & ~n1112 ;
  assign n10587 = n10586 ^ n8111 ^ 1'b0 ;
  assign n10588 = n10587 ^ n8122 ^ n2214 ;
  assign n10589 = ( n2960 & n5710 ) | ( n2960 & n6608 ) | ( n5710 & n6608 ) ;
  assign n10590 = ( ~n10585 & n10588 ) | ( ~n10585 & n10589 ) | ( n10588 & n10589 ) ;
  assign n10591 = ~n2829 & n5041 ;
  assign n10592 = n2112 | n10591 ;
  assign n10593 = n10592 ^ n6190 ^ n2598 ;
  assign n10594 = ( n916 & n2659 ) | ( n916 & n6739 ) | ( n2659 & n6739 ) ;
  assign n10595 = n6148 ^ n5759 ^ 1'b0 ;
  assign n10596 = ~n6540 & n10595 ;
  assign n10597 = n10596 ^ n8857 ^ n7021 ;
  assign n10598 = ~x230 & n10597 ;
  assign n10599 = n10413 ^ n7584 ^ n1020 ;
  assign n10600 = n10599 ^ n4018 ^ x5 ;
  assign n10601 = n2338 & ~n8757 ;
  assign n10602 = n8274 & n10601 ;
  assign n10605 = n518 | n1883 ;
  assign n10606 = n2140 & ~n10605 ;
  assign n10603 = n4128 | n6469 ;
  assign n10604 = n2350 & ~n10603 ;
  assign n10607 = n10606 ^ n10604 ^ n9754 ;
  assign n10609 = n9242 ^ n5139 ^ n4338 ;
  assign n10608 = n8904 ^ n4279 ^ 1'b0 ;
  assign n10610 = n10609 ^ n10608 ^ n4404 ;
  assign n10611 = n374 & ~n8528 ;
  assign n10618 = n3148 ^ x8 ^ 1'b0 ;
  assign n10619 = n9560 | n10618 ;
  assign n10614 = n4822 ^ n772 ^ 1'b0 ;
  assign n10615 = ~n884 & n10614 ;
  assign n10616 = n10615 ^ n3608 ^ n520 ;
  assign n10613 = ( ~n1302 & n5031 ) | ( ~n1302 & n6994 ) | ( n5031 & n6994 ) ;
  assign n10612 = n2569 ^ n888 ^ 1'b0 ;
  assign n10617 = n10616 ^ n10613 ^ n10612 ;
  assign n10620 = n10619 ^ n10617 ^ n8233 ;
  assign n10625 = n4839 ^ n780 ^ n575 ;
  assign n10621 = n8407 ^ n5470 ^ n3792 ;
  assign n10622 = n3881 & n10173 ;
  assign n10623 = n2538 & n10622 ;
  assign n10624 = n10621 & ~n10623 ;
  assign n10626 = n10625 ^ n10624 ^ 1'b0 ;
  assign n10627 = n7838 ^ n5618 ^ n4881 ;
  assign n10628 = x85 & n10627 ;
  assign n10629 = n10628 ^ n7735 ^ 1'b0 ;
  assign n10630 = ~n1449 & n4465 ;
  assign n10631 = n10630 ^ n4646 ^ 1'b0 ;
  assign n10632 = ~n4409 & n4817 ;
  assign n10633 = ( n10153 & n10631 ) | ( n10153 & ~n10632 ) | ( n10631 & ~n10632 ) ;
  assign n10634 = ( n4351 & n4499 ) | ( n4351 & ~n10092 ) | ( n4499 & ~n10092 ) ;
  assign n10635 = n4298 & ~n10634 ;
  assign n10636 = n2746 ^ n1766 ^ n828 ;
  assign n10637 = ~n9290 & n9544 ;
  assign n10638 = ~n2796 & n10637 ;
  assign n10639 = n10638 ^ n6999 ^ 1'b0 ;
  assign n10640 = ( n5531 & ~n10636 ) | ( n5531 & n10639 ) | ( ~n10636 & n10639 ) ;
  assign n10641 = n1537 & ~n6384 ;
  assign n10642 = n2751 | n4700 ;
  assign n10643 = n5885 | n10642 ;
  assign n10644 = n10641 & ~n10643 ;
  assign n10645 = ( n8086 & n10640 ) | ( n8086 & n10644 ) | ( n10640 & n10644 ) ;
  assign n10646 = n7689 ^ n4721 ^ 1'b0 ;
  assign n10647 = ~n4343 & n10646 ;
  assign n10648 = n2444 & n3586 ;
  assign n10649 = ~n10647 & n10648 ;
  assign n10650 = n10314 | n10649 ;
  assign n10651 = n3421 & ~n10650 ;
  assign n10652 = ( n2237 & n5431 ) | ( n2237 & ~n10651 ) | ( n5431 & ~n10651 ) ;
  assign n10653 = ( x170 & n818 ) | ( x170 & ~n858 ) | ( n818 & ~n858 ) ;
  assign n10654 = n8915 ^ n2832 ^ n593 ;
  assign n10655 = n1893 | n4176 ;
  assign n10656 = n10654 & ~n10655 ;
  assign n10657 = ( n7553 & n10653 ) | ( n7553 & n10656 ) | ( n10653 & n10656 ) ;
  assign n10658 = n10657 ^ x155 ^ 1'b0 ;
  assign n10659 = n7298 ^ n6327 ^ n6035 ;
  assign n10660 = n7876 ^ n3439 ^ n3064 ;
  assign n10669 = ( n1718 & n2915 ) | ( n1718 & ~n3355 ) | ( n2915 & ~n3355 ) ;
  assign n10663 = n2843 & ~n3101 ;
  assign n10664 = n7384 & n10663 ;
  assign n10665 = n1794 & n10664 ;
  assign n10666 = n5262 ^ n5115 ^ 1'b0 ;
  assign n10667 = n10665 | n10666 ;
  assign n10668 = x85 & n10667 ;
  assign n10661 = n8245 ^ n7832 ^ n5728 ;
  assign n10662 = ( n6615 & ~n10115 ) | ( n6615 & n10661 ) | ( ~n10115 & n10661 ) ;
  assign n10670 = n10669 ^ n10668 ^ n10662 ;
  assign n10671 = n5451 ^ n3885 ^ n1675 ;
  assign n10672 = ( x61 & ~n1632 ) | ( x61 & n2417 ) | ( ~n1632 & n2417 ) ;
  assign n10673 = n1703 & n10672 ;
  assign n10674 = n7631 & ~n10673 ;
  assign n10675 = n10674 ^ n10524 ^ 1'b0 ;
  assign n10676 = n10671 & ~n10675 ;
  assign n10681 = n10127 ^ n1183 ^ 1'b0 ;
  assign n10677 = n1420 & ~n4220 ;
  assign n10678 = ( n1642 & n3865 ) | ( n1642 & n4654 ) | ( n3865 & n4654 ) ;
  assign n10679 = ( ~n3640 & n10677 ) | ( ~n3640 & n10678 ) | ( n10677 & n10678 ) ;
  assign n10680 = ( n2441 & ~n4134 ) | ( n2441 & n10679 ) | ( ~n4134 & n10679 ) ;
  assign n10682 = n10681 ^ n10680 ^ 1'b0 ;
  assign n10683 = n7347 & ~n8659 ;
  assign n10684 = n6989 & ~n9182 ;
  assign n10689 = n10068 ^ n6354 ^ 1'b0 ;
  assign n10685 = ( n5799 & ~n6135 ) | ( n5799 & n6430 ) | ( ~n6135 & n6430 ) ;
  assign n10686 = n10685 ^ n2057 ^ 1'b0 ;
  assign n10687 = n3827 & ~n10686 ;
  assign n10688 = n4319 & n10687 ;
  assign n10690 = n10689 ^ n10688 ^ 1'b0 ;
  assign n10691 = n10690 ^ n765 ^ 1'b0 ;
  assign n10692 = n2467 ^ n1617 ^ 1'b0 ;
  assign n10693 = ( n8727 & n8871 ) | ( n8727 & n10692 ) | ( n8871 & n10692 ) ;
  assign n10707 = n3871 ^ n3184 ^ n701 ;
  assign n10696 = n7008 ^ n4936 ^ n2769 ;
  assign n10697 = n10696 ^ n1163 ^ 1'b0 ;
  assign n10698 = n2433 & ~n10697 ;
  assign n10699 = n10698 ^ n7722 ^ 1'b0 ;
  assign n10700 = n1064 & ~n2099 ;
  assign n10701 = n5984 & n10700 ;
  assign n10702 = n4772 ^ n3377 ^ 1'b0 ;
  assign n10703 = n7248 | n10702 ;
  assign n10704 = n10701 & ~n10703 ;
  assign n10705 = n10704 ^ n557 ^ 1'b0 ;
  assign n10706 = ~n10699 & n10705 ;
  assign n10694 = n1374 ^ n645 ^ 1'b0 ;
  assign n10695 = n9138 & ~n10694 ;
  assign n10708 = n10707 ^ n10706 ^ n10695 ;
  assign n10714 = n1831 & ~n7544 ;
  assign n10715 = ~n8117 & n10714 ;
  assign n10709 = ( ~x117 & n2171 ) | ( ~x117 & n4582 ) | ( n2171 & n4582 ) ;
  assign n10710 = ( ~n1075 & n4876 ) | ( ~n1075 & n6446 ) | ( n4876 & n6446 ) ;
  assign n10711 = n9473 | n10710 ;
  assign n10712 = n10709 & ~n10711 ;
  assign n10713 = n2679 | n10712 ;
  assign n10716 = n10715 ^ n10713 ^ n6566 ;
  assign n10717 = ( ~n3878 & n5260 ) | ( ~n3878 & n6611 ) | ( n5260 & n6611 ) ;
  assign n10718 = n10717 ^ n9926 ^ n9802 ;
  assign n10720 = n2807 ^ n1840 ^ n805 ;
  assign n10721 = ~n2213 & n7490 ;
  assign n10722 = n10720 & n10721 ;
  assign n10719 = n8591 & n9199 ;
  assign n10723 = n10722 ^ n10719 ^ 1'b0 ;
  assign n10724 = ( x228 & n4659 ) | ( x228 & ~n7618 ) | ( n4659 & ~n7618 ) ;
  assign n10725 = ( ~n2922 & n4015 ) | ( ~n2922 & n10724 ) | ( n4015 & n10724 ) ;
  assign n10726 = n3476 & ~n7537 ;
  assign n10727 = n3752 & n10726 ;
  assign n10728 = n2695 & ~n10727 ;
  assign n10729 = ~n6201 & n6806 ;
  assign n10730 = n427 & n10729 ;
  assign n10731 = n7899 ^ n852 ^ 1'b0 ;
  assign n10732 = ~n3770 & n10731 ;
  assign n10733 = n10732 ^ n7537 ^ 1'b0 ;
  assign n10734 = n9114 & ~n10507 ;
  assign n10735 = n10734 ^ n1005 ^ 1'b0 ;
  assign n10736 = n4152 ^ n1590 ^ 1'b0 ;
  assign n10737 = ( n4066 & n5507 ) | ( n4066 & n7228 ) | ( n5507 & n7228 ) ;
  assign n10738 = n10737 ^ n3750 ^ n796 ;
  assign n10739 = ( n9780 & ~n10736 ) | ( n9780 & n10738 ) | ( ~n10736 & n10738 ) ;
  assign n10740 = n6174 ^ n5085 ^ x171 ;
  assign n10741 = n5086 | n10740 ;
  assign n10742 = n10741 ^ n7640 ^ 1'b0 ;
  assign n10743 = n5411 & ~n5486 ;
  assign n10744 = n8007 ^ n2062 ^ 1'b0 ;
  assign n10745 = n1508 & n10744 ;
  assign n10746 = n10743 & n10745 ;
  assign n10747 = n2808 ^ n1626 ^ 1'b0 ;
  assign n10748 = n10746 | n10747 ;
  assign n10749 = ( n2315 & n9380 ) | ( n2315 & ~n10748 ) | ( n9380 & ~n10748 ) ;
  assign n10750 = n10742 & n10749 ;
  assign n10751 = n10750 ^ n6544 ^ 1'b0 ;
  assign n10754 = n7497 ^ n2946 ^ 1'b0 ;
  assign n10755 = n7746 & n10754 ;
  assign n10756 = n10755 ^ n4193 ^ n725 ;
  assign n10757 = ~n4885 & n10756 ;
  assign n10758 = ~n6031 & n10757 ;
  assign n10752 = ~n5370 & n7186 ;
  assign n10753 = ~n1162 & n10752 ;
  assign n10759 = n10758 ^ n10753 ^ 1'b0 ;
  assign n10760 = n4493 & n10759 ;
  assign n10761 = ( ~n2755 & n5293 ) | ( ~n2755 & n6069 ) | ( n5293 & n6069 ) ;
  assign n10762 = n10760 & n10761 ;
  assign n10763 = n10751 & n10762 ;
  assign n10764 = n4553 & n6026 ;
  assign n10765 = n5150 & n10764 ;
  assign n10766 = n10765 ^ n9053 ^ 1'b0 ;
  assign n10767 = n5663 | n10766 ;
  assign n10768 = n10767 ^ n3884 ^ 1'b0 ;
  assign n10780 = ( x66 & ~n6062 ) | ( x66 & n6423 ) | ( ~n6062 & n6423 ) ;
  assign n10781 = ~n8478 & n10780 ;
  assign n10774 = n3923 | n8754 ;
  assign n10775 = n3213 & n10774 ;
  assign n10776 = n10775 ^ n1326 ^ 1'b0 ;
  assign n10777 = ( ~n1671 & n4412 ) | ( ~n1671 & n10776 ) | ( n4412 & n10776 ) ;
  assign n10769 = ( ~n372 & n596 ) | ( ~n372 & n9467 ) | ( n596 & n9467 ) ;
  assign n10770 = ( x232 & n4876 ) | ( x232 & n9039 ) | ( n4876 & n9039 ) ;
  assign n10771 = ~n10769 & n10770 ;
  assign n10772 = n704 & n10771 ;
  assign n10773 = n10772 ^ n6817 ^ n1277 ;
  assign n10778 = n10777 ^ n10773 ^ n6103 ;
  assign n10779 = ( n4283 & n4662 ) | ( n4283 & ~n10778 ) | ( n4662 & ~n10778 ) ;
  assign n10782 = n10781 ^ n10779 ^ n6248 ;
  assign n10783 = n8059 | n9971 ;
  assign n10784 = n10783 ^ n4723 ^ 1'b0 ;
  assign n10785 = n10784 ^ n9418 ^ 1'b0 ;
  assign n10786 = ( n1028 & n1966 ) | ( n1028 & ~n10785 ) | ( n1966 & ~n10785 ) ;
  assign n10787 = n7411 ^ n4328 ^ 1'b0 ;
  assign n10788 = ( n1228 & ~n3612 ) | ( n1228 & n10787 ) | ( ~n3612 & n10787 ) ;
  assign n10792 = ~n3659 & n6399 ;
  assign n10791 = n4501 & ~n6655 ;
  assign n10793 = n10792 ^ n10791 ^ 1'b0 ;
  assign n10789 = n7018 ^ n4100 ^ n282 ;
  assign n10790 = n10789 ^ n3416 ^ n2613 ;
  assign n10794 = n10793 ^ n10790 ^ n5700 ;
  assign n10796 = n7829 ^ n1183 ^ x167 ;
  assign n10795 = n526 & n3565 ;
  assign n10797 = n10796 ^ n10795 ^ n8168 ;
  assign n10798 = n4213 ^ n4206 ^ 1'b0 ;
  assign n10799 = n3178 & ~n10798 ;
  assign n10802 = n5093 ^ n3309 ^ n624 ;
  assign n10800 = n4071 & ~n6169 ;
  assign n10801 = ( ~n6448 & n7850 ) | ( ~n6448 & n10800 ) | ( n7850 & n10800 ) ;
  assign n10803 = n10802 ^ n10801 ^ n9394 ;
  assign n10804 = n2847 ^ n1002 ^ n536 ;
  assign n10805 = n4348 ^ n812 ^ 1'b0 ;
  assign n10806 = ~n6048 & n10805 ;
  assign n10807 = ( n9911 & n10804 ) | ( n9911 & n10806 ) | ( n10804 & n10806 ) ;
  assign n10808 = n5840 ^ n2271 ^ n536 ;
  assign n10809 = ( n7525 & n9060 ) | ( n7525 & ~n10808 ) | ( n9060 & ~n10808 ) ;
  assign n10810 = n4300 & ~n5997 ;
  assign n10811 = n5347 ^ n3754 ^ 1'b0 ;
  assign n10812 = n9220 ^ n3097 ^ 1'b0 ;
  assign n10813 = n2228 | n10812 ;
  assign n10814 = ( n1311 & ~n5475 ) | ( n1311 & n10813 ) | ( ~n5475 & n10813 ) ;
  assign n10816 = n1508 & ~n7152 ;
  assign n10817 = ~x230 & n10816 ;
  assign n10818 = n10817 ^ n594 ^ 1'b0 ;
  assign n10819 = n1261 & n10818 ;
  assign n10815 = n4302 ^ n2813 ^ n2283 ;
  assign n10820 = n10819 ^ n10815 ^ n2513 ;
  assign n10821 = ( n1760 & ~n1807 ) | ( n1760 & n3266 ) | ( ~n1807 & n3266 ) ;
  assign n10822 = n10821 ^ n7718 ^ n4169 ;
  assign n10823 = ( n6408 & n10820 ) | ( n6408 & ~n10822 ) | ( n10820 & ~n10822 ) ;
  assign n10824 = ( n4061 & n9914 ) | ( n4061 & ~n10823 ) | ( n9914 & ~n10823 ) ;
  assign n10825 = ( ~n945 & n4078 ) | ( ~n945 & n4721 ) | ( n4078 & n4721 ) ;
  assign n10826 = ~n3426 & n7197 ;
  assign n10827 = n10826 ^ n6954 ^ n3261 ;
  assign n10828 = ( n2520 & n10825 ) | ( n2520 & ~n10827 ) | ( n10825 & ~n10827 ) ;
  assign n10829 = ( n10814 & n10824 ) | ( n10814 & n10828 ) | ( n10824 & n10828 ) ;
  assign n10830 = ( n688 & n1302 ) | ( n688 & ~n2043 ) | ( n1302 & ~n2043 ) ;
  assign n10831 = n8357 ^ x157 ^ 1'b0 ;
  assign n10832 = ( x29 & ~n3441 ) | ( x29 & n3770 ) | ( ~n3441 & n3770 ) ;
  assign n10833 = ( ~n497 & n8858 ) | ( ~n497 & n10832 ) | ( n8858 & n10832 ) ;
  assign n10834 = n10833 ^ n3208 ^ 1'b0 ;
  assign n10835 = ( n10830 & ~n10831 ) | ( n10830 & n10834 ) | ( ~n10831 & n10834 ) ;
  assign n10836 = ( n3374 & n4373 ) | ( n3374 & ~n7880 ) | ( n4373 & ~n7880 ) ;
  assign n10837 = ( ~n393 & n10304 ) | ( ~n393 & n10836 ) | ( n10304 & n10836 ) ;
  assign n10838 = n10837 ^ n689 ^ n317 ;
  assign n10839 = n8500 ^ n3187 ^ 1'b0 ;
  assign n10840 = ~n514 & n10839 ;
  assign n10841 = n6961 & n10840 ;
  assign n10842 = n10838 & n10841 ;
  assign n10843 = n10232 ^ n2615 ^ 1'b0 ;
  assign n10845 = ~n5284 & n5486 ;
  assign n10844 = n8170 ^ n5826 ^ x250 ;
  assign n10846 = n10845 ^ n10844 ^ n7083 ;
  assign n10853 = n1296 | n8026 ;
  assign n10854 = n5451 & ~n10853 ;
  assign n10855 = n10854 ^ n9167 ^ 1'b0 ;
  assign n10847 = n3490 & ~n5744 ;
  assign n10848 = n10847 ^ n4770 ^ 1'b0 ;
  assign n10849 = n3309 ^ n1583 ^ n819 ;
  assign n10850 = n10849 ^ n3835 ^ n3818 ;
  assign n10851 = n7729 & ~n10850 ;
  assign n10852 = n10848 & n10851 ;
  assign n10856 = n10855 ^ n10852 ^ n3468 ;
  assign n10857 = n10224 & ~n10856 ;
  assign n10858 = ~n10846 & n10857 ;
  assign n10859 = x184 & ~n4274 ;
  assign n10860 = n9258 ^ n5258 ^ 1'b0 ;
  assign n10861 = n10859 & n10860 ;
  assign n10862 = ( n2911 & n3835 ) | ( n2911 & ~n10861 ) | ( n3835 & ~n10861 ) ;
  assign n10863 = ( n969 & ~n8674 ) | ( n969 & n10862 ) | ( ~n8674 & n10862 ) ;
  assign n10864 = n8563 & ~n10454 ;
  assign n10865 = n1267 & ~n3231 ;
  assign n10866 = n10865 ^ n325 ^ 1'b0 ;
  assign n10867 = x167 & n10866 ;
  assign n10868 = n6421 ^ n6206 ^ 1'b0 ;
  assign n10869 = n4317 & n10868 ;
  assign n10870 = n3011 & n5469 ;
  assign n10871 = ( n7070 & n10869 ) | ( n7070 & n10870 ) | ( n10869 & n10870 ) ;
  assign n10872 = n10871 ^ n8229 ^ n7748 ;
  assign n10873 = ~n6655 & n10872 ;
  assign n10874 = n885 & n9463 ;
  assign n10875 = ( n1336 & n2882 ) | ( n1336 & ~n3560 ) | ( n2882 & ~n3560 ) ;
  assign n10876 = n8305 ^ n8284 ^ n3949 ;
  assign n10877 = ( n1955 & n7877 ) | ( n1955 & ~n10876 ) | ( n7877 & ~n10876 ) ;
  assign n10879 = ~n6232 & n9973 ;
  assign n10880 = n10879 ^ n1420 ^ 1'b0 ;
  assign n10878 = n5363 & ~n5551 ;
  assign n10881 = n10880 ^ n10878 ^ 1'b0 ;
  assign n10882 = n10881 ^ n8830 ^ 1'b0 ;
  assign n10883 = n8876 & n10882 ;
  assign n10884 = ( n4866 & n4950 ) | ( n4866 & n9319 ) | ( n4950 & n9319 ) ;
  assign n10885 = n10884 ^ n5342 ^ 1'b0 ;
  assign n10886 = ( ~n1046 & n9856 ) | ( ~n1046 & n10885 ) | ( n9856 & n10885 ) ;
  assign n10887 = ( n2583 & n3604 ) | ( n2583 & ~n10886 ) | ( n3604 & ~n10886 ) ;
  assign n10888 = n4627 ^ n466 ^ 1'b0 ;
  assign n10889 = ~n10887 & n10888 ;
  assign n10890 = n10463 ^ n1382 ^ 1'b0 ;
  assign n10891 = n9027 ^ n1227 ^ 1'b0 ;
  assign n10892 = n2030 | n6737 ;
  assign n10893 = n8907 ^ n7858 ^ 1'b0 ;
  assign n10894 = n9314 ^ n5168 ^ 1'b0 ;
  assign n10895 = ~n10025 & n10894 ;
  assign n10896 = n9544 ^ n8919 ^ n957 ;
  assign n10897 = n7453 | n8995 ;
  assign n10898 = ( n1246 & n4087 ) | ( n1246 & n10897 ) | ( n4087 & n10897 ) ;
  assign n10899 = n2173 ^ n640 ^ 1'b0 ;
  assign n10900 = n8002 | n10899 ;
  assign n10901 = x23 & ~n10900 ;
  assign n10902 = n10901 ^ n491 ^ 1'b0 ;
  assign n10903 = ( n10896 & ~n10898 ) | ( n10896 & n10902 ) | ( ~n10898 & n10902 ) ;
  assign n10904 = n3124 ^ n1296 ^ 1'b0 ;
  assign n10905 = n10904 ^ n7051 ^ 1'b0 ;
  assign n10906 = ( x190 & x254 ) | ( x190 & ~n10905 ) | ( x254 & ~n10905 ) ;
  assign n10907 = ~n2247 & n3363 ;
  assign n10908 = ( ~n2669 & n5665 ) | ( ~n2669 & n10907 ) | ( n5665 & n10907 ) ;
  assign n10909 = ( x136 & ~n2717 ) | ( x136 & n9233 ) | ( ~n2717 & n9233 ) ;
  assign n10915 = n3732 ^ n3089 ^ n3037 ;
  assign n10912 = n10732 ^ n9836 ^ 1'b0 ;
  assign n10913 = n7811 & n10912 ;
  assign n10910 = n4166 & ~n5593 ;
  assign n10911 = n8592 & n10910 ;
  assign n10914 = n10913 ^ n10911 ^ n6027 ;
  assign n10916 = n10915 ^ n10914 ^ n4640 ;
  assign n10920 = n9643 ^ n1706 ^ 1'b0 ;
  assign n10917 = ~n683 & n5363 ;
  assign n10918 = n10917 ^ n2432 ^ n634 ;
  assign n10919 = ( ~n2210 & n7117 ) | ( ~n2210 & n10918 ) | ( n7117 & n10918 ) ;
  assign n10921 = n10920 ^ n10919 ^ n2422 ;
  assign n10922 = n6564 | n10921 ;
  assign n10930 = ( ~n5836 & n7097 ) | ( ~n5836 & n7381 ) | ( n7097 & n7381 ) ;
  assign n10925 = n3285 | n3615 ;
  assign n10926 = n10925 ^ n8413 ^ 1'b0 ;
  assign n10927 = ( ~n4240 & n8340 ) | ( ~n4240 & n10926 ) | ( n8340 & n10926 ) ;
  assign n10928 = n10927 ^ n3823 ^ n3094 ;
  assign n10929 = n10928 ^ n6111 ^ 1'b0 ;
  assign n10923 = n6610 ^ n2574 ^ 1'b0 ;
  assign n10924 = n4533 & n10923 ;
  assign n10931 = n10930 ^ n10929 ^ n10924 ;
  assign n10932 = n8768 & ~n10931 ;
  assign n10933 = n7966 & n10932 ;
  assign n10934 = n1043 ^ x90 ^ 1'b0 ;
  assign n10935 = ~n4078 & n10934 ;
  assign n10936 = ( n1651 & n3884 ) | ( n1651 & ~n10935 ) | ( n3884 & ~n10935 ) ;
  assign n10937 = ( x220 & n303 ) | ( x220 & n10936 ) | ( n303 & n10936 ) ;
  assign n10941 = ~x136 & n2448 ;
  assign n10938 = n7270 ^ n6197 ^ 1'b0 ;
  assign n10939 = ~n3211 & n10938 ;
  assign n10940 = ~n4448 & n10939 ;
  assign n10942 = n10941 ^ n10940 ^ 1'b0 ;
  assign n10943 = n10942 ^ n5576 ^ 1'b0 ;
  assign n10944 = n6944 & n9719 ;
  assign n10945 = n10944 ^ n8888 ^ 1'b0 ;
  assign n10946 = n1216 & ~n5200 ;
  assign n10947 = n10946 ^ n9482 ^ 1'b0 ;
  assign n10948 = n10945 & ~n10947 ;
  assign n10949 = ( n1606 & n2504 ) | ( n1606 & ~n5364 ) | ( n2504 & ~n5364 ) ;
  assign n10950 = n7165 ^ n4507 ^ 1'b0 ;
  assign n10951 = n1830 & n10950 ;
  assign n10952 = n2744 | n3454 ;
  assign n10953 = n10952 ^ n5048 ^ n4418 ;
  assign n10954 = n8817 ^ n775 ^ 1'b0 ;
  assign n10955 = ~n9856 & n10954 ;
  assign n10956 = n3807 & n10955 ;
  assign n10957 = n10956 ^ n3640 ^ 1'b0 ;
  assign n10958 = ~n3264 & n10813 ;
  assign n10959 = n10958 ^ n8738 ^ 1'b0 ;
  assign n10960 = n6565 & ~n6700 ;
  assign n10961 = ( n2357 & n7477 ) | ( n2357 & n9373 ) | ( n7477 & n9373 ) ;
  assign n10962 = n7708 & n10961 ;
  assign n10963 = n10962 ^ n899 ^ 1'b0 ;
  assign n10964 = x155 & n10700 ;
  assign n10965 = n10964 ^ n3344 ^ 1'b0 ;
  assign n10966 = n9270 & ~n10965 ;
  assign n10967 = n6301 & ~n6995 ;
  assign n10968 = n10359 & n10967 ;
  assign n10969 = n10968 ^ n8206 ^ 1'b0 ;
  assign n10970 = n7810 | n10969 ;
  assign n10971 = n6312 & ~n10970 ;
  assign n10972 = n8479 ^ n4865 ^ 1'b0 ;
  assign n10973 = n1673 ^ x137 ^ 1'b0 ;
  assign n10974 = n10972 & ~n10973 ;
  assign n10975 = n10974 ^ n2195 ^ 1'b0 ;
  assign n10976 = ( n438 & n610 ) | ( n438 & n3940 ) | ( n610 & n3940 ) ;
  assign n10977 = n9573 | n10976 ;
  assign n10980 = n8212 ^ n1373 ^ 1'b0 ;
  assign n10981 = n10980 ^ n5727 ^ 1'b0 ;
  assign n10982 = n10981 ^ n1629 ^ 1'b0 ;
  assign n10983 = n6368 | n10982 ;
  assign n10984 = ( n1988 & n9138 ) | ( n1988 & n10983 ) | ( n9138 & n10983 ) ;
  assign n10985 = n6696 | n10984 ;
  assign n10986 = n10985 ^ n7705 ^ 1'b0 ;
  assign n10978 = n6159 & ~n7630 ;
  assign n10979 = n10978 ^ n5715 ^ 1'b0 ;
  assign n10987 = n10986 ^ n10979 ^ n465 ;
  assign n10988 = n10977 & ~n10987 ;
  assign n10989 = ~n5812 & n5856 ;
  assign n10990 = n10989 ^ n7971 ^ n5346 ;
  assign n10991 = n1042 ^ n1003 ^ 1'b0 ;
  assign n10992 = n8847 ^ n2233 ^ 1'b0 ;
  assign n10993 = n10992 ^ n9599 ^ n9526 ;
  assign n10994 = n10993 ^ n9989 ^ n2993 ;
  assign n10995 = n10991 & ~n10994 ;
  assign n10996 = n775 & n10995 ;
  assign n10998 = x233 & n10636 ;
  assign n10997 = ~n826 & n4204 ;
  assign n10999 = n10998 ^ n10997 ^ 1'b0 ;
  assign n11000 = n8550 ^ n1061 ^ n491 ;
  assign n11001 = n11000 ^ n941 ^ x40 ;
  assign n11002 = n1291 | n9157 ;
  assign n11003 = n11001 & ~n11002 ;
  assign n11004 = n5950 ^ n1566 ^ n1469 ;
  assign n11005 = n9246 ^ n5659 ^ 1'b0 ;
  assign n11006 = n7354 & ~n11005 ;
  assign n11010 = n9365 ^ n2553 ^ 1'b0 ;
  assign n11011 = ~n7477 & n11010 ;
  assign n11007 = n8636 ^ n1434 ^ 1'b0 ;
  assign n11008 = ~n4040 & n11007 ;
  assign n11009 = ( ~n436 & n773 ) | ( ~n436 & n11008 ) | ( n773 & n11008 ) ;
  assign n11012 = n11011 ^ n11009 ^ n4490 ;
  assign n11013 = n11012 ^ n2102 ^ n1224 ;
  assign n11014 = ~n7221 & n8794 ;
  assign n11015 = n11014 ^ n5469 ^ 1'b0 ;
  assign n11016 = ( ~n3199 & n4086 ) | ( ~n3199 & n9586 ) | ( n4086 & n9586 ) ;
  assign n11017 = n8762 & n11016 ;
  assign n11018 = n4972 ^ n1982 ^ n327 ;
  assign n11019 = n7746 | n11018 ;
  assign n11020 = n3661 | n11019 ;
  assign n11021 = n4409 ^ n2373 ^ n1830 ;
  assign n11022 = n5490 ^ n1608 ^ 1'b0 ;
  assign n11023 = n11022 ^ n10770 ^ x80 ;
  assign n11024 = ~n3701 & n11023 ;
  assign n11025 = ( n1700 & n7101 ) | ( n1700 & ~n9617 ) | ( n7101 & ~n9617 ) ;
  assign n11026 = n7799 ^ n2398 ^ n1648 ;
  assign n11027 = n7815 ^ n7069 ^ 1'b0 ;
  assign n11028 = ~n6357 & n11027 ;
  assign n11029 = n11028 ^ n7199 ^ n4326 ;
  assign n11034 = n10021 ^ n859 ^ n378 ;
  assign n11032 = n256 & ~n3203 ;
  assign n11033 = n11032 ^ x130 ^ 1'b0 ;
  assign n11035 = n11034 ^ n11033 ^ n2915 ;
  assign n11030 = n3704 ^ n1206 ^ 1'b0 ;
  assign n11031 = n7370 & ~n11030 ;
  assign n11036 = n11035 ^ n11031 ^ 1'b0 ;
  assign n11037 = ~n3132 & n11036 ;
  assign n11038 = n3452 ^ n2001 ^ x100 ;
  assign n11039 = n2167 & ~n11038 ;
  assign n11040 = n3920 ^ x158 ^ 1'b0 ;
  assign n11041 = n1969 & ~n6897 ;
  assign n11042 = n11041 ^ n7846 ^ 1'b0 ;
  assign n11043 = ~n5082 & n7366 ;
  assign n11044 = n7282 ^ n1862 ^ 1'b0 ;
  assign n11045 = ( n11042 & n11043 ) | ( n11042 & n11044 ) | ( n11043 & n11044 ) ;
  assign n11046 = ( ~n4293 & n6951 ) | ( ~n4293 & n7927 ) | ( n6951 & n7927 ) ;
  assign n11047 = n4650 ^ n2085 ^ 1'b0 ;
  assign n11048 = ~n11046 & n11047 ;
  assign n11049 = n11048 ^ n576 ^ 1'b0 ;
  assign n11050 = n6796 & ~n11049 ;
  assign n11051 = n8071 ^ n7433 ^ n3927 ;
  assign n11052 = n3080 | n11051 ;
  assign n11053 = n11052 ^ n4813 ^ 1'b0 ;
  assign n11054 = n11050 & ~n11053 ;
  assign n11055 = n10127 ^ n3470 ^ n689 ;
  assign n11056 = n11055 ^ n4797 ^ 1'b0 ;
  assign n11057 = n11056 ^ n592 ^ 1'b0 ;
  assign n11058 = n1502 ^ n748 ^ n711 ;
  assign n11059 = ( n4786 & n9265 ) | ( n4786 & n9739 ) | ( n9265 & n9739 ) ;
  assign n11060 = n799 | n9338 ;
  assign n11065 = ( n4305 & ~n6485 ) | ( n4305 & n8718 ) | ( ~n6485 & n8718 ) ;
  assign n11061 = n6227 | n7757 ;
  assign n11062 = n7838 & ~n11061 ;
  assign n11063 = n11062 ^ n1296 ^ 1'b0 ;
  assign n11064 = n9583 & n11063 ;
  assign n11066 = n11065 ^ n11064 ^ 1'b0 ;
  assign n11067 = n11066 ^ n3596 ^ 1'b0 ;
  assign n11068 = ~n11060 & n11067 ;
  assign n11069 = ( n11058 & n11059 ) | ( n11058 & ~n11068 ) | ( n11059 & ~n11068 ) ;
  assign n11073 = ( n2183 & ~n2422 ) | ( n2183 & n5075 ) | ( ~n2422 & n5075 ) ;
  assign n11074 = ( n4463 & n4807 ) | ( n4463 & n11073 ) | ( n4807 & n11073 ) ;
  assign n11070 = ~n598 & n2669 ;
  assign n11071 = ~n1599 & n11070 ;
  assign n11072 = n6208 | n11071 ;
  assign n11075 = n11074 ^ n11072 ^ 1'b0 ;
  assign n11076 = n3221 ^ n2128 ^ n344 ;
  assign n11077 = n7605 ^ n1133 ^ n803 ;
  assign n11078 = n8669 & n11077 ;
  assign n11079 = ( n4630 & n7292 ) | ( n4630 & n11078 ) | ( n7292 & n11078 ) ;
  assign n11080 = ( x29 & ~n11076 ) | ( x29 & n11079 ) | ( ~n11076 & n11079 ) ;
  assign n11083 = n992 ^ x28 ^ 1'b0 ;
  assign n11081 = n5535 | n8566 ;
  assign n11082 = n2143 & ~n11081 ;
  assign n11084 = n11083 ^ n11082 ^ n1879 ;
  assign n11085 = n1558 & n5994 ;
  assign n11086 = n11085 ^ n5946 ^ 1'b0 ;
  assign n11087 = ( ~x111 & n1023 ) | ( ~x111 & n4405 ) | ( n1023 & n4405 ) ;
  assign n11088 = n11087 ^ n3327 ^ n3036 ;
  assign n11089 = n1581 ^ n625 ^ 1'b0 ;
  assign n11090 = n11089 ^ n3507 ^ n1740 ;
  assign n11091 = ( n890 & n11088 ) | ( n890 & ~n11090 ) | ( n11088 & ~n11090 ) ;
  assign n11092 = n11086 | n11091 ;
  assign n11098 = n3105 & n3636 ;
  assign n11099 = n11098 ^ n7820 ^ 1'b0 ;
  assign n11100 = ~n647 & n11099 ;
  assign n11101 = ~n10350 & n11100 ;
  assign n11093 = n5974 ^ n5003 ^ 1'b0 ;
  assign n11094 = n4153 | n11093 ;
  assign n11095 = ( n2001 & n2110 ) | ( n2001 & ~n9541 ) | ( n2110 & ~n9541 ) ;
  assign n11096 = ( ~n1305 & n7221 ) | ( ~n1305 & n11095 ) | ( n7221 & n11095 ) ;
  assign n11097 = n11094 & n11096 ;
  assign n11102 = n11101 ^ n11097 ^ 1'b0 ;
  assign n11103 = n5578 ^ n4812 ^ 1'b0 ;
  assign n11104 = n8525 | n11103 ;
  assign n11108 = n9060 ^ n7300 ^ 1'b0 ;
  assign n11105 = n4180 & ~n10570 ;
  assign n11106 = n2556 | n7333 ;
  assign n11107 = ( n5855 & ~n11105 ) | ( n5855 & n11106 ) | ( ~n11105 & n11106 ) ;
  assign n11109 = n11108 ^ n11107 ^ n8196 ;
  assign n11110 = n2130 ^ n959 ^ 1'b0 ;
  assign n11111 = n2850 & ~n11110 ;
  assign n11112 = n11111 ^ n2627 ^ 1'b0 ;
  assign n11113 = ( ~n1597 & n4499 ) | ( ~n1597 & n11112 ) | ( n4499 & n11112 ) ;
  assign n11114 = n5939 & ~n9174 ;
  assign n11118 = n1724 & ~n8540 ;
  assign n11115 = n4495 ^ n3858 ^ n922 ;
  assign n11116 = ~n3054 & n11115 ;
  assign n11117 = ~n9056 & n11116 ;
  assign n11119 = n11118 ^ n11117 ^ n2759 ;
  assign n11120 = n9677 ^ n3343 ^ x97 ;
  assign n11121 = ( ~n2110 & n8455 ) | ( ~n2110 & n11120 ) | ( n8455 & n11120 ) ;
  assign n11122 = n11121 ^ n3565 ^ 1'b0 ;
  assign n11123 = ( n2886 & n4203 ) | ( n2886 & n4428 ) | ( n4203 & n4428 ) ;
  assign n11124 = ~n11122 & n11123 ;
  assign n11125 = n11124 ^ n6630 ^ n909 ;
  assign n11126 = n6712 ^ n2707 ^ 1'b0 ;
  assign n11127 = n10210 & n11126 ;
  assign n11128 = n10518 ^ n10106 ^ n4450 ;
  assign n11129 = n3837 & ~n8649 ;
  assign n11130 = n9385 & ~n11129 ;
  assign n11131 = n9161 & ~n11130 ;
  assign n11132 = n11131 ^ x201 ^ 1'b0 ;
  assign n11133 = ~n7415 & n8072 ;
  assign n11134 = n11133 ^ n9694 ^ 1'b0 ;
  assign n11135 = ~n437 & n4833 ;
  assign n11136 = ~n6468 & n11135 ;
  assign n11146 = n10438 ^ n8806 ^ n6962 ;
  assign n11147 = ( n1810 & ~n2667 ) | ( n1810 & n2701 ) | ( ~n2667 & n2701 ) ;
  assign n11148 = ~n11146 & n11147 ;
  assign n11149 = ~n3967 & n11148 ;
  assign n11137 = n8726 & n11008 ;
  assign n11138 = ( x59 & ~n5363 ) | ( x59 & n11137 ) | ( ~n5363 & n11137 ) ;
  assign n11139 = ( ~n4479 & n5622 ) | ( ~n4479 & n11138 ) | ( n5622 & n11138 ) ;
  assign n11140 = ~n4338 & n8903 ;
  assign n11141 = n11140 ^ n1153 ^ 1'b0 ;
  assign n11142 = n2030 | n7503 ;
  assign n11143 = n11141 & ~n11142 ;
  assign n11144 = n11139 | n11143 ;
  assign n11145 = n11144 ^ n8239 ^ 1'b0 ;
  assign n11150 = n11149 ^ n11145 ^ n7685 ;
  assign n11153 = ( n2089 & n2875 ) | ( n2089 & n5017 ) | ( n2875 & n5017 ) ;
  assign n11151 = ~n4315 & n5119 ;
  assign n11152 = ( n3582 & n4448 ) | ( n3582 & n11151 ) | ( n4448 & n11151 ) ;
  assign n11154 = n11153 ^ n11152 ^ n3236 ;
  assign n11155 = n4055 ^ n3886 ^ 1'b0 ;
  assign n11156 = n11155 ^ n5685 ^ 1'b0 ;
  assign n11157 = n1478 & ~n11156 ;
  assign n11158 = n2776 | n3046 ;
  assign n11159 = n11157 & ~n11158 ;
  assign n11160 = ~n9497 & n11159 ;
  assign n11161 = ( n5779 & n8121 ) | ( n5779 & ~n11160 ) | ( n8121 & ~n11160 ) ;
  assign n11162 = n3202 & n11161 ;
  assign n11163 = n282 & ~n4943 ;
  assign n11164 = n4001 & n11163 ;
  assign n11166 = n6615 ^ n6235 ^ 1'b0 ;
  assign n11165 = n5066 | n11143 ;
  assign n11167 = n11166 ^ n11165 ^ 1'b0 ;
  assign n11168 = ( n1486 & ~n5182 ) | ( n1486 & n10819 ) | ( ~n5182 & n10819 ) ;
  assign n11169 = n11168 ^ n2698 ^ 1'b0 ;
  assign n11170 = ~n11167 & n11169 ;
  assign n11171 = n4524 ^ n3202 ^ n3036 ;
  assign n11172 = n1472 | n11171 ;
  assign n11173 = ( n7218 & n11170 ) | ( n7218 & ~n11172 ) | ( n11170 & ~n11172 ) ;
  assign n11174 = ( ~n873 & n9437 ) | ( ~n873 & n11173 ) | ( n9437 & n11173 ) ;
  assign n11175 = ( n2686 & n4324 ) | ( n2686 & n7470 ) | ( n4324 & n7470 ) ;
  assign n11176 = n394 & ~n11175 ;
  assign n11177 = n9094 & n11176 ;
  assign n11178 = n6351 ^ n4874 ^ n4499 ;
  assign n11179 = ( n1145 & n3879 ) | ( n1145 & n11178 ) | ( n3879 & n11178 ) ;
  assign n11180 = ( ~n4000 & n10222 ) | ( ~n4000 & n11179 ) | ( n10222 & n11179 ) ;
  assign n11181 = n2794 ^ n828 ^ 1'b0 ;
  assign n11182 = n8810 | n11181 ;
  assign n11183 = n2515 & ~n11182 ;
  assign n11184 = n11180 | n11183 ;
  assign n11185 = n11184 ^ n2899 ^ 1'b0 ;
  assign n11186 = n11185 ^ n8378 ^ n4593 ;
  assign n11190 = ~n1052 & n1733 ;
  assign n11187 = n963 & n4164 ;
  assign n11188 = n11187 ^ n1621 ^ 1'b0 ;
  assign n11189 = n11188 ^ n4707 ^ n2858 ;
  assign n11191 = n11190 ^ n11189 ^ 1'b0 ;
  assign n11192 = ~n2127 & n11191 ;
  assign n11196 = x206 & ~n8442 ;
  assign n11193 = n9214 ^ n6677 ^ n3798 ;
  assign n11194 = n4876 | n5520 ;
  assign n11195 = n11193 | n11194 ;
  assign n11197 = n11196 ^ n11195 ^ 1'b0 ;
  assign n11198 = ( n6347 & ~n7125 ) | ( n6347 & n11197 ) | ( ~n7125 & n11197 ) ;
  assign n11199 = ~n2500 & n11198 ;
  assign n11200 = n11199 ^ n7905 ^ 1'b0 ;
  assign n11201 = n7077 ^ n6074 ^ n3382 ;
  assign n11202 = n2863 & ~n3236 ;
  assign n11203 = n11202 ^ n2596 ^ 1'b0 ;
  assign n11205 = n9135 ^ n2393 ^ n2051 ;
  assign n11204 = n10880 ^ n1000 ^ 1'b0 ;
  assign n11206 = n11205 ^ n11204 ^ n7551 ;
  assign n11207 = n9639 ^ n4045 ^ 1'b0 ;
  assign n11208 = ( n1028 & n11206 ) | ( n1028 & n11207 ) | ( n11206 & n11207 ) ;
  assign n11209 = n10152 ^ n4828 ^ n1473 ;
  assign n11210 = n11209 ^ n1910 ^ n1837 ;
  assign n11211 = n4848 ^ x115 ^ 1'b0 ;
  assign n11212 = n3256 | n11211 ;
  assign n11213 = n6611 ^ n5814 ^ n971 ;
  assign n11214 = n11212 | n11213 ;
  assign n11215 = n9017 & ~n11214 ;
  assign n11216 = ( ~x81 & n3042 ) | ( ~x81 & n4820 ) | ( n3042 & n4820 ) ;
  assign n11221 = n4124 ^ n3923 ^ 1'b0 ;
  assign n11220 = n7806 ^ n7579 ^ n4627 ;
  assign n11217 = ( n3162 & n3923 ) | ( n3162 & ~n9928 ) | ( n3923 & ~n9928 ) ;
  assign n11218 = n11217 ^ n4387 ^ n3047 ;
  assign n11219 = n11218 ^ n5783 ^ 1'b0 ;
  assign n11222 = n11221 ^ n11220 ^ n11219 ;
  assign n11223 = n11222 ^ n10063 ^ n8790 ;
  assign n11224 = ~n5279 & n11223 ;
  assign n11225 = ~n11216 & n11224 ;
  assign n11226 = ( n2587 & n3065 ) | ( n2587 & n4575 ) | ( n3065 & n4575 ) ;
  assign n11227 = ( n3052 & n4638 ) | ( n3052 & n11226 ) | ( n4638 & n11226 ) ;
  assign n11228 = n9643 ^ n8002 ^ 1'b0 ;
  assign n11229 = ~n2773 & n11228 ;
  assign n11230 = n4929 & n11229 ;
  assign n11231 = n11230 ^ n5779 ^ 1'b0 ;
  assign n11232 = n11227 & ~n11231 ;
  assign n11233 = n9697 ^ n353 ^ 1'b0 ;
  assign n11234 = ~n2002 & n11233 ;
  assign n11235 = n4630 ^ n1257 ^ 1'b0 ;
  assign n11236 = ~n6583 & n11235 ;
  assign n11237 = ( n6932 & n8996 ) | ( n6932 & ~n11236 ) | ( n8996 & ~n11236 ) ;
  assign n11238 = ( x99 & n11234 ) | ( x99 & ~n11237 ) | ( n11234 & ~n11237 ) ;
  assign n11239 = ( n7729 & n11232 ) | ( n7729 & ~n11238 ) | ( n11232 & ~n11238 ) ;
  assign n11240 = n1849 & ~n4883 ;
  assign n11241 = ( n3002 & ~n4317 ) | ( n3002 & n10003 ) | ( ~n4317 & n10003 ) ;
  assign n11242 = n11241 ^ n10288 ^ n4797 ;
  assign n11243 = ( ~n6349 & n7710 ) | ( ~n6349 & n11242 ) | ( n7710 & n11242 ) ;
  assign n11244 = n11243 ^ n2948 ^ 1'b0 ;
  assign n11245 = n11244 ^ n3661 ^ n1179 ;
  assign n11246 = ( n5075 & ~n11240 ) | ( n5075 & n11245 ) | ( ~n11240 & n11245 ) ;
  assign n11247 = ( n6241 & ~n10113 ) | ( n6241 & n11246 ) | ( ~n10113 & n11246 ) ;
  assign n11248 = n1797 & ~n8804 ;
  assign n11249 = ( n1981 & ~n2163 ) | ( n1981 & n5245 ) | ( ~n2163 & n5245 ) ;
  assign n11250 = ( n1370 & n9357 ) | ( n1370 & ~n11249 ) | ( n9357 & ~n11249 ) ;
  assign n11251 = n4772 ^ n3453 ^ 1'b0 ;
  assign n11252 = ( n4752 & n6500 ) | ( n4752 & ~n11251 ) | ( n6500 & ~n11251 ) ;
  assign n11253 = n3747 | n11252 ;
  assign n11254 = ( n7213 & n7234 ) | ( n7213 & ~n11253 ) | ( n7234 & ~n11253 ) ;
  assign n11255 = ( n3013 & n3459 ) | ( n3013 & ~n6497 ) | ( n3459 & ~n6497 ) ;
  assign n11256 = n11255 ^ n2906 ^ 1'b0 ;
  assign n11257 = n10067 ^ n4834 ^ n1825 ;
  assign n11258 = ( n4000 & ~n4634 ) | ( n4000 & n11257 ) | ( ~n4634 & n11257 ) ;
  assign n11259 = n11258 ^ n5845 ^ n1610 ;
  assign n11260 = n1822 & n11259 ;
  assign n11261 = ~n7278 & n11260 ;
  assign n11262 = n11261 ^ n7033 ^ 1'b0 ;
  assign n11263 = n8821 & n11262 ;
  assign n11264 = n11263 ^ n4745 ^ 1'b0 ;
  assign n11265 = n3747 | n11264 ;
  assign n11266 = n10821 ^ n5880 ^ n3955 ;
  assign n11267 = n11266 ^ x60 ^ 1'b0 ;
  assign n11268 = n9317 & n11267 ;
  assign n11269 = n6357 ^ n2543 ^ 1'b0 ;
  assign n11270 = n11269 ^ n6668 ^ n3324 ;
  assign n11271 = n4067 | n5097 ;
  assign n11272 = n3171 & n11271 ;
  assign n11273 = n11272 ^ n4764 ^ 1'b0 ;
  assign n11274 = ( n6266 & n9766 ) | ( n6266 & n11273 ) | ( n9766 & n11273 ) ;
  assign n11275 = ( n2677 & ~n2799 ) | ( n2677 & n6847 ) | ( ~n2799 & n6847 ) ;
  assign n11276 = n10772 | n11275 ;
  assign n11277 = ( n950 & n8754 ) | ( n950 & n11276 ) | ( n8754 & n11276 ) ;
  assign n11278 = n10951 & n11277 ;
  assign n11279 = n2676 & ~n11278 ;
  assign n11280 = n11279 ^ n7908 ^ 1'b0 ;
  assign n11288 = n5393 ^ n1081 ^ 1'b0 ;
  assign n11282 = n5260 & n8985 ;
  assign n11281 = n674 & ~n5467 ;
  assign n11283 = n11282 ^ n11281 ^ 1'b0 ;
  assign n11284 = x30 & n4194 ;
  assign n11285 = n11283 & n11284 ;
  assign n11286 = n11285 ^ n11000 ^ n5526 ;
  assign n11287 = n11286 ^ n4774 ^ 1'b0 ;
  assign n11289 = n11288 ^ n11287 ^ n3430 ;
  assign n11290 = n9599 ^ n8538 ^ n4660 ;
  assign n11291 = x163 | n4645 ;
  assign n11292 = n10206 ^ x253 ^ 1'b0 ;
  assign n11293 = ~n9404 & n11292 ;
  assign n11294 = ~n11291 & n11293 ;
  assign n11295 = x212 & n8614 ;
  assign n11296 = n11294 & n11295 ;
  assign n11297 = ~n1366 & n1824 ;
  assign n11298 = n11297 ^ n10159 ^ n570 ;
  assign n11299 = ~n6291 & n11298 ;
  assign n11302 = n2352 & ~n5649 ;
  assign n11303 = n11302 ^ n291 ^ 1'b0 ;
  assign n11300 = n2759 ^ n1131 ^ 1'b0 ;
  assign n11301 = ~n2034 & n11300 ;
  assign n11304 = n11303 ^ n11301 ^ n7397 ;
  assign n11305 = n10256 ^ n6387 ^ 1'b0 ;
  assign n11306 = ( n3821 & n6353 ) | ( n3821 & ~n11305 ) | ( n6353 & ~n11305 ) ;
  assign n11307 = ~n2907 & n4027 ;
  assign n11308 = n11307 ^ n9454 ^ 1'b0 ;
  assign n11309 = n4058 & ~n11308 ;
  assign n11310 = n11309 ^ n4057 ^ 1'b0 ;
  assign n11311 = ( ~n3054 & n3878 ) | ( ~n3054 & n7478 ) | ( n3878 & n7478 ) ;
  assign n11312 = n7501 ^ n5523 ^ 1'b0 ;
  assign n11313 = n11312 ^ n1404 ^ 1'b0 ;
  assign n11314 = ( ~n11310 & n11311 ) | ( ~n11310 & n11313 ) | ( n11311 & n11313 ) ;
  assign n11315 = n5277 ^ n2198 ^ 1'b0 ;
  assign n11316 = n5574 & ~n11315 ;
  assign n11317 = n5321 & ~n7440 ;
  assign n11318 = ~n11316 & n11317 ;
  assign n11319 = ( ~n6151 & n10261 ) | ( ~n6151 & n11318 ) | ( n10261 & n11318 ) ;
  assign n11320 = n10201 ^ n7013 ^ n6423 ;
  assign n11321 = n10300 & n11320 ;
  assign n11324 = n3355 & n4297 ;
  assign n11322 = n8128 ^ n459 ^ x63 ;
  assign n11323 = n6507 | n11322 ;
  assign n11325 = n11324 ^ n11323 ^ 1'b0 ;
  assign n11326 = n9596 ^ n5463 ^ n4470 ;
  assign n11327 = n9965 ^ x96 ^ 1'b0 ;
  assign n11328 = ~n6023 & n9606 ;
  assign n11329 = n11328 ^ n3495 ^ n513 ;
  assign n11330 = n1303 & n3329 ;
  assign n11331 = ~n10582 & n11330 ;
  assign n11332 = ( n6203 & ~n11329 ) | ( n6203 & n11331 ) | ( ~n11329 & n11331 ) ;
  assign n11333 = n6555 & n11332 ;
  assign n11334 = n11333 ^ n4184 ^ 1'b0 ;
  assign n11335 = ( x154 & n6174 ) | ( x154 & n8026 ) | ( n6174 & n8026 ) ;
  assign n11336 = ( n3851 & n4054 ) | ( n3851 & ~n11335 ) | ( n4054 & ~n11335 ) ;
  assign n11337 = n6941 ^ n2506 ^ 1'b0 ;
  assign n11338 = n10602 & ~n11337 ;
  assign n11339 = ~n1877 & n6329 ;
  assign n11340 = n1512 ^ n513 ^ 1'b0 ;
  assign n11341 = ~n11339 & n11340 ;
  assign n11342 = ~n4864 & n11341 ;
  assign n11343 = n10852 & n11342 ;
  assign n11344 = n11343 ^ n10607 ^ n7430 ;
  assign n11345 = n7782 | n11344 ;
  assign n11346 = n2765 | n11345 ;
  assign n11347 = n8162 ^ n2984 ^ 1'b0 ;
  assign n11348 = n1152 & n7907 ;
  assign n11349 = n2464 & n11348 ;
  assign n11350 = ( n564 & ~n7511 ) | ( n564 & n11349 ) | ( ~n7511 & n11349 ) ;
  assign n11351 = ( n3575 & n6536 ) | ( n3575 & n9517 ) | ( n6536 & n9517 ) ;
  assign n11352 = ( ~n594 & n2015 ) | ( ~n594 & n10604 ) | ( n2015 & n10604 ) ;
  assign n11366 = n8478 ^ n6659 ^ n5198 ;
  assign n11353 = n3962 & n5147 ;
  assign n11354 = n1832 ^ n1611 ^ 1'b0 ;
  assign n11355 = ~n6183 & n11354 ;
  assign n11356 = n11355 ^ n3863 ^ 1'b0 ;
  assign n11357 = n412 & n11356 ;
  assign n11358 = n11357 ^ n7217 ^ 1'b0 ;
  assign n11359 = n10293 & ~n11358 ;
  assign n11360 = n5494 & ~n7253 ;
  assign n11361 = n7436 & ~n11360 ;
  assign n11362 = n11361 ^ n6267 ^ 1'b0 ;
  assign n11363 = ~n11359 & n11362 ;
  assign n11364 = ( ~n3320 & n10905 ) | ( ~n3320 & n11363 ) | ( n10905 & n11363 ) ;
  assign n11365 = ~n11353 & n11364 ;
  assign n11367 = n11366 ^ n11365 ^ 1'b0 ;
  assign n11369 = n2146 | n2986 ;
  assign n11370 = n1708 & ~n11369 ;
  assign n11368 = n10319 ^ n2726 ^ n528 ;
  assign n11371 = n11370 ^ n11368 ^ 1'b0 ;
  assign n11372 = n940 & n11201 ;
  assign n11373 = n3518 ^ n865 ^ 1'b0 ;
  assign n11377 = n2061 | n2340 ;
  assign n11378 = n11377 ^ n1761 ^ 1'b0 ;
  assign n11379 = n11378 ^ n10432 ^ n1776 ;
  assign n11374 = n2676 | n4646 ;
  assign n11375 = ( n301 & ~n477 ) | ( n301 & n6860 ) | ( ~n477 & n6860 ) ;
  assign n11376 = ( ~n1229 & n11374 ) | ( ~n1229 & n11375 ) | ( n11374 & n11375 ) ;
  assign n11380 = n11379 ^ n11376 ^ 1'b0 ;
  assign n11381 = n5533 ^ n4925 ^ 1'b0 ;
  assign n11382 = n11381 ^ n9418 ^ x37 ;
  assign n11383 = n5172 & n6648 ;
  assign n11384 = ( x178 & n4070 ) | ( x178 & n11383 ) | ( n4070 & n11383 ) ;
  assign n11389 = ( n1908 & n2641 ) | ( n1908 & ~n4338 ) | ( n2641 & ~n4338 ) ;
  assign n11387 = ( ~n959 & n7316 ) | ( ~n959 & n9118 ) | ( n7316 & n9118 ) ;
  assign n11385 = n10446 ^ n6088 ^ 1'b0 ;
  assign n11386 = ~n10019 & n11385 ;
  assign n11388 = n11387 ^ n11386 ^ n4613 ;
  assign n11390 = n11389 ^ n11388 ^ n9513 ;
  assign n11391 = n2837 ^ n2402 ^ 1'b0 ;
  assign n11392 = x6 & ~n11391 ;
  assign n11393 = n2045 & ~n11392 ;
  assign n11394 = n7792 ^ n5101 ^ 1'b0 ;
  assign n11395 = n11393 & ~n11394 ;
  assign n11396 = n506 & n3105 ;
  assign n11397 = n11396 ^ n3107 ^ 1'b0 ;
  assign n11398 = n1023 | n11397 ;
  assign n11399 = n7072 & ~n11398 ;
  assign n11400 = ( ~n5884 & n10821 ) | ( ~n5884 & n11399 ) | ( n10821 & n11399 ) ;
  assign n11401 = n2429 ^ n1081 ^ 1'b0 ;
  assign n11402 = ~n2826 & n11401 ;
  assign n11403 = n11402 ^ n1802 ^ 1'b0 ;
  assign n11404 = n11400 | n11403 ;
  assign n11409 = ~n2010 & n3401 ;
  assign n11410 = n11409 ^ n5509 ^ 1'b0 ;
  assign n11405 = n6249 ^ n1746 ^ 1'b0 ;
  assign n11406 = ~n6074 & n11405 ;
  assign n11407 = n11406 ^ n5619 ^ 1'b0 ;
  assign n11408 = n11407 ^ n1387 ^ 1'b0 ;
  assign n11411 = n11410 ^ n11408 ^ 1'b0 ;
  assign n11413 = ( n1359 & ~n5010 ) | ( n1359 & n5549 ) | ( ~n5010 & n5549 ) ;
  assign n11412 = n3450 | n9189 ;
  assign n11414 = n11413 ^ n11412 ^ 1'b0 ;
  assign n11415 = n3953 & ~n11414 ;
  assign n11419 = ( ~n2426 & n2498 ) | ( ~n2426 & n5229 ) | ( n2498 & n5229 ) ;
  assign n11418 = n9033 | n10075 ;
  assign n11420 = n11419 ^ n11418 ^ 1'b0 ;
  assign n11416 = n9921 ^ n2325 ^ x58 ;
  assign n11417 = n11416 ^ n10438 ^ 1'b0 ;
  assign n11421 = n11420 ^ n11417 ^ n6831 ;
  assign n11422 = n11363 ^ n10315 ^ n3897 ;
  assign n11423 = n9223 ^ n6495 ^ n3982 ;
  assign n11424 = n7280 ^ n5562 ^ n4259 ;
  assign n11425 = ( n999 & ~n1056 ) | ( n999 & n4316 ) | ( ~n1056 & n4316 ) ;
  assign n11426 = n3725 & n11425 ;
  assign n11427 = n11426 ^ n11288 ^ n2471 ;
  assign n11428 = n6310 ^ n3880 ^ 1'b0 ;
  assign n11429 = n1699 | n7525 ;
  assign n11430 = ~n4771 & n7725 ;
  assign n11431 = n11430 ^ n4519 ^ 1'b0 ;
  assign n11432 = n9102 ^ n2036 ^ 1'b0 ;
  assign n11433 = ~n8896 & n11432 ;
  assign n11434 = n11433 ^ n697 ^ 1'b0 ;
  assign n11435 = ( n2832 & ~n4723 ) | ( n2832 & n6330 ) | ( ~n4723 & n6330 ) ;
  assign n11436 = ( n1286 & n5081 ) | ( n1286 & n11435 ) | ( n5081 & n11435 ) ;
  assign n11437 = ~n1474 & n11436 ;
  assign n11438 = n7862 & n11437 ;
  assign n11439 = n11438 ^ n10457 ^ n9406 ;
  assign n11440 = n7395 ^ n6235 ^ n5782 ;
  assign n11441 = n1768 | n11440 ;
  assign n11442 = n11257 ^ n3490 ^ 1'b0 ;
  assign n11443 = n4421 & n11442 ;
  assign n11444 = ~n3029 & n11443 ;
  assign n11445 = ~n11216 & n11444 ;
  assign n11446 = n2218 | n6111 ;
  assign n11447 = n504 | n9363 ;
  assign n11448 = n11446 | n11447 ;
  assign n11449 = n2313 & n8606 ;
  assign n11450 = ~n5666 & n11449 ;
  assign n11451 = n11450 ^ n5129 ^ 1'b0 ;
  assign n11456 = n3643 | n9012 ;
  assign n11457 = ~n4546 & n11456 ;
  assign n11458 = n11457 ^ n1183 ^ 1'b0 ;
  assign n11459 = n11458 ^ n5727 ^ x230 ;
  assign n11452 = n3545 ^ n1199 ^ 1'b0 ;
  assign n11453 = n8429 ^ n6434 ^ 1'b0 ;
  assign n11454 = n4778 & ~n11453 ;
  assign n11455 = ( ~n3799 & n11452 ) | ( ~n3799 & n11454 ) | ( n11452 & n11454 ) ;
  assign n11460 = n11459 ^ n11455 ^ n1160 ;
  assign n11461 = ( n2142 & n3259 ) | ( n2142 & n4985 ) | ( n3259 & n4985 ) ;
  assign n11462 = n11461 ^ n6188 ^ 1'b0 ;
  assign n11463 = n11460 & n11462 ;
  assign n11464 = n7908 ^ n1637 ^ 1'b0 ;
  assign n11465 = n11463 & ~n11464 ;
  assign n11466 = ( ~n3480 & n4883 ) | ( ~n3480 & n9506 ) | ( n4883 & n9506 ) ;
  assign n11467 = n9469 ^ n890 ^ 1'b0 ;
  assign n11468 = ( ~n787 & n11466 ) | ( ~n787 & n11467 ) | ( n11466 & n11467 ) ;
  assign n11470 = ( n1319 & ~n1567 ) | ( n1319 & n8026 ) | ( ~n1567 & n8026 ) ;
  assign n11471 = ~n2059 & n11470 ;
  assign n11472 = n6655 & n11471 ;
  assign n11469 = ~n1676 & n9399 ;
  assign n11473 = n11472 ^ n11469 ^ 1'b0 ;
  assign n11474 = n11473 ^ n10895 ^ 1'b0 ;
  assign n11475 = n6980 & n10071 ;
  assign n11476 = n6123 & n11475 ;
  assign n11477 = n7501 ^ n2871 ^ n1322 ;
  assign n11478 = ( ~x227 & n7356 ) | ( ~x227 & n10192 ) | ( n7356 & n10192 ) ;
  assign n11479 = n11477 | n11478 ;
  assign n11480 = n8742 ^ n620 ^ n416 ;
  assign n11481 = n5408 & ~n11480 ;
  assign n11482 = n11481 ^ n1588 ^ 1'b0 ;
  assign n11483 = n5320 | n8557 ;
  assign n11484 = n11483 ^ n8191 ^ 1'b0 ;
  assign n11485 = n11484 ^ n9493 ^ n589 ;
  assign n11486 = n11485 ^ n1079 ^ 1'b0 ;
  assign n11487 = n11482 & ~n11486 ;
  assign n11488 = n4659 | n6879 ;
  assign n11491 = n5745 ^ n2677 ^ 1'b0 ;
  assign n11492 = n1374 & n11491 ;
  assign n11489 = n2896 & n3307 ;
  assign n11490 = ( n5158 & ~n11466 ) | ( n5158 & n11489 ) | ( ~n11466 & n11489 ) ;
  assign n11493 = n11492 ^ n11490 ^ n6368 ;
  assign n11494 = n10541 & ~n11493 ;
  assign n11495 = n11494 ^ n501 ^ 1'b0 ;
  assign n11496 = ~n5715 & n8059 ;
  assign n11497 = n2867 | n4294 ;
  assign n11498 = n6432 ^ n2342 ^ 1'b0 ;
  assign n11499 = n11497 | n11498 ;
  assign n11500 = n11499 ^ n11250 ^ n6057 ;
  assign n11511 = n3470 & n5730 ;
  assign n11512 = n11511 ^ n10083 ^ 1'b0 ;
  assign n11506 = n2222 | n3159 ;
  assign n11507 = n1140 & ~n2737 ;
  assign n11508 = ( n1791 & ~n11506 ) | ( n1791 & n11507 ) | ( ~n11506 & n11507 ) ;
  assign n11509 = ~n5048 & n11508 ;
  assign n11510 = ( ~n6709 & n10501 ) | ( ~n6709 & n11509 ) | ( n10501 & n11509 ) ;
  assign n11502 = ~n3851 & n9451 ;
  assign n11503 = n11502 ^ n8785 ^ 1'b0 ;
  assign n11504 = n11503 ^ n10664 ^ n3440 ;
  assign n11501 = n7973 | n11012 ;
  assign n11505 = n11504 ^ n11501 ^ 1'b0 ;
  assign n11513 = n11512 ^ n11510 ^ n11505 ;
  assign n11514 = n1813 & ~n4283 ;
  assign n11515 = n11514 ^ n2293 ^ 1'b0 ;
  assign n11516 = ~n1993 & n9641 ;
  assign n11517 = n1675 ^ x2 ^ 1'b0 ;
  assign n11518 = ( n6257 & n11516 ) | ( n6257 & ~n11517 ) | ( n11516 & ~n11517 ) ;
  assign n11527 = ( n6148 & ~n7704 ) | ( n6148 & n8544 ) | ( ~n7704 & n8544 ) ;
  assign n11522 = ~n604 & n6255 ;
  assign n11523 = n11522 ^ n5544 ^ 1'b0 ;
  assign n11524 = n11523 ^ n3325 ^ n1709 ;
  assign n11525 = n11524 ^ n3134 ^ x181 ;
  assign n11519 = n2367 & ~n3290 ;
  assign n11520 = n11519 ^ n7385 ^ 1'b0 ;
  assign n11521 = n807 | n11520 ;
  assign n11526 = n11525 ^ n11521 ^ 1'b0 ;
  assign n11528 = n11527 ^ n11526 ^ n7535 ;
  assign n11529 = n2539 ^ n1915 ^ 1'b0 ;
  assign n11530 = ( n2095 & ~n10702 ) | ( n2095 & n11529 ) | ( ~n10702 & n11529 ) ;
  assign n11531 = n2736 ^ x188 ^ 1'b0 ;
  assign n11532 = ~n975 & n11531 ;
  assign n11533 = n11532 ^ n1694 ^ n310 ;
  assign n11534 = ~n11530 & n11533 ;
  assign n11535 = n9005 ^ n4348 ^ 1'b0 ;
  assign n11536 = n4941 & ~n11535 ;
  assign n11537 = ( n4089 & n6916 ) | ( n4089 & n11536 ) | ( n6916 & n11536 ) ;
  assign n11538 = ( n450 & n2619 ) | ( n450 & n4516 ) | ( n2619 & n4516 ) ;
  assign n11539 = n4526 ^ n1595 ^ 1'b0 ;
  assign n11540 = n4370 & ~n11539 ;
  assign n11541 = ( n3004 & n10673 ) | ( n3004 & n11540 ) | ( n10673 & n11540 ) ;
  assign n11542 = ( ~n1129 & n11538 ) | ( ~n1129 & n11541 ) | ( n11538 & n11541 ) ;
  assign n11543 = n11542 ^ n4320 ^ n4085 ;
  assign n11544 = n3636 | n10570 ;
  assign n11545 = n11544 ^ n2851 ^ 1'b0 ;
  assign n11546 = n11545 ^ n10850 ^ n419 ;
  assign n11547 = n5365 ^ n1793 ^ 1'b0 ;
  assign n11548 = n10991 & n11547 ;
  assign n11549 = n7662 ^ n1710 ^ 1'b0 ;
  assign n11550 = x240 & n11549 ;
  assign n11551 = n11550 ^ n6173 ^ 1'b0 ;
  assign n11552 = n7631 & ~n11551 ;
  assign n11553 = n1084 & ~n11042 ;
  assign n11554 = n6046 ^ n5707 ^ 1'b0 ;
  assign n11555 = n10021 & n11554 ;
  assign n11556 = n6368 ^ n487 ^ 1'b0 ;
  assign n11557 = n10887 ^ n9884 ^ 1'b0 ;
  assign n11558 = n11556 & ~n11557 ;
  assign n11559 = n11129 ^ n10571 ^ n5238 ;
  assign n11560 = n3790 & n5301 ;
  assign n11561 = x215 & ~n11560 ;
  assign n11562 = ~n11559 & n11561 ;
  assign n11563 = n5227 & ~n11562 ;
  assign n11564 = n5386 & n11563 ;
  assign n11565 = n5972 ^ n2706 ^ 1'b0 ;
  assign n11566 = n8555 & n11565 ;
  assign n11569 = n3577 | n5182 ;
  assign n11570 = n2348 & ~n11569 ;
  assign n11571 = n4681 | n11570 ;
  assign n11572 = x171 | n11571 ;
  assign n11567 = n1890 ^ n1403 ^ 1'b0 ;
  assign n11568 = n4522 & ~n11567 ;
  assign n11573 = n11572 ^ n11568 ^ 1'b0 ;
  assign n11576 = n324 & n9972 ;
  assign n11577 = n11576 ^ n4754 ^ 1'b0 ;
  assign n11578 = n6307 & n11577 ;
  assign n11579 = ( ~n1690 & n9946 ) | ( ~n1690 & n11578 ) | ( n9946 & n11578 ) ;
  assign n11574 = n5707 ^ n2349 ^ 1'b0 ;
  assign n11575 = ~n327 & n11574 ;
  assign n11580 = n11579 ^ n11575 ^ 1'b0 ;
  assign n11581 = x53 & n8499 ;
  assign n11582 = n11581 ^ n707 ^ 1'b0 ;
  assign n11583 = ( n1416 & n4051 ) | ( n1416 & n10694 ) | ( n4051 & n10694 ) ;
  assign n11584 = n9433 ^ n7901 ^ n4359 ;
  assign n11585 = n3670 & ~n11584 ;
  assign n11587 = x172 & n2074 ;
  assign n11588 = n11587 ^ n5036 ^ 1'b0 ;
  assign n11589 = ( n776 & ~n1722 ) | ( n776 & n1843 ) | ( ~n1722 & n1843 ) ;
  assign n11590 = ( n4307 & n5830 ) | ( n4307 & ~n11589 ) | ( n5830 & ~n11589 ) ;
  assign n11591 = ~n11588 & n11590 ;
  assign n11592 = n11591 ^ n3770 ^ 1'b0 ;
  assign n11593 = ( n563 & n752 ) | ( n563 & ~n4018 ) | ( n752 & ~n4018 ) ;
  assign n11594 = n11593 ^ n1311 ^ n953 ;
  assign n11595 = ( ~n1072 & n6859 ) | ( ~n1072 & n7117 ) | ( n6859 & n7117 ) ;
  assign n11596 = ~n11594 & n11595 ;
  assign n11597 = ~n5075 & n11596 ;
  assign n11598 = ( ~n1054 & n11592 ) | ( ~n1054 & n11597 ) | ( n11592 & n11597 ) ;
  assign n11586 = n4562 | n4871 ;
  assign n11599 = n11598 ^ n11586 ^ 1'b0 ;
  assign n11600 = n4139 ^ n1834 ^ 1'b0 ;
  assign n11601 = n11600 ^ n1733 ^ 1'b0 ;
  assign n11602 = x23 & n10677 ;
  assign n11603 = n461 & n11602 ;
  assign n11604 = n11538 ^ n7766 ^ n3055 ;
  assign n11605 = ( n408 & n1054 ) | ( n408 & n2309 ) | ( n1054 & n2309 ) ;
  assign n11606 = ( n1881 & n7965 ) | ( n1881 & ~n11605 ) | ( n7965 & ~n11605 ) ;
  assign n11607 = ( n4839 & n11604 ) | ( n4839 & n11606 ) | ( n11604 & n11606 ) ;
  assign n11608 = n11607 ^ n6241 ^ n2917 ;
  assign n11609 = n11608 ^ n9310 ^ n4103 ;
  assign n11610 = ~n11603 & n11609 ;
  assign n11611 = n11601 & n11610 ;
  assign n11612 = n10376 ^ n4584 ^ 1'b0 ;
  assign n11613 = n5617 & n11612 ;
  assign n11614 = n10483 ^ n5688 ^ n4313 ;
  assign n11617 = ( ~n1439 & n6065 ) | ( ~n1439 & n10709 ) | ( n6065 & n10709 ) ;
  assign n11616 = ( n1521 & n1598 ) | ( n1521 & n4595 ) | ( n1598 & n4595 ) ;
  assign n11618 = n11617 ^ n11616 ^ n5197 ;
  assign n11619 = n11618 ^ n10736 ^ n1965 ;
  assign n11615 = n8446 ^ n1136 ^ 1'b0 ;
  assign n11620 = n11619 ^ n11615 ^ n8326 ;
  assign n11621 = n2596 ^ n1891 ^ 1'b0 ;
  assign n11622 = n4746 & ~n11621 ;
  assign n11623 = n5432 ^ x63 ^ 1'b0 ;
  assign n11624 = n11622 & ~n11623 ;
  assign n11625 = n6237 ^ n1618 ^ 1'b0 ;
  assign n11632 = n8770 ^ n6634 ^ n2052 ;
  assign n11628 = ( x153 & n1328 ) | ( x153 & n1777 ) | ( n1328 & n1777 ) ;
  assign n11629 = n2924 | n11628 ;
  assign n11626 = ~n2039 & n2280 ;
  assign n11627 = n11626 ^ n9314 ^ 1'b0 ;
  assign n11630 = n11629 ^ n11627 ^ n4034 ;
  assign n11631 = ( n6476 & n11432 ) | ( n6476 & n11630 ) | ( n11432 & n11630 ) ;
  assign n11633 = n11632 ^ n11631 ^ x8 ;
  assign n11634 = n4881 ^ n2386 ^ n1469 ;
  assign n11635 = n11634 ^ n2978 ^ n394 ;
  assign n11636 = n11635 ^ n5225 ^ n4022 ;
  assign n11637 = ( x206 & n4571 ) | ( x206 & ~n6637 ) | ( n4571 & ~n6637 ) ;
  assign n11638 = n10935 ^ n2302 ^ n613 ;
  assign n11639 = ~n1603 & n8880 ;
  assign n11640 = n11639 ^ n6294 ^ 1'b0 ;
  assign n11641 = n11640 ^ n5168 ^ n3005 ;
  assign n11642 = ( x150 & n11638 ) | ( x150 & ~n11641 ) | ( n11638 & ~n11641 ) ;
  assign n11643 = n11642 ^ n9547 ^ n8251 ;
  assign n11644 = n9175 & ~n11643 ;
  assign n11645 = n8753 ^ n4000 ^ 1'b0 ;
  assign n11650 = n4717 ^ n3752 ^ n852 ;
  assign n11651 = ( ~n5268 & n9130 ) | ( ~n5268 & n11650 ) | ( n9130 & n11650 ) ;
  assign n11646 = n8003 ^ n1776 ^ 1'b0 ;
  assign n11647 = ( n1887 & n8848 ) | ( n1887 & n11646 ) | ( n8848 & n11646 ) ;
  assign n11648 = n11647 ^ n6838 ^ 1'b0 ;
  assign n11649 = n4833 & n11648 ;
  assign n11652 = n11651 ^ n11649 ^ n4071 ;
  assign n11656 = n5297 ^ x187 ^ 1'b0 ;
  assign n11654 = n10104 ^ n5693 ^ 1'b0 ;
  assign n11655 = n5031 & n11654 ;
  assign n11657 = n11656 ^ n11655 ^ n1513 ;
  assign n11653 = n7892 ^ n1430 ^ n917 ;
  assign n11658 = n11657 ^ n11653 ^ n3758 ;
  assign n11659 = n11658 ^ n8249 ^ n1214 ;
  assign n11660 = n7188 ^ n4943 ^ 1'b0 ;
  assign n11661 = n6761 & n11660 ;
  assign n11662 = n9635 ^ n734 ^ 1'b0 ;
  assign n11663 = n11661 & n11662 ;
  assign n11664 = ( n8920 & n11659 ) | ( n8920 & ~n11663 ) | ( n11659 & ~n11663 ) ;
  assign n11665 = n1429 ^ x58 ^ 1'b0 ;
  assign n11666 = n2139 | n11665 ;
  assign n11667 = n10281 ^ n7860 ^ n6432 ;
  assign n11668 = ( ~n2270 & n11666 ) | ( ~n2270 & n11667 ) | ( n11666 & n11667 ) ;
  assign n11669 = n5112 | n11668 ;
  assign n11670 = n4384 | n11669 ;
  assign n11671 = n3492 | n3749 ;
  assign n11672 = n4015 ^ n2015 ^ n446 ;
  assign n11673 = n11672 ^ n6925 ^ 1'b0 ;
  assign n11674 = ( n8109 & n11666 ) | ( n8109 & ~n11673 ) | ( n11666 & ~n11673 ) ;
  assign n11675 = n633 | n4532 ;
  assign n11676 = n11674 & n11675 ;
  assign n11677 = n5953 ^ n2892 ^ n1723 ;
  assign n11678 = ( ~n1790 & n4224 ) | ( ~n1790 & n11677 ) | ( n4224 & n11677 ) ;
  assign n11679 = n11678 ^ n7290 ^ n1213 ;
  assign n11680 = n8328 & n11679 ;
  assign n11686 = n11234 ^ n8781 ^ n5542 ;
  assign n11687 = n11686 ^ n6389 ^ n6293 ;
  assign n11681 = n6207 ^ n4068 ^ 1'b0 ;
  assign n11682 = n1077 & ~n1126 ;
  assign n11683 = ( ~n690 & n6935 ) | ( ~n690 & n11682 ) | ( n6935 & n11682 ) ;
  assign n11684 = ~n4847 & n11683 ;
  assign n11685 = n11681 & n11684 ;
  assign n11688 = n11687 ^ n11685 ^ n7462 ;
  assign n11689 = n1164 | n8853 ;
  assign n11690 = n4527 | n11689 ;
  assign n11691 = n11671 ^ n2450 ^ 1'b0 ;
  assign n11692 = n5547 ^ n3051 ^ n2471 ;
  assign n11693 = n1530 & ~n10765 ;
  assign n11694 = n4877 & n11693 ;
  assign n11695 = n11692 | n11694 ;
  assign n11696 = n11695 ^ n5715 ^ 1'b0 ;
  assign n11700 = n5596 & ~n7668 ;
  assign n11701 = ~n9702 & n11700 ;
  assign n11702 = ~n1543 & n11701 ;
  assign n11697 = n3935 ^ n3002 ^ n740 ;
  assign n11698 = ( x254 & n1826 ) | ( x254 & ~n11697 ) | ( n1826 & ~n11697 ) ;
  assign n11699 = n9115 & ~n11698 ;
  assign n11703 = n11702 ^ n11699 ^ 1'b0 ;
  assign n11712 = n1419 & ~n9250 ;
  assign n11713 = n9250 & n11712 ;
  assign n11704 = n5211 ^ n1621 ^ 1'b0 ;
  assign n11705 = n4229 ^ n4057 ^ n2950 ;
  assign n11706 = ( n5395 & n11704 ) | ( n5395 & n11705 ) | ( n11704 & n11705 ) ;
  assign n11707 = ~n1703 & n3245 ;
  assign n11708 = n2497 & n11707 ;
  assign n11709 = n11708 ^ n8740 ^ n2040 ;
  assign n11710 = ~n11706 & n11709 ;
  assign n11711 = n11706 & n11710 ;
  assign n11714 = n11713 ^ n11711 ^ n9136 ;
  assign n11720 = n11407 ^ n4626 ^ n598 ;
  assign n11715 = n6351 ^ n5808 ^ 1'b0 ;
  assign n11716 = n6510 ^ n5281 ^ n4209 ;
  assign n11717 = ( n673 & n7642 ) | ( n673 & ~n11716 ) | ( n7642 & ~n11716 ) ;
  assign n11718 = n11717 ^ n11594 ^ 1'b0 ;
  assign n11719 = n11715 & n11718 ;
  assign n11721 = n11720 ^ n11719 ^ n3182 ;
  assign n11722 = n6772 ^ n6177 ^ n5587 ;
  assign n11723 = ( n7510 & n11721 ) | ( n7510 & n11722 ) | ( n11721 & n11722 ) ;
  assign n11724 = ( n7433 & n8828 ) | ( n7433 & n11723 ) | ( n8828 & n11723 ) ;
  assign n11725 = n603 & n866 ;
  assign n11726 = n11725 ^ n668 ^ 1'b0 ;
  assign n11727 = n2000 ^ n1087 ^ n900 ;
  assign n11728 = ( n2446 & ~n3163 ) | ( n2446 & n4521 ) | ( ~n3163 & n4521 ) ;
  assign n11729 = n11728 ^ n5477 ^ n307 ;
  assign n11730 = ( n3845 & n6029 ) | ( n3845 & ~n11729 ) | ( n6029 & ~n11729 ) ;
  assign n11731 = ~n11727 & n11730 ;
  assign n11732 = n11731 ^ n2625 ^ 1'b0 ;
  assign n11733 = ( ~n313 & n5051 ) | ( ~n313 & n8634 ) | ( n5051 & n8634 ) ;
  assign n11735 = n1299 ^ n989 ^ 1'b0 ;
  assign n11734 = n893 | n9357 ;
  assign n11736 = n11735 ^ n11734 ^ 1'b0 ;
  assign n11737 = ( n3919 & ~n5902 ) | ( n3919 & n11736 ) | ( ~n5902 & n11736 ) ;
  assign n11738 = n1659 & ~n11737 ;
  assign n11739 = n11738 ^ n7987 ^ 1'b0 ;
  assign n11740 = n1717 & n11739 ;
  assign n11741 = n11733 & n11740 ;
  assign n11742 = ~n6027 & n11741 ;
  assign n11743 = n11732 | n11742 ;
  assign n11744 = n11726 & ~n11743 ;
  assign n11757 = ( n1103 & n8017 ) | ( n1103 & ~n11402 ) | ( n8017 & ~n11402 ) ;
  assign n11758 = n11757 ^ n9854 ^ 1'b0 ;
  assign n11752 = n1444 | n1846 ;
  assign n11753 = ~n5323 & n11752 ;
  assign n11754 = ~n935 & n11753 ;
  assign n11755 = n11754 ^ n8145 ^ n6038 ;
  assign n11756 = n5152 & n11755 ;
  assign n11745 = n9625 ^ n625 ^ 1'b0 ;
  assign n11746 = n3476 & ~n11745 ;
  assign n11747 = ( n1682 & n9804 ) | ( n1682 & n11746 ) | ( n9804 & n11746 ) ;
  assign n11748 = ~n10563 & n11747 ;
  assign n11749 = ( x188 & n4755 ) | ( x188 & n9537 ) | ( n4755 & n9537 ) ;
  assign n11750 = n11749 ^ n10068 ^ 1'b0 ;
  assign n11751 = n11748 & ~n11750 ;
  assign n11759 = n11758 ^ n11756 ^ n11751 ;
  assign n11760 = ( ~n5919 & n7285 ) | ( ~n5919 & n11205 ) | ( n7285 & n11205 ) ;
  assign n11761 = n5655 & ~n11760 ;
  assign n11762 = n6747 ^ n6025 ^ 1'b0 ;
  assign n11763 = ( n10980 & n11761 ) | ( n10980 & n11762 ) | ( n11761 & n11762 ) ;
  assign n11764 = n7766 ^ n7056 ^ 1'b0 ;
  assign n11765 = n10621 ^ n683 ^ 1'b0 ;
  assign n11766 = n4512 | n11765 ;
  assign n11767 = n8337 ^ n2707 ^ 1'b0 ;
  assign n11768 = ~n4245 & n11767 ;
  assign n11769 = n11766 & n11768 ;
  assign n11771 = ( n592 & ~n593 ) | ( n592 & n5145 ) | ( ~n593 & n5145 ) ;
  assign n11770 = x192 & ~n888 ;
  assign n11772 = n11771 ^ n11770 ^ 1'b0 ;
  assign n11773 = n6232 ^ n3586 ^ 1'b0 ;
  assign n11774 = n11773 ^ n2087 ^ n1714 ;
  assign n11775 = n6583 ^ n6407 ^ n4634 ;
  assign n11776 = n11775 ^ n901 ^ 1'b0 ;
  assign n11777 = n11774 & ~n11776 ;
  assign n11778 = n11772 & n11777 ;
  assign n11779 = ~n6186 & n11778 ;
  assign n11780 = ( ~n3109 & n4696 ) | ( ~n3109 & n11779 ) | ( n4696 & n11779 ) ;
  assign n11784 = n2380 & n5262 ;
  assign n11782 = ( n1246 & n2472 ) | ( n1246 & ~n4307 ) | ( n2472 & ~n4307 ) ;
  assign n11783 = ( n260 & ~n8032 ) | ( n260 & n11782 ) | ( ~n8032 & n11782 ) ;
  assign n11785 = n11784 ^ n11783 ^ n7477 ;
  assign n11781 = n4117 & ~n7596 ;
  assign n11786 = n11785 ^ n11781 ^ 1'b0 ;
  assign n11787 = n410 | n10153 ;
  assign n11788 = n813 | n7806 ;
  assign n11789 = ~n1747 & n5676 ;
  assign n11790 = ~n5705 & n11789 ;
  assign n11791 = ~n11788 & n11790 ;
  assign n11792 = n3365 & ~n11791 ;
  assign n11793 = n11792 ^ n3385 ^ 1'b0 ;
  assign n11794 = ( x88 & ~n2532 ) | ( x88 & n11793 ) | ( ~n2532 & n11793 ) ;
  assign n11795 = ( n10652 & ~n11180 ) | ( n10652 & n11794 ) | ( ~n11180 & n11794 ) ;
  assign n11796 = n1461 & n10499 ;
  assign n11797 = n2014 & n5264 ;
  assign n11798 = ~n459 & n11797 ;
  assign n11799 = n4415 | n11798 ;
  assign n11800 = n3593 | n11799 ;
  assign n11801 = n6167 ^ n6106 ^ 1'b0 ;
  assign n11802 = n11801 ^ n11733 ^ 1'b0 ;
  assign n11803 = n11802 ^ n8858 ^ n4191 ;
  assign n11804 = n4798 & n11359 ;
  assign n11805 = ~n4800 & n11804 ;
  assign n11806 = ( n11800 & n11803 ) | ( n11800 & n11805 ) | ( n11803 & n11805 ) ;
  assign n11807 = n2042 | n11798 ;
  assign n11808 = n2067 | n11807 ;
  assign n11811 = n10261 ^ n8843 ^ 1'b0 ;
  assign n11809 = ~n1091 & n3162 ;
  assign n11810 = n11809 ^ n11366 ^ 1'b0 ;
  assign n11812 = n11811 ^ n11810 ^ n5555 ;
  assign n11813 = n11812 ^ n9805 ^ 1'b0 ;
  assign n11814 = n5014 | n11813 ;
  assign n11815 = n4229 & n6403 ;
  assign n11816 = n6451 & n11815 ;
  assign n11817 = ( n6353 & n7664 ) | ( n6353 & n11641 ) | ( n7664 & n11641 ) ;
  assign n11818 = n8580 ^ n6297 ^ 1'b0 ;
  assign n11819 = n11818 ^ n2388 ^ 1'b0 ;
  assign n11820 = n11221 ^ n9671 ^ n3831 ;
  assign n11821 = ( x145 & n9064 ) | ( x145 & ~n11820 ) | ( n9064 & ~n11820 ) ;
  assign n11822 = ( n4524 & n11819 ) | ( n4524 & ~n11821 ) | ( n11819 & ~n11821 ) ;
  assign n11823 = n8933 ^ n5759 ^ 1'b0 ;
  assign n11832 = n433 & ~n9643 ;
  assign n11833 = n11832 ^ n9135 ^ 1'b0 ;
  assign n11834 = ( n6384 & ~n6519 ) | ( n6384 & n11833 ) | ( ~n6519 & n11833 ) ;
  assign n11835 = n3159 | n3825 ;
  assign n11836 = n11834 | n11835 ;
  assign n11831 = n9604 ^ n3891 ^ 1'b0 ;
  assign n11837 = n11836 ^ n11831 ^ n2562 ;
  assign n11830 = n3167 ^ n399 ^ 1'b0 ;
  assign n11838 = n11837 ^ n11830 ^ n8444 ;
  assign n11826 = n3629 | n5059 ;
  assign n11827 = n11826 ^ n6483 ^ 1'b0 ;
  assign n11828 = n11827 ^ n2405 ^ n774 ;
  assign n11824 = ~n1293 & n8425 ;
  assign n11825 = n975 | n11824 ;
  assign n11829 = n11828 ^ n11825 ^ 1'b0 ;
  assign n11839 = n11838 ^ n11829 ^ n8539 ;
  assign n11840 = n7480 ^ n6590 ^ n1414 ;
  assign n11841 = n11840 ^ n6954 ^ 1'b0 ;
  assign n11842 = n9328 ^ n4975 ^ n3851 ;
  assign n11843 = n3643 & ~n5277 ;
  assign n11845 = ( ~n2746 & n4206 ) | ( ~n2746 & n5392 ) | ( n4206 & n5392 ) ;
  assign n11844 = n2651 ^ x193 ^ 1'b0 ;
  assign n11846 = n11845 ^ n11844 ^ n4640 ;
  assign n11848 = n5631 ^ n3999 ^ n643 ;
  assign n11849 = ( n5709 & ~n6440 ) | ( n5709 & n11848 ) | ( ~n6440 & n11848 ) ;
  assign n11847 = ~n2592 & n11258 ;
  assign n11850 = n11849 ^ n11847 ^ 1'b0 ;
  assign n11857 = n1180 | n2298 ;
  assign n11858 = n11857 ^ n1575 ^ 1'b0 ;
  assign n11859 = ( n3247 & n4305 ) | ( n3247 & n11858 ) | ( n4305 & n11858 ) ;
  assign n11860 = ~n5469 & n11859 ;
  assign n11861 = n8979 & n11860 ;
  assign n11862 = n4113 & ~n11861 ;
  assign n11863 = n11862 ^ n1528 ^ 1'b0 ;
  assign n11853 = n10808 ^ n765 ^ 1'b0 ;
  assign n11854 = n8646 | n11853 ;
  assign n11852 = ( n865 & n4960 ) | ( n865 & n6616 ) | ( n4960 & n6616 ) ;
  assign n11851 = n4948 ^ n4469 ^ n3756 ;
  assign n11855 = n11854 ^ n11852 ^ n11851 ;
  assign n11856 = n11855 ^ n11335 ^ n9946 ;
  assign n11864 = n11863 ^ n11856 ^ 1'b0 ;
  assign n11865 = n1100 | n11864 ;
  assign n11866 = n8425 ^ n6006 ^ 1'b0 ;
  assign n11868 = ~n3606 & n4633 ;
  assign n11867 = x44 | n3055 ;
  assign n11869 = n11868 ^ n11867 ^ 1'b0 ;
  assign n11870 = ~n3567 & n11869 ;
  assign n11871 = n11866 & n11870 ;
  assign n11872 = n7303 & ~n7780 ;
  assign n11873 = n11872 ^ n5263 ^ 1'b0 ;
  assign n11874 = ( n300 & n11380 ) | ( n300 & n11873 ) | ( n11380 & n11873 ) ;
  assign n11875 = ( n2493 & n7596 ) | ( n2493 & ~n9641 ) | ( n7596 & ~n9641 ) ;
  assign n11876 = n5679 ^ n1993 ^ 1'b0 ;
  assign n11877 = n2317 | n2822 ;
  assign n11878 = n11877 ^ n4618 ^ 1'b0 ;
  assign n11879 = ~n1112 & n7832 ;
  assign n11880 = n11878 & n11879 ;
  assign n11881 = n11880 ^ n6662 ^ n5991 ;
  assign n11882 = n313 & n11881 ;
  assign n11883 = n11876 & n11882 ;
  assign n11884 = n8003 ^ n3043 ^ x246 ;
  assign n11885 = ( n3931 & n8734 ) | ( n3931 & n11884 ) | ( n8734 & n11884 ) ;
  assign n11886 = n1638 ^ n1162 ^ 1'b0 ;
  assign n11887 = ( n1015 & n1919 ) | ( n1015 & n4499 ) | ( n1919 & n4499 ) ;
  assign n11888 = n3774 | n11887 ;
  assign n11889 = n3644 & ~n11888 ;
  assign n11890 = n6169 & n11889 ;
  assign n11891 = ( ~n6767 & n11886 ) | ( ~n6767 & n11890 ) | ( n11886 & n11890 ) ;
  assign n11892 = ( n11883 & ~n11885 ) | ( n11883 & n11891 ) | ( ~n11885 & n11891 ) ;
  assign n11893 = ( ~n565 & n3933 ) | ( ~n565 & n6062 ) | ( n3933 & n6062 ) ;
  assign n11894 = n11893 ^ n5353 ^ 1'b0 ;
  assign n11895 = n7818 & n11894 ;
  assign n11896 = ( n2050 & ~n4225 ) | ( n2050 & n11895 ) | ( ~n4225 & n11895 ) ;
  assign n11897 = n11896 ^ n7052 ^ 1'b0 ;
  assign n11898 = ( ~n857 & n5317 ) | ( ~n857 & n9900 ) | ( n5317 & n9900 ) ;
  assign n11899 = x71 & ~n2064 ;
  assign n11900 = ~x239 & n11899 ;
  assign n11901 = n1886 & n4592 ;
  assign n11902 = n10004 & n11901 ;
  assign n11903 = n11900 & n11902 ;
  assign n11904 = ( n2807 & n2992 ) | ( n2807 & ~n11903 ) | ( n2992 & ~n11903 ) ;
  assign n11905 = n4379 ^ n2664 ^ 1'b0 ;
  assign n11906 = n6780 ^ n6326 ^ 1'b0 ;
  assign n11907 = n10918 & ~n11906 ;
  assign n11908 = n11905 & n11907 ;
  assign n11909 = n11904 & ~n11908 ;
  assign n11910 = n5283 & n11909 ;
  assign n11911 = n6909 ^ n3994 ^ 1'b0 ;
  assign n11912 = n6618 & n11911 ;
  assign n11913 = n4097 & n11912 ;
  assign n11914 = n11913 ^ n902 ^ 1'b0 ;
  assign n11915 = ( n1834 & n5876 ) | ( n1834 & n11914 ) | ( n5876 & n11914 ) ;
  assign n11916 = n10177 ^ n1938 ^ n1404 ;
  assign n11917 = n11916 ^ n1655 ^ 1'b0 ;
  assign n11918 = n11917 ^ n6822 ^ 1'b0 ;
  assign n11919 = n11915 & ~n11918 ;
  assign n11920 = ( n2237 & ~n2819 ) | ( n2237 & n7047 ) | ( ~n2819 & n7047 ) ;
  assign n11921 = ~n1190 & n3472 ;
  assign n11922 = ~x91 & n11921 ;
  assign n11923 = n10667 ^ n7425 ^ 1'b0 ;
  assign n11924 = n11492 ^ n7573 ^ n2217 ;
  assign n11925 = ( ~n9512 & n11283 ) | ( ~n9512 & n11924 ) | ( n11283 & n11924 ) ;
  assign n11926 = n11827 ^ n8376 ^ n6410 ;
  assign n11927 = ( x166 & n6049 ) | ( x166 & n11926 ) | ( n6049 & n11926 ) ;
  assign n11928 = x183 & n5833 ;
  assign n11929 = n8393 & n11928 ;
  assign n11930 = n2452 | n7572 ;
  assign n11931 = n4257 | n11930 ;
  assign n11932 = ( n2434 & n2871 ) | ( n2434 & ~n11931 ) | ( n2871 & ~n11931 ) ;
  assign n11933 = ( ~n9041 & n11929 ) | ( ~n9041 & n11932 ) | ( n11929 & n11932 ) ;
  assign n11934 = n7171 & ~n11933 ;
  assign n11935 = n2130 & n11934 ;
  assign n11936 = n1088 | n6925 ;
  assign n11937 = n11936 ^ n3484 ^ 1'b0 ;
  assign n11942 = n1391 & ~n10709 ;
  assign n11938 = ~n2355 & n6966 ;
  assign n11939 = n2329 & n11938 ;
  assign n11940 = n1892 | n11939 ;
  assign n11941 = n11940 ^ n355 ^ 1'b0 ;
  assign n11943 = n11942 ^ n11941 ^ n6768 ;
  assign n11944 = n8218 ^ n3516 ^ 1'b0 ;
  assign n11945 = ( n1007 & n1087 ) | ( n1007 & ~n2492 ) | ( n1087 & ~n2492 ) ;
  assign n11946 = n4063 ^ x68 ^ 1'b0 ;
  assign n11947 = n2667 & n11946 ;
  assign n11948 = n1872 & n11947 ;
  assign n11949 = n11948 ^ n5234 ^ 1'b0 ;
  assign n11950 = ( n1705 & ~n11945 ) | ( n1705 & n11949 ) | ( ~n11945 & n11949 ) ;
  assign n11951 = n11950 ^ n3692 ^ n585 ;
  assign n11952 = ( n4529 & n11944 ) | ( n4529 & n11951 ) | ( n11944 & n11951 ) ;
  assign n11953 = n2280 & n2697 ;
  assign n11954 = n11953 ^ n4972 ^ 1'b0 ;
  assign n11955 = ~n556 & n11954 ;
  assign n11956 = n8017 & n11955 ;
  assign n11957 = n11956 ^ n1334 ^ n1104 ;
  assign n11958 = n3171 & ~n10424 ;
  assign n11959 = n9278 ^ n6318 ^ 1'b0 ;
  assign n11961 = n9672 ^ n4865 ^ n802 ;
  assign n11960 = ( n1612 & n4441 ) | ( n1612 & n8475 ) | ( n4441 & n8475 ) ;
  assign n11962 = n11961 ^ n11960 ^ n5562 ;
  assign n11963 = n6760 & n7795 ;
  assign n11964 = n11962 & n11963 ;
  assign n11965 = n4309 | n11964 ;
  assign n11966 = n5519 & n8716 ;
  assign n11967 = n1984 & n10239 ;
  assign n11968 = n4722 & ~n11967 ;
  assign n11969 = n1961 & n4674 ;
  assign n11970 = ( n11966 & ~n11968 ) | ( n11966 & n11969 ) | ( ~n11968 & n11969 ) ;
  assign n11971 = ( ~n984 & n5147 ) | ( ~n984 & n5620 ) | ( n5147 & n5620 ) ;
  assign n11972 = n11971 ^ n11050 ^ 1'b0 ;
  assign n11973 = n286 & ~n11972 ;
  assign n11974 = n4800 & n6075 ;
  assign n11975 = n4500 ^ n2115 ^ 1'b0 ;
  assign n11976 = ( ~n7347 & n11974 ) | ( ~n7347 & n11975 ) | ( n11974 & n11975 ) ;
  assign n11977 = n5875 ^ n5254 ^ 1'b0 ;
  assign n11978 = n1866 | n11977 ;
  assign n11979 = n2022 | n11978 ;
  assign n11980 = n11976 | n11979 ;
  assign n11981 = n2954 ^ x18 ^ 1'b0 ;
  assign n11982 = ~n2250 & n11981 ;
  assign n11983 = n2394 & n2992 ;
  assign n11984 = ~n11982 & n11983 ;
  assign n11985 = n11984 ^ n10506 ^ n3353 ;
  assign n11986 = n11985 ^ n3955 ^ n2526 ;
  assign n11987 = ( n6204 & n10172 ) | ( n6204 & ~n10328 ) | ( n10172 & ~n10328 ) ;
  assign n11991 = n2993 ^ n676 ^ 1'b0 ;
  assign n11996 = n1580 ^ n808 ^ n806 ;
  assign n11995 = n1538 & ~n2478 ;
  assign n11992 = n2442 ^ n775 ^ n540 ;
  assign n11993 = n3159 | n11992 ;
  assign n11994 = n11993 ^ n7189 ^ 1'b0 ;
  assign n11997 = n11996 ^ n11995 ^ n11994 ;
  assign n11998 = ( n2967 & ~n11991 ) | ( n2967 & n11997 ) | ( ~n11991 & n11997 ) ;
  assign n11988 = n4064 & n8996 ;
  assign n11989 = n11988 ^ x227 ^ 1'b0 ;
  assign n11990 = ( n1140 & ~n2146 ) | ( n1140 & n11989 ) | ( ~n2146 & n11989 ) ;
  assign n11999 = n11998 ^ n11990 ^ 1'b0 ;
  assign n12000 = ( n5321 & n7309 ) | ( n5321 & n11793 ) | ( n7309 & n11793 ) ;
  assign n12001 = n12000 ^ n9132 ^ n2657 ;
  assign n12002 = ( ~x164 & n3255 ) | ( ~x164 & n4783 ) | ( n3255 & n4783 ) ;
  assign n12003 = n12002 ^ n900 ^ 1'b0 ;
  assign n12004 = n5411 & n12003 ;
  assign n12005 = n10996 & n12004 ;
  assign n12006 = n11046 & ~n12005 ;
  assign n12007 = n1226 | n2497 ;
  assign n12008 = n1166 & n4451 ;
  assign n12009 = n6844 | n12008 ;
  assign n12010 = n12007 & ~n12009 ;
  assign n12011 = n6038 ^ n1763 ^ 1'b0 ;
  assign n12012 = n3933 & n10229 ;
  assign n12013 = n298 & ~n345 ;
  assign n12014 = n12012 & n12013 ;
  assign n12032 = n5110 ^ n780 ^ x34 ;
  assign n12033 = ( ~n8119 & n10738 ) | ( ~n8119 & n12032 ) | ( n10738 & n12032 ) ;
  assign n12034 = ( n3650 & n8704 ) | ( n3650 & n12033 ) | ( n8704 & n12033 ) ;
  assign n12015 = n7708 ^ n5721 ^ n1185 ;
  assign n12023 = x132 & n2045 ;
  assign n12024 = n12023 ^ n3497 ^ 1'b0 ;
  assign n12018 = x133 & ~n6944 ;
  assign n12016 = n7036 ^ n1278 ^ 1'b0 ;
  assign n12017 = n7851 & ~n12016 ;
  assign n12019 = n12018 ^ n12017 ^ n9205 ;
  assign n12020 = x254 & ~n12019 ;
  assign n12021 = n870 & n12020 ;
  assign n12022 = ~n4375 & n12021 ;
  assign n12025 = n12024 ^ n12022 ^ 1'b0 ;
  assign n12026 = ~n7164 & n12025 ;
  assign n12027 = n2936 & n10918 ;
  assign n12028 = n12027 ^ n9938 ^ 1'b0 ;
  assign n12029 = n12028 ^ n8027 ^ 1'b0 ;
  assign n12030 = ( ~n4518 & n12026 ) | ( ~n4518 & n12029 ) | ( n12026 & n12029 ) ;
  assign n12031 = n12015 & n12030 ;
  assign n12035 = n12034 ^ n12031 ^ 1'b0 ;
  assign n12036 = ( n2736 & n2840 ) | ( n2736 & ~n5236 ) | ( n2840 & ~n5236 ) ;
  assign n12037 = n9558 ^ n7769 ^ n6702 ;
  assign n12038 = ~n12036 & n12037 ;
  assign n12048 = n1433 & ~n7683 ;
  assign n12043 = ~n900 & n8163 ;
  assign n12044 = n12043 ^ n11735 ^ 1'b0 ;
  assign n12045 = ( n2707 & ~n3486 ) | ( n2707 & n12044 ) | ( ~n3486 & n12044 ) ;
  assign n12046 = n10099 | n12045 ;
  assign n12047 = n12046 ^ n2631 ^ n1044 ;
  assign n12039 = n5732 & n8143 ;
  assign n12040 = n12039 ^ n2543 ^ 1'b0 ;
  assign n12041 = n5894 & n12040 ;
  assign n12042 = ( n1102 & n2209 ) | ( n1102 & n12041 ) | ( n2209 & n12041 ) ;
  assign n12049 = n12048 ^ n12047 ^ n12042 ;
  assign n12064 = ( n1288 & n1816 ) | ( n1288 & ~n10765 ) | ( n1816 & ~n10765 ) ;
  assign n12065 = n12064 ^ n5454 ^ n4709 ;
  assign n12058 = n1822 ^ n475 ^ 1'b0 ;
  assign n12059 = n2994 & n12058 ;
  assign n12060 = n12059 ^ n11379 ^ n472 ;
  assign n12061 = n2184 ^ n905 ^ 1'b0 ;
  assign n12062 = n12060 & ~n12061 ;
  assign n12052 = n5281 ^ n4517 ^ n1767 ;
  assign n12053 = n12052 ^ n7035 ^ 1'b0 ;
  assign n12054 = n478 & ~n7718 ;
  assign n12055 = n2657 & n12054 ;
  assign n12056 = n12055 ^ n3015 ^ 1'b0 ;
  assign n12057 = ~n12053 & n12056 ;
  assign n12050 = n788 ^ x184 ^ 1'b0 ;
  assign n12051 = n12050 ^ n6365 ^ 1'b0 ;
  assign n12063 = n12062 ^ n12057 ^ n12051 ;
  assign n12066 = n12065 ^ n12063 ^ n3569 ;
  assign n12067 = n5262 & ~n6260 ;
  assign n12068 = ~n9117 & n12067 ;
  assign n12069 = n6485 ^ n2292 ^ n1152 ;
  assign n12070 = ( n5810 & ~n8168 ) | ( n5810 & n12069 ) | ( ~n8168 & n12069 ) ;
  assign n12071 = n12070 ^ n10872 ^ n7349 ;
  assign n12073 = n2173 ^ n1536 ^ 1'b0 ;
  assign n12072 = ~n7973 & n9305 ;
  assign n12074 = n12073 ^ n12072 ^ 1'b0 ;
  assign n12075 = n9167 & ~n12074 ;
  assign n12076 = n10252 | n12075 ;
  assign n12077 = ~n6706 & n8472 ;
  assign n12078 = n12077 ^ n9461 ^ 1'b0 ;
  assign n12080 = ( x31 & ~n1097 ) | ( x31 & n1129 ) | ( ~n1097 & n1129 ) ;
  assign n12081 = n3157 & n12080 ;
  assign n12082 = ~n3234 & n12081 ;
  assign n12083 = n12082 ^ n2593 ^ 1'b0 ;
  assign n12079 = n10738 & ~n10877 ;
  assign n12084 = n12083 ^ n12079 ^ 1'b0 ;
  assign n12085 = n9069 ^ n1833 ^ n510 ;
  assign n12086 = ( ~n3532 & n9072 ) | ( ~n3532 & n10140 ) | ( n9072 & n10140 ) ;
  assign n12087 = n12086 ^ n9115 ^ 1'b0 ;
  assign n12088 = n4018 ^ n2702 ^ 1'b0 ;
  assign n12089 = ~n2610 & n12088 ;
  assign n12090 = ( n5601 & n10243 ) | ( n5601 & ~n12089 ) | ( n10243 & ~n12089 ) ;
  assign n12092 = n5390 ^ n4510 ^ 1'b0 ;
  assign n12093 = n2638 | n12092 ;
  assign n12091 = n2873 & ~n6000 ;
  assign n12094 = n12093 ^ n12091 ^ 1'b0 ;
  assign n12100 = n7354 ^ n6881 ^ n1157 ;
  assign n12097 = n1864 | n10246 ;
  assign n12095 = n9461 ^ n3544 ^ 1'b0 ;
  assign n12096 = n5643 & ~n12095 ;
  assign n12098 = n12097 ^ n12096 ^ n11820 ;
  assign n12099 = n12098 ^ n11638 ^ n9997 ;
  assign n12101 = n12100 ^ n12099 ^ 1'b0 ;
  assign n12102 = n9238 & ~n12101 ;
  assign n12103 = n10030 ^ n7125 ^ n2209 ;
  assign n12104 = n12103 ^ n8135 ^ n5346 ;
  assign n12105 = ( ~n2474 & n9460 ) | ( ~n2474 & n12104 ) | ( n9460 & n12104 ) ;
  assign n12106 = n381 & ~n8991 ;
  assign n12107 = x186 & ~n7248 ;
  assign n12108 = n12107 ^ n5317 ^ 1'b0 ;
  assign n12109 = n5732 ^ n5569 ^ n1867 ;
  assign n12110 = n260 & ~n6965 ;
  assign n12111 = ~n2325 & n12110 ;
  assign n12112 = n12109 & n12111 ;
  assign n12113 = x69 ^ x3 ^ 1'b0 ;
  assign n12114 = n3979 ^ n1358 ^ n954 ;
  assign n12115 = x88 & ~n12114 ;
  assign n12116 = ~n9394 & n12115 ;
  assign n12117 = n2817 ^ n1177 ^ x154 ;
  assign n12118 = n12117 ^ x75 ^ 1'b0 ;
  assign n12119 = ~n9752 & n12118 ;
  assign n12120 = ~n12116 & n12119 ;
  assign n12121 = ( n547 & n12113 ) | ( n547 & ~n12120 ) | ( n12113 & ~n12120 ) ;
  assign n12124 = n1829 & n6501 ;
  assign n12125 = n9167 & n12124 ;
  assign n12122 = n337 | n7186 ;
  assign n12123 = n12122 ^ n6711 ^ 1'b0 ;
  assign n12126 = n12125 ^ n12123 ^ 1'b0 ;
  assign n12127 = ~n6261 & n12126 ;
  assign n12128 = n3326 & n6413 ;
  assign n12129 = n12128 ^ n11914 ^ n7511 ;
  assign n12130 = ( n436 & n1431 ) | ( n436 & n12129 ) | ( n1431 & n12129 ) ;
  assign n12131 = n4633 ^ n3646 ^ n2914 ;
  assign n12132 = n5856 ^ n1228 ^ n443 ;
  assign n12133 = ( n7633 & n12131 ) | ( n7633 & ~n12132 ) | ( n12131 & ~n12132 ) ;
  assign n12134 = n12133 ^ n11651 ^ n6913 ;
  assign n12135 = n1370 & ~n8066 ;
  assign n12136 = n12135 ^ x185 ^ 1'b0 ;
  assign n12137 = ~n4386 & n12136 ;
  assign n12138 = n12137 ^ n10815 ^ 1'b0 ;
  assign n12139 = ~n6062 & n8307 ;
  assign n12140 = n12139 ^ n1062 ^ 1'b0 ;
  assign n12141 = n12140 ^ n10555 ^ n7306 ;
  assign n12142 = n8260 & ~n12141 ;
  assign n12143 = n6300 ^ n3620 ^ n1014 ;
  assign n12144 = ( ~n1755 & n6190 ) | ( ~n1755 & n12143 ) | ( n6190 & n12143 ) ;
  assign n12145 = n12144 ^ n10068 ^ n8762 ;
  assign n12146 = n12145 ^ n4820 ^ n678 ;
  assign n12147 = n2008 ^ n910 ^ 1'b0 ;
  assign n12148 = n5715 | n12147 ;
  assign n12149 = ( ~n3278 & n6107 ) | ( ~n3278 & n12148 ) | ( n6107 & n12148 ) ;
  assign n12150 = x198 & n3324 ;
  assign n12151 = ~n3367 & n12150 ;
  assign n12152 = ( n304 & n10512 ) | ( n304 & ~n12151 ) | ( n10512 & ~n12151 ) ;
  assign n12153 = ~n3618 & n11990 ;
  assign n12154 = n8707 ^ n2168 ^ 1'b0 ;
  assign n12155 = n8493 | n12154 ;
  assign n12156 = n8705 ^ n4926 ^ 1'b0 ;
  assign n12157 = ~n5728 & n12156 ;
  assign n12158 = n4194 & n10383 ;
  assign n12161 = ( n4873 & n10159 ) | ( n4873 & ~n11022 ) | ( n10159 & ~n11022 ) ;
  assign n12159 = ~n687 & n3280 ;
  assign n12160 = ~n3134 & n12159 ;
  assign n12162 = n12161 ^ n12160 ^ 1'b0 ;
  assign n12166 = n5676 & ~n8241 ;
  assign n12167 = n12166 ^ n7702 ^ 1'b0 ;
  assign n12163 = ( n1856 & ~n2367 ) | ( n1856 & n8853 ) | ( ~n2367 & n8853 ) ;
  assign n12164 = ( n6994 & n9548 ) | ( n6994 & ~n12144 ) | ( n9548 & ~n12144 ) ;
  assign n12165 = n12163 & ~n12164 ;
  assign n12168 = n12167 ^ n12165 ^ 1'b0 ;
  assign n12169 = n5302 & n7938 ;
  assign n12170 = n7195 ^ n462 ^ 1'b0 ;
  assign n12171 = n12169 & n12170 ;
  assign n12172 = n6696 & n8606 ;
  assign n12173 = n12172 ^ n4948 ^ 1'b0 ;
  assign n12176 = n6634 ^ n6608 ^ n5541 ;
  assign n12177 = n12176 ^ n4813 ^ n3350 ;
  assign n12174 = n4288 ^ n2680 ^ 1'b0 ;
  assign n12175 = n11530 | n12174 ;
  assign n12178 = n12177 ^ n12175 ^ 1'b0 ;
  assign n12179 = ( ~x148 & n5343 ) | ( ~x148 & n5723 ) | ( n5343 & n5723 ) ;
  assign n12180 = n12179 ^ n4971 ^ n887 ;
  assign n12181 = n12180 ^ n10159 ^ 1'b0 ;
  assign n12182 = ( n2036 & n12178 ) | ( n2036 & ~n12181 ) | ( n12178 & ~n12181 ) ;
  assign n12183 = n2648 & ~n3485 ;
  assign n12184 = ~n3798 & n12183 ;
  assign n12185 = ( n2163 & n9758 ) | ( n2163 & ~n12184 ) | ( n9758 & ~n12184 ) ;
  assign n12186 = n12185 ^ x188 ^ 1'b0 ;
  assign n12187 = n6901 | n12186 ;
  assign n12188 = ( n2369 & n3483 ) | ( n2369 & ~n6826 ) | ( n3483 & ~n6826 ) ;
  assign n12189 = n2773 | n12188 ;
  assign n12190 = n8416 & ~n12189 ;
  assign n12191 = n5992 ^ n446 ^ 1'b0 ;
  assign n12192 = n1277 & n8505 ;
  assign n12193 = ~n3231 & n12192 ;
  assign n12194 = n3043 & ~n12193 ;
  assign n12195 = ~n6554 & n10010 ;
  assign n12196 = n12195 ^ n2194 ^ 1'b0 ;
  assign n12197 = ( n1720 & ~n4210 ) | ( n1720 & n11784 ) | ( ~n4210 & n11784 ) ;
  assign n12201 = n497 | n8759 ;
  assign n12198 = ( ~n2255 & n6649 ) | ( ~n2255 & n8124 ) | ( n6649 & n8124 ) ;
  assign n12199 = n12198 ^ n6232 ^ 1'b0 ;
  assign n12200 = n12199 ^ n8187 ^ 1'b0 ;
  assign n12202 = n12201 ^ n12200 ^ n9761 ;
  assign n12203 = n12202 ^ n10928 ^ 1'b0 ;
  assign n12204 = n12197 & n12203 ;
  assign n12205 = ~n305 & n8084 ;
  assign n12206 = n12205 ^ n408 ^ 1'b0 ;
  assign n12207 = ( n3804 & n7381 ) | ( n3804 & ~n12206 ) | ( n7381 & ~n12206 ) ;
  assign n12208 = n12207 ^ n8634 ^ 1'b0 ;
  assign n12209 = ( n1756 & n2014 ) | ( n1756 & ~n8130 ) | ( n2014 & ~n8130 ) ;
  assign n12210 = n10021 ^ n4042 ^ 1'b0 ;
  assign n12211 = n5391 & n12210 ;
  assign n12212 = n6678 & n12211 ;
  assign n12213 = ~n12209 & n12212 ;
  assign n12214 = n2483 | n4137 ;
  assign n12215 = n1403 & n12214 ;
  assign n12226 = ( n734 & ~n4756 ) | ( n734 & n6234 ) | ( ~n4756 & n6234 ) ;
  assign n12227 = n12226 ^ n3895 ^ 1'b0 ;
  assign n12216 = n8492 ^ n3187 ^ n2768 ;
  assign n12217 = n9056 ^ n6966 ^ 1'b0 ;
  assign n12218 = ~n4512 & n12217 ;
  assign n12219 = n4437 & ~n12218 ;
  assign n12220 = n12219 ^ n11141 ^ n6582 ;
  assign n12221 = n8445 ^ n1755 ^ n1102 ;
  assign n12222 = ( ~x193 & n3725 ) | ( ~x193 & n12221 ) | ( n3725 & n12221 ) ;
  assign n12223 = n8411 | n12222 ;
  assign n12224 = n12220 & ~n12223 ;
  assign n12225 = n12216 & ~n12224 ;
  assign n12228 = n12227 ^ n12225 ^ 1'b0 ;
  assign n12229 = ~n3687 & n10928 ;
  assign n12230 = x34 & ~n2066 ;
  assign n12231 = n12230 ^ n5738 ^ n438 ;
  assign n12232 = ( n6099 & ~n9283 ) | ( n6099 & n12231 ) | ( ~n9283 & n12231 ) ;
  assign n12233 = n3493 ^ n1544 ^ n1014 ;
  assign n12234 = ( n2493 & n4329 ) | ( n2493 & n6883 ) | ( n4329 & n6883 ) ;
  assign n12235 = ( n6762 & ~n12233 ) | ( n6762 & n12234 ) | ( ~n12233 & n12234 ) ;
  assign n12236 = n12235 ^ n4462 ^ 1'b0 ;
  assign n12237 = n8008 ^ n6994 ^ 1'b0 ;
  assign n12238 = n10261 ^ n7636 ^ n1485 ;
  assign n12239 = n12238 ^ n4716 ^ n3825 ;
  assign n12240 = n11740 | n12239 ;
  assign n12241 = n12240 ^ n1734 ^ 1'b0 ;
  assign n12242 = n7696 & ~n12241 ;
  assign n12243 = n3259 ^ n2213 ^ n472 ;
  assign n12244 = ( n554 & n1773 ) | ( n554 & ~n12243 ) | ( n1773 & ~n12243 ) ;
  assign n12245 = n12244 ^ n9155 ^ n7936 ;
  assign n12246 = n6971 | n10480 ;
  assign n12247 = n4967 & ~n12246 ;
  assign n12248 = n12247 ^ n1351 ^ 1'b0 ;
  assign n12249 = ( x15 & n2031 ) | ( x15 & n4024 ) | ( n2031 & n4024 ) ;
  assign n12250 = n12249 ^ n2329 ^ 1'b0 ;
  assign n12251 = n2056 & ~n2794 ;
  assign n12252 = n12251 ^ n3481 ^ 1'b0 ;
  assign n12253 = ~n9167 & n10129 ;
  assign n12254 = ~n12252 & n12253 ;
  assign n12255 = ~n5784 & n12254 ;
  assign n12256 = n12250 | n12255 ;
  assign n12257 = n7904 & ~n12256 ;
  assign n12258 = n8148 & n8170 ;
  assign n12259 = n12258 ^ n10751 ^ 1'b0 ;
  assign n12261 = n3331 ^ n753 ^ 1'b0 ;
  assign n12260 = ( n2165 & n4464 ) | ( n2165 & n8113 ) | ( n4464 & n8113 ) ;
  assign n12262 = n12261 ^ n12260 ^ n8888 ;
  assign n12263 = n1330 & ~n6368 ;
  assign n12264 = n10260 | n12263 ;
  assign n12265 = ~n3439 & n8931 ;
  assign n12266 = n5393 ^ x235 ^ 1'b0 ;
  assign n12267 = n10779 ^ n9616 ^ n5055 ;
  assign n12268 = n12267 ^ n7906 ^ 1'b0 ;
  assign n12269 = ~n12266 & n12268 ;
  assign n12270 = ( ~n9531 & n11387 ) | ( ~n9531 & n12269 ) | ( n11387 & n12269 ) ;
  assign n12271 = n933 & ~n6171 ;
  assign n12272 = n12271 ^ n2962 ^ 1'b0 ;
  assign n12273 = x164 & ~n12272 ;
  assign n12274 = ~n2106 & n12273 ;
  assign n12275 = ~n4850 & n9627 ;
  assign n12276 = ( ~n5121 & n12274 ) | ( ~n5121 & n12275 ) | ( n12274 & n12275 ) ;
  assign n12279 = n9675 ^ n3406 ^ n1150 ;
  assign n12277 = n5669 ^ n3440 ^ n1433 ;
  assign n12278 = ( n4458 & ~n11791 ) | ( n4458 & n12277 ) | ( ~n11791 & n12277 ) ;
  assign n12280 = n12279 ^ n12278 ^ n4892 ;
  assign n12281 = n12280 ^ n10367 ^ 1'b0 ;
  assign n12282 = n6848 & n12281 ;
  assign n12283 = n2785 & n3261 ;
  assign n12284 = n12283 ^ n6111 ^ 1'b0 ;
  assign n12285 = n12284 ^ n2942 ^ 1'b0 ;
  assign n12286 = ( n2997 & n9101 ) | ( n2997 & ~n12285 ) | ( n9101 & ~n12285 ) ;
  assign n12287 = n7358 ^ n805 ^ 1'b0 ;
  assign n12288 = ~n7822 & n12287 ;
  assign n12289 = ( ~n6186 & n7494 ) | ( ~n6186 & n8865 ) | ( n7494 & n8865 ) ;
  assign n12290 = n994 | n12289 ;
  assign n12291 = ( ~n986 & n7384 ) | ( ~n986 & n8064 ) | ( n7384 & n8064 ) ;
  assign n12292 = ( n3793 & n6849 ) | ( n3793 & n12291 ) | ( n6849 & n12291 ) ;
  assign n12293 = n5746 & n12292 ;
  assign n12294 = ~n270 & n6250 ;
  assign n12295 = n2261 & n12294 ;
  assign n12296 = n12295 ^ n9658 ^ n5933 ;
  assign n12297 = n8319 ^ n7431 ^ x231 ;
  assign n12298 = n12297 ^ n8752 ^ n4403 ;
  assign n12299 = n11708 ^ n2434 ^ n1398 ;
  assign n12300 = n1044 & n6471 ;
  assign n12301 = n1465 & n10965 ;
  assign n12302 = n5720 ^ n4291 ^ n3003 ;
  assign n12303 = ( n10287 & n12301 ) | ( n10287 & n12302 ) | ( n12301 & n12302 ) ;
  assign n12304 = n5298 | n7206 ;
  assign n12305 = n3781 & ~n12304 ;
  assign n12306 = n12305 ^ n7638 ^ 1'b0 ;
  assign n12307 = ~n3335 & n12306 ;
  assign n12308 = n12307 ^ n2588 ^ 1'b0 ;
  assign n12309 = n12303 & n12308 ;
  assign n12310 = n3133 & ~n3755 ;
  assign n12311 = ( ~n4974 & n5687 ) | ( ~n4974 & n12310 ) | ( n5687 & n12310 ) ;
  assign n12312 = n3054 ^ n2536 ^ 1'b0 ;
  assign n12313 = n12312 ^ n9871 ^ n4714 ;
  assign n12314 = ~n2740 & n5051 ;
  assign n12315 = n12314 ^ n6846 ^ 1'b0 ;
  assign n12316 = n5541 ^ n4904 ^ 1'b0 ;
  assign n12317 = ( ~n3703 & n12315 ) | ( ~n3703 & n12316 ) | ( n12315 & n12316 ) ;
  assign n12318 = ( n12311 & ~n12313 ) | ( n12311 & n12317 ) | ( ~n12313 & n12317 ) ;
  assign n12319 = ( n3974 & ~n4556 ) | ( n3974 & n8139 ) | ( ~n4556 & n8139 ) ;
  assign n12320 = n4569 ^ n3612 ^ n2417 ;
  assign n12321 = n12188 ^ n10108 ^ n2644 ;
  assign n12327 = n3674 ^ n2124 ^ 1'b0 ;
  assign n12328 = n5172 & n12327 ;
  assign n12329 = n4752 | n12328 ;
  assign n12322 = n1814 & ~n7088 ;
  assign n12323 = n12322 ^ n4006 ^ 1'b0 ;
  assign n12324 = n12323 ^ n10709 ^ n3777 ;
  assign n12325 = n423 & n7626 ;
  assign n12326 = ( ~n9010 & n12324 ) | ( ~n9010 & n12325 ) | ( n12324 & n12325 ) ;
  assign n12330 = n12329 ^ n12326 ^ 1'b0 ;
  assign n12331 = ~n10181 & n12330 ;
  assign n12332 = n275 | n3575 ;
  assign n12333 = ~n7138 & n12332 ;
  assign n12334 = n3143 & n12333 ;
  assign n12335 = n12334 ^ n10377 ^ 1'b0 ;
  assign n12336 = n7924 & ~n12335 ;
  assign n12337 = ( ~n256 & n2750 ) | ( ~n256 & n3847 ) | ( n2750 & n3847 ) ;
  assign n12338 = ( n432 & n643 ) | ( n432 & n12337 ) | ( n643 & n12337 ) ;
  assign n12339 = n1444 | n2392 ;
  assign n12340 = n12339 ^ n7133 ^ 1'b0 ;
  assign n12341 = ( n416 & n11758 ) | ( n416 & n12340 ) | ( n11758 & n12340 ) ;
  assign n12342 = ~n12338 & n12341 ;
  assign n12344 = n1097 | n5723 ;
  assign n12343 = n4240 & n5737 ;
  assign n12345 = n12344 ^ n12343 ^ 1'b0 ;
  assign n12346 = n11666 ^ n6951 ^ 1'b0 ;
  assign n12347 = n2693 & ~n8366 ;
  assign n12348 = n12347 ^ n5245 ^ 1'b0 ;
  assign n12349 = n12346 & n12348 ;
  assign n12350 = ~n12345 & n12349 ;
  assign n12351 = n2272 ^ n745 ^ 1'b0 ;
  assign n12355 = n7079 ^ x116 ^ 1'b0 ;
  assign n12356 = ~n4375 & n12355 ;
  assign n12353 = n3467 & n6350 ;
  assign n12354 = ( ~n2138 & n6621 ) | ( ~n2138 & n12353 ) | ( n6621 & n12353 ) ;
  assign n12352 = n6773 & ~n8636 ;
  assign n12357 = n12356 ^ n12354 ^ n12352 ;
  assign n12358 = n5285 ^ n1245 ^ 1'b0 ;
  assign n12359 = n12358 ^ n9740 ^ n3142 ;
  assign n12360 = n545 & n4046 ;
  assign n12361 = n12360 ^ n5956 ^ n5825 ;
  assign n12364 = n5484 ^ n4437 ^ 1'b0 ;
  assign n12365 = n2777 | n12364 ;
  assign n12362 = n11570 ^ n7928 ^ 1'b0 ;
  assign n12363 = n12362 ^ n6525 ^ n742 ;
  assign n12366 = n12365 ^ n12363 ^ 1'b0 ;
  assign n12367 = n1311 & n2587 ;
  assign n12368 = n12367 ^ n9365 ^ 1'b0 ;
  assign n12370 = n7366 ^ n4109 ^ 1'b0 ;
  assign n12369 = n3863 & ~n4910 ;
  assign n12371 = n12370 ^ n12369 ^ 1'b0 ;
  assign n12372 = n12371 ^ n5176 ^ n3468 ;
  assign n12375 = ~n6897 & n9622 ;
  assign n12376 = n12375 ^ n4532 ^ 1'b0 ;
  assign n12377 = ( n8655 & n9871 ) | ( n8655 & ~n12376 ) | ( n9871 & ~n12376 ) ;
  assign n12373 = n3221 | n6301 ;
  assign n12374 = n12373 ^ n9682 ^ 1'b0 ;
  assign n12378 = n12377 ^ n12374 ^ 1'b0 ;
  assign n12379 = n901 | n2141 ;
  assign n12380 = n12379 ^ n11635 ^ n10602 ;
  assign n12381 = n12380 ^ n464 ^ 1'b0 ;
  assign n12382 = n350 & n12381 ;
  assign n12383 = n9672 ^ n2530 ^ 1'b0 ;
  assign n12384 = n7042 & n12383 ;
  assign n12385 = ( n3166 & ~n3749 ) | ( n3166 & n12384 ) | ( ~n3749 & n12384 ) ;
  assign n12386 = ( n8043 & n9437 ) | ( n8043 & n12385 ) | ( n9437 & n12385 ) ;
  assign n12387 = x110 & n3898 ;
  assign n12388 = ~x62 & n3081 ;
  assign n12389 = ~n1359 & n11845 ;
  assign n12390 = n7249 & n12389 ;
  assign n12391 = n12390 ^ n5097 ^ 1'b0 ;
  assign n12392 = n12388 | n12391 ;
  assign n12393 = n12392 ^ n1049 ^ 1'b0 ;
  assign n12394 = n1323 & n12393 ;
  assign n12395 = n12394 ^ n5516 ^ 1'b0 ;
  assign n12396 = ~n12387 & n12395 ;
  assign n12397 = ~n4061 & n4139 ;
  assign n12398 = ~n2696 & n12397 ;
  assign n12399 = n5153 & ~n12398 ;
  assign n12400 = n12399 ^ n10235 ^ 1'b0 ;
  assign n12401 = n4467 & n12400 ;
  assign n12402 = n2106 | n8334 ;
  assign n12403 = n6091 ^ n1895 ^ n1492 ;
  assign n12404 = n1625 & ~n11360 ;
  assign n12405 = n12403 & n12404 ;
  assign n12412 = n2739 ^ n1839 ^ n436 ;
  assign n12406 = n8740 | n12235 ;
  assign n12407 = n12406 ^ n8139 ^ 1'b0 ;
  assign n12408 = n5723 ^ n1627 ^ n1569 ;
  assign n12409 = n8733 ^ n4829 ^ n2864 ;
  assign n12410 = ~n12408 & n12409 ;
  assign n12411 = ~n12407 & n12410 ;
  assign n12413 = n12412 ^ n12411 ^ n1354 ;
  assign n12417 = n10464 ^ n6023 ^ n4416 ;
  assign n12416 = n9386 ^ n7727 ^ n5965 ;
  assign n12414 = ( n4307 & n5014 ) | ( n4307 & n7138 ) | ( n5014 & n7138 ) ;
  assign n12415 = n4433 & ~n12414 ;
  assign n12418 = n12417 ^ n12416 ^ n12415 ;
  assign n12435 = n7867 ^ n4761 ^ n2188 ;
  assign n12428 = n3986 & ~n4134 ;
  assign n12429 = ~n7477 & n12428 ;
  assign n12432 = ( n638 & n2025 ) | ( n638 & ~n3452 ) | ( n2025 & ~n3452 ) ;
  assign n12430 = n2295 & ~n7478 ;
  assign n12431 = n12430 ^ n11916 ^ n7588 ;
  assign n12433 = n12432 ^ n12431 ^ 1'b0 ;
  assign n12434 = n12429 | n12433 ;
  assign n12425 = ~n4291 & n4316 ;
  assign n12426 = n12425 ^ n6404 ^ 1'b0 ;
  assign n12419 = n3019 ^ n1284 ^ n419 ;
  assign n12420 = n395 & n4633 ;
  assign n12421 = n6956 ^ n962 ^ 1'b0 ;
  assign n12422 = n12420 & n12421 ;
  assign n12423 = ~n12419 & n12422 ;
  assign n12424 = ~n3110 & n12423 ;
  assign n12427 = n12426 ^ n12424 ^ 1'b0 ;
  assign n12436 = n12435 ^ n12434 ^ n12427 ;
  assign n12437 = ( n3532 & ~n3768 ) | ( n3532 & n6401 ) | ( ~n3768 & n6401 ) ;
  assign n12438 = n5362 & ~n7027 ;
  assign n12439 = n12438 ^ n12313 ^ n5437 ;
  assign n12440 = n1859 ^ n1302 ^ n759 ;
  assign n12441 = n12440 ^ n8915 ^ n3358 ;
  assign n12442 = n12441 ^ n10372 ^ n310 ;
  assign n12443 = n12442 ^ n11175 ^ n1487 ;
  assign n12445 = n3453 ^ n2495 ^ 1'b0 ;
  assign n12446 = n1214 & n12445 ;
  assign n12444 = n4851 | n8376 ;
  assign n12447 = n12446 ^ n12444 ^ 1'b0 ;
  assign n12448 = n12447 ^ n9464 ^ n1531 ;
  assign n12449 = n12161 ^ n2467 ^ n1421 ;
  assign n12450 = n5302 ^ n4375 ^ 1'b0 ;
  assign n12451 = ( n1680 & n6033 ) | ( n1680 & n11775 ) | ( n6033 & n11775 ) ;
  assign n12452 = n7116 | n12451 ;
  assign n12453 = n12450 & ~n12452 ;
  assign n12454 = n12416 ^ n2726 ^ 1'b0 ;
  assign n12455 = n12454 ^ n9319 ^ n2393 ;
  assign n12456 = ~n5730 & n6025 ;
  assign n12457 = n4922 | n12456 ;
  assign n12459 = x79 & ~n5704 ;
  assign n12460 = n3531 & n12459 ;
  assign n12461 = n12460 ^ n1776 ^ n499 ;
  assign n12462 = n2885 & ~n12461 ;
  assign n12463 = n8864 & n12462 ;
  assign n12458 = n2932 | n8987 ;
  assign n12464 = n12463 ^ n12458 ^ 1'b0 ;
  assign n12465 = ( ~n12455 & n12457 ) | ( ~n12455 & n12464 ) | ( n12457 & n12464 ) ;
  assign n12466 = ( n490 & n6876 ) | ( n490 & n8602 ) | ( n6876 & n8602 ) ;
  assign n12467 = n12466 ^ n7814 ^ 1'b0 ;
  assign n12468 = n5026 & n9247 ;
  assign n12469 = n12468 ^ n12052 ^ n320 ;
  assign n12470 = n1162 & ~n12469 ;
  assign n12471 = n4256 & ~n7089 ;
  assign n12472 = n8468 ^ n4983 ^ 1'b0 ;
  assign n12473 = ( n4086 & ~n12471 ) | ( n4086 & n12472 ) | ( ~n12471 & n12472 ) ;
  assign n12474 = ~n1438 & n6653 ;
  assign n12475 = ~x135 & n12474 ;
  assign n12476 = n12475 ^ n6960 ^ n3616 ;
  assign n12477 = n10222 ^ n3408 ^ 1'b0 ;
  assign n12478 = ~n8756 & n12477 ;
  assign n12479 = n12441 ^ n7590 ^ 1'b0 ;
  assign n12480 = ( n12476 & ~n12478 ) | ( n12476 & n12479 ) | ( ~n12478 & n12479 ) ;
  assign n12481 = ~n5797 & n10890 ;
  assign n12482 = ~x227 & x240 ;
  assign n12483 = ~n6528 & n12482 ;
  assign n12484 = n12483 ^ n3877 ^ 1'b0 ;
  assign n12485 = n2493 ^ n1942 ^ 1'b0 ;
  assign n12487 = ( n2978 & n6135 ) | ( n2978 & n8797 ) | ( n6135 & n8797 ) ;
  assign n12486 = n3840 & n4924 ;
  assign n12488 = n12487 ^ n12486 ^ n8942 ;
  assign n12489 = n8980 ^ n6200 ^ n707 ;
  assign n12490 = n12489 ^ n1637 ^ 1'b0 ;
  assign n12491 = n1993 & ~n12490 ;
  assign n12492 = n9761 ^ n4828 ^ 1'b0 ;
  assign n12493 = n8136 & n12492 ;
  assign n12500 = n5403 ^ n4325 ^ n575 ;
  assign n12494 = ( n582 & n3476 ) | ( n582 & ~n11859 ) | ( n3476 & ~n11859 ) ;
  assign n12495 = ( n9890 & n11666 ) | ( n9890 & n12494 ) | ( n11666 & n12494 ) ;
  assign n12496 = n3113 & ~n12495 ;
  assign n12497 = n12496 ^ n10270 ^ 1'b0 ;
  assign n12498 = ( n5838 & ~n10401 ) | ( n5838 & n12497 ) | ( ~n10401 & n12497 ) ;
  assign n12499 = ( n7042 & ~n7579 ) | ( n7042 & n12498 ) | ( ~n7579 & n12498 ) ;
  assign n12501 = n12500 ^ n12499 ^ n7022 ;
  assign n12502 = n3172 ^ x91 ^ 1'b0 ;
  assign n12503 = n10936 ^ n4421 ^ n1043 ;
  assign n12504 = ( n3579 & n4747 ) | ( n3579 & n6972 ) | ( n4747 & n6972 ) ;
  assign n12505 = n6146 ^ x126 ^ 1'b0 ;
  assign n12506 = n12504 & n12505 ;
  assign n12507 = ( n6483 & ~n12503 ) | ( n6483 & n12506 ) | ( ~n12503 & n12506 ) ;
  assign n12508 = ~n8449 & n11118 ;
  assign n12509 = n8965 ^ n6365 ^ n2316 ;
  assign n12511 = ( ~n471 & n925 ) | ( ~n471 & n6347 ) | ( n925 & n6347 ) ;
  assign n12512 = ( ~n5729 & n7674 ) | ( ~n5729 & n12511 ) | ( n7674 & n12511 ) ;
  assign n12513 = n10052 ^ n7238 ^ n2503 ;
  assign n12514 = n12513 ^ n6032 ^ n2120 ;
  assign n12515 = ( n9042 & n12512 ) | ( n9042 & ~n12514 ) | ( n12512 & ~n12514 ) ;
  assign n12510 = n343 & n1740 ;
  assign n12516 = n12515 ^ n12510 ^ n7155 ;
  assign n12517 = ( n11793 & n12509 ) | ( n11793 & ~n12516 ) | ( n12509 & ~n12516 ) ;
  assign n12518 = ( ~n9773 & n10370 ) | ( ~n9773 & n12238 ) | ( n10370 & n12238 ) ;
  assign n12519 = x24 & n4488 ;
  assign n12520 = ~n6314 & n12519 ;
  assign n12521 = n12520 ^ n4864 ^ n400 ;
  assign n12522 = ( n1236 & n2086 ) | ( n1236 & ~n12521 ) | ( n2086 & ~n12521 ) ;
  assign n12523 = ( ~n2784 & n3723 ) | ( ~n2784 & n8453 ) | ( n3723 & n8453 ) ;
  assign n12524 = n5134 | n12523 ;
  assign n12525 = n3731 & n12524 ;
  assign n12526 = x93 & n1045 ;
  assign n12527 = n12526 ^ n1096 ^ 1'b0 ;
  assign n12528 = ~n3786 & n8965 ;
  assign n12529 = n12527 & n12528 ;
  assign n12530 = n12529 ^ n4646 ^ n3869 ;
  assign n12531 = n5018 & n6293 ;
  assign n12532 = n12531 ^ n5544 ^ 1'b0 ;
  assign n12533 = ~n9070 & n12532 ;
  assign n12534 = n12533 ^ n2955 ^ 1'b0 ;
  assign n12535 = n8019 ^ n7842 ^ n6083 ;
  assign n12536 = n4538 & ~n11043 ;
  assign n12537 = ( ~n773 & n4553 ) | ( ~n773 & n5583 ) | ( n4553 & n5583 ) ;
  assign n12538 = n12537 ^ n8775 ^ n6171 ;
  assign n12539 = ( n1189 & ~n3783 ) | ( n1189 & n12538 ) | ( ~n3783 & n12538 ) ;
  assign n12543 = ( n2347 & n2551 ) | ( n2347 & n2563 ) | ( n2551 & n2563 ) ;
  assign n12544 = ( n2791 & n4000 ) | ( n2791 & n12543 ) | ( n4000 & n12543 ) ;
  assign n12540 = n11728 ^ n8649 ^ n4113 ;
  assign n12541 = ~n8899 & n12540 ;
  assign n12542 = ~n10749 & n12541 ;
  assign n12545 = n12544 ^ n12542 ^ 1'b0 ;
  assign n12546 = n8479 | n12545 ;
  assign n12547 = n1570 | n7188 ;
  assign n12548 = n12546 & ~n12547 ;
  assign n12549 = ~n630 & n5845 ;
  assign n12550 = n12549 ^ n12431 ^ n8644 ;
  assign n12552 = n5129 ^ n1845 ^ n1639 ;
  assign n12551 = ( n1500 & n4680 ) | ( n1500 & ~n10246 ) | ( n4680 & ~n10246 ) ;
  assign n12553 = n12552 ^ n12551 ^ n9727 ;
  assign n12554 = n12553 ^ n3552 ^ 1'b0 ;
  assign n12555 = n6092 & ~n12554 ;
  assign n12556 = ( ~n276 & n2348 ) | ( ~n276 & n3229 ) | ( n2348 & n3229 ) ;
  assign n12557 = n12556 ^ n4725 ^ n1863 ;
  assign n12558 = n3024 ^ n716 ^ 1'b0 ;
  assign n12559 = n12558 ^ n6911 ^ n3529 ;
  assign n12560 = n5967 | n12559 ;
  assign n12561 = n12560 ^ n2760 ^ 1'b0 ;
  assign n12562 = n12561 ^ n3595 ^ n549 ;
  assign n12563 = n12562 ^ n4022 ^ n2190 ;
  assign n12564 = ( n7855 & n12557 ) | ( n7855 & n12563 ) | ( n12557 & n12563 ) ;
  assign n12565 = n2649 & n12564 ;
  assign n12566 = n9357 ^ n4480 ^ 1'b0 ;
  assign n12568 = ( n2080 & ~n2135 ) | ( n2080 & n2780 ) | ( ~n2135 & n2780 ) ;
  assign n12569 = ~n7588 & n9635 ;
  assign n12570 = n12569 ^ n2686 ^ 1'b0 ;
  assign n12571 = n12568 & n12570 ;
  assign n12572 = n12571 ^ n8801 ^ 1'b0 ;
  assign n12573 = n12572 ^ n11205 ^ 1'b0 ;
  assign n12567 = n1518 & ~n6109 ;
  assign n12574 = n12573 ^ n12567 ^ 1'b0 ;
  assign n12575 = n2682 ^ n2250 ^ 1'b0 ;
  assign n12576 = n2210 & n12575 ;
  assign n12577 = ~n6266 & n7674 ;
  assign n12578 = ~n12576 & n12577 ;
  assign n12579 = n12578 ^ n900 ^ 1'b0 ;
  assign n12580 = ~n1138 & n9132 ;
  assign n12581 = n10892 ^ n5509 ^ 1'b0 ;
  assign n12582 = n5337 & ~n7224 ;
  assign n12583 = n12582 ^ n6255 ^ 1'b0 ;
  assign n12585 = ( ~n1026 & n1758 ) | ( ~n1026 & n2727 ) | ( n1758 & n2727 ) ;
  assign n12586 = n12585 ^ n2861 ^ n751 ;
  assign n12587 = ( ~n5093 & n9761 ) | ( ~n5093 & n10067 ) | ( n9761 & n10067 ) ;
  assign n12588 = n12586 & ~n12587 ;
  assign n12589 = ~n5828 & n12588 ;
  assign n12584 = n9765 ^ n7672 ^ n4522 ;
  assign n12590 = n12589 ^ n12584 ^ n9739 ;
  assign n12591 = ( ~x117 & n1236 ) | ( ~x117 & n1598 ) | ( n1236 & n1598 ) ;
  assign n12592 = ( n1122 & ~n2782 ) | ( n1122 & n12591 ) | ( ~n2782 & n12591 ) ;
  assign n12593 = ( n1401 & ~n11558 ) | ( n1401 & n12592 ) | ( ~n11558 & n12592 ) ;
  assign n12594 = ( n4184 & ~n5004 ) | ( n4184 & n9409 ) | ( ~n5004 & n9409 ) ;
  assign n12595 = n12594 ^ n9716 ^ n4931 ;
  assign n12596 = n6955 & n12595 ;
  assign n12597 = n4613 ^ x104 ^ 1'b0 ;
  assign n12598 = n6920 & n12597 ;
  assign n12599 = n4320 & n12598 ;
  assign n12600 = ( n1323 & ~n7314 ) | ( n1323 & n10362 ) | ( ~n7314 & n10362 ) ;
  assign n12601 = ( n859 & n3217 ) | ( n859 & n8826 ) | ( n3217 & n8826 ) ;
  assign n12602 = ( n801 & n12600 ) | ( n801 & n12601 ) | ( n12600 & n12601 ) ;
  assign n12603 = n12602 ^ n4698 ^ n981 ;
  assign n12604 = n12603 ^ n7419 ^ 1'b0 ;
  assign n12608 = n7346 ^ n6018 ^ n4570 ;
  assign n12609 = n5908 & ~n12608 ;
  assign n12605 = n786 | n1446 ;
  assign n12606 = n12605 ^ n5739 ^ n1121 ;
  assign n12607 = n12606 ^ n5830 ^ n3939 ;
  assign n12610 = n12609 ^ n12607 ^ n9154 ;
  assign n12611 = ~n3129 & n6520 ;
  assign n12612 = n1966 & n12611 ;
  assign n12613 = n12612 ^ n4674 ^ 1'b0 ;
  assign n12614 = n10850 | n12613 ;
  assign n12615 = x7 & n1246 ;
  assign n12616 = n12615 ^ n427 ^ 1'b0 ;
  assign n12617 = n4103 & n12616 ;
  assign n12618 = n10410 & n12617 ;
  assign n12619 = n12618 ^ x88 ^ 1'b0 ;
  assign n12620 = n558 & ~n12619 ;
  assign n12621 = n7345 ^ n2537 ^ n1775 ;
  assign n12622 = n7881 | n12621 ;
  assign n12623 = n10099 & ~n12622 ;
  assign n12624 = n2027 & n4051 ;
  assign n12625 = ( ~n2763 & n6763 ) | ( ~n2763 & n12624 ) | ( n6763 & n12624 ) ;
  assign n12626 = n11682 ^ n4885 ^ n4746 ;
  assign n12627 = n6097 ^ n2022 ^ 1'b0 ;
  assign n12628 = n11421 & n12627 ;
  assign n12629 = n5801 & ~n5844 ;
  assign n12630 = n4676 & n12629 ;
  assign n12631 = n12630 ^ n11051 ^ 1'b0 ;
  assign n12632 = n2308 ^ x63 ^ 1'b0 ;
  assign n12633 = n1452 | n12632 ;
  assign n12634 = ( ~n8466 & n12515 ) | ( ~n8466 & n12633 ) | ( n12515 & n12633 ) ;
  assign n12635 = ~n7895 & n12634 ;
  assign n12636 = n624 & n12635 ;
  assign n12637 = n5470 ^ n1297 ^ 1'b0 ;
  assign n12638 = n12637 ^ n5968 ^ n4542 ;
  assign n12639 = ( n7748 & n12636 ) | ( n7748 & n12638 ) | ( n12636 & n12638 ) ;
  assign n12640 = ( ~n1926 & n4402 ) | ( ~n1926 & n5792 ) | ( n4402 & n5792 ) ;
  assign n12641 = n4149 ^ n2350 ^ n1264 ;
  assign n12642 = x218 & ~n3209 ;
  assign n12643 = n12642 ^ n2666 ^ 1'b0 ;
  assign n12644 = ( n12640 & ~n12641 ) | ( n12640 & n12643 ) | ( ~n12641 & n12643 ) ;
  assign n12646 = n2627 & ~n4487 ;
  assign n12647 = n12646 ^ n469 ^ 1'b0 ;
  assign n12645 = n3592 & ~n10215 ;
  assign n12648 = n12647 ^ n12645 ^ 1'b0 ;
  assign n12649 = x125 & n10573 ;
  assign n12650 = n12649 ^ n4553 ^ 1'b0 ;
  assign n12651 = ( n536 & n767 ) | ( n536 & ~n12650 ) | ( n767 & ~n12650 ) ;
  assign n12654 = x132 & n5363 ;
  assign n12655 = n4618 | n6037 ;
  assign n12656 = n4312 | n12655 ;
  assign n12657 = n12654 & n12656 ;
  assign n12658 = ~n6314 & n12657 ;
  assign n12659 = n9304 ^ n6462 ^ x73 ;
  assign n12660 = n12658 & n12659 ;
  assign n12661 = x39 & ~n6086 ;
  assign n12662 = n7674 & n12661 ;
  assign n12663 = n12662 ^ n9589 ^ 1'b0 ;
  assign n12664 = n12660 | n12663 ;
  assign n12652 = n9437 ^ n4134 ^ n2002 ;
  assign n12653 = n3255 & n12652 ;
  assign n12665 = n12664 ^ n12653 ^ x194 ;
  assign n12670 = n11552 ^ n2771 ^ 1'b0 ;
  assign n12666 = n5781 ^ n4750 ^ 1'b0 ;
  assign n12667 = n2342 & ~n12666 ;
  assign n12668 = n12667 ^ n10986 ^ n4762 ;
  assign n12669 = ~n1561 & n12668 ;
  assign n12671 = n12670 ^ n12669 ^ 1'b0 ;
  assign n12673 = n8064 ^ n4315 ^ 1'b0 ;
  assign n12674 = ( n7085 & n9216 ) | ( n7085 & ~n12673 ) | ( n9216 & ~n12673 ) ;
  assign n12672 = n6921 & ~n7330 ;
  assign n12675 = n12674 ^ n12672 ^ 1'b0 ;
  assign n12676 = n10709 ^ n3938 ^ n2168 ;
  assign n12677 = ( n1043 & n1556 ) | ( n1043 & ~n2609 ) | ( n1556 & ~n2609 ) ;
  assign n12678 = ( n7102 & ~n12676 ) | ( n7102 & n12677 ) | ( ~n12676 & n12677 ) ;
  assign n12679 = n12678 ^ n9447 ^ n7478 ;
  assign n12680 = ( n5390 & ~n6148 ) | ( n5390 & n8558 ) | ( ~n6148 & n8558 ) ;
  assign n12681 = n1676 | n12680 ;
  assign n12682 = ( n7501 & ~n8079 ) | ( n7501 & n9196 ) | ( ~n8079 & n9196 ) ;
  assign n12683 = n3814 & n8409 ;
  assign n12684 = ( n12681 & n12682 ) | ( n12681 & ~n12683 ) | ( n12682 & ~n12683 ) ;
  assign n12685 = n12679 & n12684 ;
  assign n12686 = ( n1888 & n3626 ) | ( n1888 & ~n8691 ) | ( n3626 & ~n8691 ) ;
  assign n12687 = ( n4492 & n7539 ) | ( n4492 & ~n12686 ) | ( n7539 & ~n12686 ) ;
  assign n12693 = n4483 & n4505 ;
  assign n12694 = ~n6869 & n12693 ;
  assign n12695 = ( n1745 & ~n5856 ) | ( n1745 & n12694 ) | ( ~n5856 & n12694 ) ;
  assign n12688 = n1308 & ~n4349 ;
  assign n12689 = ~n6422 & n12688 ;
  assign n12690 = ~n12677 & n12689 ;
  assign n12691 = n12690 ^ n9523 ^ 1'b0 ;
  assign n12692 = n1994 & ~n12691 ;
  assign n12696 = n12695 ^ n12692 ^ 1'b0 ;
  assign n12697 = ( n5900 & n7118 ) | ( n5900 & ~n11667 ) | ( n7118 & ~n11667 ) ;
  assign n12698 = n12697 ^ n5066 ^ n1339 ;
  assign n12699 = n2623 ^ n602 ^ 1'b0 ;
  assign n12700 = n3475 & n12699 ;
  assign n12701 = n12700 ^ n3722 ^ n3240 ;
  assign n12702 = n9482 ^ n7129 ^ n4632 ;
  assign n12703 = n11956 & ~n12702 ;
  assign n12704 = n12701 & n12703 ;
  assign n12705 = n5092 & n7259 ;
  assign n12706 = n4829 & n5373 ;
  assign n12707 = ~n440 & n12706 ;
  assign n12708 = ~n938 & n8572 ;
  assign n12709 = n5126 | n5970 ;
  assign n12710 = n1337 ^ n386 ^ 1'b0 ;
  assign n12711 = n1528 | n2042 ;
  assign n12712 = n3867 & ~n12711 ;
  assign n12713 = n12710 & ~n12712 ;
  assign n12714 = n12713 ^ n4195 ^ 1'b0 ;
  assign n12715 = n11593 ^ n8302 ^ n5725 ;
  assign n12716 = ~n12714 & n12715 ;
  assign n12717 = n12709 & n12716 ;
  assign n12725 = n8792 ^ n6601 ^ 1'b0 ;
  assign n12726 = ~n1112 & n9645 ;
  assign n12727 = n12725 & n12726 ;
  assign n12728 = n5410 | n12727 ;
  assign n12729 = n2879 | n12728 ;
  assign n12722 = n3481 & ~n5411 ;
  assign n12718 = n9555 ^ n5041 ^ 1'b0 ;
  assign n12719 = n593 & ~n12718 ;
  assign n12720 = n9066 & n9936 ;
  assign n12721 = ~n12719 & n12720 ;
  assign n12723 = n12722 ^ n12721 ^ n2771 ;
  assign n12724 = ~n5034 & n12723 ;
  assign n12730 = n12729 ^ n12724 ^ 1'b0 ;
  assign n12731 = ( n5700 & n5911 ) | ( n5700 & ~n10802 ) | ( n5911 & ~n10802 ) ;
  assign n12732 = n5566 ^ n4662 ^ 1'b0 ;
  assign n12733 = ~n1343 & n12732 ;
  assign n12745 = n7982 ^ n5170 ^ 1'b0 ;
  assign n12746 = ~n4010 & n12745 ;
  assign n12734 = x159 & n971 ;
  assign n12735 = n10456 & n12734 ;
  assign n12736 = n1972 | n5253 ;
  assign n12737 = n8744 & ~n12736 ;
  assign n12740 = ~n7029 & n11995 ;
  assign n12738 = n1064 & n3213 ;
  assign n12739 = n1739 & n12738 ;
  assign n12741 = n12740 ^ n12739 ^ 1'b0 ;
  assign n12742 = ~n12737 & n12741 ;
  assign n12743 = ~n10152 & n12742 ;
  assign n12744 = n12735 & n12743 ;
  assign n12747 = n12746 ^ n12744 ^ n6915 ;
  assign n12750 = n11735 ^ n4220 ^ n3225 ;
  assign n12751 = n12750 ^ n9697 ^ n8797 ;
  assign n12748 = ( ~x218 & n4251 ) | ( ~x218 & n5834 ) | ( n4251 & n5834 ) ;
  assign n12749 = n7541 & ~n12748 ;
  assign n12752 = n12751 ^ n12749 ^ 1'b0 ;
  assign n12753 = ~n362 & n2653 ;
  assign n12754 = ( n876 & n9835 ) | ( n876 & n12753 ) | ( n9835 & n12753 ) ;
  assign n12755 = n12754 ^ n3969 ^ n2510 ;
  assign n12756 = ( ~n5047 & n6600 ) | ( ~n5047 & n12755 ) | ( n6600 & n12755 ) ;
  assign n12757 = ~n5923 & n9189 ;
  assign n12758 = n12757 ^ n9151 ^ 1'b0 ;
  assign n12759 = n10048 ^ n5373 ^ 1'b0 ;
  assign n12760 = n5553 ^ n5156 ^ 1'b0 ;
  assign n12761 = n5018 & ~n12760 ;
  assign n12762 = n4807 & ~n8220 ;
  assign n12763 = n12762 ^ n5640 ^ n2942 ;
  assign n12764 = n7298 & ~n11593 ;
  assign n12765 = n8944 ^ n6036 ^ 1'b0 ;
  assign n12766 = n1952 & n5297 ;
  assign n12767 = ( ~n1946 & n3703 ) | ( ~n1946 & n4365 ) | ( n3703 & n4365 ) ;
  assign n12768 = ( n5133 & n12766 ) | ( n5133 & n12767 ) | ( n12766 & n12767 ) ;
  assign n12769 = ( n12764 & n12765 ) | ( n12764 & n12768 ) | ( n12765 & n12768 ) ;
  assign n12770 = ( n432 & ~n4634 ) | ( n432 & n12769 ) | ( ~n4634 & n12769 ) ;
  assign n12771 = n10679 ^ n579 ^ 1'b0 ;
  assign n12772 = ~n7819 & n12771 ;
  assign n12773 = n12772 ^ n5950 ^ n4456 ;
  assign n12774 = ~n1614 & n5091 ;
  assign n12775 = n10395 ^ n7766 ^ n4307 ;
  assign n12776 = n4394 & n12420 ;
  assign n12777 = ~n12775 & n12776 ;
  assign n12778 = ( ~n1558 & n12598 ) | ( ~n1558 & n12777 ) | ( n12598 & n12777 ) ;
  assign n12779 = n797 & ~n9580 ;
  assign n12780 = n7672 ^ x195 ^ 1'b0 ;
  assign n12781 = n5401 | n12780 ;
  assign n12782 = n3449 & n5321 ;
  assign n12783 = n12782 ^ n12157 ^ 1'b0 ;
  assign n12784 = n12208 ^ n3369 ^ 1'b0 ;
  assign n12785 = n12783 | n12784 ;
  assign n12786 = n11638 ^ n9019 ^ n4340 ;
  assign n12787 = ( n564 & ~n9580 ) | ( n564 & n9767 ) | ( ~n9580 & n9767 ) ;
  assign n12788 = n12787 ^ n5469 ^ n2104 ;
  assign n12789 = n12788 ^ n3220 ^ 1'b0 ;
  assign n12790 = ~n12786 & n12789 ;
  assign n12791 = n9723 ^ n1783 ^ 1'b0 ;
  assign n12792 = ~n9258 & n12791 ;
  assign n12793 = ( n7510 & n9926 ) | ( n7510 & n10599 ) | ( n9926 & n10599 ) ;
  assign n12794 = n1527 & n3522 ;
  assign n12795 = n3348 ^ n2606 ^ n2149 ;
  assign n12796 = n12795 ^ n2394 ^ 1'b0 ;
  assign n12797 = ( n3417 & n4780 ) | ( n3417 & n7436 ) | ( n4780 & n7436 ) ;
  assign n12798 = ( ~x221 & n9177 ) | ( ~x221 & n12797 ) | ( n9177 & n12797 ) ;
  assign n12799 = ( n12794 & n12796 ) | ( n12794 & n12798 ) | ( n12796 & n12798 ) ;
  assign n12800 = n3230 & n10647 ;
  assign n12801 = n8806 & ~n12800 ;
  assign n12802 = ( ~n9083 & n12799 ) | ( ~n9083 & n12801 ) | ( n12799 & n12801 ) ;
  assign n12805 = ( n2670 & n3257 ) | ( n2670 & ~n10001 ) | ( n3257 & ~n10001 ) ;
  assign n12803 = ( n1411 & ~n3105 ) | ( n1411 & n8635 ) | ( ~n3105 & n8635 ) ;
  assign n12804 = n12803 ^ n3367 ^ n2592 ;
  assign n12806 = n12805 ^ n12804 ^ 1'b0 ;
  assign n12807 = n5881 & ~n12806 ;
  assign n12808 = n267 | n12807 ;
  assign n12809 = n2914 | n12808 ;
  assign n12810 = n1099 & n5420 ;
  assign n12811 = n12810 ^ n8026 ^ 1'b0 ;
  assign n12812 = n6364 | n11830 ;
  assign n12813 = ( n8451 & n12811 ) | ( n8451 & n12812 ) | ( n12811 & n12812 ) ;
  assign n12815 = x106 & ~n8507 ;
  assign n12816 = n12815 ^ n5791 ^ 1'b0 ;
  assign n12814 = n4532 | n5927 ;
  assign n12817 = n12816 ^ n12814 ^ n11546 ;
  assign n12818 = n12817 ^ n6006 ^ n1988 ;
  assign n12819 = ~n551 & n12818 ;
  assign n12820 = n12819 ^ n6334 ^ 1'b0 ;
  assign n12824 = ( ~n1994 & n9056 ) | ( ~n1994 & n9350 ) | ( n9056 & n9350 ) ;
  assign n12825 = n6646 & ~n12824 ;
  assign n12826 = n12825 ^ n5991 ^ n3256 ;
  assign n12821 = n3070 ^ n2244 ^ n1671 ;
  assign n12822 = n12821 ^ n9925 ^ 1'b0 ;
  assign n12823 = ~n12794 & n12822 ;
  assign n12827 = n12826 ^ n12823 ^ 1'b0 ;
  assign n12828 = n7501 & ~n12827 ;
  assign n12830 = n8774 ^ x88 ^ 1'b0 ;
  assign n12829 = ( n5027 & ~n8349 ) | ( n5027 & n8646 ) | ( ~n8349 & n8646 ) ;
  assign n12831 = n12830 ^ n12829 ^ n5895 ;
  assign n12832 = n2214 ^ n1246 ^ 1'b0 ;
  assign n12833 = n5617 & n6921 ;
  assign n12835 = ( n1713 & n2267 ) | ( n1713 & n2727 ) | ( n2267 & n2727 ) ;
  assign n12834 = n8445 ^ n1772 ^ x46 ;
  assign n12836 = n12835 ^ n12834 ^ 1'b0 ;
  assign n12837 = x128 & n12836 ;
  assign n12838 = ( n12832 & ~n12833 ) | ( n12832 & n12837 ) | ( ~n12833 & n12837 ) ;
  assign n12840 = n4403 ^ n4385 ^ n2040 ;
  assign n12839 = n5696 | n7994 ;
  assign n12841 = n12840 ^ n12839 ^ 1'b0 ;
  assign n12842 = n12841 ^ n11978 ^ 1'b0 ;
  assign n12843 = n8145 ^ n7692 ^ 1'b0 ;
  assign n12844 = n12843 ^ n12069 ^ n575 ;
  assign n12845 = n4015 & n12844 ;
  assign n12849 = n7597 ^ n5713 ^ n2115 ;
  assign n12850 = n12849 ^ n4768 ^ 1'b0 ;
  assign n12848 = n1716 | n5254 ;
  assign n12846 = n8015 & n11774 ;
  assign n12847 = n12846 ^ n8135 ^ 1'b0 ;
  assign n12851 = n12850 ^ n12848 ^ n12847 ;
  assign n12852 = n10049 ^ n2867 ^ n2474 ;
  assign n12858 = n9832 ^ n5618 ^ n2866 ;
  assign n12859 = n12858 ^ n7621 ^ n6887 ;
  assign n12860 = n12859 ^ n6292 ^ n1787 ;
  assign n12853 = n2547 & ~n12497 ;
  assign n12854 = ( ~n596 & n6873 ) | ( ~n596 & n9144 ) | ( n6873 & n9144 ) ;
  assign n12855 = n12854 ^ n6583 ^ n4478 ;
  assign n12856 = ( n614 & n12853 ) | ( n614 & ~n12855 ) | ( n12853 & ~n12855 ) ;
  assign n12857 = n12856 ^ x191 ^ 1'b0 ;
  assign n12861 = n12860 ^ n12857 ^ x155 ;
  assign n12862 = n12852 & n12861 ;
  assign n12863 = n12862 ^ n7646 ^ 1'b0 ;
  assign n12864 = n3470 ^ n3394 ^ 1'b0 ;
  assign n12865 = n5737 & ~n12864 ;
  assign n12867 = n4407 | n7306 ;
  assign n12868 = n12867 ^ n11954 ^ 1'b0 ;
  assign n12866 = n323 & n3935 ;
  assign n12869 = n12868 ^ n12866 ^ x1 ;
  assign n12870 = n4782 & ~n12869 ;
  assign n12871 = n12870 ^ n3925 ^ 1'b0 ;
  assign n12872 = n12870 & n12871 ;
  assign n12873 = ( ~n7430 & n12865 ) | ( ~n7430 & n12872 ) | ( n12865 & n12872 ) ;
  assign n12874 = n4622 & ~n6298 ;
  assign n12875 = ~n1330 & n12874 ;
  assign n12876 = ~n4277 & n11733 ;
  assign n12877 = n12875 & n12876 ;
  assign n12878 = n12877 ^ n1304 ^ 1'b0 ;
  assign n12879 = n12873 & n12878 ;
  assign n12884 = n3729 ^ n689 ^ 1'b0 ;
  assign n12882 = n909 ^ n734 ^ 1'b0 ;
  assign n12880 = n8158 ^ x126 ^ 1'b0 ;
  assign n12881 = n9491 | n12880 ;
  assign n12883 = n12882 ^ n12881 ^ n1772 ;
  assign n12885 = n12884 ^ n12883 ^ n3605 ;
  assign n12886 = n6940 ^ n4563 ^ n423 ;
  assign n12891 = n1653 & n3095 ;
  assign n12887 = n2111 ^ n1432 ^ 1'b0 ;
  assign n12888 = n12887 ^ n8431 ^ n3635 ;
  assign n12889 = n11101 & n12888 ;
  assign n12890 = ( n6211 & ~n8006 ) | ( n6211 & n12889 ) | ( ~n8006 & n12889 ) ;
  assign n12892 = n12891 ^ n12890 ^ n1020 ;
  assign n12896 = ( n4583 & n5317 ) | ( n4583 & ~n6139 ) | ( n5317 & ~n6139 ) ;
  assign n12897 = n2607 & ~n9292 ;
  assign n12898 = ( n686 & n916 ) | ( n686 & ~n5864 ) | ( n916 & ~n5864 ) ;
  assign n12899 = n6196 | n12898 ;
  assign n12900 = ( ~n8291 & n12897 ) | ( ~n8291 & n12899 ) | ( n12897 & n12899 ) ;
  assign n12901 = ~n12896 & n12900 ;
  assign n12902 = n12901 ^ n9801 ^ 1'b0 ;
  assign n12893 = ~x55 & n1745 ;
  assign n12894 = n4071 & n12893 ;
  assign n12895 = n4814 & ~n12894 ;
  assign n12903 = n12902 ^ n12895 ^ 1'b0 ;
  assign n12904 = n11407 ^ n6418 ^ n1305 ;
  assign n12910 = n4014 | n8316 ;
  assign n12911 = x241 & ~n8651 ;
  assign n12912 = ~n12910 & n12911 ;
  assign n12905 = ~n4216 & n8109 ;
  assign n12906 = n1657 & n12905 ;
  assign n12907 = n2676 ^ n1816 ^ 1'b0 ;
  assign n12908 = n10022 | n12907 ;
  assign n12909 = ( n4024 & n12906 ) | ( n4024 & ~n12908 ) | ( n12906 & ~n12908 ) ;
  assign n12913 = n12912 ^ n12909 ^ 1'b0 ;
  assign n12918 = n4866 ^ n2841 ^ 1'b0 ;
  assign n12919 = n4746 & n12918 ;
  assign n12916 = n11058 ^ n645 ^ 1'b0 ;
  assign n12914 = n8700 ^ n748 ^ 1'b0 ;
  assign n12915 = n12914 ^ n6275 ^ 1'b0 ;
  assign n12917 = n12916 ^ n12915 ^ n5258 ;
  assign n12920 = n12919 ^ n12917 ^ 1'b0 ;
  assign n12921 = n2265 ^ n2228 ^ 1'b0 ;
  assign n12922 = ~n8366 & n12921 ;
  assign n12923 = n11836 ^ n2204 ^ 1'b0 ;
  assign n12924 = n12923 ^ n1905 ^ 1'b0 ;
  assign n12925 = n2951 | n12924 ;
  assign n12926 = n6323 ^ n3959 ^ 1'b0 ;
  assign n12927 = n4905 & n12926 ;
  assign n12928 = n5085 & n12927 ;
  assign n12929 = n1141 | n2993 ;
  assign n12930 = ( x186 & n1164 ) | ( x186 & ~n1587 ) | ( n1164 & ~n1587 ) ;
  assign n12931 = ( n2809 & n5363 ) | ( n2809 & n5989 ) | ( n5363 & n5989 ) ;
  assign n12932 = ( n5883 & n12930 ) | ( n5883 & ~n12931 ) | ( n12930 & ~n12931 ) ;
  assign n12933 = n8007 | n12932 ;
  assign n12934 = n1362 & ~n12933 ;
  assign n12935 = ( n10930 & n12929 ) | ( n10930 & n12934 ) | ( n12929 & n12934 ) ;
  assign n12936 = n4351 | n12935 ;
  assign n12937 = n12532 ^ n1567 ^ 1'b0 ;
  assign n12938 = n2401 ^ n2212 ^ n331 ;
  assign n12939 = n12938 ^ n5375 ^ n572 ;
  assign n12940 = ( n775 & n7780 ) | ( n775 & n12939 ) | ( n7780 & n12939 ) ;
  assign n12941 = n12940 ^ n3497 ^ n2206 ;
  assign n12942 = n9319 & ~n10483 ;
  assign n12943 = n6653 ^ n3255 ^ 1'b0 ;
  assign n12944 = n12943 ^ n2887 ^ n2880 ;
  assign n12945 = n2498 & n4342 ;
  assign n12946 = ( n1141 & n2080 ) | ( n1141 & ~n5125 ) | ( n2080 & ~n5125 ) ;
  assign n12947 = n4310 ^ n783 ^ n504 ;
  assign n12948 = n12947 ^ n807 ^ 1'b0 ;
  assign n12949 = n12946 | n12948 ;
  assign n12950 = n7722 | n12949 ;
  assign n12951 = n10781 ^ n5349 ^ 1'b0 ;
  assign n12952 = n12951 ^ n8389 ^ n562 ;
  assign n12953 = n11513 ^ n1666 ^ 1'b0 ;
  assign n12954 = n10505 & ~n12953 ;
  assign n12956 = n6428 ^ n6179 ^ 1'b0 ;
  assign n12957 = n9486 | n12956 ;
  assign n12955 = n9170 & n12586 ;
  assign n12958 = n12957 ^ n12955 ^ n11430 ;
  assign n12959 = n10428 ^ n4259 ^ 1'b0 ;
  assign n12960 = n8307 ^ n6889 ^ n4782 ;
  assign n12961 = ( n1205 & n12959 ) | ( n1205 & n12960 ) | ( n12959 & n12960 ) ;
  assign n12962 = n12026 ^ n7350 ^ x125 ;
  assign n12963 = n8109 & n9167 ;
  assign n12964 = n12963 ^ n2104 ^ 1'b0 ;
  assign n12965 = n12964 ^ n4728 ^ n1738 ;
  assign n12966 = n10874 ^ n6868 ^ 1'b0 ;
  assign n12967 = n12965 & ~n12966 ;
  assign n12968 = n12967 ^ n3462 ^ 1'b0 ;
  assign n12969 = n7928 ^ n5294 ^ 1'b0 ;
  assign n12970 = n2855 & ~n12969 ;
  assign n12971 = n4489 ^ n2640 ^ n1318 ;
  assign n12972 = n8109 ^ n6450 ^ 1'b0 ;
  assign n12973 = n1158 | n3555 ;
  assign n12974 = n3148 & ~n12973 ;
  assign n12975 = ( n1723 & ~n2036 ) | ( n1723 & n5956 ) | ( ~n2036 & n5956 ) ;
  assign n12976 = ( ~n4602 & n12974 ) | ( ~n4602 & n12975 ) | ( n12974 & n12975 ) ;
  assign n12977 = n12976 ^ n5231 ^ 1'b0 ;
  assign n12978 = n12972 & ~n12977 ;
  assign n12979 = n12971 & n12978 ;
  assign n12980 = n12970 & n12979 ;
  assign n12982 = n3979 ^ n2575 ^ x157 ;
  assign n12983 = ( n3199 & n3259 ) | ( n3199 & ~n12982 ) | ( n3259 & ~n12982 ) ;
  assign n12981 = x76 & ~n11249 ;
  assign n12984 = n12983 ^ n12981 ^ 1'b0 ;
  assign n12985 = n12984 ^ n7579 ^ n2373 ;
  assign n12986 = ~n8648 & n12985 ;
  assign n12987 = n12980 & n12986 ;
  assign n12988 = n4774 | n7739 ;
  assign n12989 = ( n7042 & ~n7550 ) | ( n7042 & n12988 ) | ( ~n7550 & n12988 ) ;
  assign n12990 = n10229 | n12989 ;
  assign n12991 = n781 & n2701 ;
  assign n12992 = n5767 & ~n12991 ;
  assign n12993 = n12992 ^ n2610 ^ 1'b0 ;
  assign n12994 = ( n3884 & n8855 ) | ( n3884 & ~n12993 ) | ( n8855 & ~n12993 ) ;
  assign n12996 = n8493 ^ n1984 ^ 1'b0 ;
  assign n12995 = n7446 ^ n3878 ^ n3350 ;
  assign n12997 = n12996 ^ n12995 ^ n4508 ;
  assign n12999 = n7120 ^ n2986 ^ 1'b0 ;
  assign n12998 = n4702 ^ n4494 ^ n1930 ;
  assign n13000 = n12999 ^ n12998 ^ n5860 ;
  assign n13001 = ~n1880 & n7531 ;
  assign n13002 = n13001 ^ n4724 ^ 1'b0 ;
  assign n13003 = ( ~n7702 & n8111 ) | ( ~n7702 & n13002 ) | ( n8111 & n13002 ) ;
  assign n13006 = n9089 ^ n6907 ^ n3169 ;
  assign n13004 = n9136 ^ n4926 ^ n401 ;
  assign n13005 = n6102 & ~n13004 ;
  assign n13007 = n13006 ^ n13005 ^ n6105 ;
  assign n13008 = n4351 & n11719 ;
  assign n13009 = n13008 ^ n3043 ^ 1'b0 ;
  assign n13010 = n1542 & ~n10772 ;
  assign n13011 = n13010 ^ n6456 ^ n2514 ;
  assign n13012 = ( n7950 & ~n9418 ) | ( n7950 & n11670 ) | ( ~n9418 & n11670 ) ;
  assign n13013 = n10495 ^ n9206 ^ 1'b0 ;
  assign n13014 = n2943 & ~n13013 ;
  assign n13015 = x98 & ~n9845 ;
  assign n13016 = n13015 ^ n2409 ^ 1'b0 ;
  assign n13017 = n9262 & n11775 ;
  assign n13018 = n7989 ^ n7094 ^ 1'b0 ;
  assign n13019 = n12377 ^ n2607 ^ 1'b0 ;
  assign n13020 = ( n1632 & ~n2342 ) | ( n1632 & n3097 ) | ( ~n2342 & n3097 ) ;
  assign n13021 = n13020 ^ n1693 ^ n646 ;
  assign n13022 = n13021 ^ n8580 ^ n5310 ;
  assign n13023 = n9436 & ~n13022 ;
  assign n13024 = ~n8250 & n13023 ;
  assign n13026 = n2946 & n3025 ;
  assign n13027 = n1818 & n13026 ;
  assign n13025 = ( ~n602 & n2272 ) | ( ~n602 & n5026 ) | ( n2272 & n5026 ) ;
  assign n13028 = n13027 ^ n13025 ^ n266 ;
  assign n13029 = n5066 | n12014 ;
  assign n13030 = n12559 ^ n1863 ^ 1'b0 ;
  assign n13031 = n2259 & n13030 ;
  assign n13038 = ( x127 & n1445 ) | ( x127 & n4042 ) | ( n1445 & n4042 ) ;
  assign n13032 = n6723 ^ n1351 ^ 1'b0 ;
  assign n13033 = x99 & ~n13032 ;
  assign n13034 = ~n2143 & n13033 ;
  assign n13035 = n13034 ^ n7053 ^ 1'b0 ;
  assign n13036 = ~x174 & n7746 ;
  assign n13037 = n13035 & n13036 ;
  assign n13039 = n13038 ^ n13037 ^ 1'b0 ;
  assign n13040 = ~n13031 & n13039 ;
  assign n13041 = ~n6947 & n13040 ;
  assign n13042 = n891 | n6347 ;
  assign n13043 = n2006 ^ x117 ^ 1'b0 ;
  assign n13044 = n12299 & n13043 ;
  assign n13045 = ~n13042 & n13044 ;
  assign n13046 = n5782 ^ n3031 ^ 1'b0 ;
  assign n13047 = n13046 ^ n10004 ^ n2546 ;
  assign n13048 = ~n2885 & n8996 ;
  assign n13049 = n13048 ^ n8442 ^ n5939 ;
  assign n13050 = n13049 ^ n2906 ^ 1'b0 ;
  assign n13051 = n3951 | n13050 ;
  assign n13052 = ( n631 & n3257 ) | ( n631 & ~n9635 ) | ( n3257 & ~n9635 ) ;
  assign n13053 = ( ~n3233 & n9380 ) | ( ~n3233 & n13052 ) | ( n9380 & n13052 ) ;
  assign n13054 = ( x187 & n11308 ) | ( x187 & ~n13053 ) | ( n11308 & ~n13053 ) ;
  assign n13055 = ( n1830 & n3368 ) | ( n1830 & n10054 ) | ( n3368 & n10054 ) ;
  assign n13056 = n13055 ^ n5773 ^ n5347 ;
  assign n13057 = ( n6806 & n12570 ) | ( n6806 & n13056 ) | ( n12570 & n13056 ) ;
  assign n13058 = ( ~n279 & n4418 ) | ( ~n279 & n6702 ) | ( n4418 & n6702 ) ;
  assign n13059 = ( ~n3552 & n8522 ) | ( ~n3552 & n13058 ) | ( n8522 & n13058 ) ;
  assign n13060 = n5532 & ~n8979 ;
  assign n13061 = n13060 ^ n2937 ^ 1'b0 ;
  assign n13062 = n2761 & ~n5873 ;
  assign n13063 = n550 & n13062 ;
  assign n13064 = ( ~n662 & n12339 ) | ( ~n662 & n13063 ) | ( n12339 & n13063 ) ;
  assign n13065 = n13064 ^ x8 ^ 1'b0 ;
  assign n13066 = n13061 & ~n13065 ;
  assign n13067 = ( ~n5446 & n13059 ) | ( ~n5446 & n13066 ) | ( n13059 & n13066 ) ;
  assign n13071 = n6992 ^ n5956 ^ 1'b0 ;
  assign n13072 = n3655 & n13071 ;
  assign n13069 = n4128 ^ n1083 ^ 1'b0 ;
  assign n13070 = ( n3801 & n4653 ) | ( n3801 & n13069 ) | ( n4653 & n13069 ) ;
  assign n13073 = n13072 ^ n13070 ^ 1'b0 ;
  assign n13074 = n4451 & ~n13073 ;
  assign n13075 = ( x49 & n1787 ) | ( x49 & ~n5973 ) | ( n1787 & ~n5973 ) ;
  assign n13076 = n13075 ^ n5992 ^ 1'b0 ;
  assign n13077 = n13074 & ~n13076 ;
  assign n13068 = n8147 ^ n2209 ^ 1'b0 ;
  assign n13078 = n13077 ^ n13068 ^ n9059 ;
  assign n13080 = ~n4328 & n11204 ;
  assign n13079 = n4165 & ~n9303 ;
  assign n13081 = n13080 ^ n13079 ^ 1'b0 ;
  assign n13082 = n11635 ^ n7753 ^ 1'b0 ;
  assign n13083 = n7878 & ~n13082 ;
  assign n13084 = n3033 & n13083 ;
  assign n13085 = n505 & ~n9816 ;
  assign n13086 = n10450 ^ n10425 ^ 1'b0 ;
  assign n13087 = ~n13085 & n13086 ;
  assign n13094 = ( n5099 & n6247 ) | ( n5099 & n7539 ) | ( n6247 & n7539 ) ;
  assign n13088 = n2865 & n4533 ;
  assign n13089 = n807 | n3204 ;
  assign n13090 = n3013 & ~n13089 ;
  assign n13091 = n13090 ^ n5200 ^ 1'b0 ;
  assign n13092 = ~n13088 & n13091 ;
  assign n13093 = n13092 ^ n8274 ^ n4384 ;
  assign n13095 = n13094 ^ n13093 ^ 1'b0 ;
  assign n13097 = ~n2160 & n4027 ;
  assign n13098 = n12344 ^ n434 ^ 1'b0 ;
  assign n13099 = n13097 & ~n13098 ;
  assign n13100 = n13099 ^ n5648 ^ n1639 ;
  assign n13096 = n12412 ^ n3544 ^ 1'b0 ;
  assign n13101 = n13100 ^ n13096 ^ n10439 ;
  assign n13102 = ( n946 & n5290 ) | ( n946 & ~n8951 ) | ( n5290 & ~n8951 ) ;
  assign n13103 = ( ~n4322 & n6884 ) | ( ~n4322 & n10021 ) | ( n6884 & n10021 ) ;
  assign n13104 = n7253 & ~n13103 ;
  assign n13105 = ~n8817 & n13104 ;
  assign n13112 = ( n3739 & ~n5305 ) | ( n3739 & n11634 ) | ( ~n5305 & n11634 ) ;
  assign n13113 = n4083 ^ n704 ^ 1'b0 ;
  assign n13114 = n13113 ^ n7110 ^ n4906 ;
  assign n13115 = ( n594 & n13112 ) | ( n594 & ~n13114 ) | ( n13112 & ~n13114 ) ;
  assign n13110 = n3522 ^ n1449 ^ 1'b0 ;
  assign n13106 = n1153 & n1589 ;
  assign n13107 = n2560 & n13106 ;
  assign n13108 = n4076 | n8759 ;
  assign n13109 = n13107 & ~n13108 ;
  assign n13111 = n13110 ^ n13109 ^ n3656 ;
  assign n13116 = n13115 ^ n13111 ^ n9385 ;
  assign n13117 = ( ~x176 & n2376 ) | ( ~x176 & n2448 ) | ( n2376 & n2448 ) ;
  assign n13118 = n4428 | n13117 ;
  assign n13119 = n13118 ^ n2611 ^ 1'b0 ;
  assign n13122 = n8960 ^ n2232 ^ n1264 ;
  assign n13123 = n13122 ^ n1261 ^ 1'b0 ;
  assign n13120 = n2018 | n5160 ;
  assign n13121 = ( ~n4275 & n5314 ) | ( ~n4275 & n13120 ) | ( n5314 & n13120 ) ;
  assign n13124 = n13123 ^ n13121 ^ 1'b0 ;
  assign n13125 = n7855 ^ n4085 ^ 1'b0 ;
  assign n13126 = n12357 ^ n8489 ^ n6314 ;
  assign n13127 = n10139 ^ n2928 ^ n2541 ;
  assign n13128 = ( n6113 & n7219 ) | ( n6113 & n13127 ) | ( n7219 & n13127 ) ;
  assign n13129 = n7213 ^ n1376 ^ 1'b0 ;
  assign n13130 = x155 & ~n6084 ;
  assign n13136 = n567 & ~n2114 ;
  assign n13137 = n13136 ^ n1796 ^ 1'b0 ;
  assign n13138 = n13137 ^ n6097 ^ 1'b0 ;
  assign n13135 = n12431 ^ n10495 ^ n2076 ;
  assign n13131 = n8917 ^ n5364 ^ 1'b0 ;
  assign n13132 = n9944 ^ n6469 ^ n4234 ;
  assign n13133 = n13132 ^ n6769 ^ 1'b0 ;
  assign n13134 = ~n13131 & n13133 ;
  assign n13139 = n13138 ^ n13135 ^ n13134 ;
  assign n13146 = ( n943 & n2691 ) | ( n943 & n6146 ) | ( n2691 & n6146 ) ;
  assign n13140 = x3 & ~n10499 ;
  assign n13141 = n13140 ^ n1675 ^ 1'b0 ;
  assign n13142 = ( n1791 & n2755 ) | ( n1791 & n13141 ) | ( n2755 & n13141 ) ;
  assign n13143 = n1064 & n13142 ;
  assign n13144 = n13143 ^ n11763 ^ 1'b0 ;
  assign n13145 = n12243 & ~n13144 ;
  assign n13147 = n13146 ^ n13145 ^ 1'b0 ;
  assign n13148 = ~n6118 & n6170 ;
  assign n13149 = n8701 ^ n1527 ^ n436 ;
  assign n13150 = ( n3523 & n8177 ) | ( n3523 & ~n13149 ) | ( n8177 & ~n13149 ) ;
  assign n13151 = n13150 ^ n1826 ^ 1'b0 ;
  assign n13152 = ~n13148 & n13151 ;
  assign n13153 = n8164 ^ n6474 ^ n2571 ;
  assign n13154 = n4176 ^ n3016 ^ n2206 ;
  assign n13155 = n13154 ^ n1935 ^ 1'b0 ;
  assign n13158 = n5372 ^ n5303 ^ 1'b0 ;
  assign n13156 = n6855 ^ n2676 ^ 1'b0 ;
  assign n13157 = n13156 ^ n10668 ^ n10599 ;
  assign n13159 = n13158 ^ n13157 ^ n1138 ;
  assign n13160 = n13155 & n13159 ;
  assign n13161 = n13153 | n13160 ;
  assign n13162 = ~n4340 & n13161 ;
  assign n13163 = ~n13152 & n13162 ;
  assign n13164 = n4408 ^ n2800 ^ n638 ;
  assign n13165 = n5556 | n13164 ;
  assign n13167 = n1430 | n10504 ;
  assign n13166 = ( n752 & ~n1257 ) | ( n752 & n5277 ) | ( ~n1257 & n5277 ) ;
  assign n13168 = n13167 ^ n13166 ^ n2913 ;
  assign n13169 = n13165 | n13168 ;
  assign n13170 = n6373 ^ n1883 ^ 1'b0 ;
  assign n13171 = n595 & ~n13170 ;
  assign n13172 = n13171 ^ n1366 ^ 1'b0 ;
  assign n13173 = n8605 & ~n13172 ;
  assign n13174 = n13173 ^ n5776 ^ 1'b0 ;
  assign n13175 = ( n3351 & n4087 ) | ( n3351 & n4985 ) | ( n4087 & n4985 ) ;
  assign n13176 = ~n10888 & n13175 ;
  assign n13177 = ( ~n1937 & n7114 ) | ( ~n1937 & n13176 ) | ( n7114 & n13176 ) ;
  assign n13178 = n13177 ^ n6114 ^ 1'b0 ;
  assign n13179 = n2025 & ~n13178 ;
  assign n13183 = ( n2222 & n4293 ) | ( n2222 & n9534 ) | ( n4293 & n9534 ) ;
  assign n13180 = n3398 ^ n1399 ^ 1'b0 ;
  assign n13181 = n435 & n13180 ;
  assign n13182 = ~n4759 & n13181 ;
  assign n13184 = n13183 ^ n13182 ^ 1'b0 ;
  assign n13185 = n3863 & n9052 ;
  assign n13186 = n13185 ^ n5724 ^ 1'b0 ;
  assign n13187 = n2732 & n2988 ;
  assign n13188 = n13187 ^ n1665 ^ 1'b0 ;
  assign n13189 = n1373 | n5713 ;
  assign n13190 = n13189 ^ n4809 ^ 1'b0 ;
  assign n13191 = n13188 & n13190 ;
  assign n13192 = n13191 ^ n3472 ^ 1'b0 ;
  assign n13193 = n2561 ^ n746 ^ 1'b0 ;
  assign n13194 = n7030 & n13193 ;
  assign n13195 = n13194 ^ n4428 ^ n4285 ;
  assign n13196 = n13195 ^ n7379 ^ n3986 ;
  assign n13197 = ~n13192 & n13196 ;
  assign n13198 = n13197 ^ n300 ^ 1'b0 ;
  assign n13199 = n4654 & ~n7558 ;
  assign n13200 = n13199 ^ n8619 ^ n5217 ;
  assign n13201 = n10259 ^ n6248 ^ n1067 ;
  assign n13202 = ( n7362 & ~n9468 ) | ( n7362 & n9565 ) | ( ~n9468 & n9565 ) ;
  assign n13203 = ( n10589 & ~n13201 ) | ( n10589 & n13202 ) | ( ~n13201 & n13202 ) ;
  assign n13204 = n6608 ^ n5024 ^ n1780 ;
  assign n13205 = n13204 ^ n8323 ^ n818 ;
  assign n13206 = n5486 & ~n10753 ;
  assign n13207 = n13206 ^ n2549 ^ 1'b0 ;
  assign n13208 = n13207 ^ n5907 ^ n1108 ;
  assign n13209 = ( x139 & ~n6668 ) | ( x139 & n13208 ) | ( ~n6668 & n13208 ) ;
  assign n13210 = n10425 ^ n6716 ^ n3353 ;
  assign n13211 = n13210 ^ n3124 ^ n1759 ;
  assign n13213 = n545 & ~n3912 ;
  assign n13214 = ~x201 & n13213 ;
  assign n13215 = ( ~n7630 & n8073 ) | ( ~n7630 & n13214 ) | ( n8073 & n13214 ) ;
  assign n13212 = n5788 ^ n3536 ^ n1682 ;
  assign n13216 = n13215 ^ n13212 ^ n3707 ;
  assign n13217 = n13216 ^ n7547 ^ n4244 ;
  assign n13218 = n1217 & ~n2584 ;
  assign n13219 = n13218 ^ n11173 ^ 1'b0 ;
  assign n13220 = ( n534 & n11635 ) | ( n534 & n13219 ) | ( n11635 & n13219 ) ;
  assign n13221 = ( ~n2409 & n2667 ) | ( ~n2409 & n7019 ) | ( n2667 & n7019 ) ;
  assign n13222 = n2324 & n6007 ;
  assign n13223 = n13222 ^ n11536 ^ 1'b0 ;
  assign n13228 = n2522 ^ n1462 ^ 1'b0 ;
  assign n13229 = ~n4960 & n13228 ;
  assign n13230 = ( n3848 & ~n6431 ) | ( n3848 & n13229 ) | ( ~n6431 & n13229 ) ;
  assign n13231 = n1182 & n13230 ;
  assign n13232 = n13231 ^ n5339 ^ n5036 ;
  assign n13224 = n8455 | n12143 ;
  assign n13225 = ~n589 & n11618 ;
  assign n13226 = n5800 & n13225 ;
  assign n13227 = n13224 & n13226 ;
  assign n13233 = n13232 ^ n13227 ^ n12650 ;
  assign n13234 = n11686 ^ n1184 ^ 1'b0 ;
  assign n13235 = n13233 | n13234 ;
  assign n13236 = n12087 ^ n2947 ^ n2071 ;
  assign n13237 = ( n797 & ~n6661 ) | ( n797 & n9836 ) | ( ~n6661 & n9836 ) ;
  assign n13239 = n1376 ^ n1358 ^ 1'b0 ;
  assign n13240 = n1897 | n13239 ;
  assign n13241 = n13240 ^ n7973 ^ n4938 ;
  assign n13238 = n12505 ^ n7658 ^ n2263 ;
  assign n13242 = n13241 ^ n13238 ^ 1'b0 ;
  assign n13243 = n9130 ^ n4297 ^ 1'b0 ;
  assign n13244 = ( n3925 & n13002 ) | ( n3925 & ~n13243 ) | ( n13002 & ~n13243 ) ;
  assign n13245 = ~n7390 & n13244 ;
  assign n13247 = n1761 & ~n9724 ;
  assign n13246 = n1551 ^ n692 ^ 1'b0 ;
  assign n13248 = n13247 ^ n13246 ^ n3073 ;
  assign n13249 = n2706 & n6067 ;
  assign n13250 = n13249 ^ n13123 ^ n8795 ;
  assign n13251 = n5310 ^ n2928 ^ n725 ;
  assign n13252 = ( n1836 & ~n6628 ) | ( n1836 & n8407 ) | ( ~n6628 & n8407 ) ;
  assign n13253 = ( ~n1518 & n7197 ) | ( ~n1518 & n7286 ) | ( n7197 & n7286 ) ;
  assign n13254 = ( n3425 & ~n8995 ) | ( n3425 & n13253 ) | ( ~n8995 & n13253 ) ;
  assign n13255 = n13254 ^ n8123 ^ 1'b0 ;
  assign n13256 = n13252 & ~n13255 ;
  assign n13257 = n13132 ^ n3314 ^ n1746 ;
  assign n13258 = ( n7147 & ~n7482 ) | ( n7147 & n13257 ) | ( ~n7482 & n13257 ) ;
  assign n13259 = n13258 ^ n1241 ^ 1'b0 ;
  assign n13264 = n4834 ^ n2970 ^ 1'b0 ;
  assign n13263 = ( ~n5809 & n5823 ) | ( ~n5809 & n12591 ) | ( n5823 & n12591 ) ;
  assign n13260 = n1303 & ~n1825 ;
  assign n13261 = n3161 & n13260 ;
  assign n13262 = n13261 ^ n7521 ^ 1'b0 ;
  assign n13265 = n13264 ^ n13263 ^ n13262 ;
  assign n13266 = n8190 ^ n3573 ^ x14 ;
  assign n13267 = ( n7511 & n10242 ) | ( n7511 & ~n12422 ) | ( n10242 & ~n12422 ) ;
  assign n13268 = n11793 ^ n5938 ^ 1'b0 ;
  assign n13269 = n3613 & n10038 ;
  assign n13270 = n7805 & n13269 ;
  assign n13271 = n13270 ^ n2480 ^ 1'b0 ;
  assign n13272 = n6198 ^ n500 ^ 1'b0 ;
  assign n13273 = ( n708 & ~n4738 ) | ( n708 & n13272 ) | ( ~n4738 & n13272 ) ;
  assign n13274 = ( n1997 & n3479 ) | ( n1997 & n9206 ) | ( n3479 & n9206 ) ;
  assign n13276 = ~n1425 & n2631 ;
  assign n13277 = n1022 & n13276 ;
  assign n13275 = n2754 ^ n866 ^ 1'b0 ;
  assign n13278 = n13277 ^ n13275 ^ n12295 ;
  assign n13279 = ~n13274 & n13278 ;
  assign n13280 = ( n13271 & n13273 ) | ( n13271 & n13279 ) | ( n13273 & n13279 ) ;
  assign n13285 = ( n2594 & n5501 ) | ( n2594 & ~n8320 ) | ( n5501 & ~n8320 ) ;
  assign n13286 = n13285 ^ n3254 ^ n3070 ;
  assign n13287 = n4858 & ~n13286 ;
  assign n13281 = n2732 & ~n3195 ;
  assign n13282 = n13281 ^ n2269 ^ 1'b0 ;
  assign n13283 = n5239 | n13282 ;
  assign n13284 = n13283 ^ n8134 ^ 1'b0 ;
  assign n13288 = n13287 ^ n13284 ^ n1683 ;
  assign n13290 = n6585 | n7845 ;
  assign n13291 = ( ~n2066 & n8987 ) | ( ~n2066 & n13290 ) | ( n8987 & n13290 ) ;
  assign n13292 = n13291 ^ n4247 ^ n3821 ;
  assign n13289 = n10794 ^ n4464 ^ n2374 ;
  assign n13293 = n13292 ^ n13289 ^ n7005 ;
  assign n13294 = n10452 ^ n6162 ^ n5494 ;
  assign n13295 = n13294 ^ n405 ^ n260 ;
  assign n13297 = n1543 & n6365 ;
  assign n13298 = ~n1411 & n13297 ;
  assign n13299 = n2112 ^ n724 ^ 1'b0 ;
  assign n13300 = ( ~n10424 & n13298 ) | ( ~n10424 & n13299 ) | ( n13298 & n13299 ) ;
  assign n13296 = ( n5208 & ~n8654 ) | ( n5208 & n11755 ) | ( ~n8654 & n11755 ) ;
  assign n13301 = n13300 ^ n13296 ^ 1'b0 ;
  assign n13302 = n6976 | n13301 ;
  assign n13303 = ( ~n5133 & n12442 ) | ( ~n5133 & n13302 ) | ( n12442 & n13302 ) ;
  assign n13304 = n5522 | n13011 ;
  assign n13305 = x190 & ~n7097 ;
  assign n13306 = n6023 | n13305 ;
  assign n13307 = n11465 & ~n13306 ;
  assign n13308 = n11694 & n13307 ;
  assign n13309 = n10410 ^ n9240 ^ 1'b0 ;
  assign n13310 = n4734 & n6907 ;
  assign n13311 = ~n13309 & n13310 ;
  assign n13312 = n3457 & n3644 ;
  assign n13313 = ( n5079 & n9476 ) | ( n5079 & n9522 ) | ( n9476 & n9522 ) ;
  assign n13314 = ( ~n8409 & n12157 ) | ( ~n8409 & n13313 ) | ( n12157 & n13313 ) ;
  assign n13315 = n13312 | n13314 ;
  assign n13316 = n7714 ^ n3362 ^ 1'b0 ;
  assign n13319 = n7089 ^ n2035 ^ n959 ;
  assign n13317 = n4586 ^ n695 ^ x0 ;
  assign n13318 = n13317 ^ n10593 ^ 1'b0 ;
  assign n13320 = n13319 ^ n13318 ^ n7203 ;
  assign n13321 = n7136 ^ n523 ^ 1'b0 ;
  assign n13322 = ( n3409 & ~n5499 ) | ( n3409 & n13321 ) | ( ~n5499 & n13321 ) ;
  assign n13323 = ( ~n2511 & n7360 ) | ( ~n2511 & n9126 ) | ( n7360 & n9126 ) ;
  assign n13324 = n3294 & ~n5527 ;
  assign n13325 = n13324 ^ n9101 ^ n953 ;
  assign n13327 = n2700 | n11627 ;
  assign n13328 = n7463 & ~n13327 ;
  assign n13329 = ~n924 & n13328 ;
  assign n13330 = n13329 ^ n9144 ^ 1'b0 ;
  assign n13331 = n13330 ^ n9928 ^ 1'b0 ;
  assign n13332 = n2417 & n13331 ;
  assign n13333 = n13332 ^ n6222 ^ n5166 ;
  assign n13326 = n3899 | n10880 ;
  assign n13334 = n13333 ^ n13326 ^ 1'b0 ;
  assign n13335 = n10124 ^ n2127 ^ 1'b0 ;
  assign n13336 = n10258 ^ n6693 ^ n1701 ;
  assign n13337 = n13336 ^ n3503 ^ n2187 ;
  assign n13338 = ( ~n3435 & n13093 ) | ( ~n3435 & n13337 ) | ( n13093 & n13337 ) ;
  assign n13340 = n9677 ^ n8507 ^ n4257 ;
  assign n13339 = n6720 & ~n12304 ;
  assign n13341 = n13340 ^ n13339 ^ 1'b0 ;
  assign n13342 = n12297 | n12964 ;
  assign n13343 = ( n3453 & ~n11954 ) | ( n3453 & n12112 ) | ( ~n11954 & n12112 ) ;
  assign n13344 = n12883 ^ n4196 ^ 1'b0 ;
  assign n13345 = ~n1826 & n2641 ;
  assign n13346 = ( n10501 & n11603 ) | ( n10501 & ~n13345 ) | ( n11603 & ~n13345 ) ;
  assign n13347 = n5662 & ~n8301 ;
  assign n13348 = n13277 ^ n7219 ^ n4350 ;
  assign n13349 = n13348 ^ n11819 ^ 1'b0 ;
  assign n13350 = n13347 | n13349 ;
  assign n13351 = n2008 ^ n1041 ^ 1'b0 ;
  assign n13352 = n12606 & ~n13351 ;
  assign n13353 = ( ~n6869 & n9802 ) | ( ~n6869 & n10656 ) | ( n9802 & n10656 ) ;
  assign n13354 = n1359 | n13353 ;
  assign n13355 = ~n13352 & n13354 ;
  assign n13356 = n5599 ^ n3678 ^ 1'b0 ;
  assign n13357 = n1519 ^ n1399 ^ 1'b0 ;
  assign n13358 = n11716 & n13357 ;
  assign n13359 = n894 & n13358 ;
  assign n13360 = ~n5522 & n13359 ;
  assign n13361 = ( ~n10669 & n13356 ) | ( ~n10669 & n13360 ) | ( n13356 & n13360 ) ;
  assign n13362 = n2828 | n9924 ;
  assign n13363 = n13362 ^ n9208 ^ 1'b0 ;
  assign n13364 = n13363 ^ n13033 ^ n385 ;
  assign n13365 = n3450 ^ n2402 ^ 1'b0 ;
  assign n13366 = n2623 & ~n13365 ;
  assign n13367 = ( n4989 & n9694 ) | ( n4989 & ~n13366 ) | ( n9694 & ~n13366 ) ;
  assign n13368 = ( n9530 & n13364 ) | ( n9530 & ~n13367 ) | ( n13364 & ~n13367 ) ;
  assign n13369 = n13368 ^ n13358 ^ 1'b0 ;
  assign n13370 = n10828 & n13369 ;
  assign n13372 = n1349 ^ n387 ^ x154 ;
  assign n13371 = ~n1505 & n7201 ;
  assign n13373 = n13372 ^ n13371 ^ x250 ;
  assign n13374 = ( n2652 & ~n7217 ) | ( n2652 & n12766 ) | ( ~n7217 & n12766 ) ;
  assign n13375 = x49 & n1851 ;
  assign n13376 = ~n13374 & n13375 ;
  assign n13377 = ( ~n362 & n1045 ) | ( ~n362 & n6244 ) | ( n1045 & n6244 ) ;
  assign n13378 = n1274 | n4956 ;
  assign n13379 = n1007 & ~n13378 ;
  assign n13380 = ( n3793 & n13377 ) | ( n3793 & n13379 ) | ( n13377 & n13379 ) ;
  assign n13381 = n11240 ^ n1770 ^ 1'b0 ;
  assign n13382 = n13113 ^ n5711 ^ 1'b0 ;
  assign n13383 = n10481 ^ n7378 ^ 1'b0 ;
  assign n13384 = ~n11959 & n13383 ;
  assign n13388 = n2226 & n9125 ;
  assign n13389 = n5087 & ~n13388 ;
  assign n13390 = n5266 & n13389 ;
  assign n13385 = n12461 ^ n7596 ^ n3608 ;
  assign n13386 = n13385 ^ n7122 ^ 1'b0 ;
  assign n13387 = n5229 & n13386 ;
  assign n13391 = n13390 ^ n13387 ^ n10499 ;
  assign n13392 = n10344 | n11533 ;
  assign n13393 = n13392 ^ n573 ^ 1'b0 ;
  assign n13394 = n2355 | n2613 ;
  assign n13396 = n3113 | n6146 ;
  assign n13395 = n4825 & n9655 ;
  assign n13397 = n13396 ^ n13395 ^ 1'b0 ;
  assign n13398 = ( n950 & n13394 ) | ( n950 & n13397 ) | ( n13394 & n13397 ) ;
  assign n13403 = n599 & n895 ;
  assign n13404 = ~n8785 & n13403 ;
  assign n13399 = n1706 & n7931 ;
  assign n13400 = n7723 ^ n2325 ^ n1909 ;
  assign n13401 = n13399 | n13400 ;
  assign n13402 = n5251 & ~n13401 ;
  assign n13405 = n13404 ^ n13402 ^ n9491 ;
  assign n13406 = n8206 & ~n12344 ;
  assign n13407 = n13406 ^ n5054 ^ n3590 ;
  assign n13412 = n4495 & ~n8939 ;
  assign n13413 = ~n6592 & n13412 ;
  assign n13408 = n6169 ^ n2285 ^ 1'b0 ;
  assign n13409 = n13408 ^ n9040 ^ 1'b0 ;
  assign n13410 = n7038 & ~n13409 ;
  assign n13411 = n13410 ^ n12486 ^ x196 ;
  assign n13414 = n13413 ^ n13411 ^ 1'b0 ;
  assign n13415 = n11429 ^ n8007 ^ 1'b0 ;
  assign n13416 = n489 & ~n3658 ;
  assign n13417 = ~n489 & n13416 ;
  assign n13418 = x128 & n5284 ;
  assign n13419 = ~n9434 & n13418 ;
  assign n13420 = n13417 | n13419 ;
  assign n13421 = n13417 & ~n13420 ;
  assign n13422 = ( x195 & ~n2128 ) | ( x195 & n6581 ) | ( ~n2128 & n6581 ) ;
  assign n13423 = ( ~n684 & n3785 ) | ( ~n684 & n13422 ) | ( n3785 & n13422 ) ;
  assign n13424 = n13423 ^ n10415 ^ 1'b0 ;
  assign n13425 = ~n2965 & n6647 ;
  assign n13426 = ~n3675 & n13425 ;
  assign n13427 = n4524 | n7244 ;
  assign n13428 = ~n13426 & n13427 ;
  assign n13429 = n5653 ^ n5651 ^ 1'b0 ;
  assign n13430 = ~n4365 & n8907 ;
  assign n13431 = n5804 | n13430 ;
  assign n13432 = n13431 ^ n4055 ^ 1'b0 ;
  assign n13433 = ( n11805 & ~n13429 ) | ( n11805 & n13432 ) | ( ~n13429 & n13432 ) ;
  assign n13434 = n10996 ^ n4747 ^ 1'b0 ;
  assign n13435 = n8900 & n13434 ;
  assign n13436 = ( n1990 & ~n7566 ) | ( n1990 & n7849 ) | ( ~n7566 & n7849 ) ;
  assign n13437 = ( ~n1093 & n3466 ) | ( ~n1093 & n13436 ) | ( n3466 & n13436 ) ;
  assign n13438 = ( ~n6180 & n6500 ) | ( ~n6180 & n10559 ) | ( n6500 & n10559 ) ;
  assign n13439 = n3871 ^ n3217 ^ 1'b0 ;
  assign n13440 = n2224 | n13439 ;
  assign n13441 = n13440 ^ n11672 ^ n10844 ;
  assign n13442 = ( ~n2898 & n3968 ) | ( ~n2898 & n5305 ) | ( n3968 & n5305 ) ;
  assign n13443 = n13442 ^ n4012 ^ 1'b0 ;
  assign n13444 = n10468 & n13443 ;
  assign n13445 = n12954 & n13444 ;
  assign n13446 = n13445 ^ n7049 ^ 1'b0 ;
  assign n13447 = n13165 ^ n8537 ^ n7099 ;
  assign n13448 = n13447 ^ n11633 ^ n11461 ;
  assign n13449 = n1537 & ~n5522 ;
  assign n13450 = ~x31 & n13449 ;
  assign n13451 = n13450 ^ n10297 ^ 1'b0 ;
  assign n13452 = ( n636 & n692 ) | ( n636 & n2970 ) | ( n692 & n2970 ) ;
  assign n13453 = n13452 ^ n6718 ^ 1'b0 ;
  assign n13454 = n6070 & n6532 ;
  assign n13455 = n13454 ^ n2883 ^ 1'b0 ;
  assign n13456 = ( n273 & n1197 ) | ( n273 & n9363 ) | ( n1197 & n9363 ) ;
  assign n13457 = n4385 & ~n13456 ;
  assign n13458 = n3746 & n13457 ;
  assign n13459 = ~n4123 & n4929 ;
  assign n13460 = n13458 & n13459 ;
  assign n13467 = n4756 & ~n10475 ;
  assign n13468 = ~n8019 & n13467 ;
  assign n13461 = ( ~n1798 & n1897 ) | ( ~n1798 & n4079 ) | ( n1897 & n4079 ) ;
  assign n13462 = n2330 & n6683 ;
  assign n13463 = x113 & n9739 ;
  assign n13464 = n13463 ^ n6950 ^ 1'b0 ;
  assign n13465 = ( ~n13461 & n13462 ) | ( ~n13461 & n13464 ) | ( n13462 & n13464 ) ;
  assign n13466 = n5007 & n13465 ;
  assign n13469 = n13468 ^ n13466 ^ 1'b0 ;
  assign n13470 = n13469 ^ n4239 ^ 1'b0 ;
  assign n13471 = n1791 ^ n1743 ^ 1'b0 ;
  assign n13472 = ~n5076 & n13471 ;
  assign n13473 = ( n1646 & ~n5521 ) | ( n1646 & n13472 ) | ( ~n5521 & n13472 ) ;
  assign n13478 = ~n1439 & n6285 ;
  assign n13476 = ( ~n948 & n8595 ) | ( ~n948 & n10284 ) | ( n8595 & n10284 ) ;
  assign n13477 = n6959 | n13476 ;
  assign n13479 = n13478 ^ n13477 ^ 1'b0 ;
  assign n13474 = n412 & n10617 ;
  assign n13475 = n13474 ^ n3365 ^ 1'b0 ;
  assign n13480 = n13479 ^ n13475 ^ n13058 ;
  assign n13481 = ( n3480 & n3896 ) | ( n3480 & ~n13480 ) | ( n3896 & ~n13480 ) ;
  assign n13482 = n4869 & n5221 ;
  assign n13483 = ( n10737 & n11771 ) | ( n10737 & n12640 ) | ( n11771 & n12640 ) ;
  assign n13484 = ( n2255 & n2680 ) | ( n2255 & ~n10744 ) | ( n2680 & ~n10744 ) ;
  assign n13485 = ~n6802 & n13484 ;
  assign n13486 = n13485 ^ n5686 ^ 1'b0 ;
  assign n13487 = n13486 ^ n6327 ^ 1'b0 ;
  assign n13488 = n6246 & n7990 ;
  assign n13489 = n13488 ^ n3756 ^ 1'b0 ;
  assign n13490 = ( n4697 & ~n12399 ) | ( n4697 & n13489 ) | ( ~n12399 & n13489 ) ;
  assign n13491 = n9538 ^ n5637 ^ 1'b0 ;
  assign n13492 = n10029 & n13491 ;
  assign n13493 = n13492 ^ n2103 ^ n492 ;
  assign n13494 = ( n8472 & ~n13490 ) | ( n8472 & n13493 ) | ( ~n13490 & n13493 ) ;
  assign n13495 = ( n329 & ~n2022 ) | ( n329 & n2748 ) | ( ~n2022 & n2748 ) ;
  assign n13496 = n13495 ^ n6802 ^ n4785 ;
  assign n13505 = n12475 ^ n7189 ^ 1'b0 ;
  assign n13500 = n3927 ^ n2863 ^ 1'b0 ;
  assign n13501 = n1004 & n13500 ;
  assign n13502 = n13501 ^ n2425 ^ 1'b0 ;
  assign n13497 = n3052 ^ n2809 ^ n2765 ;
  assign n13498 = n1659 & n13497 ;
  assign n13499 = n13498 ^ n5589 ^ 1'b0 ;
  assign n13503 = n13502 ^ n13499 ^ 1'b0 ;
  assign n13504 = n5355 & n13503 ;
  assign n13506 = n13505 ^ n13504 ^ 1'b0 ;
  assign n13507 = n7907 & n13506 ;
  assign n13508 = n13507 ^ n10081 ^ 1'b0 ;
  assign n13509 = n13508 ^ n4816 ^ n3531 ;
  assign n13510 = n13509 ^ n5776 ^ n1192 ;
  assign n13511 = n7915 ^ n1028 ^ 1'b0 ;
  assign n13512 = n5873 | n13511 ;
  assign n13513 = ( n9223 & n12974 ) | ( n9223 & n13512 ) | ( n12974 & n13512 ) ;
  assign n13514 = n13513 ^ n2018 ^ 1'b0 ;
  assign n13515 = n6450 & n13514 ;
  assign n13516 = n6007 & n13515 ;
  assign n13517 = n13516 ^ n8748 ^ 1'b0 ;
  assign n13518 = n9832 ^ x240 ^ 1'b0 ;
  assign n13519 = n11715 & ~n13518 ;
  assign n13520 = n2976 ^ n2280 ^ 1'b0 ;
  assign n13521 = ~n2607 & n13520 ;
  assign n13522 = ( n7696 & n11249 ) | ( n7696 & n13521 ) | ( n11249 & n13521 ) ;
  assign n13523 = n3448 | n13522 ;
  assign n13524 = n2711 & n13523 ;
  assign n13525 = ~n13519 & n13524 ;
  assign n13526 = n13525 ^ n10533 ^ n3523 ;
  assign n13527 = n5910 & n7671 ;
  assign n13528 = n12667 & n13527 ;
  assign n13529 = n2506 | n13528 ;
  assign n13530 = n5580 | n13529 ;
  assign n13531 = n13530 ^ x188 ^ 1'b0 ;
  assign n13532 = n13531 ^ n8380 ^ 1'b0 ;
  assign n13539 = n12441 ^ n11494 ^ n2666 ;
  assign n13533 = n4625 ^ n3398 ^ 1'b0 ;
  assign n13534 = n5353 | n13533 ;
  assign n13535 = ( n2639 & ~n3294 ) | ( n2639 & n4627 ) | ( ~n3294 & n4627 ) ;
  assign n13536 = n5472 | n13535 ;
  assign n13537 = n13534 & ~n13536 ;
  assign n13538 = n13537 ^ n8903 ^ n4651 ;
  assign n13540 = n13539 ^ n13538 ^ 1'b0 ;
  assign n13541 = ~n1643 & n5522 ;
  assign n13542 = n3591 | n6925 ;
  assign n13543 = n13542 ^ n2843 ^ 1'b0 ;
  assign n13544 = ~n547 & n13543 ;
  assign n13545 = n13544 ^ n6005 ^ 1'b0 ;
  assign n13546 = n2903 & n4824 ;
  assign n13547 = ( n6622 & n12833 ) | ( n6622 & n13546 ) | ( n12833 & n13546 ) ;
  assign n13548 = n5026 ^ n2481 ^ 1'b0 ;
  assign n13549 = n4848 & ~n13548 ;
  assign n13550 = n368 & n5595 ;
  assign n13551 = ~n7598 & n13550 ;
  assign n13552 = n1969 & ~n9635 ;
  assign n13553 = n7504 | n13552 ;
  assign n13554 = n13553 ^ n1697 ^ 1'b0 ;
  assign n13562 = n6004 ^ n1154 ^ 1'b0 ;
  assign n13563 = x186 & n13562 ;
  assign n13561 = n3006 | n5372 ;
  assign n13564 = n13563 ^ n13561 ^ 1'b0 ;
  assign n13559 = n3997 ^ n2695 ^ n1815 ;
  assign n13555 = n2806 | n5340 ;
  assign n13556 = n2987 & n13555 ;
  assign n13557 = n2434 & n13556 ;
  assign n13558 = ( n8198 & n9491 ) | ( n8198 & n13557 ) | ( n9491 & n13557 ) ;
  assign n13560 = n13559 ^ n13558 ^ 1'b0 ;
  assign n13565 = n13564 ^ n13560 ^ n8955 ;
  assign n13567 = n3522 ^ n308 ^ 1'b0 ;
  assign n13566 = n8284 ^ n2900 ^ n1431 ;
  assign n13568 = n13567 ^ n13566 ^ n5516 ;
  assign n13569 = n13568 ^ n4489 ^ x111 ;
  assign n13570 = n5695 ^ n4011 ^ n787 ;
  assign n13571 = n1885 & n13570 ;
  assign n13572 = n13571 ^ n8531 ^ 1'b0 ;
  assign n13573 = n7008 ^ n2350 ^ 1'b0 ;
  assign n13574 = n11655 | n13573 ;
  assign n13575 = n12148 ^ n2751 ^ 1'b0 ;
  assign n13576 = n3750 & n13575 ;
  assign n13577 = ( n1431 & n13574 ) | ( n1431 & ~n13576 ) | ( n13574 & ~n13576 ) ;
  assign n13594 = n12219 ^ n7277 ^ n2384 ;
  assign n13578 = n8007 ^ n5222 ^ n3339 ;
  assign n13580 = ~n1924 & n5253 ;
  assign n13579 = n3484 & ~n3992 ;
  assign n13581 = n13580 ^ n13579 ^ 1'b0 ;
  assign n13589 = n12328 ^ n2737 ^ n2138 ;
  assign n13582 = x113 & n4430 ;
  assign n13583 = n890 & n13582 ;
  assign n13584 = n13583 ^ n3655 ^ n666 ;
  assign n13585 = x159 & n13584 ;
  assign n13586 = n13585 ^ n2365 ^ 1'b0 ;
  assign n13587 = ( n2546 & n2584 ) | ( n2546 & n13586 ) | ( n2584 & n13586 ) ;
  assign n13588 = n9555 & n13587 ;
  assign n13590 = n13589 ^ n13588 ^ 1'b0 ;
  assign n13591 = n13590 ^ n3470 ^ n1971 ;
  assign n13592 = n13581 | n13591 ;
  assign n13593 = n13578 | n13592 ;
  assign n13595 = n13594 ^ n13593 ^ 1'b0 ;
  assign n13596 = ( n1032 & n2691 ) | ( n1032 & ~n3303 ) | ( n2691 & ~n3303 ) ;
  assign n13597 = n3214 & n13596 ;
  assign n13598 = ~n1258 & n5071 ;
  assign n13599 = n7317 & n13598 ;
  assign n13600 = n13599 ^ n11737 ^ 1'b0 ;
  assign n13601 = n12844 & ~n13600 ;
  assign n13602 = n2594 & ~n7588 ;
  assign n13603 = ~n1198 & n13602 ;
  assign n13604 = ( ~n1609 & n9742 ) | ( ~n1609 & n13603 ) | ( n9742 & n13603 ) ;
  assign n13607 = n5092 & n5646 ;
  assign n13608 = n1802 & n13607 ;
  assign n13609 = n13608 ^ n4403 ^ 1'b0 ;
  assign n13605 = n1004 & ~n3774 ;
  assign n13606 = n13605 ^ n6385 ^ 1'b0 ;
  assign n13610 = n13609 ^ n13606 ^ n13320 ;
  assign n13612 = n6899 ^ n4046 ^ 1'b0 ;
  assign n13611 = n10897 ^ n6569 ^ n1527 ;
  assign n13613 = n13612 ^ n13611 ^ 1'b0 ;
  assign n13614 = ( n2955 & n10093 ) | ( n2955 & ~n12686 ) | ( n10093 & ~n12686 ) ;
  assign n13615 = n13614 ^ n12556 ^ n3939 ;
  assign n13618 = n2367 & n2421 ;
  assign n13616 = ( n300 & n843 ) | ( n300 & n1635 ) | ( n843 & n1635 ) ;
  assign n13617 = n13616 ^ n3948 ^ 1'b0 ;
  assign n13619 = n13618 ^ n13617 ^ 1'b0 ;
  assign n13620 = n13110 & ~n13619 ;
  assign n13621 = ~n1934 & n13620 ;
  assign n13622 = ~n13615 & n13621 ;
  assign n13623 = n5524 & n13622 ;
  assign n13624 = n13623 ^ n5874 ^ 1'b0 ;
  assign n13625 = n1662 | n3325 ;
  assign n13626 = n6378 & ~n13625 ;
  assign n13627 = n13626 ^ n12841 ^ 1'b0 ;
  assign n13628 = x76 & n13489 ;
  assign n13629 = n9188 & n13628 ;
  assign n13630 = ( ~n4040 & n13627 ) | ( ~n4040 & n13629 ) | ( n13627 & n13629 ) ;
  assign n13631 = n10761 ^ n9375 ^ n2348 ;
  assign n13632 = n9583 & n10118 ;
  assign n13633 = n11320 ^ n10449 ^ 1'b0 ;
  assign n13635 = n1807 | n3212 ;
  assign n13634 = n432 & n11366 ;
  assign n13636 = n13635 ^ n13634 ^ n4613 ;
  assign n13637 = ( n1173 & ~n13633 ) | ( n1173 & n13636 ) | ( ~n13633 & n13636 ) ;
  assign n13638 = n12756 ^ n5504 ^ n3897 ;
  assign n13640 = n5539 ^ n3961 ^ n3666 ;
  assign n13639 = ~n647 & n8859 ;
  assign n13641 = n13640 ^ n13639 ^ n6498 ;
  assign n13642 = n10744 ^ n8173 ^ 1'b0 ;
  assign n13643 = n13642 ^ n11589 ^ 1'b0 ;
  assign n13644 = ~n1203 & n13643 ;
  assign n13645 = n5712 ^ n1784 ^ 1'b0 ;
  assign n13646 = n6976 & ~n8700 ;
  assign n13647 = ~n533 & n12055 ;
  assign n13648 = n13647 ^ n2278 ^ n1112 ;
  assign n13651 = n3880 ^ n3271 ^ 1'b0 ;
  assign n13649 = n9599 ^ n2723 ^ 1'b0 ;
  assign n13650 = n11868 & n13649 ;
  assign n13652 = n13651 ^ n13650 ^ 1'b0 ;
  assign n13653 = n8656 ^ n6006 ^ 1'b0 ;
  assign n13654 = n6796 & n13653 ;
  assign n13655 = n13654 ^ n778 ^ 1'b0 ;
  assign n13656 = n13583 ^ n3776 ^ x2 ;
  assign n13657 = n13656 ^ n13275 ^ n7264 ;
  assign n13658 = ( ~n322 & n2526 ) | ( ~n322 & n3978 ) | ( n2526 & n3978 ) ;
  assign n13659 = ~n11831 & n13658 ;
  assign n13660 = n13659 ^ n8893 ^ 1'b0 ;
  assign n13661 = ( n1230 & n2528 ) | ( n1230 & ~n11366 ) | ( n2528 & ~n11366 ) ;
  assign n13662 = n7752 ^ n2316 ^ 1'b0 ;
  assign n13663 = ~n1802 & n13662 ;
  assign n13664 = ( n4978 & ~n6061 ) | ( n4978 & n7490 ) | ( ~n6061 & n7490 ) ;
  assign n13665 = n13663 & ~n13664 ;
  assign n13666 = n13661 & ~n13665 ;
  assign n13667 = n13666 ^ n10652 ^ 1'b0 ;
  assign n13669 = n3633 | n7582 ;
  assign n13670 = n13669 ^ n9770 ^ 1'b0 ;
  assign n13668 = ~n1648 & n13190 ;
  assign n13671 = n13670 ^ n13668 ^ 1'b0 ;
  assign n13672 = ( n10004 & n10685 ) | ( n10004 & n13671 ) | ( n10685 & n13671 ) ;
  assign n13673 = n8040 ^ n6966 ^ 1'b0 ;
  assign n13674 = ( n1849 & n7112 ) | ( n1849 & ~n13673 ) | ( n7112 & ~n13673 ) ;
  assign n13675 = ( n3567 & n13617 ) | ( n3567 & n13674 ) | ( n13617 & n13674 ) ;
  assign n13676 = n5323 ^ n761 ^ 1'b0 ;
  assign n13677 = ~n6704 & n13676 ;
  assign n13678 = ( n1398 & ~n5340 ) | ( n1398 & n9784 ) | ( ~n5340 & n9784 ) ;
  assign n13679 = n4775 ^ n3845 ^ 1'b0 ;
  assign n13680 = n2920 | n12408 ;
  assign n13681 = n13679 | n13680 ;
  assign n13682 = n2649 & ~n13681 ;
  assign n13683 = ( ~n10592 & n13678 ) | ( ~n10592 & n13682 ) | ( n13678 & n13682 ) ;
  assign n13684 = n9386 ^ x128 ^ 1'b0 ;
  assign n13685 = n3381 & n6741 ;
  assign n13686 = n7774 | n10708 ;
  assign n13687 = n12063 | n13686 ;
  assign n13688 = ( n710 & n1274 ) | ( n710 & n2851 ) | ( n1274 & n2851 ) ;
  assign n13689 = ( n1294 & n4136 ) | ( n1294 & n13688 ) | ( n4136 & n13688 ) ;
  assign n13690 = ~n3200 & n13689 ;
  assign n13691 = ~n5321 & n13690 ;
  assign n13692 = n8943 ^ n2257 ^ n741 ;
  assign n13693 = n13692 ^ n4980 ^ n4670 ;
  assign n13695 = n3694 & ~n5600 ;
  assign n13694 = n9026 ^ n528 ^ x219 ;
  assign n13696 = n13695 ^ n13694 ^ n4574 ;
  assign n13697 = n13693 | n13696 ;
  assign n13698 = n13691 & ~n13697 ;
  assign n13699 = n10151 ^ n9912 ^ n3918 ;
  assign n13700 = ( n2476 & n4251 ) | ( n2476 & ~n13699 ) | ( n4251 & ~n13699 ) ;
  assign n13701 = ( ~n2946 & n8350 ) | ( ~n2946 & n10099 ) | ( n8350 & n10099 ) ;
  assign n13702 = ( ~n2097 & n6737 ) | ( ~n2097 & n9544 ) | ( n6737 & n9544 ) ;
  assign n13703 = ( n7731 & n10550 ) | ( n7731 & ~n13702 ) | ( n10550 & ~n13702 ) ;
  assign n13704 = n4775 ^ x89 ^ 1'b0 ;
  assign n13705 = n7782 | n13704 ;
  assign n13706 = n4405 | n13705 ;
  assign n13707 = n3694 & n13706 ;
  assign n13708 = n7862 ^ n4082 ^ n3601 ;
  assign n13716 = n8703 ^ n4056 ^ 1'b0 ;
  assign n13717 = ( ~n1680 & n2991 ) | ( ~n1680 & n3674 ) | ( n2991 & n3674 ) ;
  assign n13718 = n13716 & ~n13717 ;
  assign n13712 = n10302 ^ n4028 ^ n1588 ;
  assign n13713 = n13712 ^ n10337 ^ n1282 ;
  assign n13714 = n5435 | n13713 ;
  assign n13715 = n9242 & ~n13714 ;
  assign n13709 = n1366 & ~n12206 ;
  assign n13710 = n9385 & n13709 ;
  assign n13711 = n13710 ^ n13618 ^ 1'b0 ;
  assign n13719 = n13718 ^ n13715 ^ n13711 ;
  assign n13720 = ( n1828 & ~n3518 ) | ( n1828 & n10058 ) | ( ~n3518 & n10058 ) ;
  assign n13721 = n6096 ^ n589 ^ 1'b0 ;
  assign n13722 = n707 | n13721 ;
  assign n13723 = ( n8062 & n13720 ) | ( n8062 & n13722 ) | ( n13720 & n13722 ) ;
  assign n13728 = n6207 ^ n1010 ^ n977 ;
  assign n13724 = n4373 ^ n716 ^ n491 ;
  assign n13725 = n13724 ^ n5561 ^ n1516 ;
  assign n13726 = ( ~n5665 & n12339 ) | ( ~n5665 & n13725 ) | ( n12339 & n13725 ) ;
  assign n13727 = n8101 & n13726 ;
  assign n13729 = n13728 ^ n13727 ^ 1'b0 ;
  assign n13730 = ( n710 & ~n13342 ) | ( n710 & n13729 ) | ( ~n13342 & n13729 ) ;
  assign n13731 = ~n4201 & n8406 ;
  assign n13732 = n13731 ^ n8744 ^ n3787 ;
  assign n13733 = n6282 & n6946 ;
  assign n13734 = n10359 & ~n13733 ;
  assign n13735 = n13734 ^ n8429 ^ 1'b0 ;
  assign n13736 = ( ~n2526 & n2812 ) | ( ~n2526 & n2900 ) | ( n2812 & n2900 ) ;
  assign n13737 = n13736 ^ n7824 ^ n4798 ;
  assign n13738 = n13557 ^ n10254 ^ n1943 ;
  assign n13739 = n13738 ^ n10136 ^ 1'b0 ;
  assign n13740 = n9176 ^ n7568 ^ 1'b0 ;
  assign n13741 = ( ~n13737 & n13739 ) | ( ~n13737 & n13740 ) | ( n13739 & n13740 ) ;
  assign n13742 = n3024 & ~n6456 ;
  assign n13743 = n13610 & ~n13742 ;
  assign n13744 = n13743 ^ n5572 ^ 1'b0 ;
  assign n13745 = ~n2185 & n2634 ;
  assign n13746 = n13745 ^ n1246 ^ 1'b0 ;
  assign n13747 = n13586 ^ n5236 ^ n1949 ;
  assign n13748 = n12331 & ~n13747 ;
  assign n13749 = n13748 ^ n5671 ^ 1'b0 ;
  assign n13750 = n13749 ^ n7139 ^ 1'b0 ;
  assign n13751 = ~n13746 & n13750 ;
  assign n13752 = ( n4476 & ~n9317 ) | ( n4476 & n9655 ) | ( ~n9317 & n9655 ) ;
  assign n13759 = n5418 ^ n5322 ^ 1'b0 ;
  assign n13760 = n13759 ^ n11073 ^ n10606 ;
  assign n13753 = n9721 ^ n786 ^ 1'b0 ;
  assign n13754 = n8138 & n13753 ;
  assign n13756 = n3962 & ~n12887 ;
  assign n13755 = ( n8617 & n8696 ) | ( n8617 & n9662 ) | ( n8696 & n9662 ) ;
  assign n13757 = n13756 ^ n13755 ^ 1'b0 ;
  assign n13758 = n13754 & n13757 ;
  assign n13761 = n13760 ^ n13758 ^ 1'b0 ;
  assign n13762 = x48 & n13761 ;
  assign n13763 = n10090 ^ n8215 ^ 1'b0 ;
  assign n13764 = n2853 & ~n13763 ;
  assign n13765 = n5156 & n12059 ;
  assign n13766 = n5992 & n13765 ;
  assign n13767 = n13766 ^ n7854 ^ n2183 ;
  assign n13768 = ( n2764 & n4888 ) | ( n2764 & ~n13767 ) | ( n4888 & ~n13767 ) ;
  assign n13769 = n3213 & ~n13768 ;
  assign n13770 = ( ~n2560 & n13565 ) | ( ~n2560 & n13769 ) | ( n13565 & n13769 ) ;
  assign n13774 = ~n5880 & n8536 ;
  assign n13775 = n13774 ^ n6395 ^ 1'b0 ;
  assign n13773 = ~n8805 & n9779 ;
  assign n13771 = n1967 & ~n3033 ;
  assign n13772 = n13771 ^ n10833 ^ 1'b0 ;
  assign n13776 = n13775 ^ n13773 ^ n13772 ;
  assign n13777 = n3917 & n5992 ;
  assign n13778 = n5800 ^ n4999 ^ 1'b0 ;
  assign n13780 = ( n495 & n3226 ) | ( n495 & ~n4866 ) | ( n3226 & ~n4866 ) ;
  assign n13779 = ~n2053 & n3042 ;
  assign n13781 = n13780 ^ n13779 ^ 1'b0 ;
  assign n13782 = ( n2434 & n13778 ) | ( n2434 & ~n13781 ) | ( n13778 & ~n13781 ) ;
  assign n13790 = x90 & ~n924 ;
  assign n13791 = n3051 & n13790 ;
  assign n13789 = n384 | n11113 ;
  assign n13792 = n13791 ^ n13789 ^ 1'b0 ;
  assign n13783 = n5449 | n8754 ;
  assign n13784 = n13783 ^ n6962 ^ 1'b0 ;
  assign n13785 = ( ~n7387 & n8438 ) | ( ~n7387 & n10929 ) | ( n8438 & n10929 ) ;
  assign n13786 = ( n2877 & n13784 ) | ( n2877 & ~n13785 ) | ( n13784 & ~n13785 ) ;
  assign n13787 = ~n11076 & n13786 ;
  assign n13788 = ~n2369 & n13787 ;
  assign n13793 = n13792 ^ n13788 ^ n4201 ;
  assign n13794 = ( n1850 & ~n1874 ) | ( n1850 & n2425 ) | ( ~n1874 & n2425 ) ;
  assign n13795 = ( ~n844 & n1767 ) | ( ~n844 & n10132 ) | ( n1767 & n10132 ) ;
  assign n13796 = ( n1673 & n2402 ) | ( n1673 & n13795 ) | ( n2402 & n13795 ) ;
  assign n13797 = n13796 ^ n6761 ^ n6546 ;
  assign n13798 = n13797 ^ n13259 ^ 1'b0 ;
  assign n13799 = n13794 & n13798 ;
  assign n13800 = n3988 | n5404 ;
  assign n13801 = n13800 ^ n9548 ^ 1'b0 ;
  assign n13802 = n13801 ^ n5733 ^ 1'b0 ;
  assign n13803 = ( ~n9942 & n10208 ) | ( ~n9942 & n13802 ) | ( n10208 & n13802 ) ;
  assign n13804 = n7810 ^ n516 ^ 1'b0 ;
  assign n13805 = ( ~n2285 & n3220 ) | ( ~n2285 & n12931 ) | ( n3220 & n12931 ) ;
  assign n13806 = n2690 ^ n1014 ^ 1'b0 ;
  assign n13807 = ( n1347 & ~n10277 ) | ( n1347 & n13806 ) | ( ~n10277 & n13806 ) ;
  assign n13808 = n13807 ^ n12275 ^ n305 ;
  assign n13809 = n5713 | n8574 ;
  assign n13810 = n7563 & ~n13809 ;
  assign n13811 = ( n4958 & n11873 ) | ( n4958 & n13810 ) | ( n11873 & n13810 ) ;
  assign n13812 = n13811 ^ n3499 ^ n1067 ;
  assign n13813 = n11818 ^ n4777 ^ 1'b0 ;
  assign n13814 = ( ~n6176 & n6527 ) | ( ~n6176 & n13813 ) | ( n6527 & n13813 ) ;
  assign n13819 = n6857 ^ n6492 ^ n1892 ;
  assign n13815 = n4415 ^ n2641 ^ 1'b0 ;
  assign n13816 = n13815 ^ n3884 ^ n443 ;
  assign n13817 = n4683 & n8107 ;
  assign n13818 = n13816 & n13817 ;
  assign n13820 = n13819 ^ n13818 ^ 1'b0 ;
  assign n13821 = n2555 & ~n3760 ;
  assign n13822 = n4152 & n13821 ;
  assign n13823 = n13822 ^ n6695 ^ 1'b0 ;
  assign n13824 = ( n7220 & n7280 ) | ( n7220 & n13823 ) | ( n7280 & n13823 ) ;
  assign n13825 = n13824 ^ n7471 ^ 1'b0 ;
  assign n13826 = n11145 ^ n3595 ^ 1'b0 ;
  assign n13827 = n7716 & n13826 ;
  assign n13828 = ( n1466 & n3161 ) | ( n1466 & ~n13611 ) | ( n3161 & ~n13611 ) ;
  assign n13829 = n13573 | n13768 ;
  assign n13830 = n1671 | n10805 ;
  assign n13831 = n6509 ^ n358 ^ x178 ;
  assign n13835 = n7265 ^ n6704 ^ n1125 ;
  assign n13836 = ( ~n1107 & n4204 ) | ( ~n1107 & n13835 ) | ( n4204 & n13835 ) ;
  assign n13832 = ~n4830 & n8881 ;
  assign n13833 = ~n6727 & n13832 ;
  assign n13834 = n13190 & ~n13833 ;
  assign n13837 = n13836 ^ n13834 ^ 1'b0 ;
  assign n13838 = ( ~n1304 & n13831 ) | ( ~n1304 & n13837 ) | ( n13831 & n13837 ) ;
  assign n13839 = ( n9773 & ~n10086 ) | ( n9773 & n13838 ) | ( ~n10086 & n13838 ) ;
  assign n13840 = n1897 | n10820 ;
  assign n13841 = n7766 | n13840 ;
  assign n13842 = ~n8090 & n13841 ;
  assign n13843 = n13842 ^ n873 ^ 1'b0 ;
  assign n13854 = n2619 & ~n13379 ;
  assign n13855 = n7506 & n13854 ;
  assign n13844 = n807 ^ n296 ^ 1'b0 ;
  assign n13845 = ~n3664 & n13844 ;
  assign n13847 = n5106 ^ n2572 ^ x82 ;
  assign n13846 = n826 & ~n5074 ;
  assign n13848 = n13847 ^ n13846 ^ n1940 ;
  assign n13849 = n13848 ^ n11692 ^ n1784 ;
  assign n13850 = ( n5789 & ~n11196 ) | ( n5789 & n13849 ) | ( ~n11196 & n13849 ) ;
  assign n13851 = ( n8059 & n9154 ) | ( n8059 & n13850 ) | ( n9154 & n13850 ) ;
  assign n13852 = n13851 ^ n13109 ^ 1'b0 ;
  assign n13853 = n13845 & n13852 ;
  assign n13856 = n13855 ^ n13853 ^ 1'b0 ;
  assign n13857 = n6752 ^ n2803 ^ x173 ;
  assign n13858 = n13857 ^ n6286 ^ n2097 ;
  assign n13859 = ( n712 & n6255 ) | ( n712 & n13858 ) | ( n6255 & n13858 ) ;
  assign n13862 = n6434 ^ n4184 ^ n801 ;
  assign n13863 = ( n7097 & n7927 ) | ( n7097 & ~n13862 ) | ( n7927 & ~n13862 ) ;
  assign n13864 = n13863 ^ n8164 ^ 1'b0 ;
  assign n13860 = ( x194 & n4998 ) | ( x194 & ~n12974 ) | ( n4998 & ~n12974 ) ;
  assign n13861 = ~n12475 & n13860 ;
  assign n13865 = n13864 ^ n13861 ^ 1'b0 ;
  assign n13866 = ( n8417 & ~n13859 ) | ( n8417 & n13865 ) | ( ~n13859 & n13865 ) ;
  assign n13867 = ( ~n7919 & n10299 ) | ( ~n7919 & n11145 ) | ( n10299 & n11145 ) ;
  assign n13868 = ( n565 & n2374 ) | ( n565 & n6468 ) | ( n2374 & n6468 ) ;
  assign n13869 = n4209 & n13868 ;
  assign n13870 = n13869 ^ n10151 ^ 1'b0 ;
  assign n13871 = n13870 ^ n8311 ^ 1'b0 ;
  assign n13872 = n9444 | n13871 ;
  assign n13873 = n10871 ^ n6701 ^ n465 ;
  assign n13874 = ( n2406 & n2615 ) | ( n2406 & ~n9291 ) | ( n2615 & ~n9291 ) ;
  assign n13875 = n4155 & n13874 ;
  assign n13876 = n13873 & ~n13875 ;
  assign n13877 = n13872 & n13876 ;
  assign n13878 = n13336 ^ n9547 ^ 1'b0 ;
  assign n13879 = ( ~n6136 & n13877 ) | ( ~n6136 & n13878 ) | ( n13877 & n13878 ) ;
  assign n13880 = n5063 | n12523 ;
  assign n13881 = n13880 ^ n2312 ^ 1'b0 ;
  assign n13882 = n10438 ^ n5801 ^ 1'b0 ;
  assign n13883 = n10315 | n11327 ;
  assign n13884 = n4279 & ~n8965 ;
  assign n13885 = n4477 | n13884 ;
  assign n13886 = n13885 ^ n3214 ^ n435 ;
  assign n13887 = x235 & n13886 ;
  assign n13888 = ~n6793 & n13887 ;
  assign n13889 = ( n6190 & n12434 ) | ( n6190 & ~n13888 ) | ( n12434 & ~n13888 ) ;
  assign n13890 = n7498 ^ n5231 ^ 1'b0 ;
  assign n13891 = n13890 ^ n11436 ^ n10469 ;
  assign n13892 = n8548 | n13891 ;
  assign n13893 = n829 & ~n2326 ;
  assign n13894 = n4837 ^ n1927 ^ n860 ;
  assign n13895 = n8136 ^ n6577 ^ n5729 ;
  assign n13896 = ( ~n6630 & n10993 ) | ( ~n6630 & n13895 ) | ( n10993 & n13895 ) ;
  assign n13897 = n7053 | n13896 ;
  assign n13898 = n13894 & ~n13897 ;
  assign n13901 = n12370 ^ n6961 ^ 1'b0 ;
  assign n13902 = n1271 & n13901 ;
  assign n13899 = n10019 ^ n1570 ^ 1'b0 ;
  assign n13900 = n13899 ^ n11239 ^ n8763 ;
  assign n13903 = n13902 ^ n13900 ^ n13211 ;
  assign n13904 = n6887 ^ n2918 ^ n2362 ;
  assign n13905 = ~n12097 & n13904 ;
  assign n13906 = n13905 ^ n2247 ^ 1'b0 ;
  assign n13907 = n13906 ^ n1793 ^ n478 ;
  assign n13908 = ~n2922 & n3897 ;
  assign n13909 = n13908 ^ n2863 ^ 1'b0 ;
  assign n13910 = n6507 | n13909 ;
  assign n13911 = n13907 | n13910 ;
  assign n13912 = n1690 & n7110 ;
  assign n13913 = n13912 ^ n7588 ^ 1'b0 ;
  assign n13914 = n7964 ^ n7456 ^ 1'b0 ;
  assign n13915 = ( n11301 & ~n13913 ) | ( n11301 & n13914 ) | ( ~n13913 & n13914 ) ;
  assign n13916 = n4577 | n13915 ;
  assign n13917 = ( n10019 & n11376 ) | ( n10019 & n13916 ) | ( n11376 & n13916 ) ;
  assign n13918 = n3817 ^ n3190 ^ n2881 ;
  assign n13919 = ( n646 & n2593 ) | ( n646 & n13918 ) | ( n2593 & n13918 ) ;
  assign n13920 = n5631 ^ n1987 ^ 1'b0 ;
  assign n13921 = ~n3285 & n13920 ;
  assign n13922 = ( ~n4073 & n13919 ) | ( ~n4073 & n13921 ) | ( n13919 & n13921 ) ;
  assign n13923 = ~n3867 & n13922 ;
  assign n13924 = n13923 ^ n1022 ^ 1'b0 ;
  assign n13925 = n9652 & n13924 ;
  assign n13926 = n5456 ^ n4156 ^ x20 ;
  assign n13927 = n13926 ^ n10432 ^ n6035 ;
  assign n13928 = n4997 ^ x177 ^ 1'b0 ;
  assign n13929 = n11205 | n13928 ;
  assign n13930 = n13929 ^ n10252 ^ 1'b0 ;
  assign n13931 = ~n6681 & n13930 ;
  assign n13932 = n13410 ^ n2494 ^ 1'b0 ;
  assign n13933 = n6001 & ~n10880 ;
  assign n13934 = n10994 & n13933 ;
  assign n13935 = ( ~n946 & n13760 ) | ( ~n946 & n13934 ) | ( n13760 & n13934 ) ;
  assign n13936 = n1962 & ~n13935 ;
  assign n13937 = x110 & n11031 ;
  assign n13938 = n6791 | n7843 ;
  assign n13939 = n13937 | n13938 ;
  assign n13948 = ~n5756 & n9365 ;
  assign n13949 = n5377 & n13948 ;
  assign n13950 = n13949 ^ n10191 ^ 1'b0 ;
  assign n13940 = n4519 & ~n8886 ;
  assign n13941 = ~n1323 & n13940 ;
  assign n13943 = n10405 ^ n4836 ^ n1804 ;
  assign n13942 = ( ~n1590 & n5478 ) | ( ~n1590 & n6932 ) | ( n5478 & n6932 ) ;
  assign n13944 = n13943 ^ n13942 ^ n5976 ;
  assign n13945 = ~n13941 & n13944 ;
  assign n13946 = n13945 ^ n9275 ^ 1'b0 ;
  assign n13947 = n4770 | n13946 ;
  assign n13951 = n13950 ^ n13947 ^ 1'b0 ;
  assign n13952 = ~n6362 & n9740 ;
  assign n13953 = n4193 & n13952 ;
  assign n13954 = n13953 ^ n3258 ^ x159 ;
  assign n13955 = ( ~n2641 & n5104 ) | ( ~n2641 & n5432 ) | ( n5104 & n5432 ) ;
  assign n13956 = n7535 & ~n13955 ;
  assign n13957 = ~n542 & n7727 ;
  assign n13958 = n13957 ^ x191 ^ 1'b0 ;
  assign n13959 = n8704 & ~n13958 ;
  assign n13960 = n13959 ^ n4868 ^ 1'b0 ;
  assign n13961 = ( n2478 & n8509 ) | ( n2478 & n13960 ) | ( n8509 & n13960 ) ;
  assign n13962 = n13961 ^ n4983 ^ 1'b0 ;
  assign n13963 = ( n7268 & ~n7543 ) | ( n7268 & n8087 ) | ( ~n7543 & n8087 ) ;
  assign n13964 = n923 & ~n13851 ;
  assign n13965 = n10444 & n13964 ;
  assign n13966 = n4602 | n11962 ;
  assign n13967 = n8017 & ~n13966 ;
  assign n13968 = ( n6668 & n10544 ) | ( n6668 & n13002 ) | ( n10544 & n13002 ) ;
  assign n13969 = ( n3784 & n4010 ) | ( n3784 & ~n4521 ) | ( n4010 & ~n4521 ) ;
  assign n13970 = n5815 ^ x222 ^ 1'b0 ;
  assign n13971 = ~n4333 & n13970 ;
  assign n13972 = ( n9779 & n13969 ) | ( n9779 & n13971 ) | ( n13969 & n13971 ) ;
  assign n13973 = n4601 & ~n7597 ;
  assign n13974 = n13973 ^ n6667 ^ 1'b0 ;
  assign n13975 = n9936 & ~n13974 ;
  assign n13976 = n13972 & n13975 ;
  assign n13981 = n6242 ^ n1307 ^ n851 ;
  assign n13982 = n550 | n13981 ;
  assign n13983 = n13982 ^ n4762 ^ 1'b0 ;
  assign n13984 = n13983 ^ n2691 ^ 1'b0 ;
  assign n13977 = n4582 & n4626 ;
  assign n13978 = n9136 ^ n5150 ^ n3625 ;
  assign n13979 = n6562 | n13978 ;
  assign n13980 = ( ~n4795 & n13977 ) | ( ~n4795 & n13979 ) | ( n13977 & n13979 ) ;
  assign n13985 = n13984 ^ n13980 ^ n2155 ;
  assign n13986 = n13985 ^ n10072 ^ n553 ;
  assign n13987 = ( n6070 & n13976 ) | ( n6070 & n13986 ) | ( n13976 & n13986 ) ;
  assign n13988 = ( n604 & n3908 ) | ( n604 & n7637 ) | ( n3908 & n7637 ) ;
  assign n13989 = n5158 ^ n2478 ^ 1'b0 ;
  assign n13990 = ( n4783 & ~n13988 ) | ( n4783 & n13989 ) | ( ~n13988 & n13989 ) ;
  assign n13991 = n13990 ^ n7258 ^ n3906 ;
  assign n13992 = n12388 ^ n2592 ^ n898 ;
  assign n13993 = n13992 ^ n7612 ^ 1'b0 ;
  assign n13994 = ~n13991 & n13993 ;
  assign n13995 = n1442 | n3024 ;
  assign n13996 = n13995 ^ n332 ^ 1'b0 ;
  assign n13997 = n2896 & n8933 ;
  assign n13998 = ~n6183 & n9205 ;
  assign n13999 = n13998 ^ n13717 ^ 1'b0 ;
  assign n14000 = n13999 ^ n3452 ^ 1'b0 ;
  assign n14001 = ~n13997 & n14000 ;
  assign n14002 = ( n9938 & n10953 ) | ( n9938 & n13366 ) | ( n10953 & n13366 ) ;
  assign n14003 = ~n470 & n10897 ;
  assign n14004 = n14003 ^ n7645 ^ n2682 ;
  assign n14005 = ~n285 & n7271 ;
  assign n14006 = ( n3141 & n5223 ) | ( n3141 & n7076 ) | ( n5223 & n7076 ) ;
  assign n14007 = n14006 ^ n13729 ^ n556 ;
  assign n14008 = ( ~n12536 & n14005 ) | ( ~n12536 & n14007 ) | ( n14005 & n14007 ) ;
  assign n14009 = ( n1442 & n5032 ) | ( n1442 & ~n9220 ) | ( n5032 & ~n9220 ) ;
  assign n14010 = n14009 ^ n7280 ^ n4305 ;
  assign n14011 = ( n4927 & n10920 ) | ( n4927 & n13404 ) | ( n10920 & n13404 ) ;
  assign n14023 = ( n1176 & n2785 ) | ( n1176 & n4279 ) | ( n2785 & n4279 ) ;
  assign n14020 = n4514 ^ n450 ^ 1'b0 ;
  assign n14021 = n708 & n14020 ;
  assign n14016 = n3146 & ~n7269 ;
  assign n14017 = ~x198 & n14016 ;
  assign n14014 = n11867 ^ n8678 ^ 1'b0 ;
  assign n14015 = n1323 & n14014 ;
  assign n14018 = n14017 ^ n14015 ^ 1'b0 ;
  assign n14019 = n8361 & ~n14018 ;
  assign n14022 = n14021 ^ n14019 ^ n11388 ;
  assign n14012 = n1862 ^ x54 ^ 1'b0 ;
  assign n14013 = n8661 & ~n14012 ;
  assign n14024 = n14023 ^ n14022 ^ n14013 ;
  assign n14025 = ( n4305 & n5086 ) | ( n4305 & ~n12970 ) | ( n5086 & ~n12970 ) ;
  assign n14026 = n14025 ^ n3049 ^ 1'b0 ;
  assign n14027 = n13222 | n14026 ;
  assign n14028 = n10769 ^ n5101 ^ 1'b0 ;
  assign n14029 = ( n5799 & ~n6114 ) | ( n5799 & n11757 ) | ( ~n6114 & n11757 ) ;
  assign n14030 = n1858 | n14029 ;
  assign n14031 = n14030 ^ n10555 ^ 1'b0 ;
  assign n14039 = x196 & ~n2120 ;
  assign n14040 = n14039 ^ n8785 ^ 1'b0 ;
  assign n14041 = ( n2543 & ~n7108 ) | ( n2543 & n14040 ) | ( ~n7108 & n14040 ) ;
  assign n14042 = ( n582 & ~n842 ) | ( n582 & n14041 ) | ( ~n842 & n14041 ) ;
  assign n14032 = ( n3673 & ~n7801 ) | ( n3673 & n9890 ) | ( ~n7801 & n9890 ) ;
  assign n14035 = ( ~n1122 & n5352 ) | ( ~n1122 & n7610 ) | ( n5352 & n7610 ) ;
  assign n14036 = n14035 ^ n8584 ^ n5325 ;
  assign n14033 = ( ~n1589 & n4850 ) | ( ~n1589 & n11709 ) | ( n4850 & n11709 ) ;
  assign n14034 = n9025 & ~n14033 ;
  assign n14037 = n14036 ^ n14034 ^ 1'b0 ;
  assign n14038 = n14032 & ~n14037 ;
  assign n14043 = n14042 ^ n14038 ^ 1'b0 ;
  assign n14044 = n14043 ^ n10485 ^ n9684 ;
  assign n14045 = n7839 & n13112 ;
  assign n14046 = n7329 & ~n11408 ;
  assign n14049 = n12993 ^ n2478 ^ n1551 ;
  assign n14047 = n3070 | n6510 ;
  assign n14048 = n5424 | n14047 ;
  assign n14050 = n14049 ^ n14048 ^ 1'b0 ;
  assign n14051 = n1705 ^ n1507 ^ 1'b0 ;
  assign n14052 = n14051 ^ n5346 ^ n4433 ;
  assign n14053 = n6727 ^ n4079 ^ 1'b0 ;
  assign n14054 = ( ~n3109 & n5145 ) | ( ~n3109 & n14053 ) | ( n5145 & n14053 ) ;
  assign n14055 = ~n1561 & n14054 ;
  assign n14056 = n1270 & ~n2923 ;
  assign n14057 = n14055 & n14056 ;
  assign n14058 = n3626 ^ n1188 ^ 1'b0 ;
  assign n14059 = n1300 | n14058 ;
  assign n14060 = n13678 | n14059 ;
  assign n14061 = ( ~n4483 & n14057 ) | ( ~n4483 & n14060 ) | ( n14057 & n14060 ) ;
  assign n14062 = n14061 ^ n5038 ^ n562 ;
  assign n14063 = ( n6376 & n14052 ) | ( n6376 & ~n14062 ) | ( n14052 & ~n14062 ) ;
  assign n14064 = n10942 ^ n6611 ^ n1836 ;
  assign n14065 = ~n1573 & n5470 ;
  assign n14066 = ~n3699 & n5516 ;
  assign n14067 = n14066 ^ n9720 ^ 1'b0 ;
  assign n14068 = ( n1885 & n6496 ) | ( n1885 & n14067 ) | ( n6496 & n14067 ) ;
  assign n14076 = n10785 ^ n934 ^ 1'b0 ;
  assign n14074 = n11046 ^ n1431 ^ 1'b0 ;
  assign n14071 = n6965 ^ n6534 ^ x14 ;
  assign n14072 = x33 & ~n14071 ;
  assign n14073 = n905 & n14072 ;
  assign n14069 = n3368 ^ n1717 ^ n295 ;
  assign n14070 = n12045 & n14069 ;
  assign n14075 = n14074 ^ n14073 ^ n14070 ;
  assign n14077 = n14076 ^ n14075 ^ n2884 ;
  assign n14078 = n3511 | n5671 ;
  assign n14079 = n14078 ^ n8531 ^ n1279 ;
  assign n14080 = ~n2200 & n14079 ;
  assign n14081 = n2693 ^ n1296 ^ x36 ;
  assign n14082 = n14081 ^ n12694 ^ 1'b0 ;
  assign n14083 = ( n883 & n12544 ) | ( n883 & n12550 ) | ( n12544 & n12550 ) ;
  assign n14084 = n4645 | n6184 ;
  assign n14087 = n12045 ^ n8579 ^ 1'b0 ;
  assign n14085 = n5567 & n12511 ;
  assign n14086 = n14085 ^ n6458 ^ n2365 ;
  assign n14088 = n14087 ^ n14086 ^ 1'b0 ;
  assign n14089 = n9938 & ~n14088 ;
  assign n14090 = n14089 ^ n959 ^ 1'b0 ;
  assign n14091 = n11303 ^ n10517 ^ n483 ;
  assign n14092 = n12623 ^ n9464 ^ 1'b0 ;
  assign n14093 = n1130 & n14092 ;
  assign n14094 = ( ~n7547 & n8354 ) | ( ~n7547 & n13841 ) | ( n8354 & n13841 ) ;
  assign n14095 = n13568 ^ n567 ^ x163 ;
  assign n14098 = ( n2042 & ~n3046 ) | ( n2042 & n12676 ) | ( ~n3046 & n12676 ) ;
  assign n14096 = ( x89 & n2845 ) | ( x89 & ~n12591 ) | ( n2845 & ~n12591 ) ;
  assign n14097 = n14096 ^ n3190 ^ n3156 ;
  assign n14099 = n14098 ^ n14097 ^ n9802 ;
  assign n14103 = n10103 ^ n351 ^ x225 ;
  assign n14100 = n9537 ^ n4516 ^ 1'b0 ;
  assign n14101 = n6391 ^ n2376 ^ 1'b0 ;
  assign n14102 = ( n11011 & n14100 ) | ( n11011 & ~n14101 ) | ( n14100 & ~n14101 ) ;
  assign n14104 = n14103 ^ n14102 ^ n3949 ;
  assign n14105 = n2105 & n4124 ;
  assign n14106 = n14105 ^ n781 ^ 1'b0 ;
  assign n14107 = n14106 ^ n6950 ^ n1692 ;
  assign n14108 = n5616 ^ n1277 ^ 1'b0 ;
  assign n14109 = n10058 ^ n1826 ^ 1'b0 ;
  assign n14110 = n14109 ^ n7722 ^ 1'b0 ;
  assign n14111 = ~n14108 & n14110 ;
  assign n14112 = ~n520 & n7901 ;
  assign n14113 = ~n8694 & n14112 ;
  assign n14114 = n10886 ^ n1209 ^ x87 ;
  assign n14116 = n1804 ^ n1050 ^ 1'b0 ;
  assign n14115 = n3831 | n12125 ;
  assign n14117 = n14116 ^ n14115 ^ 1'b0 ;
  assign n14118 = n4779 & ~n5184 ;
  assign n14119 = n7392 | n11538 ;
  assign n14120 = n14118 | n14119 ;
  assign n14121 = n14117 & ~n14120 ;
  assign n14122 = ( n6626 & n7521 ) | ( n6626 & ~n14121 ) | ( n7521 & ~n14121 ) ;
  assign n14125 = ( n2664 & ~n4085 ) | ( n2664 & n5676 ) | ( ~n4085 & n5676 ) ;
  assign n14123 = n4987 & ~n7999 ;
  assign n14124 = n471 & ~n14123 ;
  assign n14126 = n14125 ^ n14124 ^ 1'b0 ;
  assign n14127 = n5906 | n14126 ;
  assign n14128 = n12003 ^ n2084 ^ 1'b0 ;
  assign n14129 = ( ~n260 & n3499 ) | ( ~n260 & n5008 ) | ( n3499 & n5008 ) ;
  assign n14130 = ( n9216 & n14128 ) | ( n9216 & ~n14129 ) | ( n14128 & ~n14129 ) ;
  assign n14131 = x27 & ~n4291 ;
  assign n14132 = ( n10532 & n11380 ) | ( n10532 & ~n12348 ) | ( n11380 & ~n12348 ) ;
  assign n14133 = n13149 ^ n5216 ^ 1'b0 ;
  assign n14134 = n7706 | n14133 ;
  assign n14135 = n675 & n14134 ;
  assign n14136 = ~n4570 & n12313 ;
  assign n14137 = ( n1784 & n10517 ) | ( n1784 & n14136 ) | ( n10517 & n14136 ) ;
  assign n14138 = ~n704 & n3185 ;
  assign n14139 = n14138 ^ n6564 ^ 1'b0 ;
  assign n14140 = n8867 ^ n6430 ^ n5682 ;
  assign n14141 = ~n7147 & n14140 ;
  assign n14142 = n14141 ^ n2951 ^ 1'b0 ;
  assign n14143 = n9460 & ~n14142 ;
  assign n14144 = ~n7722 & n14143 ;
  assign n14145 = n10625 & ~n14144 ;
  assign n14146 = n14139 & n14145 ;
  assign n14147 = ~n7337 & n12243 ;
  assign n14148 = n5388 ^ n2318 ^ 1'b0 ;
  assign n14149 = n7475 ^ n521 ^ 1'b0 ;
  assign n14150 = n14148 & n14149 ;
  assign n14151 = n10140 ^ n8956 ^ x60 ;
  assign n14152 = n8272 & ~n14151 ;
  assign n14153 = n14150 & n14152 ;
  assign n14159 = n5302 ^ n2104 ^ n368 ;
  assign n14160 = n9922 | n14159 ;
  assign n14161 = n14160 ^ n9996 ^ 1'b0 ;
  assign n14154 = n1197 & n3532 ;
  assign n14155 = n14154 ^ n5520 ^ 1'b0 ;
  assign n14156 = ( ~n7606 & n9816 ) | ( ~n7606 & n10152 ) | ( n9816 & n10152 ) ;
  assign n14157 = n14156 ^ n5947 ^ 1'b0 ;
  assign n14158 = n14155 & ~n14157 ;
  assign n14162 = n14161 ^ n14158 ^ 1'b0 ;
  assign n14163 = ~n14153 & n14162 ;
  assign n14164 = ( ~x181 & n1532 ) | ( ~x181 & n3193 ) | ( n1532 & n3193 ) ;
  assign n14165 = n14164 ^ n443 ^ 1'b0 ;
  assign n14166 = ~n1884 & n5809 ;
  assign n14167 = ~n2427 & n14166 ;
  assign n14168 = n14019 ^ n10831 ^ n1597 ;
  assign n14169 = n6520 ^ n2260 ^ 1'b0 ;
  assign n14170 = n14169 ^ n10919 ^ n6847 ;
  assign n14171 = ~n4086 & n14170 ;
  assign n14172 = ~n14168 & n14171 ;
  assign n14173 = ( ~n14165 & n14167 ) | ( ~n14165 & n14172 ) | ( n14167 & n14172 ) ;
  assign n14174 = n5767 & n8294 ;
  assign n14175 = n1393 ^ n901 ^ 1'b0 ;
  assign n14176 = n14175 ^ n2097 ^ n733 ;
  assign n14177 = n5421 & n14176 ;
  assign n14178 = ~n572 & n14177 ;
  assign n14179 = n1657 | n2212 ;
  assign n14180 = n579 | n14179 ;
  assign n14181 = ( n10541 & ~n14178 ) | ( n10541 & n14180 ) | ( ~n14178 & n14180 ) ;
  assign n14182 = n279 & n14181 ;
  assign n14183 = ( n1820 & n4801 ) | ( n1820 & ~n6655 ) | ( n4801 & ~n6655 ) ;
  assign n14184 = n9962 & n14183 ;
  assign n14185 = ~n4204 & n14184 ;
  assign n14188 = ~n895 & n2381 ;
  assign n14189 = ( n11975 & ~n12097 ) | ( n11975 & n14188 ) | ( ~n12097 & n14188 ) ;
  assign n14186 = ( n1831 & n1926 ) | ( n1831 & n6989 ) | ( n1926 & n6989 ) ;
  assign n14187 = x65 & ~n14186 ;
  assign n14190 = n14189 ^ n14187 ^ 1'b0 ;
  assign n14191 = ( n5664 & ~n13472 ) | ( n5664 & n14190 ) | ( ~n13472 & n14190 ) ;
  assign n14192 = ( n6186 & n11287 ) | ( n6186 & ~n14191 ) | ( n11287 & ~n14191 ) ;
  assign n14193 = ( n12772 & n14185 ) | ( n12772 & n14192 ) | ( n14185 & n14192 ) ;
  assign n14194 = n14193 ^ n7669 ^ 1'b0 ;
  assign n14195 = ( n689 & ~n3763 ) | ( n689 & n4261 ) | ( ~n3763 & n4261 ) ;
  assign n14196 = n8231 ^ n448 ^ 1'b0 ;
  assign n14197 = ~n14195 & n14196 ;
  assign n14198 = ~n6146 & n14197 ;
  assign n14199 = n14198 ^ n10585 ^ 1'b0 ;
  assign n14200 = ~n11537 & n14199 ;
  assign n14201 = n14200 ^ n10704 ^ 1'b0 ;
  assign n14207 = n5640 ^ n3785 ^ 1'b0 ;
  assign n14208 = n14207 ^ n11275 ^ 1'b0 ;
  assign n14209 = n14208 ^ n4811 ^ 1'b0 ;
  assign n14210 = n11523 & ~n14209 ;
  assign n14202 = n8987 ^ n7395 ^ n6589 ;
  assign n14203 = n14202 ^ n14148 ^ n8895 ;
  assign n14204 = n1264 & ~n14203 ;
  assign n14205 = n14204 ^ n13408 ^ 1'b0 ;
  assign n14206 = ( n3163 & n11922 ) | ( n3163 & n14205 ) | ( n11922 & n14205 ) ;
  assign n14211 = n14210 ^ n14206 ^ n11482 ;
  assign n14212 = n4357 & n5180 ;
  assign n14213 = n14212 ^ n6659 ^ 1'b0 ;
  assign n14218 = n425 & ~n5673 ;
  assign n14219 = ~n10377 & n14218 ;
  assign n14220 = n14219 ^ n10281 ^ n4524 ;
  assign n14221 = n14220 ^ n12614 ^ 1'b0 ;
  assign n14214 = ( n1107 & n2460 ) | ( n1107 & n10884 ) | ( n2460 & n10884 ) ;
  assign n14215 = ( n395 & ~n6981 ) | ( n395 & n14214 ) | ( ~n6981 & n14214 ) ;
  assign n14216 = n13410 ^ n7265 ^ 1'b0 ;
  assign n14217 = n14215 | n14216 ;
  assign n14222 = n14221 ^ n14217 ^ 1'b0 ;
  assign n14223 = n12198 ^ n11749 ^ n8580 ;
  assign n14224 = ( n640 & ~n10352 ) | ( n640 & n14223 ) | ( ~n10352 & n14223 ) ;
  assign n14226 = n5946 ^ n3801 ^ 1'b0 ;
  assign n14227 = ~n2793 & n14226 ;
  assign n14225 = n3626 & ~n7120 ;
  assign n14228 = n14227 ^ n14225 ^ 1'b0 ;
  assign n14229 = ~n7993 & n14228 ;
  assign n14230 = n14229 ^ n11304 ^ 1'b0 ;
  assign n14233 = n10672 ^ n3507 ^ 1'b0 ;
  assign n14234 = n14233 ^ n320 ^ 1'b0 ;
  assign n14231 = n1643 & ~n3445 ;
  assign n14232 = n14231 ^ n6185 ^ 1'b0 ;
  assign n14235 = n14234 ^ n14232 ^ n6959 ;
  assign n14236 = ( n6384 & ~n8286 ) | ( n6384 & n14235 ) | ( ~n8286 & n14235 ) ;
  assign n14237 = ( n1886 & ~n5278 ) | ( n1886 & n14236 ) | ( ~n5278 & n14236 ) ;
  assign n14243 = n11721 & n11809 ;
  assign n14238 = n10941 | n12365 ;
  assign n14239 = n661 | n14238 ;
  assign n14240 = n14239 ^ n9362 ^ 1'b0 ;
  assign n14241 = n5908 & n14240 ;
  assign n14242 = n1367 & n14241 ;
  assign n14244 = n14243 ^ n14242 ^ 1'b0 ;
  assign n14245 = ( n5195 & n6069 ) | ( n5195 & n14244 ) | ( n6069 & n14244 ) ;
  assign n14246 = n7605 ^ n1836 ^ n1404 ;
  assign n14247 = n14246 ^ n8109 ^ 1'b0 ;
  assign n14248 = x114 & n997 ;
  assign n14249 = n7440 & n14248 ;
  assign n14250 = n14249 ^ n8438 ^ 1'b0 ;
  assign n14251 = n14250 ^ n6608 ^ 1'b0 ;
  assign n14252 = n6540 | n14251 ;
  assign n14253 = ( x187 & n7320 ) | ( x187 & n14252 ) | ( n7320 & n14252 ) ;
  assign n14254 = n604 | n7083 ;
  assign n14255 = n1294 | n14254 ;
  assign n14256 = n8900 ^ n3398 ^ n2555 ;
  assign n14257 = ( ~n3148 & n10063 ) | ( ~n3148 & n12681 ) | ( n10063 & n12681 ) ;
  assign n14259 = n8257 ^ n5320 ^ 1'b0 ;
  assign n14258 = ( ~n3317 & n4399 ) | ( ~n3317 & n9375 ) | ( n4399 & n9375 ) ;
  assign n14260 = n14259 ^ n14258 ^ 1'b0 ;
  assign n14261 = n11056 & ~n14260 ;
  assign n14262 = ( n9911 & n14257 ) | ( n9911 & ~n14261 ) | ( n14257 & ~n14261 ) ;
  assign n14263 = ~n401 & n6105 ;
  assign n14264 = n9620 & n14263 ;
  assign n14265 = ( ~n450 & n1861 ) | ( ~n450 & n14264 ) | ( n1861 & n14264 ) ;
  assign n14266 = ~n4024 & n4521 ;
  assign n14267 = ~n609 & n14266 ;
  assign n14268 = x99 | n6351 ;
  assign n14269 = x83 & ~n603 ;
  assign n14270 = n3689 & ~n3911 ;
  assign n14271 = ( ~n1914 & n3615 ) | ( ~n1914 & n14270 ) | ( n3615 & n14270 ) ;
  assign n14272 = n5033 ^ n4094 ^ n1167 ;
  assign n14273 = n7229 | n14272 ;
  assign n14274 = n14271 & ~n14273 ;
  assign n14276 = n10617 ^ n8882 ^ n2478 ;
  assign n14275 = n1924 | n5593 ;
  assign n14277 = n14276 ^ n14275 ^ 1'b0 ;
  assign n14278 = n5055 | n14277 ;
  assign n14279 = n7605 ^ n2807 ^ n636 ;
  assign n14280 = n12082 ^ n10777 ^ n7397 ;
  assign n14281 = n14279 & ~n14280 ;
  assign n14282 = n13867 ^ n5082 ^ 1'b0 ;
  assign n14283 = ~n9402 & n14282 ;
  assign n14285 = n7448 ^ n6767 ^ 1'b0 ;
  assign n14284 = n3464 & ~n9614 ;
  assign n14286 = n14285 ^ n14284 ^ 1'b0 ;
  assign n14287 = n4522 & ~n14286 ;
  assign n14288 = n2798 ^ n2438 ^ 1'b0 ;
  assign n14289 = n14288 ^ n3557 ^ 1'b0 ;
  assign n14290 = n7985 & ~n14289 ;
  assign n14291 = n14287 & ~n14290 ;
  assign n14297 = n2584 & n9039 ;
  assign n14292 = n10075 ^ n6691 ^ n3481 ;
  assign n14293 = n2233 ^ n1827 ^ x251 ;
  assign n14294 = n14292 | n14293 ;
  assign n14295 = ( n4413 & n7203 ) | ( n4413 & n10881 ) | ( n7203 & n10881 ) ;
  assign n14296 = ( n937 & n14294 ) | ( n937 & ~n14295 ) | ( n14294 & ~n14295 ) ;
  assign n14298 = n14297 ^ n14296 ^ n2999 ;
  assign n14299 = n5003 ^ n3145 ^ n317 ;
  assign n14300 = n789 & ~n14299 ;
  assign n14301 = n14300 ^ n13502 ^ n1182 ;
  assign n14302 = n14301 ^ n11485 ^ n3437 ;
  assign n14304 = ~n1569 & n8224 ;
  assign n14305 = n14304 ^ n4453 ^ 1'b0 ;
  assign n14303 = ( n271 & ~n5933 ) | ( n271 & n6329 ) | ( ~n5933 & n6329 ) ;
  assign n14306 = n14305 ^ n14303 ^ n13847 ;
  assign n14307 = n5268 ^ n4681 ^ 1'b0 ;
  assign n14308 = ~n2773 & n12057 ;
  assign n14309 = ~n1737 & n14308 ;
  assign n14310 = n12510 ^ n9778 ^ n847 ;
  assign n14311 = ( n6404 & n9043 ) | ( n6404 & ~n14254 ) | ( n9043 & ~n14254 ) ;
  assign n14312 = ( n9448 & n14310 ) | ( n9448 & n14311 ) | ( n14310 & n14311 ) ;
  assign n14313 = n11290 ^ n8566 ^ x36 ;
  assign n14316 = n11389 ^ n8903 ^ n6795 ;
  assign n14314 = ( n746 & ~n3448 ) | ( n746 & n11653 ) | ( ~n3448 & n11653 ) ;
  assign n14315 = n14314 ^ n8466 ^ n5704 ;
  assign n14317 = n14316 ^ n14315 ^ 1'b0 ;
  assign n14318 = ( n1313 & n2066 ) | ( n1313 & ~n10979 ) | ( n2066 & ~n10979 ) ;
  assign n14322 = n5937 ^ n4479 ^ 1'b0 ;
  assign n14323 = n5783 ^ n562 ^ 1'b0 ;
  assign n14324 = ~n14322 & n14323 ;
  assign n14325 = n327 & n14324 ;
  assign n14326 = ( ~n1227 & n2939 ) | ( ~n1227 & n14325 ) | ( n2939 & n14325 ) ;
  assign n14327 = n4524 ^ n1671 ^ 1'b0 ;
  assign n14328 = n14326 & ~n14327 ;
  assign n14321 = ( ~n2766 & n4857 ) | ( ~n2766 & n11034 ) | ( n4857 & n11034 ) ;
  assign n14319 = n1138 & n6320 ;
  assign n14320 = ( n4275 & ~n13529 ) | ( n4275 & n14319 ) | ( ~n13529 & n14319 ) ;
  assign n14329 = n14328 ^ n14321 ^ n14320 ;
  assign n14330 = ( n5132 & n7406 ) | ( n5132 & ~n12301 ) | ( n7406 & ~n12301 ) ;
  assign n14331 = n11784 & ~n14330 ;
  assign n14332 = n11895 | n14331 ;
  assign n14333 = n2428 & ~n3101 ;
  assign n14334 = ~n14170 & n14333 ;
  assign n14335 = n11120 & ~n14334 ;
  assign n14336 = ~n14332 & n14335 ;
  assign n14337 = n11489 ^ n9132 ^ n3948 ;
  assign n14338 = n4697 & n14337 ;
  assign n14339 = n12621 ^ n4632 ^ n308 ;
  assign n14340 = ( ~n596 & n6998 ) | ( ~n596 & n14339 ) | ( n6998 & n14339 ) ;
  assign n14341 = ( n3567 & ~n3864 ) | ( n3567 & n4394 ) | ( ~n3864 & n4394 ) ;
  assign n14342 = ( n5588 & ~n11493 ) | ( n5588 & n14341 ) | ( ~n11493 & n14341 ) ;
  assign n14343 = n1975 & ~n5946 ;
  assign n14344 = n2984 & n14343 ;
  assign n14345 = n14344 ^ n6517 ^ 1'b0 ;
  assign n14346 = n4966 & n14345 ;
  assign n14347 = ( n2602 & ~n2986 ) | ( n2602 & n5057 ) | ( ~n2986 & n5057 ) ;
  assign n14348 = n14347 ^ n12487 ^ 1'b0 ;
  assign n14349 = n8334 ^ n3092 ^ x142 ;
  assign n14350 = n2686 & ~n3236 ;
  assign n14351 = n14350 ^ n5958 ^ 1'b0 ;
  assign n14352 = n14351 ^ n4800 ^ 1'b0 ;
  assign n14353 = ( n2614 & n12296 ) | ( n2614 & ~n14352 ) | ( n12296 & ~n14352 ) ;
  assign n14354 = ( ~n6267 & n14349 ) | ( ~n6267 & n14353 ) | ( n14349 & n14353 ) ;
  assign n14355 = ( n929 & n1152 ) | ( n929 & ~n1326 ) | ( n1152 & ~n1326 ) ;
  assign n14356 = n8157 ^ n1189 ^ 1'b0 ;
  assign n14357 = n14355 & n14356 ;
  assign n14358 = n14357 ^ n1440 ^ 1'b0 ;
  assign n14359 = n2466 & n8607 ;
  assign n14360 = n14359 ^ n9983 ^ 1'b0 ;
  assign n14361 = ( n5329 & n10677 ) | ( n5329 & ~n14360 ) | ( n10677 & ~n14360 ) ;
  assign n14362 = ~n14358 & n14361 ;
  assign n14363 = n13548 & n14362 ;
  assign n14364 = n512 & n14173 ;
  assign n14365 = ( n1526 & ~n8882 ) | ( n1526 & n12921 ) | ( ~n8882 & n12921 ) ;
  assign n14366 = n14365 ^ n9530 ^ 1'b0 ;
  assign n14367 = n8740 | n14366 ;
  assign n14368 = n1906 & ~n2278 ;
  assign n14369 = n14368 ^ n7645 ^ 1'b0 ;
  assign n14370 = ( ~n8795 & n14367 ) | ( ~n8795 & n14369 ) | ( n14367 & n14369 ) ;
  assign n14371 = n4680 ^ n2670 ^ 1'b0 ;
  assign n14372 = n1374 & ~n7065 ;
  assign n14373 = n14372 ^ n4518 ^ 1'b0 ;
  assign n14374 = ( n11138 & ~n11964 ) | ( n11138 & n14373 ) | ( ~n11964 & n14373 ) ;
  assign n14375 = n2324 | n5170 ;
  assign n14376 = n2829 | n8676 ;
  assign n14377 = n14375 | n14376 ;
  assign n14378 = n14377 ^ n11724 ^ 1'b0 ;
  assign n14379 = n11440 & n14378 ;
  assign n14381 = n4465 & ~n9973 ;
  assign n14380 = n6968 & n8834 ;
  assign n14382 = n14381 ^ n14380 ^ n4387 ;
  assign n14383 = n4559 & ~n14382 ;
  assign n14385 = ( n946 & ~n3221 ) | ( n946 & n4530 ) | ( ~n3221 & n4530 ) ;
  assign n14384 = ( n10800 & n12177 ) | ( n10800 & ~n12829 ) | ( n12177 & ~n12829 ) ;
  assign n14386 = n14385 ^ n14384 ^ n3730 ;
  assign n14387 = ( x180 & n3218 ) | ( x180 & n5404 ) | ( n3218 & n5404 ) ;
  assign n14388 = n7200 ^ n6123 ^ 1'b0 ;
  assign n14389 = n8673 | n14388 ;
  assign n14390 = ~n10118 & n12938 ;
  assign n14391 = n14389 & n14390 ;
  assign n14392 = ( n10420 & n14387 ) | ( n10420 & ~n14391 ) | ( n14387 & ~n14391 ) ;
  assign n14393 = ~n4145 & n7556 ;
  assign n14394 = ( n2084 & ~n7521 ) | ( n2084 & n10993 ) | ( ~n7521 & n10993 ) ;
  assign n14395 = ~n4622 & n14394 ;
  assign n14396 = n10662 & n14395 ;
  assign n14397 = ( n3381 & n14393 ) | ( n3381 & n14396 ) | ( n14393 & n14396 ) ;
  assign n14398 = ( n1463 & n3590 ) | ( n1463 & n4431 ) | ( n3590 & n4431 ) ;
  assign n14399 = n13385 & n14398 ;
  assign n14400 = n13109 ^ n9277 ^ 1'b0 ;
  assign n14401 = n14399 & ~n14400 ;
  assign n14402 = n3878 | n14401 ;
  assign n14406 = ( n984 & n13275 ) | ( n984 & ~n13543 ) | ( n13275 & ~n13543 ) ;
  assign n14407 = n14406 ^ n5666 ^ n3044 ;
  assign n14403 = n4195 & ~n6763 ;
  assign n14404 = n14403 ^ n2025 ^ 1'b0 ;
  assign n14405 = ~n8638 & n14404 ;
  assign n14408 = n14407 ^ n14405 ^ n1108 ;
  assign n14409 = n11103 ^ n1784 ^ 1'b0 ;
  assign n14410 = n4239 & n14409 ;
  assign n14411 = n14410 ^ n8661 ^ 1'b0 ;
  assign n14412 = ~n5212 & n14411 ;
  assign n14413 = ( ~n660 & n5912 ) | ( ~n660 & n8803 ) | ( n5912 & n8803 ) ;
  assign n14414 = n13319 ^ n5170 ^ 1'b0 ;
  assign n14415 = n14414 ^ n4301 ^ 1'b0 ;
  assign n14416 = n14415 ^ n9506 ^ n1408 ;
  assign n14417 = n308 | n6456 ;
  assign n14418 = n14416 & ~n14417 ;
  assign n14419 = ( n11967 & n14413 ) | ( n11967 & ~n14418 ) | ( n14413 & ~n14418 ) ;
  assign n14426 = n12676 ^ n12198 ^ 1'b0 ;
  assign n14420 = n4422 | n8082 ;
  assign n14421 = n5262 ^ n1058 ^ 1'b0 ;
  assign n14422 = n3587 | n14421 ;
  assign n14423 = n9066 & n14422 ;
  assign n14424 = n14420 & ~n14423 ;
  assign n14425 = n14424 ^ n2750 ^ 1'b0 ;
  assign n14427 = n14426 ^ n14425 ^ 1'b0 ;
  assign n14428 = n1802 & ~n14427 ;
  assign n14429 = ( n14412 & n14419 ) | ( n14412 & n14428 ) | ( n14419 & n14428 ) ;
  assign n14430 = n900 | n6462 ;
  assign n14431 = n13072 | n14430 ;
  assign n14432 = ~n4343 & n6139 ;
  assign n14433 = n477 & ~n10417 ;
  assign n14434 = n14432 & ~n14433 ;
  assign n14435 = ~n14431 & n14434 ;
  assign n14436 = n14435 ^ n8378 ^ n4596 ;
  assign n14437 = n6134 ^ n5065 ^ n4497 ;
  assign n14438 = ( n8457 & n13250 ) | ( n8457 & ~n14437 ) | ( n13250 & ~n14437 ) ;
  assign n14439 = n14197 ^ n10377 ^ 1'b0 ;
  assign n14440 = n14439 ^ n10261 ^ n1880 ;
  assign n14441 = n13506 ^ n13147 ^ n512 ;
  assign n14442 = x132 & ~n1669 ;
  assign n14443 = n14442 ^ n1384 ^ 1'b0 ;
  assign n14444 = n14443 ^ n3452 ^ n1510 ;
  assign n14445 = n2539 & n14444 ;
  assign n14446 = ~n6006 & n14445 ;
  assign n14447 = n613 & ~n7425 ;
  assign n14448 = n14446 | n14447 ;
  assign n14449 = n8994 | n14448 ;
  assign n14458 = x133 & n12199 ;
  assign n14459 = n10281 & n14458 ;
  assign n14452 = ( n2694 & n2737 ) | ( n2694 & ~n11589 ) | ( n2737 & ~n11589 ) ;
  assign n14453 = ~n6596 & n11271 ;
  assign n14454 = n14453 ^ n12476 ^ 1'b0 ;
  assign n14455 = ( n3608 & n14452 ) | ( n3608 & n14454 ) | ( n14452 & n14454 ) ;
  assign n14450 = n3833 & ~n4632 ;
  assign n14451 = n13002 & n14450 ;
  assign n14456 = n14455 ^ n14451 ^ 1'b0 ;
  assign n14457 = n10022 | n14456 ;
  assign n14460 = n14459 ^ n14457 ^ 1'b0 ;
  assign n14464 = ~n4618 & n5268 ;
  assign n14465 = n2874 & n14464 ;
  assign n14466 = n14465 ^ n5554 ^ n5518 ;
  assign n14467 = ~n9431 & n14466 ;
  assign n14468 = n14467 ^ n14250 ^ 1'b0 ;
  assign n14469 = ( x220 & ~n3647 ) | ( x220 & n14468 ) | ( ~n3647 & n14468 ) ;
  assign n14461 = ~n6100 & n7962 ;
  assign n14462 = n14461 ^ n10186 ^ n10120 ;
  assign n14463 = n6997 & ~n14462 ;
  assign n14470 = n14469 ^ n14463 ^ 1'b0 ;
  assign n14471 = n7605 ^ n5950 ^ 1'b0 ;
  assign n14472 = ( n4584 & ~n5912 ) | ( n4584 & n6613 ) | ( ~n5912 & n6613 ) ;
  assign n14473 = n14471 & ~n14472 ;
  assign n14474 = ~n5465 & n9404 ;
  assign n14475 = n4224 | n4401 ;
  assign n14476 = n6410 | n14475 ;
  assign n14477 = ~n3307 & n14476 ;
  assign n14478 = ( n1438 & ~n14474 ) | ( n1438 & n14477 ) | ( ~n14474 & n14477 ) ;
  assign n14479 = n14478 ^ n11167 ^ 1'b0 ;
  assign n14480 = n1828 | n9738 ;
  assign n14481 = n14480 ^ n5014 ^ 1'b0 ;
  assign n14482 = n8644 & ~n14481 ;
  assign n14483 = n4210 & n14482 ;
  assign n14484 = n12457 ^ n6850 ^ n940 ;
  assign n14485 = n10103 ^ n3531 ^ n343 ;
  assign n14486 = n14485 ^ n11542 ^ n4886 ;
  assign n14494 = ~n4501 & n8389 ;
  assign n14487 = n9919 ^ n6956 ^ 1'b0 ;
  assign n14488 = n5329 ^ n1301 ^ 1'b0 ;
  assign n14489 = n14487 & ~n14488 ;
  assign n14490 = n5345 ^ n598 ^ 1'b0 ;
  assign n14491 = ~n8103 & n14490 ;
  assign n14492 = n14491 ^ n5708 ^ n1544 ;
  assign n14493 = n14489 & ~n14492 ;
  assign n14495 = n14494 ^ n14493 ^ 1'b0 ;
  assign n14496 = n6209 & ~n14495 ;
  assign n14501 = n3946 & ~n4642 ;
  assign n14502 = n14501 ^ n6944 ^ 1'b0 ;
  assign n14503 = n1023 | n14502 ;
  assign n14499 = n1915 | n7988 ;
  assign n14500 = n14499 ^ n1826 ^ 1'b0 ;
  assign n14504 = n14503 ^ n14500 ^ n6477 ;
  assign n14497 = n11227 ^ n2494 ^ n1779 ;
  assign n14498 = n7748 & n14497 ;
  assign n14505 = n14504 ^ n14498 ^ 1'b0 ;
  assign n14507 = ~n1097 & n9974 ;
  assign n14508 = ~n1284 & n4734 ;
  assign n14509 = n14507 & n14508 ;
  assign n14506 = ( n495 & n4282 ) | ( n495 & ~n9282 ) | ( n4282 & ~n9282 ) ;
  assign n14510 = n14509 ^ n14506 ^ n5886 ;
  assign n14511 = ( ~n5826 & n6028 ) | ( ~n5826 & n13440 ) | ( n6028 & n13440 ) ;
  assign n14512 = n13223 | n14511 ;
  assign n14518 = n879 & ~n9790 ;
  assign n14519 = ~n13862 & n14518 ;
  assign n14520 = n14519 ^ n7559 ^ 1'b0 ;
  assign n14516 = ( n959 & n2759 ) | ( n959 & ~n4466 ) | ( n2759 & ~n4466 ) ;
  assign n14513 = n10468 ^ n1014 ^ 1'b0 ;
  assign n14514 = n3535 & n14513 ;
  assign n14515 = n14514 ^ n10977 ^ n3643 ;
  assign n14517 = n14516 ^ n14515 ^ n7044 ;
  assign n14521 = n14520 ^ n14517 ^ 1'b0 ;
  assign n14522 = ~n3666 & n14521 ;
  assign n14523 = ( ~n310 & n2320 ) | ( ~n310 & n7780 ) | ( n2320 & n7780 ) ;
  assign n14524 = ( n702 & n13728 ) | ( n702 & ~n14523 ) | ( n13728 & ~n14523 ) ;
  assign n14525 = n1969 & ~n13506 ;
  assign n14526 = n3775 & n14525 ;
  assign n14527 = n14526 ^ n948 ^ 1'b0 ;
  assign n14528 = n6440 & ~n14527 ;
  assign n14529 = n6973 & n14528 ;
  assign n14530 = n5003 ^ n1627 ^ 1'b0 ;
  assign n14531 = n11746 & n14530 ;
  assign n14532 = n394 & n5129 ;
  assign n14533 = n14532 ^ n5980 ^ 1'b0 ;
  assign n14534 = n2169 ^ n1319 ^ n577 ;
  assign n14535 = n12420 & ~n14534 ;
  assign n14536 = ~n3329 & n14535 ;
  assign n14537 = n6486 & n14536 ;
  assign n14540 = ( n2948 & ~n8904 ) | ( n2948 & n8907 ) | ( ~n8904 & n8907 ) ;
  assign n14538 = n4488 ^ n297 ^ 1'b0 ;
  assign n14539 = n7658 | n14538 ;
  assign n14541 = n14540 ^ n14539 ^ 1'b0 ;
  assign n14542 = ( n981 & ~n4387 ) | ( n981 & n4942 ) | ( ~n4387 & n4942 ) ;
  assign n14543 = n14542 ^ n3290 ^ 1'b0 ;
  assign n14544 = ( n1136 & n7954 ) | ( n1136 & ~n14543 ) | ( n7954 & ~n14543 ) ;
  assign n14551 = ~n437 & n5005 ;
  assign n14552 = ~n2149 & n14551 ;
  assign n14545 = n8587 ^ n7862 ^ n3827 ;
  assign n14546 = n4058 & n8309 ;
  assign n14547 = n5283 & n14546 ;
  assign n14548 = n14547 ^ n2025 ^ n1460 ;
  assign n14549 = n14545 & ~n14548 ;
  assign n14550 = ~n11482 & n14549 ;
  assign n14553 = n14552 ^ n14550 ^ n3013 ;
  assign n14554 = ( n7442 & ~n14544 ) | ( n7442 & n14553 ) | ( ~n14544 & n14553 ) ;
  assign n14555 = n8017 ^ n4022 ^ 1'b0 ;
  assign n14556 = n14555 ^ n286 ^ 1'b0 ;
  assign n14557 = n2896 & n14556 ;
  assign n14558 = n3835 & n14557 ;
  assign n14559 = n4571 & n14558 ;
  assign n14560 = n2895 ^ n1537 ^ n599 ;
  assign n14561 = n14560 ^ n11516 ^ n11121 ;
  assign n14562 = ( n838 & n2296 ) | ( n838 & ~n5651 ) | ( n2296 & ~n5651 ) ;
  assign n14563 = n14562 ^ n2801 ^ 1'b0 ;
  assign n14564 = n436 | n1139 ;
  assign n14565 = n14564 ^ n5397 ^ 1'b0 ;
  assign n14566 = n693 & n6555 ;
  assign n14567 = ~n14565 & n14566 ;
  assign n14568 = n3335 & ~n14567 ;
  assign n14580 = n14322 ^ n4866 ^ n4305 ;
  assign n14569 = n3591 ^ n2541 ^ 1'b0 ;
  assign n14570 = n14140 ^ n3252 ^ 1'b0 ;
  assign n14571 = n14569 & ~n14570 ;
  assign n14572 = ( n3919 & n5102 ) | ( n3919 & n6422 ) | ( n5102 & n6422 ) ;
  assign n14573 = n5231 | n7887 ;
  assign n14574 = n14573 ^ n1235 ^ 1'b0 ;
  assign n14575 = ~n14572 & n14574 ;
  assign n14576 = ~n14571 & n14575 ;
  assign n14577 = n3527 ^ n3210 ^ 1'b0 ;
  assign n14578 = n7920 & ~n14577 ;
  assign n14579 = n14576 & n14578 ;
  assign n14581 = n14580 ^ n14579 ^ n8487 ;
  assign n14582 = n3142 ^ x189 ^ 1'b0 ;
  assign n14583 = ~n6889 & n14582 ;
  assign n14584 = n2737 & n14583 ;
  assign n14585 = ~n1061 & n14584 ;
  assign n14588 = n14585 ^ n4659 ^ n2252 ;
  assign n14586 = n10208 ^ n8232 ^ n4020 ;
  assign n14587 = ( n954 & n14585 ) | ( n954 & ~n14586 ) | ( n14585 & ~n14586 ) ;
  assign n14589 = n14588 ^ n14587 ^ 1'b0 ;
  assign n14590 = n1012 ^ x118 ^ 1'b0 ;
  assign n14591 = ~n13212 & n14590 ;
  assign n14592 = n9681 | n14591 ;
  assign n14593 = ( ~n2592 & n3129 ) | ( ~n2592 & n7358 ) | ( n3129 & n7358 ) ;
  assign n14594 = ( n4103 & n10859 ) | ( n4103 & n14593 ) | ( n10859 & n14593 ) ;
  assign n14595 = n14543 ^ n5501 ^ n3983 ;
  assign n14596 = n14595 ^ n1560 ^ 1'b0 ;
  assign n14597 = n3200 | n10191 ;
  assign n14598 = n4345 & ~n14597 ;
  assign n14605 = n6673 ^ n5127 ^ n644 ;
  assign n14606 = n2117 | n14605 ;
  assign n14607 = n9314 | n14606 ;
  assign n14608 = n13117 ^ n4809 ^ 1'b0 ;
  assign n14609 = n14607 & ~n14608 ;
  assign n14599 = n9577 ^ n4286 ^ 1'b0 ;
  assign n14600 = n3426 & ~n14599 ;
  assign n14601 = ~n7459 & n14600 ;
  assign n14602 = n14601 ^ n9022 ^ 1'b0 ;
  assign n14603 = n11009 ^ n4936 ^ n3671 ;
  assign n14604 = ~n14602 & n14603 ;
  assign n14610 = n14609 ^ n14604 ^ 1'b0 ;
  assign n14611 = n12046 ^ n1280 ^ 1'b0 ;
  assign n14612 = n3851 & ~n12337 ;
  assign n14613 = n12147 ^ n4564 ^ n3095 ;
  assign n14614 = n5184 ^ n1077 ^ n673 ;
  assign n14615 = n11619 ^ n7964 ^ 1'b0 ;
  assign n14616 = n7497 & ~n14615 ;
  assign n14617 = n14614 & n14616 ;
  assign n14618 = ~n4785 & n14617 ;
  assign n14619 = n11010 ^ n5645 ^ n2675 ;
  assign n14620 = ( ~x7 & n6682 ) | ( ~x7 & n14619 ) | ( n6682 & n14619 ) ;
  assign n14621 = n4619 | n14620 ;
  assign n14622 = n11243 ^ n1395 ^ n1050 ;
  assign n14624 = n1544 | n9265 ;
  assign n14623 = n2690 & ~n12916 ;
  assign n14625 = n14624 ^ n14623 ^ 1'b0 ;
  assign n14626 = ( n10272 & ~n14622 ) | ( n10272 & n14625 ) | ( ~n14622 & n14625 ) ;
  assign n14627 = n14626 ^ n5726 ^ n3808 ;
  assign n14628 = n4754 & ~n14627 ;
  assign n14629 = ( n3729 & n4754 ) | ( n3729 & ~n14223 ) | ( n4754 & ~n14223 ) ;
  assign n14630 = ~n2014 & n6118 ;
  assign n14631 = n1239 | n2196 ;
  assign n14632 = n14631 ^ n924 ^ 1'b0 ;
  assign n14633 = n5316 & ~n14632 ;
  assign n14634 = n14633 ^ n6695 ^ n5673 ;
  assign n14635 = ( ~n6837 & n10385 ) | ( ~n6837 & n13490 ) | ( n10385 & n13490 ) ;
  assign n14636 = n4757 ^ x68 ^ 1'b0 ;
  assign n14637 = ~n3502 & n6003 ;
  assign n14638 = n8657 & n14637 ;
  assign n14639 = n14638 ^ n14081 ^ n10869 ;
  assign n14640 = n2091 | n2722 ;
  assign n14641 = n14639 | n14640 ;
  assign n14642 = n14636 & ~n14641 ;
  assign n14647 = ~n3562 & n5966 ;
  assign n14648 = n4880 & n14647 ;
  assign n14649 = n13006 & ~n14648 ;
  assign n14650 = n14649 ^ n1643 ^ 1'b0 ;
  assign n14643 = n10315 ^ n6850 ^ 1'b0 ;
  assign n14644 = n8926 | n14643 ;
  assign n14645 = n3615 & ~n14644 ;
  assign n14646 = x55 | n14645 ;
  assign n14651 = n14650 ^ n14646 ^ 1'b0 ;
  assign n14652 = n2305 | n3550 ;
  assign n14653 = n5889 & ~n14652 ;
  assign n14654 = n14653 ^ n900 ^ 1'b0 ;
  assign n14655 = n9985 ^ n1747 ^ 1'b0 ;
  assign n14656 = n14654 & n14655 ;
  assign n14657 = x66 & n14656 ;
  assign n14658 = ~n3436 & n7390 ;
  assign n14659 = ~n8079 & n14658 ;
  assign n14660 = n14659 ^ n13039 ^ n341 ;
  assign n14661 = n3142 & ~n13131 ;
  assign n14662 = ~n3019 & n13074 ;
  assign n14663 = n4728 & n14662 ;
  assign n14664 = n2670 & ~n4315 ;
  assign n14666 = ~n3934 & n4746 ;
  assign n14665 = n7708 ^ n3494 ^ n818 ;
  assign n14667 = n14666 ^ n14665 ^ n12416 ;
  assign n14668 = n14667 ^ n12304 ^ 1'b0 ;
  assign n14669 = ( n3804 & n8110 ) | ( n3804 & n14668 ) | ( n8110 & n14668 ) ;
  assign n14682 = n8199 ^ n6558 ^ n3961 ;
  assign n14679 = n7214 ^ n2172 ^ 1'b0 ;
  assign n14680 = n14679 ^ n5208 ^ 1'b0 ;
  assign n14676 = n2637 ^ n668 ^ 1'b0 ;
  assign n14677 = ~n3346 & n14676 ;
  assign n14678 = ~n1815 & n14677 ;
  assign n14681 = n14680 ^ n14678 ^ 1'b0 ;
  assign n14683 = n14682 ^ n14681 ^ n2782 ;
  assign n14671 = ( n3388 & n3563 ) | ( n3388 & n4056 ) | ( n3563 & n4056 ) ;
  assign n14672 = x154 & ~n14671 ;
  assign n14673 = n14672 ^ n5004 ^ 1'b0 ;
  assign n14674 = n14673 ^ n3413 ^ n2015 ;
  assign n14670 = n7576 ^ n5720 ^ 1'b0 ;
  assign n14675 = n14674 ^ n14670 ^ 1'b0 ;
  assign n14684 = n14683 ^ n14675 ^ n12029 ;
  assign n14685 = n9665 ^ n7131 ^ n1886 ;
  assign n14686 = ( ~n12508 & n13025 ) | ( ~n12508 & n14685 ) | ( n13025 & n14685 ) ;
  assign n14687 = n13157 ^ n8537 ^ 1'b0 ;
  assign n14688 = n13404 | n14687 ;
  assign n14689 = n2931 & ~n14688 ;
  assign n14690 = n6196 & n14689 ;
  assign n14691 = n9558 ^ n8876 ^ 1'b0 ;
  assign n14692 = ~n14690 & n14691 ;
  assign n14693 = n9656 ^ n2232 ^ 1'b0 ;
  assign n14694 = x32 & ~n1721 ;
  assign n14695 = ~n2448 & n14694 ;
  assign n14696 = n14695 ^ n13871 ^ n5924 ;
  assign n14697 = n6003 ^ n2874 ^ 1'b0 ;
  assign n14698 = n6521 & ~n11079 ;
  assign n14699 = n1415 & n14698 ;
  assign n14700 = n14697 & n14699 ;
  assign n14701 = n14700 ^ n9911 ^ 1'b0 ;
  assign n14702 = n14696 | n14701 ;
  assign n14703 = ~n10196 & n11774 ;
  assign n14704 = n14702 & n14703 ;
  assign n14705 = n3525 | n11782 ;
  assign n14706 = n14705 ^ n5033 ^ 1'b0 ;
  assign n14707 = ~n1734 & n2973 ;
  assign n14708 = n3073 & n14707 ;
  assign n14709 = n14706 & n14708 ;
  assign n14710 = n14709 ^ n1856 ^ 1'b0 ;
  assign n14711 = n5465 ^ n1076 ^ 1'b0 ;
  assign n14712 = n10946 ^ n4681 ^ n2664 ;
  assign n14713 = n14712 ^ n11257 ^ n6916 ;
  assign n14714 = ( ~n2157 & n3779 ) | ( ~n2157 & n6808 ) | ( n3779 & n6808 ) ;
  assign n14715 = ~n5365 & n8586 ;
  assign n14716 = n14715 ^ n6637 ^ 1'b0 ;
  assign n14720 = ~n3861 & n4249 ;
  assign n14721 = n7376 & n14720 ;
  assign n14722 = n2632 | n13583 ;
  assign n14723 = n4756 | n14722 ;
  assign n14724 = ( n1832 & ~n7399 ) | ( n1832 & n14723 ) | ( ~n7399 & n14723 ) ;
  assign n14725 = ( ~n7474 & n14721 ) | ( ~n7474 & n14724 ) | ( n14721 & n14724 ) ;
  assign n14717 = n2835 & n5624 ;
  assign n14718 = n14717 ^ x97 ^ 1'b0 ;
  assign n14719 = n1841 & n14718 ;
  assign n14726 = n14725 ^ n14719 ^ 1'b0 ;
  assign n14727 = n14716 | n14726 ;
  assign n14728 = n729 & n3274 ;
  assign n14729 = ( n5482 & n11779 ) | ( n5482 & n14728 ) | ( n11779 & n14728 ) ;
  assign n14730 = ( n1777 & n1836 ) | ( n1777 & n4268 ) | ( n1836 & n4268 ) ;
  assign n14731 = n14155 & ~n14730 ;
  assign n14732 = ~n9630 & n14731 ;
  assign n14733 = n6388 ^ n2579 ^ 1'b0 ;
  assign n14734 = ~n9658 & n14733 ;
  assign n14735 = n7316 ^ n2655 ^ 1'b0 ;
  assign n14736 = n12931 ^ n5797 ^ 1'b0 ;
  assign n14737 = ~n4577 & n14736 ;
  assign n14738 = n1048 | n5443 ;
  assign n14739 = n7894 & ~n14738 ;
  assign n14740 = ~n4191 & n6509 ;
  assign n14741 = n14740 ^ n14665 ^ n11101 ;
  assign n14742 = ( n14737 & n14739 ) | ( n14737 & ~n14741 ) | ( n14739 & ~n14741 ) ;
  assign n14748 = ( ~n567 & n6726 ) | ( ~n567 & n7297 ) | ( n6726 & n7297 ) ;
  assign n14743 = ~n7676 & n8143 ;
  assign n14744 = n14743 ^ n2291 ^ 1'b0 ;
  assign n14745 = ( x227 & n1548 ) | ( x227 & ~n8533 ) | ( n1548 & ~n8533 ) ;
  assign n14746 = n14744 | n14745 ;
  assign n14747 = n14746 ^ n12120 ^ 1'b0 ;
  assign n14749 = n14748 ^ n14747 ^ 1'b0 ;
  assign n14750 = ( ~x147 & n2918 ) | ( ~x147 & n9569 ) | ( n2918 & n9569 ) ;
  assign n14751 = n14750 ^ n11322 ^ n10915 ;
  assign n14752 = n14751 ^ n5069 ^ n3206 ;
  assign n14753 = n5470 & ~n6214 ;
  assign n14754 = n14753 ^ x222 ^ 1'b0 ;
  assign n14755 = ( n12160 & n13584 ) | ( n12160 & n14754 ) | ( n13584 & n14754 ) ;
  assign n14756 = ~n1465 & n5316 ;
  assign n14757 = n3036 ^ n717 ^ x186 ;
  assign n14758 = n14756 | n14757 ;
  assign n14759 = n14758 ^ n7072 ^ 1'b0 ;
  assign n14760 = n13424 & n14759 ;
  assign n14761 = n14760 ^ n8299 ^ 1'b0 ;
  assign n14762 = ~n3370 & n7669 ;
  assign n14763 = n14762 ^ n2576 ^ 1'b0 ;
  assign n14764 = ( n4927 & n9092 ) | ( n4927 & n12558 ) | ( n9092 & n12558 ) ;
  assign n14765 = n13519 ^ n8666 ^ 1'b0 ;
  assign n14766 = n4980 & n14765 ;
  assign n14767 = n14766 ^ n4613 ^ 1'b0 ;
  assign n14768 = n14767 ^ n7591 ^ 1'b0 ;
  assign n14769 = ( ~n991 & n12606 ) | ( ~n991 & n13934 ) | ( n12606 & n13934 ) ;
  assign n14780 = n1189 & n2417 ;
  assign n14781 = n14780 ^ n554 ^ 1'b0 ;
  assign n14782 = ~n2010 & n6355 ;
  assign n14783 = n14781 & n14782 ;
  assign n14784 = n14783 ^ n11773 ^ n280 ;
  assign n14772 = n3624 ^ n2503 ^ n962 ;
  assign n14771 = n3790 & n4385 ;
  assign n14773 = n14772 ^ n14771 ^ 1'b0 ;
  assign n14774 = ~n6704 & n9647 ;
  assign n14775 = n14774 ^ n6411 ^ 1'b0 ;
  assign n14776 = ( n10869 & ~n14773 ) | ( n10869 & n14775 ) | ( ~n14773 & n14775 ) ;
  assign n14770 = ( n1109 & ~n2433 ) | ( n1109 & n9887 ) | ( ~n2433 & n9887 ) ;
  assign n14777 = n14776 ^ n14770 ^ n4617 ;
  assign n14778 = n2438 & ~n14777 ;
  assign n14779 = n10560 & ~n14778 ;
  assign n14785 = n14784 ^ n14779 ^ 1'b0 ;
  assign n14786 = n1172 ^ n332 ^ 1'b0 ;
  assign n14787 = x0 & n14786 ;
  assign n14788 = n4639 & n14787 ;
  assign n14789 = n9990 & ~n14788 ;
  assign n14790 = n14789 ^ n5077 ^ 1'b0 ;
  assign n14791 = ( n4244 & ~n4975 ) | ( n4244 & n14790 ) | ( ~n4975 & n14790 ) ;
  assign n14798 = n11752 ^ n6917 ^ n2476 ;
  assign n14792 = n3233 & n6618 ;
  assign n14793 = ~n4381 & n14792 ;
  assign n14794 = n5595 & ~n9971 ;
  assign n14795 = ~x140 & n14794 ;
  assign n14796 = n4412 & ~n14795 ;
  assign n14797 = n14793 & n14796 ;
  assign n14799 = n14798 ^ n14797 ^ n2114 ;
  assign n14800 = n1026 & ~n2310 ;
  assign n14801 = ( n2791 & ~n13096 ) | ( n2791 & n14800 ) | ( ~n13096 & n14800 ) ;
  assign n14802 = n6501 & n6502 ;
  assign n14803 = n14801 & n14802 ;
  assign n14804 = ~n2190 & n14803 ;
  assign n14805 = n1449 & n2167 ;
  assign n14806 = n14805 ^ n6106 ^ 1'b0 ;
  assign n14807 = ( ~n5906 & n10099 ) | ( ~n5906 & n13932 ) | ( n10099 & n13932 ) ;
  assign n14810 = n1195 | n2574 ;
  assign n14811 = n14810 ^ n3989 ^ 1'b0 ;
  assign n14808 = n1993 ^ n1943 ^ 1'b0 ;
  assign n14809 = ~n6317 & n14808 ;
  assign n14812 = n14811 ^ n14809 ^ n11028 ;
  assign n14813 = ( ~n2020 & n6014 ) | ( ~n2020 & n11099 ) | ( n6014 & n11099 ) ;
  assign n14814 = n3154 & n6997 ;
  assign n14815 = ( n4385 & n14813 ) | ( n4385 & ~n14814 ) | ( n14813 & ~n14814 ) ;
  assign n14816 = n14815 ^ n5140 ^ n2360 ;
  assign n14821 = n8876 ^ n5411 ^ n2662 ;
  assign n14822 = ( n3392 & n4398 ) | ( n3392 & ~n5076 ) | ( n4398 & ~n5076 ) ;
  assign n14823 = n14822 ^ n2779 ^ n1495 ;
  assign n14824 = ~n14821 & n14823 ;
  assign n14817 = n11137 ^ x15 ^ 1'b0 ;
  assign n14818 = n11009 & ~n14817 ;
  assign n14819 = ( n6984 & n10078 ) | ( n6984 & n14818 ) | ( n10078 & n14818 ) ;
  assign n14820 = n14819 ^ n854 ^ 1'b0 ;
  assign n14825 = n14824 ^ n14820 ^ n2422 ;
  assign n14826 = n6338 ^ n2472 ^ n1953 ;
  assign n14827 = ( n1254 & n5539 ) | ( n1254 & ~n10077 ) | ( n5539 & ~n10077 ) ;
  assign n14828 = n14827 ^ n9238 ^ n3945 ;
  assign n14829 = ( ~n6393 & n14826 ) | ( ~n6393 & n14828 ) | ( n14826 & n14828 ) ;
  assign n14830 = ( n2776 & n3300 ) | ( n2776 & n7976 ) | ( n3300 & n7976 ) ;
  assign n14831 = n14830 ^ n3064 ^ 1'b0 ;
  assign n14835 = n2690 & n4312 ;
  assign n14836 = ~n1909 & n14835 ;
  assign n14837 = n14836 ^ n3494 ^ 1'b0 ;
  assign n14832 = ( n1647 & n4551 ) | ( n1647 & n8792 ) | ( n4551 & n8792 ) ;
  assign n14833 = n14832 ^ n3518 ^ n1479 ;
  assign n14834 = n14833 ^ n6413 ^ n1998 ;
  assign n14838 = n14837 ^ n14834 ^ n6888 ;
  assign n14839 = ~n5923 & n11115 ;
  assign n14840 = n14839 ^ n599 ^ 1'b0 ;
  assign n14841 = x54 | n7850 ;
  assign n14842 = ( n3958 & n14840 ) | ( n3958 & ~n14841 ) | ( n14840 & ~n14841 ) ;
  assign n14843 = n3295 ^ n1627 ^ 1'b0 ;
  assign n14844 = n12658 | n14843 ;
  assign n14845 = n8216 ^ n5867 ^ 1'b0 ;
  assign n14846 = ~n609 & n14845 ;
  assign n14847 = n14844 & n14846 ;
  assign n14848 = n11844 ^ n11011 ^ n6457 ;
  assign n14849 = n7378 & n14848 ;
  assign n14850 = n10820 ^ n1791 ^ 1'b0 ;
  assign n14851 = n10020 | n14850 ;
  assign n14852 = n9892 ^ n3413 ^ n2492 ;
  assign n14853 = n14814 & n14852 ;
  assign n14854 = n14853 ^ x7 ^ 1'b0 ;
  assign n14855 = n8389 & ~n14854 ;
  assign n14856 = n7719 & n14855 ;
  assign n14857 = ( n4480 & n7403 ) | ( n4480 & ~n14856 ) | ( n7403 & ~n14856 ) ;
  assign n14858 = n14857 ^ n14279 ^ n11833 ;
  assign n14860 = ( n518 & n3449 ) | ( n518 & ~n4660 ) | ( n3449 & ~n4660 ) ;
  assign n14861 = ( n7349 & n11034 ) | ( n7349 & ~n14860 ) | ( n11034 & ~n14860 ) ;
  assign n14859 = ( ~n1491 & n4067 ) | ( ~n1491 & n10621 ) | ( n4067 & n10621 ) ;
  assign n14862 = n14861 ^ n14859 ^ 1'b0 ;
  assign n14863 = n6532 & ~n14862 ;
  assign n14864 = n14627 & n14863 ;
  assign n14865 = ~n6180 & n14864 ;
  assign n14866 = n3404 & ~n9671 ;
  assign n14867 = n1157 & n14866 ;
  assign n14868 = ~n10649 & n14867 ;
  assign n14869 = ~n5069 & n6932 ;
  assign n14870 = ~n14868 & n14869 ;
  assign n14871 = n13427 | n14870 ;
  assign n14876 = n1690 & ~n3292 ;
  assign n14877 = n14876 ^ n6611 ^ 1'b0 ;
  assign n14878 = n1524 | n4846 ;
  assign n14879 = n14878 ^ n835 ^ 1'b0 ;
  assign n14880 = ( ~n9299 & n14877 ) | ( ~n9299 & n14879 ) | ( n14877 & n14879 ) ;
  assign n14873 = ( x46 & ~n534 ) | ( x46 & n4722 ) | ( ~n534 & n4722 ) ;
  assign n14872 = ~n2793 & n8224 ;
  assign n14874 = n14873 ^ n14872 ^ 1'b0 ;
  assign n14875 = ( n4020 & n4804 ) | ( n4020 & n14874 ) | ( n4804 & n14874 ) ;
  assign n14881 = n14880 ^ n14875 ^ n2141 ;
  assign n14882 = n8206 & ~n12520 ;
  assign n14883 = n14882 ^ n4043 ^ 1'b0 ;
  assign n14884 = ( n1101 & n6139 ) | ( n1101 & n14883 ) | ( n6139 & n14883 ) ;
  assign n14885 = n12344 ^ n779 ^ n329 ;
  assign n14886 = ( ~x86 & n5007 ) | ( ~x86 & n14885 ) | ( n5007 & n14885 ) ;
  assign n14887 = ~n8897 & n14886 ;
  assign n14888 = n8724 ^ n4006 ^ 1'b0 ;
  assign n14889 = ~n14887 & n14888 ;
  assign n14890 = n10488 ^ n10136 ^ n1081 ;
  assign n14891 = ( ~x218 & n8743 ) | ( ~x218 & n12040 ) | ( n8743 & n12040 ) ;
  assign n14892 = ( ~n7179 & n14890 ) | ( ~n7179 & n14891 ) | ( n14890 & n14891 ) ;
  assign n14893 = ( n9654 & ~n11112 ) | ( n9654 & n14892 ) | ( ~n11112 & n14892 ) ;
  assign n14894 = n4594 | n7233 ;
  assign n14895 = n14894 ^ n10454 ^ 1'b0 ;
  assign n14896 = n9201 ^ n7763 ^ n4157 ;
  assign n14897 = n14896 ^ n6553 ^ 1'b0 ;
  assign n14898 = ~n10140 & n14897 ;
  assign n14899 = ~n4884 & n8763 ;
  assign n14900 = n4927 & n14899 ;
  assign n14901 = ( ~n1391 & n5718 ) | ( ~n1391 & n11275 ) | ( n5718 & n11275 ) ;
  assign n14902 = ( ~n9842 & n14900 ) | ( ~n9842 & n14901 ) | ( n14900 & n14901 ) ;
  assign n14903 = n6871 & ~n11867 ;
  assign n14904 = n11242 ^ n2639 ^ 1'b0 ;
  assign n14905 = n14904 ^ n12576 ^ n5424 ;
  assign n14906 = ( n14902 & ~n14903 ) | ( n14902 & n14905 ) | ( ~n14903 & n14905 ) ;
  assign n14907 = n8452 ^ n5085 ^ 1'b0 ;
  assign n14908 = n673 & n14907 ;
  assign n14909 = n6424 & n14908 ;
  assign n14911 = ~n1635 & n7669 ;
  assign n14912 = n9273 & n14911 ;
  assign n14910 = x174 & ~n12463 ;
  assign n14913 = n14912 ^ n14910 ^ 1'b0 ;
  assign n14914 = ~n5311 & n14913 ;
  assign n14915 = n4262 ^ n2661 ^ 1'b0 ;
  assign n14916 = n14914 & ~n14915 ;
  assign n14917 = n465 ^ x251 ^ 1'b0 ;
  assign n14918 = n4516 ^ n1710 ^ 1'b0 ;
  assign n14919 = n1721 | n14918 ;
  assign n14920 = ( n8512 & n14917 ) | ( n8512 & n14919 ) | ( n14917 & n14919 ) ;
  assign n14921 = ( n4367 & n9050 ) | ( n4367 & n9700 ) | ( n9050 & n9700 ) ;
  assign n14922 = ( n912 & n4348 ) | ( n912 & n11887 ) | ( n4348 & n11887 ) ;
  assign n14923 = ~n1588 & n9677 ;
  assign n14924 = n10667 ^ n3340 ^ n859 ;
  assign n14925 = x104 & n1260 ;
  assign n14926 = n4396 & n14925 ;
  assign n14927 = ( ~n447 & n5609 ) | ( ~n447 & n12840 ) | ( n5609 & n12840 ) ;
  assign n14928 = n5965 ^ n2885 ^ 1'b0 ;
  assign n14929 = ( n2917 & n8136 ) | ( n2917 & n14928 ) | ( n8136 & n14928 ) ;
  assign n14930 = n5236 | n7582 ;
  assign n14931 = n14930 ^ n8616 ^ 1'b0 ;
  assign n14932 = n14783 | n14931 ;
  assign n14933 = n14929 | n14932 ;
  assign n14934 = ( n7011 & n14927 ) | ( n7011 & ~n14933 ) | ( n14927 & ~n14933 ) ;
  assign n14935 = n14926 & n14934 ;
  assign n14936 = n13999 ^ n13984 ^ n5581 ;
  assign n14937 = n6267 ^ n1841 ^ n1005 ;
  assign n14938 = n6726 ^ n733 ^ n467 ;
  assign n14939 = ( ~n4696 & n8103 ) | ( ~n4696 & n11440 ) | ( n8103 & n11440 ) ;
  assign n14940 = ( ~n9990 & n14938 ) | ( ~n9990 & n14939 ) | ( n14938 & n14939 ) ;
  assign n14942 = n1858 | n4251 ;
  assign n14941 = n9116 ^ n2671 ^ n696 ;
  assign n14943 = n14942 ^ n14941 ^ n14653 ;
  assign n14944 = ( n363 & n7821 ) | ( n363 & ~n14185 ) | ( n7821 & ~n14185 ) ;
  assign n14945 = n14944 ^ n2495 ^ 1'b0 ;
  assign n14946 = x25 & n11574 ;
  assign n14947 = n2426 ^ x93 ^ 1'b0 ;
  assign n14948 = n14946 & ~n14947 ;
  assign n14949 = n14164 ^ n3585 ^ 1'b0 ;
  assign n14950 = n5044 & ~n14949 ;
  assign n14951 = x21 | n303 ;
  assign n14952 = n14951 ^ n12586 ^ n8887 ;
  assign n14953 = n14950 & n14952 ;
  assign n14954 = n14953 ^ n3740 ^ 1'b0 ;
  assign n14955 = x222 & n14954 ;
  assign n14956 = ~n8394 & n14955 ;
  assign n14957 = ~n2997 & n5559 ;
  assign n14958 = ~n4065 & n14957 ;
  assign n14959 = n14958 ^ n1703 ^ 1'b0 ;
  assign n14960 = n2027 | n14959 ;
  assign n14961 = n7600 & n14960 ;
  assign n14962 = ( ~n3246 & n4340 ) | ( ~n3246 & n5234 ) | ( n4340 & n5234 ) ;
  assign n14963 = ~n5010 & n14962 ;
  assign n14964 = n14963 ^ n1419 ^ 1'b0 ;
  assign n14965 = n8615 & ~n14964 ;
  assign n14968 = n5699 & n5934 ;
  assign n14969 = ~n7845 & n14968 ;
  assign n14970 = ~n6389 & n14969 ;
  assign n14966 = n8342 ^ n3761 ^ 1'b0 ;
  assign n14967 = n14966 ^ n740 ^ 1'b0 ;
  assign n14971 = n14970 ^ n14967 ^ n8494 ;
  assign n14983 = n2727 & n9662 ;
  assign n14984 = n14983 ^ n2796 ^ 1'b0 ;
  assign n14982 = n2409 & n6197 ;
  assign n14985 = n14984 ^ n14982 ^ 1'b0 ;
  assign n14979 = n8877 ^ n7772 ^ 1'b0 ;
  assign n14980 = n285 | n14979 ;
  assign n14972 = n5733 | n14891 ;
  assign n14973 = n14972 ^ n10337 ^ 1'b0 ;
  assign n14974 = n14973 ^ n6621 ^ 1'b0 ;
  assign n14975 = n11249 | n14974 ;
  assign n14976 = ( n2779 & n7355 ) | ( n2779 & ~n10766 ) | ( n7355 & ~n10766 ) ;
  assign n14977 = ( n7306 & n13348 ) | ( n7306 & ~n14976 ) | ( n13348 & ~n14976 ) ;
  assign n14978 = ( n6061 & ~n14975 ) | ( n6061 & n14977 ) | ( ~n14975 & n14977 ) ;
  assign n14981 = n14980 ^ n14978 ^ n1773 ;
  assign n14986 = n14985 ^ n14981 ^ n10226 ;
  assign n14987 = n6076 & n7117 ;
  assign n14988 = n14987 ^ n8336 ^ n816 ;
  assign n14989 = n3747 & n14988 ;
  assign n14990 = n3234 & ~n6838 ;
  assign n14991 = n14990 ^ n5470 ^ 1'b0 ;
  assign n14992 = n14991 ^ n11354 ^ x66 ;
  assign n14993 = n14992 ^ n9596 ^ 1'b0 ;
  assign n14994 = ( n335 & n5765 ) | ( n335 & n10645 ) | ( n5765 & n10645 ) ;
  assign n14995 = n14994 ^ n9579 ^ n5332 ;
  assign n14996 = n12633 ^ n1304 ^ n489 ;
  assign n14997 = n2398 & n3593 ;
  assign n14998 = n14997 ^ n4348 ^ 1'b0 ;
  assign n14999 = n7470 ^ n2108 ^ 1'b0 ;
  assign n15000 = n14998 | n14999 ;
  assign n15001 = n3383 & n4680 ;
  assign n15002 = ( ~n14996 & n15000 ) | ( ~n14996 & n15001 ) | ( n15000 & n15001 ) ;
  assign n15003 = n9101 & n9875 ;
  assign n15004 = ~n12540 & n15003 ;
  assign n15005 = n15004 ^ n1995 ^ 1'b0 ;
  assign n15006 = n2930 | n15005 ;
  assign n15007 = n2374 & ~n13371 ;
  assign n15008 = n15007 ^ n12376 ^ 1'b0 ;
  assign n15009 = n15008 ^ n14819 ^ n12106 ;
  assign n15010 = ( ~n1138 & n6076 ) | ( ~n1138 & n15009 ) | ( n6076 & n15009 ) ;
  assign n15011 = n1696 & ~n4042 ;
  assign n15012 = n15011 ^ n8942 ^ 1'b0 ;
  assign n15013 = ( n1173 & n1220 ) | ( n1173 & n5598 ) | ( n1220 & n5598 ) ;
  assign n15014 = ( n10380 & ~n15012 ) | ( n10380 & n15013 ) | ( ~n15012 & n15013 ) ;
  assign n15015 = ( n8119 & ~n9879 ) | ( n8119 & n15014 ) | ( ~n9879 & n15014 ) ;
  assign n15016 = ~n744 & n15015 ;
  assign n15017 = ( n885 & ~n5991 ) | ( n885 & n9275 ) | ( ~n5991 & n9275 ) ;
  assign n15018 = ~n7815 & n15017 ;
  assign n15019 = n15018 ^ n1662 ^ 1'b0 ;
  assign n15020 = n4902 & ~n15019 ;
  assign n15025 = n7491 ^ n6248 ^ 1'b0 ;
  assign n15026 = x118 & ~n15025 ;
  assign n15022 = n5269 ^ n2304 ^ n994 ;
  assign n15023 = n7406 | n15022 ;
  assign n15021 = n8849 ^ n407 ^ 1'b0 ;
  assign n15024 = n15023 ^ n15021 ^ n4830 ;
  assign n15027 = n15026 ^ n15024 ^ n14195 ;
  assign n15028 = n8473 ^ n5741 ^ 1'b0 ;
  assign n15029 = ~n7322 & n15028 ;
  assign n15030 = n7542 | n15029 ;
  assign n15031 = n13724 & ~n15030 ;
  assign n15032 = ( ~n2247 & n5986 ) | ( ~n2247 & n15031 ) | ( n5986 & n15031 ) ;
  assign n15033 = ( n8374 & n10160 ) | ( n8374 & n12640 ) | ( n10160 & n12640 ) ;
  assign n15034 = ( n3813 & n10197 ) | ( n3813 & n12537 ) | ( n10197 & n12537 ) ;
  assign n15035 = n15034 ^ n12013 ^ n2260 ;
  assign n15036 = ( n9332 & n15033 ) | ( n9332 & ~n15035 ) | ( n15033 & ~n15035 ) ;
  assign n15037 = n6622 ^ n5033 ^ n1023 ;
  assign n15038 = n10344 ^ n9928 ^ 1'b0 ;
  assign n15039 = n11642 & n15038 ;
  assign n15040 = n15039 ^ n4227 ^ n2608 ;
  assign n15041 = n15040 ^ n10191 ^ 1'b0 ;
  assign n15042 = ( n6401 & n15037 ) | ( n6401 & n15041 ) | ( n15037 & n15041 ) ;
  assign n15043 = n15036 & n15042 ;
  assign n15044 = n11367 & n15043 ;
  assign n15045 = ( x139 & n2425 ) | ( x139 & n4989 ) | ( n2425 & n4989 ) ;
  assign n15046 = n788 | n15045 ;
  assign n15049 = n2155 | n3400 ;
  assign n15050 = n15049 ^ n4693 ^ 1'b0 ;
  assign n15047 = n5329 & n5955 ;
  assign n15048 = ~n9346 & n15047 ;
  assign n15051 = n15050 ^ n15048 ^ n8563 ;
  assign n15052 = n2576 ^ n1146 ^ 1'b0 ;
  assign n15053 = n1990 & ~n15052 ;
  assign n15054 = ( n1158 & ~n1881 ) | ( n1158 & n15053 ) | ( ~n1881 & n15053 ) ;
  assign n15055 = ~n723 & n3644 ;
  assign n15057 = ( n5341 & ~n6450 ) | ( n5341 & n6857 ) | ( ~n6450 & n6857 ) ;
  assign n15058 = n307 & ~n6625 ;
  assign n15059 = ~n15057 & n15058 ;
  assign n15056 = n9027 ^ n1203 ^ 1'b0 ;
  assign n15060 = n15059 ^ n15056 ^ n11363 ;
  assign n15061 = n7911 ^ n6612 ^ 1'b0 ;
  assign n15062 = ~n6868 & n15061 ;
  assign n15063 = n1333 | n15062 ;
  assign n15064 = ( ~n3474 & n5745 ) | ( ~n3474 & n10012 ) | ( n5745 & n10012 ) ;
  assign n15065 = ( n1998 & n10631 ) | ( n1998 & ~n15064 ) | ( n10631 & ~n15064 ) ;
  assign n15066 = n1994 & ~n11106 ;
  assign n15067 = n15066 ^ n8924 ^ 1'b0 ;
  assign n15068 = ( n15063 & n15065 ) | ( n15063 & n15067 ) | ( n15065 & n15067 ) ;
  assign n15069 = n7646 | n12291 ;
  assign n15070 = n15069 ^ n9885 ^ 1'b0 ;
  assign n15071 = n15070 ^ n824 ^ 1'b0 ;
  assign n15072 = n15071 ^ n8052 ^ 1'b0 ;
  assign n15073 = x13 & n6862 ;
  assign n15074 = n4774 & n15073 ;
  assign n15075 = ( n2012 & ~n2055 ) | ( n2012 & n14818 ) | ( ~n2055 & n14818 ) ;
  assign n15076 = n15075 ^ n11275 ^ 1'b0 ;
  assign n15077 = ( ~n3987 & n15074 ) | ( ~n3987 & n15076 ) | ( n15074 & n15076 ) ;
  assign n15078 = ~n3364 & n6220 ;
  assign n15079 = ( ~n1935 & n10090 ) | ( ~n1935 & n15078 ) | ( n10090 & n15078 ) ;
  assign n15080 = n15077 & n15079 ;
  assign n15081 = n5935 & n15080 ;
  assign n15082 = n6114 & ~n11961 ;
  assign n15083 = n15082 ^ n3962 ^ 1'b0 ;
  assign n15085 = x23 & ~n6193 ;
  assign n15086 = ~n12221 & n15085 ;
  assign n15084 = n8732 ^ n6990 ^ n3411 ;
  assign n15087 = n15086 ^ n15084 ^ n4155 ;
  assign n15088 = ( n5197 & n15083 ) | ( n5197 & n15087 ) | ( n15083 & n15087 ) ;
  assign n15089 = n10229 ^ n8978 ^ n4360 ;
  assign n15090 = n12739 | n15089 ;
  assign n15091 = ~n11961 & n15090 ;
  assign n15092 = n15091 ^ n343 ^ 1'b0 ;
  assign n15093 = n11054 & n15092 ;
  assign n15094 = ~n8899 & n13918 ;
  assign n15095 = ~n4162 & n15094 ;
  assign n15096 = n5856 & ~n15095 ;
  assign n15097 = n15096 ^ n7023 ^ 1'b0 ;
  assign n15098 = n454 & n2628 ;
  assign n15099 = n12858 ^ n2324 ^ 1'b0 ;
  assign n15100 = n2765 & ~n6635 ;
  assign n15101 = n15100 ^ n13423 ^ 1'b0 ;
  assign n15102 = ~n1912 & n15101 ;
  assign n15104 = n13190 ^ n6086 ^ n4288 ;
  assign n15105 = ( x62 & n11436 ) | ( x62 & n15104 ) | ( n11436 & n15104 ) ;
  assign n15103 = ~n7605 & n9719 ;
  assign n15106 = n15105 ^ n15103 ^ 1'b0 ;
  assign n15107 = n11786 | n15106 ;
  assign n15108 = n11190 & ~n15107 ;
  assign n15113 = n6934 ^ n6867 ^ 1'b0 ;
  assign n15114 = n13497 & n15113 ;
  assign n15109 = n3833 & ~n4488 ;
  assign n15110 = n4844 & n5025 ;
  assign n15111 = ~n9291 & n15110 ;
  assign n15112 = n15109 | n15111 ;
  assign n15115 = n15114 ^ n15112 ^ n534 ;
  assign n15116 = ( n735 & ~n14302 ) | ( n735 & n15115 ) | ( ~n14302 & n15115 ) ;
  assign n15117 = n12765 ^ n1442 ^ 1'b0 ;
  assign n15118 = n8764 ^ n2123 ^ 1'b0 ;
  assign n15119 = n2698 & ~n4950 ;
  assign n15120 = n15119 ^ n7442 ^ 1'b0 ;
  assign n15121 = ( n1334 & n8755 ) | ( n1334 & ~n15120 ) | ( n8755 & ~n15120 ) ;
  assign n15122 = n6088 & ~n15121 ;
  assign n15123 = ~n2770 & n6186 ;
  assign n15124 = n4003 & n15123 ;
  assign n15125 = n9996 ^ n9409 ^ 1'b0 ;
  assign n15126 = n13188 & ~n15125 ;
  assign n15127 = n15126 ^ n9692 ^ n6781 ;
  assign n15128 = n14902 ^ n6366 ^ 1'b0 ;
  assign n15129 = ~n8973 & n15128 ;
  assign n15130 = ~n10099 & n15129 ;
  assign n15131 = n12221 ^ n7453 ^ n2387 ;
  assign n15132 = n5723 & n15131 ;
  assign n15133 = n15132 ^ n2406 ^ 1'b0 ;
  assign n15134 = n2142 & n15133 ;
  assign n15135 = ( n539 & n7951 ) | ( n539 & n15134 ) | ( n7951 & n15134 ) ;
  assign n15136 = n765 & ~n11255 ;
  assign n15137 = ( ~n2063 & n7487 ) | ( ~n2063 & n9767 ) | ( n7487 & n9767 ) ;
  assign n15138 = ( n6355 & n14900 ) | ( n6355 & n15137 ) | ( n14900 & n15137 ) ;
  assign n15139 = ( ~x244 & n3605 ) | ( ~x244 & n10467 ) | ( n3605 & n10467 ) ;
  assign n15140 = n10292 ^ n10121 ^ 1'b0 ;
  assign n15141 = n14049 & ~n15140 ;
  assign n15142 = ~n15139 & n15141 ;
  assign n15148 = n7654 ^ n6842 ^ 1'b0 ;
  assign n15143 = n4716 & ~n7870 ;
  assign n15144 = ~n3931 & n15143 ;
  assign n15145 = n15144 ^ n6138 ^ 1'b0 ;
  assign n15146 = ~n2592 & n15145 ;
  assign n15147 = ~n11429 & n15146 ;
  assign n15149 = n15148 ^ n15147 ^ n2362 ;
  assign n15150 = n7640 & n14426 ;
  assign n15151 = n15150 ^ n13385 ^ 1'b0 ;
  assign n15152 = n15151 ^ n12473 ^ 1'b0 ;
  assign n15153 = n10696 & n15152 ;
  assign n15154 = ( x183 & n13529 ) | ( x183 & n15153 ) | ( n13529 & n15153 ) ;
  assign n15155 = n8484 ^ n4313 ^ 1'b0 ;
  assign n15156 = n13113 ^ n2085 ^ 1'b0 ;
  assign n15157 = n10206 & ~n15156 ;
  assign n15158 = n15157 ^ n1877 ^ 1'b0 ;
  assign n15159 = n10368 & n15158 ;
  assign n15160 = n15159 ^ n14493 ^ 1'b0 ;
  assign n15161 = ~n15155 & n15160 ;
  assign n15162 = ( n2069 & ~n8287 ) | ( n2069 & n13232 ) | ( ~n8287 & n13232 ) ;
  assign n15163 = ( n11242 & ~n14478 ) | ( n11242 & n15162 ) | ( ~n14478 & n15162 ) ;
  assign n15164 = n10727 ^ n8452 ^ n3178 ;
  assign n15165 = n15164 ^ n12754 ^ 1'b0 ;
  assign n15166 = n15165 ^ n3537 ^ 1'b0 ;
  assign n15167 = n15163 & n15166 ;
  assign n15168 = n3433 & ~n7710 ;
  assign n15169 = n15168 ^ n10633 ^ n9851 ;
  assign n15170 = n12508 & n15169 ;
  assign n15171 = n14116 ^ n5759 ^ n1747 ;
  assign n15172 = ( n374 & n5383 ) | ( n374 & ~n6193 ) | ( n5383 & ~n6193 ) ;
  assign n15174 = ( n3625 & ~n4498 ) | ( n3625 & n7308 ) | ( ~n4498 & n7308 ) ;
  assign n15173 = n2934 & ~n13529 ;
  assign n15175 = n15174 ^ n15173 ^ 1'b0 ;
  assign n15176 = n15175 ^ n346 ^ 1'b0 ;
  assign n15177 = n15172 & n15176 ;
  assign n15178 = n5313 & ~n11972 ;
  assign n15179 = ~n4737 & n15178 ;
  assign n15180 = ( x224 & n536 ) | ( x224 & n2541 ) | ( n536 & n2541 ) ;
  assign n15183 = n12797 ^ n12046 ^ 1'b0 ;
  assign n15181 = ( ~n1948 & n3621 ) | ( ~n1948 & n6696 ) | ( n3621 & n6696 ) ;
  assign n15182 = ( n4368 & ~n6829 ) | ( n4368 & n15181 ) | ( ~n6829 & n15181 ) ;
  assign n15184 = n15183 ^ n15182 ^ n5467 ;
  assign n15185 = ( n7181 & n15180 ) | ( n7181 & ~n15184 ) | ( n15180 & ~n15184 ) ;
  assign n15186 = n13815 ^ n9770 ^ n6398 ;
  assign n15187 = n15186 ^ n7782 ^ 1'b0 ;
  assign n15188 = ( ~n13379 & n15185 ) | ( ~n13379 & n15187 ) | ( n15185 & n15187 ) ;
  assign n15189 = ( ~n2029 & n2146 ) | ( ~n2029 & n6389 ) | ( n2146 & n6389 ) ;
  assign n15191 = n13192 ^ x168 ^ 1'b0 ;
  assign n15190 = n12551 ^ n2111 ^ 1'b0 ;
  assign n15192 = n15191 ^ n15190 ^ 1'b0 ;
  assign n15193 = n13815 & ~n15192 ;
  assign n15194 = ~n4501 & n7085 ;
  assign n15195 = n1423 & ~n15194 ;
  assign n15196 = n15195 ^ n10606 ^ 1'b0 ;
  assign n15197 = ~n8424 & n15196 ;
  assign n15198 = ~n13955 & n15197 ;
  assign n15203 = ( n6735 & n8530 ) | ( n6735 & ~n10377 ) | ( n8530 & ~n10377 ) ;
  assign n15199 = n6826 & n11392 ;
  assign n15200 = ~n2182 & n15199 ;
  assign n15201 = ( n11556 & n13622 ) | ( n11556 & ~n15200 ) | ( n13622 & ~n15200 ) ;
  assign n15202 = n15201 ^ n8087 ^ n2192 ;
  assign n15204 = n15203 ^ n15202 ^ n9409 ;
  assign n15205 = n15088 ^ n9604 ^ 1'b0 ;
  assign n15206 = ~n15204 & n15205 ;
  assign n15214 = ( ~n4046 & n12549 ) | ( ~n4046 & n14497 ) | ( n12549 & n14497 ) ;
  assign n15207 = n2215 & n2500 ;
  assign n15208 = n15207 ^ n4661 ^ 1'b0 ;
  assign n15209 = n3333 & ~n15208 ;
  assign n15210 = n15209 ^ n7096 ^ n1561 ;
  assign n15211 = n15210 ^ n11510 ^ n1187 ;
  assign n15212 = n3353 | n15211 ;
  assign n15213 = n15212 ^ n11068 ^ 1'b0 ;
  assign n15215 = n15214 ^ n15213 ^ 1'b0 ;
  assign n15216 = n11383 ^ n10500 ^ 1'b0 ;
  assign n15217 = n12456 ^ n11942 ^ n11525 ;
  assign n15218 = n15217 ^ n8217 ^ x83 ;
  assign n15219 = ( n895 & n3517 ) | ( n895 & n8942 ) | ( n3517 & n8942 ) ;
  assign n15220 = n11972 ^ n2117 ^ 1'b0 ;
  assign n15221 = ( n3529 & n3896 ) | ( n3529 & ~n12057 ) | ( n3896 & ~n12057 ) ;
  assign n15222 = n14854 ^ n8895 ^ 1'b0 ;
  assign n15223 = n15221 & n15222 ;
  assign n15224 = n6223 ^ x135 ^ 1'b0 ;
  assign n15229 = ( n1293 & n11672 ) | ( n1293 & ~n12252 ) | ( n11672 & ~n12252 ) ;
  assign n15225 = n11060 ^ n4775 ^ n2478 ;
  assign n15226 = ( n2126 & n2793 ) | ( n2126 & ~n6712 ) | ( n2793 & ~n6712 ) ;
  assign n15227 = n3585 & n15226 ;
  assign n15228 = ~n15225 & n15227 ;
  assign n15230 = n15229 ^ n15228 ^ n349 ;
  assign n15231 = n3426 & ~n14228 ;
  assign n15232 = n15231 ^ n575 ^ 1'b0 ;
  assign n15239 = n15041 ^ n14015 ^ 1'b0 ;
  assign n15240 = ~n11239 & n15239 ;
  assign n15234 = n9220 ^ n3057 ^ n1702 ;
  assign n15233 = n5145 | n9885 ;
  assign n15235 = n15234 ^ n15233 ^ 1'b0 ;
  assign n15236 = n7398 & ~n15235 ;
  assign n15237 = ~n6315 & n15236 ;
  assign n15238 = n8723 & ~n15237 ;
  assign n15241 = n15240 ^ n15238 ^ 1'b0 ;
  assign n15242 = ~n11001 & n13472 ;
  assign n15243 = n11514 ^ n3379 ^ n1734 ;
  assign n15244 = n6373 ^ n4824 ^ n2218 ;
  assign n15245 = n6080 & n15244 ;
  assign n15246 = n13353 ^ n8577 ^ 1'b0 ;
  assign n15247 = n15246 ^ n7929 ^ n1798 ;
  assign n15251 = n3379 & n6286 ;
  assign n15252 = ~n5149 & n15251 ;
  assign n15248 = n2838 | n4129 ;
  assign n15249 = n7900 & ~n15248 ;
  assign n15250 = n15249 ^ n8350 ^ n2718 ;
  assign n15253 = n15252 ^ n15250 ^ n2960 ;
  assign n15256 = ( x207 & n7783 ) | ( x207 & ~n8606 ) | ( n7783 & ~n8606 ) ;
  assign n15257 = n1113 & n15256 ;
  assign n15258 = n15257 ^ x107 ^ 1'b0 ;
  assign n15254 = n3257 & n7372 ;
  assign n15255 = n15254 ^ n2131 ^ 1'b0 ;
  assign n15259 = n15258 ^ n15255 ^ n999 ;
  assign n15260 = ( n5399 & n6334 ) | ( n5399 & n10304 ) | ( n6334 & n10304 ) ;
  assign n15261 = n15260 ^ n4209 ^ n779 ;
  assign n15263 = n8217 ^ n2731 ^ 1'b0 ;
  assign n15264 = n15263 ^ n6585 ^ n6360 ;
  assign n15262 = n10635 ^ n332 ^ 1'b0 ;
  assign n15265 = n15264 ^ n15262 ^ 1'b0 ;
  assign n15266 = n15261 | n15265 ;
  assign n15267 = n15266 ^ n2357 ^ 1'b0 ;
  assign n15268 = n2351 | n7524 ;
  assign n15269 = n15268 ^ n4991 ^ 1'b0 ;
  assign n15270 = n15269 ^ n15207 ^ n5297 ;
  assign n15271 = n8847 & ~n9723 ;
  assign n15272 = n15271 ^ n4815 ^ 1'b0 ;
  assign n15273 = n15270 | n15272 ;
  assign n15274 = n15273 ^ n9259 ^ 1'b0 ;
  assign n15275 = n6216 & n15274 ;
  assign n15276 = n12640 ^ n609 ^ x39 ;
  assign n15277 = ( n311 & ~n3853 ) | ( n311 & n15276 ) | ( ~n3853 & n15276 ) ;
  assign n15278 = n11767 | n15277 ;
  assign n15279 = ~n9143 & n15278 ;
  assign n15280 = n2107 & ~n12912 ;
  assign n15281 = n15280 ^ n2811 ^ 1'b0 ;
  assign n15282 = n5500 & n5760 ;
  assign n15283 = n780 | n6872 ;
  assign n15284 = n15282 & ~n15283 ;
  assign n15285 = n12766 ^ n11151 ^ n10444 ;
  assign n15286 = n11881 ^ n10104 ^ n2183 ;
  assign n15287 = n15286 ^ n4500 ^ 1'b0 ;
  assign n15288 = n7435 ^ n3722 ^ 1'b0 ;
  assign n15289 = ( n10761 & n11830 ) | ( n10761 & n15288 ) | ( n11830 & n15288 ) ;
  assign n15290 = n15289 ^ n10383 ^ n6734 ;
  assign n15291 = n15290 ^ n10012 ^ 1'b0 ;
  assign n15292 = n10920 ^ n3031 ^ n1583 ;
  assign n15293 = n14648 ^ n4505 ^ 1'b0 ;
  assign n15294 = n15292 | n15293 ;
  assign n15295 = n2882 & ~n15294 ;
  assign n15296 = n15295 ^ x231 ^ 1'b0 ;
  assign n15297 = n13722 | n15207 ;
  assign n15298 = n15297 ^ n9159 ^ n7932 ;
  assign n15299 = n14762 ^ n11011 ^ 1'b0 ;
  assign n15300 = n8861 ^ n3557 ^ n2309 ;
  assign n15301 = n5321 ^ n730 ^ n556 ;
  assign n15302 = ( n11071 & n15300 ) | ( n11071 & n15301 ) | ( n15300 & n15301 ) ;
  assign n15303 = ~n3716 & n13097 ;
  assign n15304 = n15303 ^ n3904 ^ 1'b0 ;
  assign n15305 = ( n2950 & ~n3906 ) | ( n2950 & n4257 ) | ( ~n3906 & n4257 ) ;
  assign n15306 = n15304 | n15305 ;
  assign n15307 = n15302 & ~n15306 ;
  assign n15308 = n4251 & ~n15307 ;
  assign n15309 = n15308 ^ n10061 ^ 1'b0 ;
  assign n15310 = n13877 | n15309 ;
  assign n15311 = n9974 & ~n15310 ;
  assign n15312 = n13154 ^ n6200 ^ n2027 ;
  assign n15313 = n1575 ^ n1156 ^ 1'b0 ;
  assign n15314 = n7827 ^ n5747 ^ 1'b0 ;
  assign n15315 = n15314 ^ n7944 ^ 1'b0 ;
  assign n15316 = n2278 | n15315 ;
  assign n15317 = ( n2851 & n15313 ) | ( n2851 & ~n15316 ) | ( n15313 & ~n15316 ) ;
  assign n15318 = n10244 ^ n7325 ^ 1'b0 ;
  assign n15319 = ( n3470 & n6242 ) | ( n3470 & ~n15318 ) | ( n6242 & ~n15318 ) ;
  assign n15320 = n15319 ^ n13971 ^ 1'b0 ;
  assign n15321 = n368 & ~n15320 ;
  assign n15322 = n15321 ^ n9496 ^ n6633 ;
  assign n15323 = n4671 ^ n1000 ^ 1'b0 ;
  assign n15324 = n15323 ^ x92 ^ 1'b0 ;
  assign n15325 = n5791 ^ n4776 ^ 1'b0 ;
  assign n15326 = ( n2131 & n3849 ) | ( n2131 & n15325 ) | ( n3849 & n15325 ) ;
  assign n15327 = n15326 ^ n2472 ^ 1'b0 ;
  assign n15328 = ~n7213 & n15327 ;
  assign n15329 = n11265 ^ n6338 ^ 1'b0 ;
  assign n15330 = n9693 & ~n15329 ;
  assign n15331 = ~n10191 & n14466 ;
  assign n15332 = ~n6435 & n15331 ;
  assign n15333 = n3249 & ~n11736 ;
  assign n15334 = ~n6993 & n15333 ;
  assign n15335 = n15334 ^ n8996 ^ n286 ;
  assign n15336 = n15335 ^ n14823 ^ n11110 ;
  assign n15337 = ~n15332 & n15336 ;
  assign n15338 = n12052 ^ n10292 ^ 1'b0 ;
  assign n15339 = n5847 ^ n2152 ^ 1'b0 ;
  assign n15340 = ~n733 & n15339 ;
  assign n15341 = n15338 | n15340 ;
  assign n15342 = n8653 ^ n4552 ^ 1'b0 ;
  assign n15343 = n8391 & n15342 ;
  assign n15344 = n11219 & n11492 ;
  assign n15345 = n15344 ^ n4613 ^ 1'b0 ;
  assign n15346 = n2200 | n13030 ;
  assign n15347 = n15346 ^ n12442 ^ n9857 ;
  assign n15348 = n15347 ^ n4441 ^ 1'b0 ;
  assign n15349 = ~n8751 & n15348 ;
  assign n15350 = n15349 ^ n495 ^ 1'b0 ;
  assign n15351 = n4129 | n9290 ;
  assign n15352 = n10917 ^ n5412 ^ n4234 ;
  assign n15353 = ( n2250 & n7752 ) | ( n2250 & n14671 ) | ( n7752 & n14671 ) ;
  assign n15354 = n15353 ^ n6784 ^ n4884 ;
  assign n15355 = n15354 ^ n13216 ^ 1'b0 ;
  assign n15356 = n14660 | n15355 ;
  assign n15357 = n13617 ^ n5396 ^ 1'b0 ;
  assign n15358 = ~n816 & n13627 ;
  assign n15359 = n15358 ^ n1935 ^ 1'b0 ;
  assign n15360 = n12605 ^ n4104 ^ n429 ;
  assign n15361 = n4464 & ~n15360 ;
  assign n15362 = n15361 ^ n13192 ^ 1'b0 ;
  assign n15364 = n12959 ^ n9570 ^ 1'b0 ;
  assign n15363 = ( ~n2187 & n3367 ) | ( ~n2187 & n6728 ) | ( n3367 & n6728 ) ;
  assign n15365 = n15364 ^ n15363 ^ 1'b0 ;
  assign n15366 = ( x72 & n10654 ) | ( x72 & n10820 ) | ( n10654 & n10820 ) ;
  assign n15367 = n2970 ^ n1319 ^ 1'b0 ;
  assign n15368 = n8309 & n15367 ;
  assign n15369 = n370 | n3985 ;
  assign n15370 = n15369 ^ n7846 ^ 1'b0 ;
  assign n15371 = n15368 & n15370 ;
  assign n15372 = n15366 & n15371 ;
  assign n15373 = n7207 ^ n5512 ^ n526 ;
  assign n15374 = ( n2376 & n14653 ) | ( n2376 & ~n14730 ) | ( n14653 & ~n14730 ) ;
  assign n15375 = n15374 ^ n11884 ^ n3721 ;
  assign n15376 = ( n3459 & n15373 ) | ( n3459 & n15375 ) | ( n15373 & n15375 ) ;
  assign n15377 = n8195 | n11082 ;
  assign n15378 = n4396 ^ n1026 ^ 1'b0 ;
  assign n15379 = n15378 ^ n9531 ^ n3996 ;
  assign n15380 = n15379 ^ n3283 ^ n2480 ;
  assign n15381 = n1442 | n2591 ;
  assign n15382 = n15381 ^ n4569 ^ 1'b0 ;
  assign n15383 = n12332 ^ n10238 ^ n6214 ;
  assign n15384 = n15383 ^ x108 ^ 1'b0 ;
  assign n15385 = n13292 & n14385 ;
  assign n15386 = n15385 ^ n11492 ^ 1'b0 ;
  assign n15387 = x202 | n1538 ;
  assign n15399 = x62 & n333 ;
  assign n15400 = ~n5417 & n15399 ;
  assign n15401 = n15400 ^ n3433 ^ n1883 ;
  assign n15402 = n15401 ^ n13974 ^ n12431 ;
  assign n15394 = n3208 ^ n1368 ^ 1'b0 ;
  assign n15395 = ( ~n1681 & n14481 ) | ( ~n1681 & n15394 ) | ( n14481 & n15394 ) ;
  assign n15396 = ( n4624 & n5523 ) | ( n4624 & n8371 ) | ( n5523 & n8371 ) ;
  assign n15397 = n15396 ^ n7217 ^ 1'b0 ;
  assign n15398 = n15395 | n15397 ;
  assign n15388 = n4425 ^ n1651 ^ 1'b0 ;
  assign n15389 = n10550 & ~n15388 ;
  assign n15390 = n15389 ^ n1045 ^ 1'b0 ;
  assign n15391 = n15390 ^ n13077 ^ n1777 ;
  assign n15392 = n11517 ^ n10429 ^ 1'b0 ;
  assign n15393 = n15391 & ~n15392 ;
  assign n15403 = n15402 ^ n15398 ^ n15393 ;
  assign n15404 = n8078 & ~n15403 ;
  assign n15405 = n10212 & n15404 ;
  assign n15406 = n10060 & n10063 ;
  assign n15409 = n7638 ^ n1767 ^ 1'b0 ;
  assign n15407 = n5048 ^ n4275 ^ 1'b0 ;
  assign n15408 = ( n937 & n3543 ) | ( n937 & n15407 ) | ( n3543 & n15407 ) ;
  assign n15410 = n15409 ^ n15408 ^ n8183 ;
  assign n15411 = ( n4365 & ~n15406 ) | ( n4365 & n15410 ) | ( ~n15406 & n15410 ) ;
  assign n15416 = n440 & ~n7483 ;
  assign n15417 = ~n2847 & n15416 ;
  assign n15418 = ~n8877 & n15417 ;
  assign n15419 = ( n7433 & n15057 ) | ( n7433 & n15418 ) | ( n15057 & n15418 ) ;
  assign n15413 = ( ~n3262 & n5693 ) | ( ~n3262 & n6783 ) | ( n5693 & n6783 ) ;
  assign n15414 = n12432 ^ n6668 ^ 1'b0 ;
  assign n15415 = ( ~n11595 & n15413 ) | ( ~n11595 & n15414 ) | ( n15413 & n15414 ) ;
  assign n15412 = ~n2497 & n14446 ;
  assign n15420 = n15419 ^ n15415 ^ n15412 ;
  assign n15421 = x106 & x246 ;
  assign n15422 = ~n1838 & n15421 ;
  assign n15423 = ( ~n1047 & n2528 ) | ( ~n1047 & n15422 ) | ( n2528 & n15422 ) ;
  assign n15424 = ( n2841 & n7463 ) | ( n2841 & n15423 ) | ( n7463 & n15423 ) ;
  assign n15425 = n13594 ^ n9948 ^ n7812 ;
  assign n15426 = n9213 ^ n4980 ^ n2553 ;
  assign n15427 = n15426 ^ n327 ^ x208 ;
  assign n15428 = n15425 & n15427 ;
  assign n15429 = n15428 ^ n14355 ^ n11086 ;
  assign n15434 = ~n2218 & n11622 ;
  assign n15435 = n10529 | n15434 ;
  assign n15436 = n15435 ^ n14624 ^ 1'b0 ;
  assign n15430 = n12378 ^ n8145 ^ 1'b0 ;
  assign n15431 = ~n4952 & n15430 ;
  assign n15432 = n15401 & n15431 ;
  assign n15433 = ~n380 & n15432 ;
  assign n15437 = n15436 ^ n15433 ^ 1'b0 ;
  assign n15438 = n15429 | n15437 ;
  assign n15439 = n10185 | n11056 ;
  assign n15440 = n6800 ^ n2640 ^ 1'b0 ;
  assign n15441 = n6829 | n15440 ;
  assign n15442 = n15441 ^ n2178 ^ 1'b0 ;
  assign n15443 = n15442 ^ n9583 ^ 1'b0 ;
  assign n15444 = ( n1213 & n6048 ) | ( n1213 & ~n8257 ) | ( n6048 & ~n8257 ) ;
  assign n15445 = n15396 & n15444 ;
  assign n15446 = n15443 | n15445 ;
  assign n15447 = ~n1510 & n11117 ;
  assign n15448 = n15447 ^ n14088 ^ n5636 ;
  assign n15449 = n3437 ^ n2198 ^ 1'b0 ;
  assign n15450 = ( n5600 & n6092 ) | ( n5600 & n11020 ) | ( n6092 & n11020 ) ;
  assign n15451 = ( n7232 & ~n15449 ) | ( n7232 & n15450 ) | ( ~n15449 & n15450 ) ;
  assign n15452 = ( n1293 & n14823 ) | ( n1293 & ~n15451 ) | ( n14823 & ~n15451 ) ;
  assign n15453 = ~n5385 & n7573 ;
  assign n15454 = n6329 & n15453 ;
  assign n15455 = ~n4313 & n15454 ;
  assign n15456 = n4925 & n11155 ;
  assign n15457 = n13846 & ~n15456 ;
  assign n15458 = n9887 ^ n9375 ^ n3359 ;
  assign n15459 = ~n2997 & n15458 ;
  assign n15460 = n15459 ^ n3892 ^ 1'b0 ;
  assign n15461 = ( n1125 & ~n5257 ) | ( n1125 & n6610 ) | ( ~n5257 & n6610 ) ;
  assign n15462 = n15460 & ~n15461 ;
  assign n15463 = n1410 & n15462 ;
  assign n15464 = n11298 ^ n10681 ^ n2014 ;
  assign n15465 = n9842 ^ n4624 ^ 1'b0 ;
  assign n15466 = ( n15463 & n15464 ) | ( n15463 & n15465 ) | ( n15464 & n15465 ) ;
  assign n15467 = ( n508 & n4448 ) | ( n508 & ~n4978 ) | ( n4448 & ~n4978 ) ;
  assign n15468 = n15467 ^ n10578 ^ 1'b0 ;
  assign n15469 = n2071 | n15468 ;
  assign n15470 = n15469 ^ n8228 ^ 1'b0 ;
  assign n15471 = n15470 ^ n14773 ^ n6993 ;
  assign n15472 = n4613 ^ n3329 ^ x129 ;
  assign n15473 = n15472 ^ n13555 ^ n6318 ;
  assign n15474 = n8939 ^ n2733 ^ n1002 ;
  assign n15475 = ( ~n2248 & n8482 ) | ( ~n2248 & n15427 ) | ( n8482 & n15427 ) ;
  assign n15476 = n5963 & n15475 ;
  assign n15477 = n3325 ^ n1068 ^ 1'b0 ;
  assign n15478 = n15476 | n15477 ;
  assign n15479 = ( n544 & n8581 ) | ( n544 & ~n13692 ) | ( n8581 & ~n13692 ) ;
  assign n15480 = ( n10371 & ~n15478 ) | ( n10371 & n15479 ) | ( ~n15478 & n15479 ) ;
  assign n15482 = n8733 ^ n2942 ^ 1'b0 ;
  assign n15481 = ( n2250 & ~n2820 ) | ( n2250 & n6520 ) | ( ~n2820 & n6520 ) ;
  assign n15483 = n15482 ^ n15481 ^ n3765 ;
  assign n15484 = n5670 | n9527 ;
  assign n15485 = ( n3297 & n7466 ) | ( n3297 & ~n15484 ) | ( n7466 & ~n15484 ) ;
  assign n15492 = n3482 ^ n1783 ^ 1'b0 ;
  assign n15493 = ~n8193 & n15492 ;
  assign n15494 = n15493 ^ n5595 ^ 1'b0 ;
  assign n15495 = n4547 ^ n1294 ^ n1278 ;
  assign n15496 = ( n3499 & ~n15494 ) | ( n3499 & n15495 ) | ( ~n15494 & n15495 ) ;
  assign n15486 = n5628 ^ n4752 ^ n3138 ;
  assign n15487 = n14773 ^ n2474 ^ 1'b0 ;
  assign n15488 = ( n6773 & n15486 ) | ( n6773 & n15487 ) | ( n15486 & n15487 ) ;
  assign n15489 = n15441 ^ n8852 ^ n5446 ;
  assign n15490 = n15489 ^ n13141 ^ 1'b0 ;
  assign n15491 = n15488 & ~n15490 ;
  assign n15497 = n15496 ^ n15491 ^ 1'b0 ;
  assign n15498 = n11301 ^ n2808 ^ x108 ;
  assign n15499 = n15498 ^ n9884 ^ n5342 ;
  assign n15500 = ( n5895 & ~n7075 ) | ( n5895 & n10150 ) | ( ~n7075 & n10150 ) ;
  assign n15501 = n15500 ^ n10534 ^ 1'b0 ;
  assign n15502 = n7702 ^ n6040 ^ n2372 ;
  assign n15503 = n322 | n10855 ;
  assign n15504 = n15503 ^ n6092 ^ n4022 ;
  assign n15505 = n15504 ^ n5714 ^ n1314 ;
  assign n15506 = n11192 & n15505 ;
  assign n15507 = ( n5723 & ~n15502 ) | ( n5723 & n15506 ) | ( ~n15502 & n15506 ) ;
  assign n15508 = n4325 & ~n11239 ;
  assign n15509 = x66 & n799 ;
  assign n15510 = ( x198 & x232 ) | ( x198 & ~n2584 ) | ( x232 & ~n2584 ) ;
  assign n15511 = n15510 ^ n5984 ^ 1'b0 ;
  assign n15512 = n14285 ^ x117 ^ 1'b0 ;
  assign n15513 = n3065 & n15512 ;
  assign n15514 = n15513 ^ n1736 ^ 1'b0 ;
  assign n15515 = n2511 | n7265 ;
  assign n15516 = n11901 | n15515 ;
  assign n15517 = n5665 & ~n10808 ;
  assign n15518 = n7428 ^ n6198 ^ n2347 ;
  assign n15519 = n15518 ^ n11155 ^ n6472 ;
  assign n15520 = ~n920 & n15519 ;
  assign n15521 = ~n15517 & n15520 ;
  assign n15522 = ~n13240 & n15521 ;
  assign n15523 = ( n9139 & n15516 ) | ( n9139 & n15522 ) | ( n15516 & n15522 ) ;
  assign n15524 = n8408 | n8501 ;
  assign n15525 = x2 & ~n8987 ;
  assign n15526 = n15525 ^ n8587 ^ 1'b0 ;
  assign n15527 = n15526 ^ n15353 ^ x197 ;
  assign n15528 = n12890 & ~n15527 ;
  assign n15529 = ~n1034 & n15528 ;
  assign n15530 = n15524 & n15529 ;
  assign n15531 = ( n880 & ~n2346 ) | ( n880 & n3554 ) | ( ~n2346 & n3554 ) ;
  assign n15532 = n15289 | n15531 ;
  assign n15533 = n15532 ^ n6148 ^ 1'b0 ;
  assign n15539 = n2644 ^ n1305 ^ n732 ;
  assign n15537 = n3268 | n7614 ;
  assign n15538 = n15537 ^ n1036 ^ 1'b0 ;
  assign n15540 = n15539 ^ n15538 ^ n751 ;
  assign n15534 = n6408 & ~n9724 ;
  assign n15535 = n15534 ^ n11798 ^ 1'b0 ;
  assign n15536 = ~n10898 & n15535 ;
  assign n15541 = n15540 ^ n15536 ^ 1'b0 ;
  assign n15542 = n15078 ^ n10440 ^ n3046 ;
  assign n15543 = ( n1894 & n13823 ) | ( n1894 & n15542 ) | ( n13823 & n15542 ) ;
  assign n15544 = n15543 ^ n4222 ^ n1105 ;
  assign n15550 = n1765 & n1836 ;
  assign n15551 = ( n2027 & ~n5349 ) | ( n2027 & n15550 ) | ( ~n5349 & n15550 ) ;
  assign n15552 = n15551 ^ n13030 ^ n9334 ;
  assign n15549 = n6626 & ~n11087 ;
  assign n15546 = n13397 ^ n8524 ^ n7578 ;
  assign n15547 = n15546 ^ n2405 ^ 1'b0 ;
  assign n15548 = n4771 & n15547 ;
  assign n15553 = n15552 ^ n15549 ^ n15548 ;
  assign n15545 = n12198 ^ n7093 ^ 1'b0 ;
  assign n15554 = n15553 ^ n15545 ^ n8791 ;
  assign n15555 = n10258 ^ n8486 ^ n4705 ;
  assign n15556 = ( n1103 & ~n9033 ) | ( n1103 & n14478 ) | ( ~n9033 & n14478 ) ;
  assign n15557 = n15556 ^ n7780 ^ 1'b0 ;
  assign n15558 = ~n4745 & n9896 ;
  assign n15559 = ~n14394 & n15558 ;
  assign n15560 = ~n4794 & n12766 ;
  assign n15561 = ( n1284 & n7023 ) | ( n1284 & ~n15560 ) | ( n7023 & ~n15560 ) ;
  assign n15562 = n13082 ^ n9185 ^ n2348 ;
  assign n15563 = n15562 ^ n6480 ^ 1'b0 ;
  assign n15564 = n15561 | n15563 ;
  assign n15567 = ( ~n1422 & n4139 ) | ( ~n1422 & n5675 ) | ( n4139 & n5675 ) ;
  assign n15565 = n6860 & n12931 ;
  assign n15566 = ~n4966 & n15565 ;
  assign n15568 = n15567 ^ n15566 ^ n1667 ;
  assign n15569 = ( n2933 & n7779 ) | ( n2933 & n15568 ) | ( n7779 & n15568 ) ;
  assign n15570 = ~x130 & n2620 ;
  assign n15571 = n2994 ^ n2651 ^ n2110 ;
  assign n15572 = ~n10400 & n15571 ;
  assign n15573 = n15572 ^ n917 ^ 1'b0 ;
  assign n15574 = ~n13150 & n15573 ;
  assign n15575 = n3638 ^ n2686 ^ x111 ;
  assign n15576 = n15575 ^ n12370 ^ n2433 ;
  assign n15577 = ( n3219 & n7736 ) | ( n3219 & ~n15576 ) | ( n7736 & ~n15576 ) ;
  assign n15578 = n8742 ^ n5097 ^ 1'b0 ;
  assign n15579 = n15577 & n15578 ;
  assign n15580 = n11982 ^ n4512 ^ 1'b0 ;
  assign n15581 = n15580 ^ n8954 ^ 1'b0 ;
  assign n15582 = n15579 & ~n15581 ;
  assign n15586 = n2960 ^ n625 ^ n401 ;
  assign n15583 = n7234 & ~n13430 ;
  assign n15584 = n15583 ^ n14051 ^ 1'b0 ;
  assign n15585 = n15584 ^ n6209 ^ n6129 ;
  assign n15587 = n15586 ^ n15585 ^ n5163 ;
  assign n15589 = n7827 ^ n493 ^ 1'b0 ;
  assign n15588 = n12238 ^ n8000 ^ n3770 ;
  assign n15590 = n15589 ^ n15588 ^ n13289 ;
  assign n15591 = ( n2393 & n3791 ) | ( n2393 & n7250 ) | ( n3791 & n7250 ) ;
  assign n15592 = n15591 ^ n14873 ^ n7162 ;
  assign n15593 = n15592 ^ n3662 ^ 1'b0 ;
  assign n15594 = n598 | n9282 ;
  assign n15595 = n15594 ^ n11597 ^ 1'b0 ;
  assign n15596 = n2293 & n3364 ;
  assign n15597 = n15596 ^ n10876 ^ n9404 ;
  assign n15598 = ( n4595 & n14507 ) | ( n4595 & ~n15597 ) | ( n14507 & ~n15597 ) ;
  assign n15599 = n12387 ^ n10247 ^ 1'b0 ;
  assign n15600 = n15598 & ~n15599 ;
  assign n15608 = n8945 ^ n5313 ^ n2283 ;
  assign n15607 = n1473 & ~n8338 ;
  assign n15609 = n15608 ^ n15607 ^ n12591 ;
  assign n15610 = n15609 ^ n8459 ^ n1323 ;
  assign n15601 = n11320 ^ n4641 ^ n1692 ;
  assign n15602 = ~n15294 & n15601 ;
  assign n15603 = n15602 ^ n3110 ^ 1'b0 ;
  assign n15604 = n9770 & ~n15603 ;
  assign n15605 = n2790 & n15604 ;
  assign n15606 = n14962 & ~n15605 ;
  assign n15611 = n15610 ^ n15606 ^ 1'b0 ;
  assign n15614 = ( n3419 & ~n4477 ) | ( n3419 & n4990 ) | ( ~n4477 & n4990 ) ;
  assign n15615 = n8334 ^ n5262 ^ n4111 ;
  assign n15616 = ( n6664 & ~n15614 ) | ( n6664 & n15615 ) | ( ~n15614 & n15615 ) ;
  assign n15612 = ( ~n528 & n6803 ) | ( ~n528 & n7747 ) | ( n6803 & n7747 ) ;
  assign n15613 = ( n8509 & n9261 ) | ( n8509 & n15612 ) | ( n9261 & n15612 ) ;
  assign n15617 = n15616 ^ n15613 ^ n601 ;
  assign n15618 = ( n4932 & n6526 ) | ( n4932 & ~n11661 ) | ( n6526 & ~n11661 ) ;
  assign n15619 = n4210 & ~n15618 ;
  assign n15620 = n15074 & n15619 ;
  assign n15621 = ( n710 & n14815 ) | ( n710 & n15620 ) | ( n14815 & n15620 ) ;
  assign n15622 = ( n3764 & n4401 ) | ( n3764 & n6114 ) | ( n4401 & n6114 ) ;
  assign n15623 = n14673 ^ n2474 ^ n2209 ;
  assign n15624 = n15622 & n15623 ;
  assign n15625 = n13919 ^ n2311 ^ 1'b0 ;
  assign n15626 = n15624 | n15625 ;
  assign n15627 = ~n1743 & n6711 ;
  assign n15628 = n3991 | n15627 ;
  assign n15629 = n2631 & n2975 ;
  assign n15630 = n15629 ^ n3925 ^ 1'b0 ;
  assign n15631 = n719 ^ n702 ^ 1'b0 ;
  assign n15632 = ( n1841 & n4519 ) | ( n1841 & n15631 ) | ( n4519 & n15631 ) ;
  assign n15633 = n4297 | n5487 ;
  assign n15634 = n15632 | n15633 ;
  assign n15635 = ~n15630 & n15634 ;
  assign n15636 = ~n1064 & n15635 ;
  assign n15637 = ( ~n5237 & n15435 ) | ( ~n5237 & n15636 ) | ( n15435 & n15636 ) ;
  assign n15638 = ( ~n710 & n1205 ) | ( ~n710 & n12202 ) | ( n1205 & n12202 ) ;
  assign n15639 = n4317 & ~n15638 ;
  assign n15640 = n12332 ^ n9839 ^ 1'b0 ;
  assign n15641 = n8475 ^ n6843 ^ n6437 ;
  assign n15642 = ( x241 & n3517 ) | ( x241 & ~n5238 ) | ( n3517 & ~n5238 ) ;
  assign n15643 = n15642 ^ n8960 ^ 1'b0 ;
  assign n15644 = n15641 | n15643 ;
  assign n15645 = n15482 ^ n10919 ^ n10673 ;
  assign n15648 = n14466 ^ n12231 ^ 1'b0 ;
  assign n15646 = ~n834 & n5688 ;
  assign n15647 = n12097 & ~n15646 ;
  assign n15649 = n15648 ^ n15647 ^ 1'b0 ;
  assign n15652 = n3835 & ~n5066 ;
  assign n15653 = n15652 ^ n8983 ^ 1'b0 ;
  assign n15654 = n15653 ^ n3501 ^ n2316 ;
  assign n15650 = n10844 ^ n9342 ^ 1'b0 ;
  assign n15651 = n15650 ^ n1101 ^ n833 ;
  assign n15655 = n15654 ^ n15651 ^ n1806 ;
  assign n15656 = n4552 ^ n3206 ^ 1'b0 ;
  assign n15657 = n2053 | n15656 ;
  assign n15660 = ( n3263 & ~n3311 ) | ( n3263 & n5804 ) | ( ~n3311 & n5804 ) ;
  assign n15658 = x57 & ~n4060 ;
  assign n15659 = n15658 ^ n1422 ^ 1'b0 ;
  assign n15661 = n15660 ^ n15659 ^ n2492 ;
  assign n15662 = n3071 ^ n1190 ^ 1'b0 ;
  assign n15663 = n15661 | n15662 ;
  assign n15664 = ~n15657 & n15663 ;
  assign n15665 = n6850 ^ n6304 ^ 1'b0 ;
  assign n15669 = n5573 ^ n5269 ^ n4530 ;
  assign n15667 = ( n2690 & n14284 ) | ( n2690 & ~n14912 ) | ( n14284 & ~n14912 ) ;
  assign n15668 = ( n2722 & ~n10755 ) | ( n2722 & n15667 ) | ( ~n10755 & n15667 ) ;
  assign n15666 = n8055 | n10445 ;
  assign n15670 = n15669 ^ n15668 ^ n15666 ;
  assign n15671 = ( n3848 & n6062 ) | ( n3848 & n15670 ) | ( n6062 & n15670 ) ;
  assign n15680 = n1840 & ~n2115 ;
  assign n15681 = n15680 ^ n7133 ^ 1'b0 ;
  assign n15672 = ~n539 & n15580 ;
  assign n15673 = n15672 ^ n4827 ^ 1'b0 ;
  assign n15674 = ( n2302 & n4228 ) | ( n2302 & n10585 ) | ( n4228 & n10585 ) ;
  assign n15675 = n15674 ^ n7518 ^ 1'b0 ;
  assign n15676 = ~n8824 & n15675 ;
  assign n15677 = ( n5931 & ~n15673 ) | ( n5931 & n15676 ) | ( ~n15673 & n15676 ) ;
  assign n15678 = ( n1197 & ~n2089 ) | ( n1197 & n15677 ) | ( ~n2089 & n15677 ) ;
  assign n15679 = n15678 ^ n10249 ^ 1'b0 ;
  assign n15682 = n15681 ^ n15679 ^ 1'b0 ;
  assign n15684 = n3986 & ~n6056 ;
  assign n15685 = ~n5049 & n15684 ;
  assign n15683 = ~n772 & n2325 ;
  assign n15686 = n15685 ^ n15683 ^ n5051 ;
  assign n15687 = n15686 ^ n12512 ^ n4209 ;
  assign n15688 = ( ~n554 & n5557 ) | ( ~n554 & n10780 ) | ( n5557 & n10780 ) ;
  assign n15689 = ( n786 & n4317 ) | ( n786 & n15688 ) | ( n4317 & n15688 ) ;
  assign n15690 = ~n14568 & n15689 ;
  assign n15691 = n7597 & n15690 ;
  assign n15692 = ~n530 & n8015 ;
  assign n15693 = n11667 & ~n15692 ;
  assign n15694 = n11479 | n13183 ;
  assign n15695 = ~n10897 & n15694 ;
  assign n15696 = n15695 ^ n8429 ^ 1'b0 ;
  assign n15697 = ( n8287 & ~n10223 ) | ( n8287 & n14270 ) | ( ~n10223 & n14270 ) ;
  assign n15698 = n15697 ^ n2536 ^ 1'b0 ;
  assign n15699 = ( n8420 & n11186 ) | ( n8420 & ~n15698 ) | ( n11186 & ~n15698 ) ;
  assign n15700 = n6353 & ~n7612 ;
  assign n15701 = n1045 & n13611 ;
  assign n15702 = n15034 ^ n3202 ^ n1243 ;
  assign n15703 = ( ~n11800 & n14420 ) | ( ~n11800 & n15702 ) | ( n14420 & n15702 ) ;
  assign n15704 = n15703 ^ n13273 ^ 1'b0 ;
  assign n15705 = n432 & n4693 ;
  assign n15706 = ~n13584 & n15705 ;
  assign n15707 = ~n2134 & n15706 ;
  assign n15708 = n851 ^ x99 ^ 1'b0 ;
  assign n15709 = n9546 ^ n4141 ^ 1'b0 ;
  assign n15710 = n2255 & ~n15709 ;
  assign n15711 = n15300 ^ n12045 ^ 1'b0 ;
  assign n15712 = n11170 & n15711 ;
  assign n15713 = ~n3080 & n11863 ;
  assign n15714 = n6237 & n15713 ;
  assign n15715 = n3601 ^ n448 ^ 1'b0 ;
  assign n15716 = n15714 | n15715 ;
  assign n15717 = ( n14471 & n15712 ) | ( n14471 & n15716 ) | ( n15712 & n15716 ) ;
  assign n15718 = n12530 ^ n4929 ^ 1'b0 ;
  assign n15719 = n1095 & n4972 ;
  assign n15720 = n8324 & n15719 ;
  assign n15721 = n15720 ^ n13224 ^ 1'b0 ;
  assign n15722 = n13865 ^ n6028 ^ 1'b0 ;
  assign n15723 = n539 & n3814 ;
  assign n15724 = n7688 | n9089 ;
  assign n15725 = n15724 ^ n2545 ^ 1'b0 ;
  assign n15726 = ( n4403 & ~n15723 ) | ( n4403 & n15725 ) | ( ~n15723 & n15725 ) ;
  assign n15727 = n1908 ^ n1798 ^ 1'b0 ;
  assign n15728 = ~n5543 & n15727 ;
  assign n15729 = n1123 | n15728 ;
  assign n15730 = n15729 ^ n11925 ^ n1122 ;
  assign n15731 = n11084 & ~n15730 ;
  assign n15732 = n15726 & n15731 ;
  assign n15733 = n15522 ^ n10574 ^ n467 ;
  assign n15734 = n12967 ^ n10206 ^ n579 ;
  assign n15735 = n9437 ^ n3559 ^ n1797 ;
  assign n15736 = n9331 | n15735 ;
  assign n15737 = ( n6917 & n8066 ) | ( n6917 & n9688 ) | ( n8066 & n9688 ) ;
  assign n15738 = n15737 ^ n14241 ^ n8301 ;
  assign n15739 = ( n1184 & ~n4527 ) | ( n1184 & n10606 ) | ( ~n4527 & n10606 ) ;
  assign n15740 = n4477 ^ n4316 ^ n3231 ;
  assign n15741 = n3653 & n15740 ;
  assign n15742 = n15741 ^ n2999 ^ 1'b0 ;
  assign n15743 = n15742 ^ n15451 ^ 1'b0 ;
  assign n15744 = n15739 | n15743 ;
  assign n15745 = n8216 ^ n5910 ^ n1620 ;
  assign n15746 = ( n3427 & n8237 ) | ( n3427 & ~n15745 ) | ( n8237 & ~n15745 ) ;
  assign n15747 = n9506 | n15746 ;
  assign n15748 = n15744 & ~n15747 ;
  assign n15749 = n14474 ^ n9156 ^ 1'b0 ;
  assign n15750 = n1428 | n15749 ;
  assign n15751 = ( n4042 & ~n6565 ) | ( n4042 & n15750 ) | ( ~n6565 & n15750 ) ;
  assign n15752 = n15751 ^ n2640 ^ 1'b0 ;
  assign n15753 = ( n559 & n1043 ) | ( n559 & ~n14757 ) | ( n1043 & ~n14757 ) ;
  assign n15754 = ( n3059 & ~n14087 ) | ( n3059 & n15753 ) | ( ~n14087 & n15753 ) ;
  assign n15755 = ~n1096 & n15754 ;
  assign n15756 = n4051 & ~n8211 ;
  assign n15757 = n15756 ^ n14865 ^ 1'b0 ;
  assign n15758 = n10534 ^ n2279 ^ n1442 ;
  assign n15759 = n15083 | n15758 ;
  assign n15760 = n15759 ^ n7995 ^ 1'b0 ;
  assign n15761 = n11174 ^ n1880 ^ 1'b0 ;
  assign n15762 = n4726 & ~n15761 ;
  assign n15766 = n9637 ^ n1107 ^ n883 ;
  assign n15767 = ( n11322 & ~n11834 ) | ( n11322 & n15766 ) | ( ~n11834 & n15766 ) ;
  assign n15763 = ~n5727 & n7554 ;
  assign n15764 = n15763 ^ n477 ^ 1'b0 ;
  assign n15765 = ~n14894 & n15764 ;
  assign n15768 = n15767 ^ n15765 ^ n10115 ;
  assign n15769 = ( x8 & ~n4634 ) | ( x8 & n8943 ) | ( ~n4634 & n8943 ) ;
  assign n15770 = ( n7417 & n13548 ) | ( n7417 & n15769 ) | ( n13548 & n15769 ) ;
  assign n15771 = n526 & ~n1703 ;
  assign n15772 = n15771 ^ n2147 ^ 1'b0 ;
  assign n15773 = ( ~n7645 & n15770 ) | ( ~n7645 & n15772 ) | ( n15770 & n15772 ) ;
  assign n15774 = n14382 ^ n8522 ^ n7929 ;
  assign n15775 = n6601 ^ n4936 ^ 1'b0 ;
  assign n15776 = n753 & n15775 ;
  assign n15777 = n13578 & ~n15776 ;
  assign n15778 = ~n13558 & n15777 ;
  assign n15779 = n15778 ^ n10456 ^ 1'b0 ;
  assign n15780 = n12493 ^ n1163 ^ 1'b0 ;
  assign n15781 = n1889 ^ n1555 ^ 1'b0 ;
  assign n15782 = n15781 ^ n2716 ^ 1'b0 ;
  assign n15783 = n2485 | n15360 ;
  assign n15784 = n15783 ^ n6025 ^ n3886 ;
  assign n15785 = n12537 ^ n7871 ^ n3458 ;
  assign n15786 = n3177 ^ n1491 ^ 1'b0 ;
  assign n15787 = ~n15785 & n15786 ;
  assign n15788 = n11606 & ~n12674 ;
  assign n15789 = ( n6491 & ~n8817 ) | ( n6491 & n15788 ) | ( ~n8817 & n15788 ) ;
  assign n15790 = ( n6392 & n15787 ) | ( n6392 & n15789 ) | ( n15787 & n15789 ) ;
  assign n15791 = n12052 ^ n10229 ^ 1'b0 ;
  assign n15792 = n15791 ^ n3875 ^ 1'b0 ;
  assign n15793 = ~n3101 & n15792 ;
  assign n15794 = n10161 ^ n4073 ^ 1'b0 ;
  assign n15795 = n12722 | n15794 ;
  assign n15796 = ( ~n884 & n8952 ) | ( ~n884 & n15795 ) | ( n8952 & n15795 ) ;
  assign n15797 = n400 & n15305 ;
  assign n15798 = n10452 ^ n4122 ^ 1'b0 ;
  assign n15799 = n6712 ^ n6573 ^ n5114 ;
  assign n15800 = n15164 | n15799 ;
  assign n15801 = n15798 & ~n15800 ;
  assign n15802 = ~n1388 & n2050 ;
  assign n15803 = n15802 ^ n9438 ^ 1'b0 ;
  assign n15804 = ~n15500 & n15803 ;
  assign n15813 = n3209 ^ n3169 ^ 1'b0 ;
  assign n15812 = ( n690 & n1166 ) | ( n690 & n2315 ) | ( n1166 & n2315 ) ;
  assign n15814 = n15813 ^ n15812 ^ 1'b0 ;
  assign n15809 = n1320 & n10016 ;
  assign n15810 = ~n4053 & n15809 ;
  assign n15811 = ( n4197 & n7358 ) | ( n4197 & ~n15810 ) | ( n7358 & ~n15810 ) ;
  assign n15815 = n15814 ^ n15811 ^ 1'b0 ;
  assign n15816 = n7908 | n15815 ;
  assign n15805 = n7490 & n13543 ;
  assign n15806 = n15805 ^ n2401 ^ 1'b0 ;
  assign n15807 = n1652 & n15806 ;
  assign n15808 = n1507 | n15807 ;
  assign n15817 = n15816 ^ n15808 ^ 1'b0 ;
  assign n15818 = n8106 & n11642 ;
  assign n15819 = n3219 & n15818 ;
  assign n15820 = n1128 | n3767 ;
  assign n15821 = n12175 ^ n8472 ^ n3653 ;
  assign n15822 = n2191 | n15821 ;
  assign n15823 = n5547 ^ n3366 ^ 1'b0 ;
  assign n15824 = n15822 | n15823 ;
  assign n15825 = n4487 ^ n2354 ^ 1'b0 ;
  assign n15826 = n13614 | n15825 ;
  assign n15827 = n15826 ^ n9688 ^ 1'b0 ;
  assign n15828 = ~n10315 & n15827 ;
  assign n15829 = n3398 | n7644 ;
  assign n15830 = n15829 ^ n6162 ^ n5659 ;
  assign n15835 = n4814 ^ n2273 ^ n1163 ;
  assign n15831 = ~n1826 & n8032 ;
  assign n15832 = n15831 ^ n3069 ^ 1'b0 ;
  assign n15833 = n4206 & n15832 ;
  assign n15834 = n15833 ^ n1609 ^ n1602 ;
  assign n15836 = n15835 ^ n15834 ^ n9277 ;
  assign n15837 = n11600 & n15836 ;
  assign n15839 = n12825 ^ n9261 ^ x162 ;
  assign n15840 = n15301 ^ n12440 ^ n3184 ;
  assign n15841 = n15840 ^ n1274 ^ 1'b0 ;
  assign n15842 = n15839 & ~n15841 ;
  assign n15838 = ~n13943 & n14639 ;
  assign n15843 = n15842 ^ n15838 ^ 1'b0 ;
  assign n15844 = n1031 | n4101 ;
  assign n15845 = n15844 ^ n13423 ^ n3256 ;
  assign n15846 = ( n1138 & ~n8164 ) | ( n1138 & n15845 ) | ( ~n8164 & n15845 ) ;
  assign n15847 = ~n15423 & n15846 ;
  assign n15848 = n13990 | n15847 ;
  assign n15849 = n9396 ^ n1018 ^ n510 ;
  assign n15850 = n13874 ^ n3814 ^ 1'b0 ;
  assign n15851 = n7003 ^ n5028 ^ n3066 ;
  assign n15852 = n15851 ^ n6158 ^ 1'b0 ;
  assign n15853 = n15852 ^ n8276 ^ 1'b0 ;
  assign n15854 = ~n15850 & n15853 ;
  assign n15855 = n2155 | n2584 ;
  assign n15856 = ( n15849 & ~n15854 ) | ( n15849 & n15855 ) | ( ~n15854 & n15855 ) ;
  assign n15857 = n15856 ^ n9013 ^ 1'b0 ;
  assign n15859 = ( n7642 & n11103 ) | ( n7642 & n11642 ) | ( n11103 & n11642 ) ;
  assign n15858 = n2057 | n5477 ;
  assign n15860 = n15859 ^ n15858 ^ 1'b0 ;
  assign n15861 = n3295 | n4632 ;
  assign n15862 = n15861 ^ n3877 ^ 1'b0 ;
  assign n15863 = n15862 ^ n3824 ^ n1028 ;
  assign n15864 = n15863 ^ n7847 ^ 1'b0 ;
  assign n15865 = n8721 ^ n6084 ^ 1'b0 ;
  assign n15866 = ~n4346 & n15865 ;
  assign n15867 = ~n3567 & n9911 ;
  assign n15868 = n15867 ^ n6696 ^ 1'b0 ;
  assign n15869 = n15866 & n15868 ;
  assign n15870 = n13298 ^ n4137 ^ n1022 ;
  assign n15871 = ~n11991 & n12426 ;
  assign n15872 = n15871 ^ n5028 ^ 1'b0 ;
  assign n15873 = n10193 ^ n6913 ^ 1'b0 ;
  assign n15874 = x194 & n15873 ;
  assign n15878 = n6795 ^ n5299 ^ 1'b0 ;
  assign n15879 = n7504 & ~n15878 ;
  assign n15880 = n15879 ^ n11240 ^ n8757 ;
  assign n15881 = n14900 & ~n15880 ;
  assign n15876 = n8779 ^ n654 ^ 1'b0 ;
  assign n15875 = n5052 ^ n4656 ^ 1'b0 ;
  assign n15877 = n15876 ^ n15875 ^ n15294 ;
  assign n15882 = n15881 ^ n15877 ^ n9147 ;
  assign n15884 = n12972 ^ n9697 ^ 1'b0 ;
  assign n15885 = n15884 ^ n9240 ^ n707 ;
  assign n15883 = n9606 | n13088 ;
  assign n15886 = n15885 ^ n15883 ^ n755 ;
  assign n15887 = n15886 ^ n12264 ^ 1'b0 ;
  assign n15888 = n7366 & n13522 ;
  assign n15889 = n7087 ^ n2217 ^ 1'b0 ;
  assign n15890 = ( n10609 & n11641 ) | ( n10609 & ~n15889 ) | ( n11641 & ~n15889 ) ;
  assign n15891 = n8260 & ~n15890 ;
  assign n15892 = n15891 ^ n12065 ^ 1'b0 ;
  assign n15893 = ( n14730 & n15888 ) | ( n14730 & n15892 ) | ( n15888 & n15892 ) ;
  assign n15894 = n401 | n965 ;
  assign n15895 = n12712 & ~n15894 ;
  assign n15896 = n11980 & ~n15895 ;
  assign n15897 = n15896 ^ n7514 ^ 1'b0 ;
  assign n15899 = n10826 & n11076 ;
  assign n15900 = ( ~n1237 & n13620 ) | ( ~n1237 & n15899 ) | ( n13620 & n15899 ) ;
  assign n15898 = ~n261 & n1646 ;
  assign n15901 = n15900 ^ n15898 ^ n3979 ;
  assign n15902 = ( n1163 & n7390 ) | ( n1163 & n13238 ) | ( n7390 & n13238 ) ;
  assign n15903 = n9621 ^ n3399 ^ 1'b0 ;
  assign n15904 = n10023 | n15903 ;
  assign n15905 = n15904 ^ n7327 ^ n5769 ;
  assign n15906 = n5810 ^ n4634 ^ 1'b0 ;
  assign n15909 = n12556 ^ n9671 ^ n4937 ;
  assign n15907 = ~n683 & n1034 ;
  assign n15908 = n5435 & n15907 ;
  assign n15910 = n15909 ^ n15908 ^ n11490 ;
  assign n15911 = n15910 ^ n3052 ^ 1'b0 ;
  assign n15912 = ~n15906 & n15911 ;
  assign n15916 = n9530 ^ n8945 ^ 1'b0 ;
  assign n15917 = n13042 & n15916 ;
  assign n15913 = n1728 & n4389 ;
  assign n15914 = n9188 ^ n3591 ^ n689 ;
  assign n15915 = ~n15913 & n15914 ;
  assign n15918 = n15917 ^ n15915 ^ 1'b0 ;
  assign n15919 = n9727 ^ n7285 ^ 1'b0 ;
  assign n15920 = n15918 & ~n15919 ;
  assign n15921 = ( n7976 & ~n8111 ) | ( n7976 & n13273 ) | ( ~n8111 & n13273 ) ;
  assign n15922 = n15921 ^ n6416 ^ n5585 ;
  assign n15925 = n6797 ^ n4893 ^ 1'b0 ;
  assign n15923 = n7988 & ~n8256 ;
  assign n15924 = n3762 & n15923 ;
  assign n15926 = n15925 ^ n15924 ^ n624 ;
  assign n15927 = ( x130 & n389 ) | ( x130 & ~n3128 ) | ( n389 & ~n3128 ) ;
  assign n15928 = n1028 & ~n1739 ;
  assign n15929 = n15928 ^ n3845 ^ 1'b0 ;
  assign n15930 = n15929 ^ n14917 ^ n13456 ;
  assign n15931 = n15927 | n15930 ;
  assign n15932 = ( n9575 & ~n12147 ) | ( n9575 & n15931 ) | ( ~n12147 & n15931 ) ;
  assign n15933 = n15932 ^ n14654 ^ n2726 ;
  assign n15935 = ~n2110 & n3195 ;
  assign n15934 = n798 & ~n9303 ;
  assign n15936 = n15935 ^ n15934 ^ 1'b0 ;
  assign n15937 = n8672 & n15936 ;
  assign n15938 = n10497 ^ n2760 ^ 1'b0 ;
  assign n15944 = n5792 & ~n13583 ;
  assign n15945 = n15944 ^ n3357 ^ 1'b0 ;
  assign n15946 = n15945 ^ n5908 ^ n1277 ;
  assign n15939 = n1362 ^ n470 ^ 1'b0 ;
  assign n15940 = n7196 & ~n9856 ;
  assign n15941 = ~n15939 & n15940 ;
  assign n15942 = n15941 ^ n2808 ^ n1581 ;
  assign n15943 = n15942 ^ x127 ^ 1'b0 ;
  assign n15947 = n15946 ^ n15943 ^ n10796 ;
  assign n15948 = n10994 ^ n3803 ^ n2638 ;
  assign n15950 = n14249 ^ n6959 ^ n2055 ;
  assign n15949 = n5172 & n10756 ;
  assign n15951 = n15950 ^ n15949 ^ 1'b0 ;
  assign n15952 = ~n3856 & n5896 ;
  assign n15953 = n15952 ^ n2474 ^ 1'b0 ;
  assign n15954 = n15953 ^ n6521 ^ 1'b0 ;
  assign n15955 = ( n683 & n7157 ) | ( n683 & ~n15954 ) | ( n7157 & ~n15954 ) ;
  assign n15956 = n15955 ^ n4499 ^ 1'b0 ;
  assign n15957 = n11906 ^ n4003 ^ 1'b0 ;
  assign n15958 = ~n750 & n15957 ;
  assign n15959 = n15958 ^ n5412 ^ n2922 ;
  assign n15960 = n15959 ^ n2885 ^ 1'b0 ;
  assign n15965 = n7884 ^ n7097 ^ 1'b0 ;
  assign n15966 = ~n6485 & n14234 ;
  assign n15967 = n4208 | n15966 ;
  assign n15968 = n15965 & ~n15967 ;
  assign n15962 = n2382 & n4466 ;
  assign n15961 = ~n2973 & n10907 ;
  assign n15963 = n15962 ^ n15961 ^ 1'b0 ;
  assign n15964 = n15963 ^ n7327 ^ n6257 ;
  assign n15969 = n15968 ^ n15964 ^ n7633 ;
  assign n15970 = ( n2727 & ~n4494 ) | ( n2727 & n4784 ) | ( ~n4494 & n4784 ) ;
  assign n15971 = n3869 | n6230 ;
  assign n15974 = n3281 | n8024 ;
  assign n15972 = n1019 & ~n1040 ;
  assign n15973 = ~n9555 & n15972 ;
  assign n15975 = n15974 ^ n15973 ^ n9033 ;
  assign n15980 = x211 & n15137 ;
  assign n15981 = ~n2217 & n15980 ;
  assign n15979 = n14322 ^ n4248 ^ n1457 ;
  assign n15976 = ( n6045 & n6474 ) | ( n6045 & n14550 ) | ( n6474 & n14550 ) ;
  assign n15977 = n15463 ^ n7854 ^ 1'b0 ;
  assign n15978 = n15976 & ~n15977 ;
  assign n15982 = n15981 ^ n15979 ^ n15978 ;
  assign n15983 = n1461 | n2813 ;
  assign n15984 = n15983 ^ n15378 ^ 1'b0 ;
  assign n15985 = n8145 ^ n7003 ^ 1'b0 ;
  assign n15986 = ( n7571 & n15984 ) | ( n7571 & n15985 ) | ( n15984 & n15985 ) ;
  assign n15987 = n15986 ^ n10181 ^ 1'b0 ;
  assign n15988 = ~n2718 & n8883 ;
  assign n15989 = n15988 ^ n8886 ^ 1'b0 ;
  assign n15990 = n6676 & ~n15989 ;
  assign n15991 = ( n6064 & n6104 ) | ( n6064 & n9516 ) | ( n6104 & n9516 ) ;
  assign n15992 = n11346 ^ n8731 ^ 1'b0 ;
  assign n16001 = n13905 ^ n7029 ^ n6106 ;
  assign n15999 = n11226 ^ n4082 ^ 1'b0 ;
  assign n16000 = n5530 | n15999 ;
  assign n15993 = ~n2871 & n5318 ;
  assign n15994 = n7805 ^ n1636 ^ 1'b0 ;
  assign n15995 = n15993 | n15994 ;
  assign n15996 = n15995 ^ n9061 ^ 1'b0 ;
  assign n15997 = ~n1837 & n9944 ;
  assign n15998 = ~n15996 & n15997 ;
  assign n16002 = n16001 ^ n16000 ^ n15998 ;
  assign n16003 = ~n1000 & n10368 ;
  assign n16004 = ~n16002 & n16003 ;
  assign n16005 = n10103 ^ n5014 ^ 1'b0 ;
  assign n16006 = n2256 | n7119 ;
  assign n16007 = n16006 ^ n270 ^ 1'b0 ;
  assign n16008 = ( n1353 & ~n15465 ) | ( n1353 & n16007 ) | ( ~n15465 & n16007 ) ;
  assign n16009 = n5391 ^ n4506 ^ 1'b0 ;
  assign n16010 = n14176 & ~n16009 ;
  assign n16011 = x116 & ~n4493 ;
  assign n16012 = n13578 & ~n16011 ;
  assign n16013 = n1098 & n16012 ;
  assign n16016 = ( n2777 & ~n4071 ) | ( n2777 & n9551 ) | ( ~n4071 & n9551 ) ;
  assign n16014 = n2194 & n5569 ;
  assign n16015 = n16014 ^ n3154 ^ 1'b0 ;
  assign n16017 = n16016 ^ n16015 ^ n7901 ;
  assign n16018 = ( n7016 & n10577 ) | ( n7016 & n10848 ) | ( n10577 & n10848 ) ;
  assign n16023 = ( ~n3811 & n4776 ) | ( ~n3811 & n8059 ) | ( n4776 & n8059 ) ;
  assign n16019 = n3126 ^ n1990 ^ 1'b0 ;
  assign n16020 = n1484 ^ n1031 ^ x166 ;
  assign n16021 = n16020 ^ n1077 ^ n668 ;
  assign n16022 = ( n3255 & n16019 ) | ( n3255 & n16021 ) | ( n16019 & n16021 ) ;
  assign n16024 = n16023 ^ n16022 ^ 1'b0 ;
  assign n16031 = n1657 ^ n1191 ^ 1'b0 ;
  assign n16032 = n5726 | n16031 ;
  assign n16029 = n2889 ^ n1485 ^ n1411 ;
  assign n16030 = n2238 & ~n16029 ;
  assign n16033 = n16032 ^ n16030 ^ n2510 ;
  assign n16025 = n4613 | n10140 ;
  assign n16026 = n16025 ^ n13692 ^ 1'b0 ;
  assign n16027 = n14665 ^ n12069 ^ 1'b0 ;
  assign n16028 = n16026 & n16027 ;
  assign n16034 = n16033 ^ n16028 ^ n15391 ;
  assign n16035 = n15881 ^ n2580 ^ 1'b0 ;
  assign n16036 = n16034 & n16035 ;
  assign n16037 = ~n7108 & n14381 ;
  assign n16044 = n5970 ^ n2021 ^ 1'b0 ;
  assign n16045 = n7606 | n16044 ;
  assign n16046 = n16045 ^ n6842 ^ 1'b0 ;
  assign n16047 = ( ~n489 & n6765 ) | ( ~n489 & n10869 ) | ( n6765 & n10869 ) ;
  assign n16048 = n6092 & n9016 ;
  assign n16049 = ( n14616 & n15045 ) | ( n14616 & n16048 ) | ( n15045 & n16048 ) ;
  assign n16050 = ( ~n14656 & n16047 ) | ( ~n14656 & n16049 ) | ( n16047 & n16049 ) ;
  assign n16051 = ( n1091 & n16046 ) | ( n1091 & n16050 ) | ( n16046 & n16050 ) ;
  assign n16052 = n12478 & n16051 ;
  assign n16041 = n13552 ^ n11244 ^ n10776 ;
  assign n16042 = ( n10269 & n14032 ) | ( n10269 & ~n16041 ) | ( n14032 & ~n16041 ) ;
  assign n16043 = n16042 ^ n12525 ^ n3446 ;
  assign n16038 = ~n4691 & n5149 ;
  assign n16039 = n6345 & n16038 ;
  assign n16040 = ( n2840 & ~n14393 ) | ( n2840 & n16039 ) | ( ~n14393 & n16039 ) ;
  assign n16053 = n16052 ^ n16043 ^ n16040 ;
  assign n16054 = n966 & n8798 ;
  assign n16055 = n15735 ^ n15423 ^ n7645 ;
  assign n16056 = n8156 ^ n310 ^ 1'b0 ;
  assign n16057 = ~n716 & n16056 ;
  assign n16058 = ( n16054 & n16055 ) | ( n16054 & n16057 ) | ( n16055 & n16057 ) ;
  assign n16062 = n13006 ^ n9673 ^ 1'b0 ;
  assign n16063 = n6720 & ~n16062 ;
  assign n16059 = n8797 ^ n1639 ^ 1'b0 ;
  assign n16060 = x211 & ~n16059 ;
  assign n16061 = n6584 & n16060 ;
  assign n16064 = n16063 ^ n16061 ^ 1'b0 ;
  assign n16065 = n16064 ^ n5263 ^ n557 ;
  assign n16066 = ~n2776 & n8921 ;
  assign n16067 = n894 & n3081 ;
  assign n16068 = n16067 ^ n13868 ^ 1'b0 ;
  assign n16069 = n6161 ^ n2603 ^ 1'b0 ;
  assign n16070 = n4966 & ~n16069 ;
  assign n16071 = n16068 & n16070 ;
  assign n16072 = n13438 | n16071 ;
  assign n16073 = n16066 | n16072 ;
  assign n16074 = ~n6705 & n8621 ;
  assign n16075 = ( n9220 & n9451 ) | ( n9220 & n15779 ) | ( n9451 & n15779 ) ;
  assign n16078 = ( n4315 & n5482 ) | ( n4315 & n10129 ) | ( n5482 & n10129 ) ;
  assign n16077 = n13069 ^ n12292 ^ 1'b0 ;
  assign n16076 = n3929 ^ n2396 ^ 1'b0 ;
  assign n16079 = n16078 ^ n16077 ^ n16076 ;
  assign n16080 = n6263 | n11673 ;
  assign n16081 = n16080 ^ n7899 ^ n2178 ;
  assign n16083 = x44 & n345 ;
  assign n16084 = n16083 ^ n1722 ^ 1'b0 ;
  assign n16082 = ( x25 & ~x214 ) | ( x25 & n7721 ) | ( ~x214 & n7721 ) ;
  assign n16085 = n16084 ^ n16082 ^ 1'b0 ;
  assign n16086 = n5075 & n16085 ;
  assign n16087 = ~n2322 & n16086 ;
  assign n16088 = n7908 ^ n7201 ^ 1'b0 ;
  assign n16089 = ( ~n2426 & n5342 ) | ( ~n2426 & n6010 ) | ( n5342 & n6010 ) ;
  assign n16090 = n13670 & ~n16089 ;
  assign n16091 = n3333 & n9055 ;
  assign n16092 = n16091 ^ n4030 ^ 1'b0 ;
  assign n16093 = n8923 & n16092 ;
  assign n16094 = n11397 ^ n10020 ^ 1'b0 ;
  assign n16095 = ~n14215 & n16094 ;
  assign n16096 = n16095 ^ n12267 ^ 1'b0 ;
  assign n16097 = n3093 | n16096 ;
  assign n16098 = n2848 & ~n6859 ;
  assign n16099 = ( n298 & ~n4750 ) | ( n298 & n16098 ) | ( ~n4750 & n16098 ) ;
  assign n16100 = n14404 ^ n13126 ^ n1903 ;
  assign n16101 = n914 & n8539 ;
  assign n16102 = n1164 & n2842 ;
  assign n16103 = n16102 ^ n595 ^ 1'b0 ;
  assign n16104 = n16103 ^ n11514 ^ 1'b0 ;
  assign n16109 = n7966 ^ n3015 ^ n661 ;
  assign n16110 = n16109 ^ n6887 ^ n1311 ;
  assign n16111 = n16110 ^ n9765 ^ n4582 ;
  assign n16105 = ( ~n737 & n4014 ) | ( ~n737 & n5241 ) | ( n4014 & n5241 ) ;
  assign n16106 = n5354 & ~n7005 ;
  assign n16107 = n16106 ^ n4086 ^ 1'b0 ;
  assign n16108 = n16105 | n16107 ;
  assign n16112 = n16111 ^ n16108 ^ 1'b0 ;
  assign n16113 = n787 & ~n4775 ;
  assign n16114 = ( n8325 & ~n11510 ) | ( n8325 & n16113 ) | ( ~n11510 & n16113 ) ;
  assign n16115 = ( n13121 & n15503 ) | ( n13121 & ~n16114 ) | ( n15503 & ~n16114 ) ;
  assign n16116 = n11001 ^ n10784 ^ 1'b0 ;
  assign n16117 = n8979 | n16116 ;
  assign n16118 = n12601 | n16117 ;
  assign n16119 = n16118 ^ n5206 ^ n3679 ;
  assign n16120 = n7332 ^ n2195 ^ 1'b0 ;
  assign n16121 = n5055 & n16120 ;
  assign n16122 = ( n3829 & ~n7827 ) | ( n3829 & n16121 ) | ( ~n7827 & n16121 ) ;
  assign n16123 = ( ~x17 & n1400 ) | ( ~x17 & n13229 ) | ( n1400 & n13229 ) ;
  assign n16124 = n5235 ^ n4908 ^ 1'b0 ;
  assign n16125 = n16123 & ~n16124 ;
  assign n16126 = n11919 ^ n5290 ^ n349 ;
  assign n16127 = n16126 ^ n603 ^ 1'b0 ;
  assign n16128 = n16125 & ~n16127 ;
  assign n16129 = n9652 ^ n8725 ^ n4391 ;
  assign n16130 = x237 & ~n16129 ;
  assign n16131 = n16130 ^ n9450 ^ 1'b0 ;
  assign n16132 = n16131 ^ n4418 ^ 1'b0 ;
  assign n16133 = ~n13222 & n16132 ;
  assign n16134 = n5695 ^ n5395 ^ n4119 ;
  assign n16135 = n11556 | n13291 ;
  assign n16136 = ( n3718 & n16134 ) | ( n3718 & ~n16135 ) | ( n16134 & ~n16135 ) ;
  assign n16137 = n5708 & ~n16136 ;
  assign n16138 = ( n729 & ~n2799 ) | ( n729 & n10505 ) | ( ~n2799 & n10505 ) ;
  assign n16139 = ( ~n1344 & n6088 ) | ( ~n1344 & n8851 ) | ( n6088 & n8851 ) ;
  assign n16140 = n16139 ^ n10530 ^ 1'b0 ;
  assign n16141 = x86 & n8777 ;
  assign n16142 = n7175 ^ n1949 ^ 1'b0 ;
  assign n16143 = n7367 ^ n5248 ^ n4397 ;
  assign n16144 = n16143 ^ n6484 ^ 1'b0 ;
  assign n16145 = n9719 & n16144 ;
  assign n16146 = n16145 ^ n15134 ^ n1293 ;
  assign n16147 = n6662 & ~n15955 ;
  assign n16148 = ~n13184 & n16147 ;
  assign n16149 = n14128 ^ n6791 ^ n5984 ;
  assign n16150 = n4460 | n16149 ;
  assign n16151 = n16150 ^ n3591 ^ 1'b0 ;
  assign n16152 = n16151 ^ n4453 ^ 1'b0 ;
  assign n16153 = n3785 & n4888 ;
  assign n16154 = ~n1761 & n16153 ;
  assign n16156 = n2588 | n7801 ;
  assign n16155 = n12219 ^ n1812 ^ n755 ;
  assign n16157 = n16156 ^ n16155 ^ n3176 ;
  assign n16158 = ( n1028 & n3542 ) | ( n1028 & n4328 ) | ( n3542 & n4328 ) ;
  assign n16159 = ( n7592 & n7664 ) | ( n7592 & n16158 ) | ( n7664 & n16158 ) ;
  assign n16162 = n6037 & ~n14071 ;
  assign n16163 = n14503 & n16162 ;
  assign n16160 = n7964 ^ n4339 ^ 1'b0 ;
  assign n16161 = n16160 ^ n8523 ^ n6736 ;
  assign n16164 = n16163 ^ n16161 ^ n14167 ;
  assign n16165 = ~n16159 & n16164 ;
  assign n16166 = ~n11789 & n16165 ;
  assign n16167 = ~n4536 & n6190 ;
  assign n16168 = n7128 & n16167 ;
  assign n16169 = n3678 | n16168 ;
  assign n16170 = n14669 & n16169 ;
  assign n16171 = n9516 ^ n8542 ^ 1'b0 ;
  assign n16172 = ~n7838 & n16171 ;
  assign n16173 = ~n693 & n16172 ;
  assign n16174 = n13916 ^ n10288 ^ n3758 ;
  assign n16175 = n5402 & ~n5864 ;
  assign n16176 = n16175 ^ n4182 ^ 1'b0 ;
  assign n16177 = ( n899 & n3931 ) | ( n899 & n4635 ) | ( n3931 & n4635 ) ;
  assign n16178 = n11059 ^ n5123 ^ 1'b0 ;
  assign n16179 = ~n14547 & n16178 ;
  assign n16180 = n16177 & n16179 ;
  assign n16181 = ~n16176 & n16180 ;
  assign n16182 = n16174 & ~n16181 ;
  assign n16183 = n13744 ^ n1005 ^ 1'b0 ;
  assign n16184 = n5184 ^ n435 ^ 1'b0 ;
  assign n16185 = n7868 ^ n851 ^ 1'b0 ;
  assign n16186 = n16185 ^ n7771 ^ n2331 ;
  assign n16187 = n16186 ^ n8617 ^ 1'b0 ;
  assign n16188 = n2641 | n16169 ;
  assign n16189 = ( ~n16184 & n16187 ) | ( ~n16184 & n16188 ) | ( n16187 & n16188 ) ;
  assign n16190 = n8782 | n13482 ;
  assign n16191 = n10751 ^ n6858 ^ 1'b0 ;
  assign n16192 = ~n4379 & n16191 ;
  assign n16193 = n11113 | n16192 ;
  assign n16194 = n6919 & n13288 ;
  assign n16195 = ~n16193 & n16194 ;
  assign n16197 = n6908 & ~n13048 ;
  assign n16198 = n16197 ^ n14745 ^ 1'b0 ;
  assign n16199 = n16198 ^ n14150 ^ 1'b0 ;
  assign n16196 = n5622 | n9980 ;
  assign n16200 = n16199 ^ n16196 ^ 1'b0 ;
  assign n16201 = n761 & ~n16200 ;
  assign n16203 = n9793 ^ n3502 ^ 1'b0 ;
  assign n16204 = n6904 & n16203 ;
  assign n16202 = n10950 ^ n7377 ^ n3419 ;
  assign n16205 = n16204 ^ n16202 ^ n4384 ;
  assign n16206 = n16205 ^ n6287 ^ 1'b0 ;
  assign n16207 = n1587 & ~n12630 ;
  assign n16208 = n16207 ^ n3875 ^ 1'b0 ;
  assign n16212 = n943 | n3368 ;
  assign n16213 = n3068 & ~n16212 ;
  assign n16214 = n4775 ^ n3723 ^ 1'b0 ;
  assign n16215 = x7 & n16214 ;
  assign n16216 = ~n4348 & n16215 ;
  assign n16217 = n16213 | n16216 ;
  assign n16209 = ( n11124 & n12140 ) | ( n11124 & ~n15441 ) | ( n12140 & ~n15441 ) ;
  assign n16210 = ~n3040 & n16209 ;
  assign n16211 = n16210 ^ n12332 ^ 1'b0 ;
  assign n16218 = n16217 ^ n16211 ^ 1'b0 ;
  assign n16225 = n2504 ^ n1478 ^ n1224 ;
  assign n16224 = n5888 & n7016 ;
  assign n16226 = n16225 ^ n16224 ^ 1'b0 ;
  assign n16221 = n2796 ^ n1297 ^ 1'b0 ;
  assign n16222 = ~n10013 & n13868 ;
  assign n16223 = ~n16221 & n16222 ;
  assign n16227 = n16226 ^ n16223 ^ 1'b0 ;
  assign n16219 = n7077 ^ n4006 ^ x124 ;
  assign n16220 = n16219 ^ n9856 ^ n9629 ;
  assign n16228 = n16227 ^ n16220 ^ n12412 ;
  assign n16229 = n16228 ^ n15954 ^ n6862 ;
  assign n16230 = n1288 & n5241 ;
  assign n16231 = n2520 ^ n1208 ^ n733 ;
  assign n16232 = n16231 ^ n1454 ^ 1'b0 ;
  assign n16233 = ( n3308 & n16230 ) | ( n3308 & n16232 ) | ( n16230 & n16232 ) ;
  assign n16236 = n8588 ^ n6713 ^ n2097 ;
  assign n16237 = n16236 ^ n13042 ^ n7681 ;
  assign n16234 = ( n5697 & n8817 ) | ( n5697 & n14772 ) | ( n8817 & n14772 ) ;
  assign n16235 = n1231 & ~n16234 ;
  assign n16238 = n16237 ^ n16235 ^ 1'b0 ;
  assign n16239 = ~n1622 & n3520 ;
  assign n16240 = ( n3329 & ~n7385 ) | ( n3329 & n16239 ) | ( ~n7385 & n16239 ) ;
  assign n16241 = n8830 | n16240 ;
  assign n16254 = n4035 | n6364 ;
  assign n16255 = n16254 ^ n1623 ^ 1'b0 ;
  assign n16253 = ~n5008 & n16123 ;
  assign n16256 = n16255 ^ n16253 ^ 1'b0 ;
  assign n16252 = ~n10438 & n13082 ;
  assign n16257 = n16256 ^ n16252 ^ n2547 ;
  assign n16258 = x123 & ~n16257 ;
  assign n16259 = n16258 ^ n2069 ^ 1'b0 ;
  assign n16242 = ( ~n3190 & n4283 ) | ( ~n3190 & n6232 ) | ( n4283 & n6232 ) ;
  assign n16243 = ( n2785 & ~n5535 ) | ( n2785 & n16242 ) | ( ~n5535 & n16242 ) ;
  assign n16244 = n1163 ^ n918 ^ n541 ;
  assign n16245 = n7766 & n16244 ;
  assign n16246 = n8739 ^ n4937 ^ 1'b0 ;
  assign n16247 = n8665 & ~n16246 ;
  assign n16248 = ~n4725 & n16247 ;
  assign n16249 = n12304 & n16248 ;
  assign n16250 = ( n3124 & ~n16245 ) | ( n3124 & n16249 ) | ( ~n16245 & n16249 ) ;
  assign n16251 = ( n13141 & ~n16243 ) | ( n13141 & n16250 ) | ( ~n16243 & n16250 ) ;
  assign n16260 = n16259 ^ n16251 ^ 1'b0 ;
  assign n16261 = n10240 & ~n11637 ;
  assign n16262 = n2076 & n16261 ;
  assign n16263 = ~n4791 & n12861 ;
  assign n16264 = n9613 ^ n2538 ^ 1'b0 ;
  assign n16265 = ~n14031 & n16264 ;
  assign n16266 = ( ~x119 & n7136 ) | ( ~x119 & n9438 ) | ( n7136 & n9438 ) ;
  assign n16267 = ( n5576 & ~n8386 ) | ( n5576 & n16266 ) | ( ~n8386 & n16266 ) ;
  assign n16268 = n16267 ^ n13460 ^ n10424 ;
  assign n16269 = n9850 | n11570 ;
  assign n16270 = n16268 & ~n16269 ;
  assign n16271 = n12751 ^ n4319 ^ n521 ;
  assign n16272 = x136 & n16047 ;
  assign n16273 = n14789 ^ n11755 ^ 1'b0 ;
  assign n16274 = ( n2267 & ~n8010 ) | ( n2267 & n16273 ) | ( ~n8010 & n16273 ) ;
  assign n16275 = n5531 & ~n6918 ;
  assign n16276 = ( n13193 & n16274 ) | ( n13193 & ~n16275 ) | ( n16274 & ~n16275 ) ;
  assign n16277 = ( n16271 & ~n16272 ) | ( n16271 & n16276 ) | ( ~n16272 & n16276 ) ;
  assign n16278 = ( x38 & n3773 ) | ( x38 & n10150 ) | ( n3773 & n10150 ) ;
  assign n16279 = n1802 | n5454 ;
  assign n16280 = n14149 ^ n8301 ^ 1'b0 ;
  assign n16281 = n8247 ^ n3881 ^ n1087 ;
  assign n16282 = n5786 ^ n4846 ^ n2551 ;
  assign n16283 = ( n6789 & ~n11640 ) | ( n6789 & n16282 ) | ( ~n11640 & n16282 ) ;
  assign n16284 = n13156 ^ n6867 ^ n5215 ;
  assign n16285 = ( ~n10136 & n15167 ) | ( ~n10136 & n16284 ) | ( n15167 & n16284 ) ;
  assign n16286 = n6642 ^ n6160 ^ n934 ;
  assign n16287 = ( ~n5754 & n9078 ) | ( ~n5754 & n12291 ) | ( n9078 & n12291 ) ;
  assign n16288 = n12755 ^ n8226 ^ n646 ;
  assign n16289 = n2669 & n10584 ;
  assign n16290 = ( n16287 & n16288 ) | ( n16287 & ~n16289 ) | ( n16288 & ~n16289 ) ;
  assign n16292 = n6219 ^ n3188 ^ 1'b0 ;
  assign n16291 = n3261 & n15975 ;
  assign n16293 = n16292 ^ n16291 ^ 1'b0 ;
  assign n16294 = n5750 ^ n4681 ^ 1'b0 ;
  assign n16295 = ~n6557 & n16294 ;
  assign n16296 = n3627 | n13722 ;
  assign n16297 = ( n4240 & n14867 ) | ( n4240 & n16296 ) | ( n14867 & n16296 ) ;
  assign n16298 = ( n11682 & n16295 ) | ( n11682 & ~n16297 ) | ( n16295 & ~n16297 ) ;
  assign n16299 = n362 | n9064 ;
  assign n16300 = n16299 ^ n13635 ^ 1'b0 ;
  assign n16301 = n15476 ^ n3582 ^ n3347 ;
  assign n16302 = n7772 ^ n6737 ^ 1'b0 ;
  assign n16303 = n3837 & n16302 ;
  assign n16304 = n5361 ^ n295 ^ 1'b0 ;
  assign n16305 = n11788 & n16304 ;
  assign n16306 = n7051 ^ n2508 ^ 1'b0 ;
  assign n16307 = ( x8 & ~n8329 ) | ( x8 & n9872 ) | ( ~n8329 & n9872 ) ;
  assign n16308 = n16307 ^ n6713 ^ n6023 ;
  assign n16309 = ( n9969 & n11880 ) | ( n9969 & ~n16308 ) | ( n11880 & ~n16308 ) ;
  assign n16310 = n13815 ^ n8859 ^ n7136 ;
  assign n16311 = n16310 ^ n5246 ^ n3290 ;
  assign n16312 = ( n5634 & ~n9905 ) | ( n5634 & n16311 ) | ( ~n9905 & n16311 ) ;
  assign n16313 = n2708 | n4707 ;
  assign n16314 = n1135 | n16313 ;
  assign n16315 = n4284 & ~n8257 ;
  assign n16316 = ~n16314 & n16315 ;
  assign n16317 = ( ~n2749 & n2778 ) | ( ~n2749 & n5996 ) | ( n2778 & n5996 ) ;
  assign n16318 = ( n6061 & n6446 ) | ( n6061 & n16317 ) | ( n6446 & n16317 ) ;
  assign n16319 = n16318 ^ n8463 ^ 1'b0 ;
  assign n16320 = ~n16316 & n16319 ;
  assign n16321 = n4937 ^ n3339 ^ n2522 ;
  assign n16322 = n2840 | n16321 ;
  assign n16323 = ( n2970 & ~n6700 ) | ( n2970 & n12605 ) | ( ~n6700 & n12605 ) ;
  assign n16324 = ( n2962 & n3068 ) | ( n2962 & ~n5238 ) | ( n3068 & ~n5238 ) ;
  assign n16325 = ~n1221 & n14426 ;
  assign n16326 = n16325 ^ n7935 ^ 1'b0 ;
  assign n16327 = ( n4189 & n10410 ) | ( n4189 & n16326 ) | ( n10410 & n16326 ) ;
  assign n16328 = ( n1291 & n4425 ) | ( n1291 & ~n16327 ) | ( n4425 & ~n16327 ) ;
  assign n16329 = ( x186 & n1039 ) | ( x186 & ~n2034 ) | ( n1039 & ~n2034 ) ;
  assign n16330 = ( ~n3092 & n4007 ) | ( ~n3092 & n16329 ) | ( n4007 & n16329 ) ;
  assign n16331 = n834 | n3320 ;
  assign n16332 = n16330 & ~n16331 ;
  assign n16333 = ( n2168 & ~n7605 ) | ( n2168 & n9984 ) | ( ~n7605 & n9984 ) ;
  assign n16334 = ( n14246 & n16332 ) | ( n14246 & n16333 ) | ( n16332 & n16333 ) ;
  assign n16335 = n2600 & ~n16334 ;
  assign n16336 = n16328 & n16335 ;
  assign n16339 = n9023 ^ n4707 ^ 1'b0 ;
  assign n16337 = ~n10850 & n12340 ;
  assign n16338 = ( n2550 & n12419 ) | ( n2550 & ~n16337 ) | ( n12419 & ~n16337 ) ;
  assign n16340 = n16339 ^ n16338 ^ n2234 ;
  assign n16341 = n7056 | n7612 ;
  assign n16342 = n16341 ^ n14789 ^ n829 ;
  assign n16355 = n4581 ^ n3741 ^ 1'b0 ;
  assign n16356 = n4768 & n16355 ;
  assign n16354 = n7442 ^ n1872 ^ n1712 ;
  assign n16353 = ( n342 & n10223 ) | ( n342 & n13440 ) | ( n10223 & n13440 ) ;
  assign n16357 = n16356 ^ n16354 ^ n16353 ;
  assign n16343 = n13440 ^ n11536 ^ 1'b0 ;
  assign n16348 = ( n933 & ~n2340 ) | ( n933 & n4073 ) | ( ~n2340 & n4073 ) ;
  assign n16346 = ~n7799 & n8807 ;
  assign n16347 = n16346 ^ n3110 ^ 1'b0 ;
  assign n16344 = n4210 & ~n4981 ;
  assign n16345 = n7487 & n16344 ;
  assign n16349 = n16348 ^ n16347 ^ n16345 ;
  assign n16350 = ~n16343 & n16349 ;
  assign n16351 = ~n7021 & n16350 ;
  assign n16352 = n16351 ^ n13531 ^ 1'b0 ;
  assign n16358 = n16357 ^ n16352 ^ n9741 ;
  assign n16359 = n4160 ^ n4041 ^ x12 ;
  assign n16360 = n11190 ^ n10900 ^ n10352 ;
  assign n16361 = n16360 ^ n15066 ^ n14650 ;
  assign n16362 = ~n16359 & n16361 ;
  assign n16363 = n16362 ^ n2237 ^ 1'b0 ;
  assign n16364 = n3516 ^ n3000 ^ 1'b0 ;
  assign n16365 = n16364 ^ n10662 ^ 1'b0 ;
  assign n16366 = ~n5426 & n16365 ;
  assign n16368 = n7209 ^ n598 ^ 1'b0 ;
  assign n16369 = n4446 & n16368 ;
  assign n16370 = n7480 ^ n6570 ^ 1'b0 ;
  assign n16371 = n16369 & n16370 ;
  assign n16367 = n12013 ^ n692 ^ 1'b0 ;
  assign n16372 = n16371 ^ n16367 ^ n8898 ;
  assign n16373 = n16372 ^ n10149 ^ 1'b0 ;
  assign n16374 = ( n1108 & n1116 ) | ( n1108 & n6184 ) | ( n1116 & n6184 ) ;
  assign n16375 = n4877 | n6325 ;
  assign n16376 = n16375 ^ n11942 ^ n4555 ;
  assign n16377 = n16376 ^ n11008 ^ n3448 ;
  assign n16378 = ( n2209 & n6381 ) | ( n2209 & ~n11153 ) | ( n6381 & ~n11153 ) ;
  assign n16379 = n10076 & n16378 ;
  assign n16380 = ~n9055 & n16379 ;
  assign n16381 = n6396 ^ n1022 ^ 1'b0 ;
  assign n16382 = n3663 | n16381 ;
  assign n16383 = n6006 & n16382 ;
  assign n16384 = n12739 & n16383 ;
  assign n16385 = ( n910 & n6600 ) | ( n910 & n11335 ) | ( n6600 & n11335 ) ;
  assign n16386 = n2121 & n8371 ;
  assign n16387 = n1633 & ~n16386 ;
  assign n16389 = n12370 ^ n593 ^ 1'b0 ;
  assign n16390 = n7393 & n16389 ;
  assign n16388 = n1266 ^ n257 ^ 1'b0 ;
  assign n16391 = n16390 ^ n16388 ^ n14466 ;
  assign n16392 = n7022 ^ n6926 ^ 1'b0 ;
  assign n16393 = n12384 ^ n3178 ^ x21 ;
  assign n16394 = n6966 & ~n16393 ;
  assign n16395 = n5667 & n16394 ;
  assign n16396 = n16395 ^ n10424 ^ 1'b0 ;
  assign n16397 = ~n16392 & n16396 ;
  assign n16398 = n16397 ^ n15435 ^ 1'b0 ;
  assign n16399 = n15929 ^ n13156 ^ 1'b0 ;
  assign n16400 = n16399 ^ n11562 ^ 1'b0 ;
  assign n16401 = ( n3037 & ~n15372 ) | ( n3037 & n16400 ) | ( ~n15372 & n16400 ) ;
  assign n16408 = n7083 ^ n1282 ^ 1'b0 ;
  assign n16402 = n8209 ^ n1201 ^ 1'b0 ;
  assign n16403 = n10030 & n16402 ;
  assign n16404 = n13154 ^ n2986 ^ 1'b0 ;
  assign n16405 = ~n4691 & n16404 ;
  assign n16406 = n1793 & n16405 ;
  assign n16407 = ~n16403 & n16406 ;
  assign n16409 = n16408 ^ n16407 ^ 1'b0 ;
  assign n16410 = n1558 & n9775 ;
  assign n16411 = ( ~n4580 & n7492 ) | ( ~n4580 & n16410 ) | ( n7492 & n16410 ) ;
  assign n16412 = n16411 ^ n11950 ^ n10766 ;
  assign n16413 = n258 & n6677 ;
  assign n16414 = n16412 & n16413 ;
  assign n16415 = n16414 ^ n7072 ^ 1'b0 ;
  assign n16416 = n5933 & n16415 ;
  assign n16417 = ( ~n4884 & n11906 ) | ( ~n4884 & n12274 ) | ( n11906 & n12274 ) ;
  assign n16418 = ~n2889 & n12686 ;
  assign n16419 = n16417 & n16418 ;
  assign n16420 = n6056 | n16419 ;
  assign n16421 = ~n4398 & n12686 ;
  assign n16422 = ~n2714 & n16421 ;
  assign n16423 = ( n5042 & n6938 ) | ( n5042 & n16422 ) | ( n6938 & n16422 ) ;
  assign n16424 = n16423 ^ n14347 ^ n2490 ;
  assign n16425 = n16424 ^ n8699 ^ 1'b0 ;
  assign n16426 = n16420 | n16425 ;
  assign n16427 = n5110 ^ x42 ^ 1'b0 ;
  assign n16428 = n4373 & n16427 ;
  assign n16429 = n796 | n4077 ;
  assign n16430 = n16428 | n16429 ;
  assign n16431 = ( n1466 & ~n8139 ) | ( n1466 & n16430 ) | ( ~n8139 & n16430 ) ;
  assign n16432 = n12505 ^ n8579 ^ x124 ;
  assign n16433 = n4846 ^ n4373 ^ 1'b0 ;
  assign n16434 = ~n2120 & n16433 ;
  assign n16435 = n821 | n16434 ;
  assign n16436 = n16435 ^ n9176 ^ 1'b0 ;
  assign n16437 = ( n3383 & ~n16347 ) | ( n3383 & n16436 ) | ( ~n16347 & n16436 ) ;
  assign n16438 = n7988 & ~n16437 ;
  assign n16439 = n3627 & n5948 ;
  assign n16442 = n16221 ^ n14562 ^ 1'b0 ;
  assign n16440 = n11640 & ~n15256 ;
  assign n16441 = n16440 ^ n2187 ^ 1'b0 ;
  assign n16443 = n16442 ^ n16441 ^ n2625 ;
  assign n16445 = n5424 ^ n1643 ^ x231 ;
  assign n16444 = ~n11051 & n11732 ;
  assign n16446 = n16445 ^ n16444 ^ 1'b0 ;
  assign n16447 = ~n9366 & n16446 ;
  assign n16448 = n2512 & n10638 ;
  assign n16449 = n10832 ^ x210 ^ 1'b0 ;
  assign n16450 = n325 | n5424 ;
  assign n16451 = n16449 & ~n16450 ;
  assign n16452 = n16451 ^ n2067 ^ 1'b0 ;
  assign n16453 = n6994 | n16452 ;
  assign n16454 = n16448 & ~n16453 ;
  assign n16455 = n10029 & ~n16454 ;
  assign n16456 = n6585 & n16455 ;
  assign n16457 = n16390 ^ n16020 ^ n8514 ;
  assign n16458 = n16457 ^ n11964 ^ n2498 ;
  assign n16459 = n6723 | n16458 ;
  assign n16460 = n16459 ^ n8254 ^ 1'b0 ;
  assign n16461 = n16460 ^ n9761 ^ n2031 ;
  assign n16462 = ( n443 & ~n2376 ) | ( n443 & n12416 ) | ( ~n2376 & n12416 ) ;
  assign n16463 = n16462 ^ n13806 ^ n13351 ;
  assign n16464 = n15104 ^ n5420 ^ n2547 ;
  assign n16465 = ( x252 & n16463 ) | ( x252 & ~n16464 ) | ( n16463 & ~n16464 ) ;
  assign n16466 = ~n5034 & n16369 ;
  assign n16467 = n16466 ^ n6762 ^ 1'b0 ;
  assign n16468 = n7310 ^ n4316 ^ 1'b0 ;
  assign n16469 = n13847 ^ n11446 ^ 1'b0 ;
  assign n16470 = n10760 & n16469 ;
  assign n16471 = n264 & n1428 ;
  assign n16472 = n15468 ^ n11810 ^ n698 ;
  assign n16473 = ( ~n12940 & n16471 ) | ( ~n12940 & n16472 ) | ( n16471 & n16472 ) ;
  assign n16474 = n16473 ^ n2756 ^ 1'b0 ;
  assign n16475 = ( n4179 & ~n4952 ) | ( n4179 & n12509 ) | ( ~n4952 & n12509 ) ;
  assign n16476 = n16475 ^ n2456 ^ 1'b0 ;
  assign n16477 = n5411 & n16476 ;
  assign n16478 = ( n1922 & n10597 ) | ( n1922 & n11932 ) | ( n10597 & n11932 ) ;
  assign n16479 = ~n320 & n735 ;
  assign n16480 = ~n16478 & n16479 ;
  assign n16481 = n4057 ^ n1595 ^ n1086 ;
  assign n16482 = n16481 ^ n8619 ^ n1393 ;
  assign n16483 = n16482 ^ n6053 ^ n3435 ;
  assign n16486 = ~n1723 & n6242 ;
  assign n16487 = n16486 ^ n16464 ^ x119 ;
  assign n16484 = n9509 ^ n1881 ^ 1'b0 ;
  assign n16485 = n11407 | n16484 ;
  assign n16488 = n16487 ^ n16485 ^ 1'b0 ;
  assign n16489 = n16488 ^ n13430 ^ n9342 ;
  assign n16490 = ~n2771 & n6893 ;
  assign n16491 = n16490 ^ n6075 ^ n2964 ;
  assign n16492 = n16491 ^ n9311 ^ n6588 ;
  assign n16493 = n12801 ^ n7688 ^ 1'b0 ;
  assign n16495 = n5063 | n9796 ;
  assign n16496 = n16495 ^ n3437 ^ 1'b0 ;
  assign n16494 = n7004 ^ n5150 ^ n4780 ;
  assign n16497 = n16496 ^ n16494 ^ n15395 ;
  assign n16498 = n16497 ^ n10495 ^ 1'b0 ;
  assign n16499 = n1203 | n10374 ;
  assign n16500 = n16498 | n16499 ;
  assign n16501 = n14734 ^ n11099 ^ n1756 ;
  assign n16502 = n16501 ^ n8373 ^ n7979 ;
  assign n16503 = n14677 ^ n3114 ^ x68 ;
  assign n16504 = n16503 ^ n6245 ^ n4012 ;
  assign n16505 = x23 & n7709 ;
  assign n16506 = n16505 ^ n7753 ^ 1'b0 ;
  assign n16507 = ( n5588 & n16504 ) | ( n5588 & n16506 ) | ( n16504 & n16506 ) ;
  assign n16508 = n4619 ^ n3759 ^ n3200 ;
  assign n16509 = n2052 & n16508 ;
  assign n16510 = ~n4974 & n16509 ;
  assign n16511 = n16507 & n16510 ;
  assign n16512 = ( ~n4439 & n6196 ) | ( ~n4439 & n6803 ) | ( n6196 & n6803 ) ;
  assign n16513 = n11112 ^ n2320 ^ 1'b0 ;
  assign n16514 = n16512 | n16513 ;
  assign n16515 = n16514 ^ n2210 ^ 1'b0 ;
  assign n16516 = n16515 ^ n9232 ^ 1'b0 ;
  assign n16517 = n6029 ^ x65 ^ 1'b0 ;
  assign n16518 = ~n12138 & n16517 ;
  assign n16519 = ( n5179 & n14545 ) | ( n5179 & ~n14914 ) | ( n14545 & ~n14914 ) ;
  assign n16520 = n12946 ^ n8699 ^ 1'b0 ;
  assign n16521 = x77 & n16520 ;
  assign n16522 = n1906 & ~n16521 ;
  assign n16523 = n3067 & ~n7030 ;
  assign n16524 = ~n8449 & n16523 ;
  assign n16528 = n12921 ^ n12676 ^ n3949 ;
  assign n16525 = n3333 & ~n4814 ;
  assign n16526 = ~n12110 & n16525 ;
  assign n16527 = ( n7712 & ~n11593 ) | ( n7712 & n16526 ) | ( ~n11593 & n16526 ) ;
  assign n16529 = n16528 ^ n16527 ^ n15588 ;
  assign n16530 = ( n5737 & ~n6856 ) | ( n5737 & n13027 ) | ( ~n6856 & n13027 ) ;
  assign n16531 = n3466 ^ n3230 ^ 1'b0 ;
  assign n16532 = n2661 & ~n16531 ;
  assign n16533 = n13181 ^ n3740 ^ 1'b0 ;
  assign n16534 = n16532 & ~n16533 ;
  assign n16535 = ~n16530 & n16534 ;
  assign n16536 = n4673 ^ n3113 ^ 1'b0 ;
  assign n16537 = n5637 | n16536 ;
  assign n16538 = ( n6240 & ~n7401 ) | ( n6240 & n16537 ) | ( ~n7401 & n16537 ) ;
  assign n16539 = ~n418 & n16442 ;
  assign n16540 = ( ~n326 & n3781 ) | ( ~n326 & n11588 ) | ( n3781 & n11588 ) ;
  assign n16541 = ( ~n1634 & n5246 ) | ( ~n1634 & n9924 ) | ( n5246 & n9924 ) ;
  assign n16542 = n4720 | n16541 ;
  assign n16543 = n16542 ^ n7084 ^ 1'b0 ;
  assign n16544 = ( n4351 & n16540 ) | ( n4351 & ~n16543 ) | ( n16540 & ~n16543 ) ;
  assign n16545 = n16544 ^ n14241 ^ n9371 ;
  assign n16548 = n2874 ^ n2557 ^ 1'b0 ;
  assign n16546 = n13070 ^ n2977 ^ 1'b0 ;
  assign n16547 = ( n3659 & ~n16077 ) | ( n3659 & n16546 ) | ( ~n16077 & n16546 ) ;
  assign n16549 = n16548 ^ n16547 ^ n8933 ;
  assign n16550 = ( n2729 & n9633 ) | ( n2729 & n10165 ) | ( n9633 & n10165 ) ;
  assign n16551 = n5160 | n8180 ;
  assign n16552 = n16551 ^ n13299 ^ n5006 ;
  assign n16553 = n16552 ^ n4261 ^ n1648 ;
  assign n16554 = n5765 & ~n16553 ;
  assign n16555 = ( n2759 & n5834 ) | ( n2759 & n9786 ) | ( n5834 & n9786 ) ;
  assign n16556 = n12454 ^ n10423 ^ 1'b0 ;
  assign n16557 = ( ~n2707 & n2778 ) | ( ~n2707 & n16556 ) | ( n2778 & n16556 ) ;
  assign n16561 = n8222 ^ n5258 ^ n2220 ;
  assign n16562 = n7817 ^ n858 ^ 1'b0 ;
  assign n16563 = ~n16561 & n16562 ;
  assign n16564 = n16563 ^ n16045 ^ n8886 ;
  assign n16558 = n3426 ^ n3329 ^ 1'b0 ;
  assign n16559 = ~n1545 & n16558 ;
  assign n16560 = n16559 ^ n10958 ^ 1'b0 ;
  assign n16565 = n16564 ^ n16560 ^ n4848 ;
  assign n16566 = n16565 ^ n13231 ^ n9761 ;
  assign n16567 = ~n1666 & n11028 ;
  assign n16568 = n16567 ^ n11968 ^ x186 ;
  assign n16569 = n10695 ^ n9263 ^ n5685 ;
  assign n16570 = n5426 ^ n4456 ^ 1'b0 ;
  assign n16571 = ( n4049 & n8415 ) | ( n4049 & n16570 ) | ( n8415 & n16570 ) ;
  assign n16572 = n11788 ^ n6437 ^ 1'b0 ;
  assign n16573 = n12881 ^ n9235 ^ n7258 ;
  assign n16574 = n2765 & ~n16573 ;
  assign n16575 = ~x117 & n16574 ;
  assign n16576 = n16575 ^ n12730 ^ 1'b0 ;
  assign n16577 = ~n2365 & n16576 ;
  assign n16578 = n16577 ^ n14606 ^ n5715 ;
  assign n16585 = x154 & n7079 ;
  assign n16586 = ( n1039 & n3835 ) | ( n1039 & n16585 ) | ( n3835 & n16585 ) ;
  assign n16587 = ( n7448 & n10494 ) | ( n7448 & n14020 ) | ( n10494 & n14020 ) ;
  assign n16588 = ~n16586 & n16587 ;
  assign n16589 = n16588 ^ n12608 ^ n9357 ;
  assign n16582 = n841 & n11297 ;
  assign n16583 = ~n5227 & n16582 ;
  assign n16579 = n7577 ^ n3219 ^ 1'b0 ;
  assign n16580 = n6038 | n16579 ;
  assign n16581 = ( n6775 & n12307 ) | ( n6775 & n16580 ) | ( n12307 & n16580 ) ;
  assign n16584 = n16583 ^ n16581 ^ 1'b0 ;
  assign n16590 = n16589 ^ n16584 ^ n15790 ;
  assign n16591 = n4173 | n13442 ;
  assign n16592 = ( n9969 & n14856 ) | ( n9969 & ~n16591 ) | ( n14856 & ~n16591 ) ;
  assign n16595 = n2528 & n3138 ;
  assign n16593 = n8785 ^ n698 ^ 1'b0 ;
  assign n16594 = n6704 & n16593 ;
  assign n16596 = n16595 ^ n16594 ^ n8411 ;
  assign n16597 = n3522 & n9930 ;
  assign n16598 = n1692 | n16597 ;
  assign n16599 = n5297 & ~n16598 ;
  assign n16600 = n12821 & n16599 ;
  assign n16602 = n6907 ^ n1176 ^ n606 ;
  assign n16603 = n7707 & n16602 ;
  assign n16604 = n4551 & ~n16603 ;
  assign n16601 = n1953 ^ n1537 ^ 1'b0 ;
  assign n16605 = n16604 ^ n16601 ^ 1'b0 ;
  assign n16606 = n12543 & n16605 ;
  assign n16607 = ~n13115 & n16606 ;
  assign n16608 = n15305 | n16004 ;
  assign n16609 = n16608 ^ n3314 ^ 1'b0 ;
  assign n16610 = n6287 ^ n1713 ^ 1'b0 ;
  assign n16611 = n13773 ^ n4441 ^ 1'b0 ;
  assign n16614 = n2314 ^ n433 ^ 1'b0 ;
  assign n16615 = n1693 | n16614 ;
  assign n16613 = ( ~n3484 & n7763 ) | ( ~n3484 & n9233 ) | ( n7763 & n9233 ) ;
  assign n16616 = n16615 ^ n16613 ^ n11914 ;
  assign n16617 = n6349 ^ n978 ^ 1'b0 ;
  assign n16618 = n16616 & ~n16617 ;
  assign n16612 = n4788 & ~n11450 ;
  assign n16619 = n16618 ^ n16612 ^ 1'b0 ;
  assign n16620 = n4034 | n11521 ;
  assign n16621 = n9483 | n13616 ;
  assign n16622 = ~n2810 & n7702 ;
  assign n16623 = n16622 ^ n10727 ^ n3785 ;
  assign n16624 = ( n368 & ~n15219 ) | ( n368 & n16623 ) | ( ~n15219 & n16623 ) ;
  assign n16625 = ( n923 & n1731 ) | ( n923 & n5359 ) | ( n1731 & n5359 ) ;
  assign n16626 = n16625 ^ n16160 ^ n7572 ;
  assign n16627 = n6613 & ~n13317 ;
  assign n16628 = n16627 ^ n3587 ^ 1'b0 ;
  assign n16629 = n7904 & n16352 ;
  assign n16630 = n13718 ^ n10992 ^ n10383 ;
  assign n16631 = n10664 ^ n7639 ^ 1'b0 ;
  assign n16632 = n16630 | n16631 ;
  assign n16634 = ~n1394 & n3110 ;
  assign n16633 = n12906 | n15104 ;
  assign n16635 = n16634 ^ n16633 ^ n1914 ;
  assign n16636 = ( n9513 & ~n16632 ) | ( n9513 & n16635 ) | ( ~n16632 & n16635 ) ;
  assign n16637 = ( n3823 & n9203 ) | ( n3823 & ~n10594 ) | ( n9203 & ~n10594 ) ;
  assign n16638 = n13059 ^ n6618 ^ 1'b0 ;
  assign n16639 = n10107 & ~n16638 ;
  assign n16640 = ( x139 & n2510 ) | ( x139 & ~n4707 ) | ( n2510 & ~n4707 ) ;
  assign n16641 = n15053 & n16640 ;
  assign n16642 = ~n3896 & n16641 ;
  assign n16643 = ( n662 & n16639 ) | ( n662 & n16642 ) | ( n16639 & n16642 ) ;
  assign n16644 = n11705 ^ n7388 ^ 1'b0 ;
  assign n16645 = n4871 ^ n3799 ^ n2892 ;
  assign n16646 = n5367 & n16049 ;
  assign n16647 = ~n16645 & n16646 ;
  assign n16648 = n16647 ^ n8438 ^ 1'b0 ;
  assign n16649 = n4582 | n5241 ;
  assign n16650 = n16649 ^ n1545 ^ 1'b0 ;
  assign n16651 = n16648 & ~n16650 ;
  assign n16652 = ~n16644 & n16651 ;
  assign n16656 = ~n4877 & n7659 ;
  assign n16653 = n1840 & ~n2410 ;
  assign n16654 = n16653 ^ n3994 ^ 1'b0 ;
  assign n16655 = x42 | n16654 ;
  assign n16657 = n16656 ^ n16655 ^ n6969 ;
  assign n16658 = n7958 & ~n9892 ;
  assign n16659 = n3374 & n16658 ;
  assign n16662 = ~n7795 & n10337 ;
  assign n16660 = ~n1108 & n13767 ;
  assign n16661 = n8919 & ~n16660 ;
  assign n16663 = n16662 ^ n16661 ^ 1'b0 ;
  assign n16664 = n16663 ^ n14170 ^ 1'b0 ;
  assign n16665 = ( n301 & ~n16659 ) | ( n301 & n16664 ) | ( ~n16659 & n16664 ) ;
  assign n16666 = n4884 ^ n4489 ^ 1'b0 ;
  assign n16667 = n5792 & n16666 ;
  assign n16668 = n393 & n7932 ;
  assign n16669 = n9254 & ~n16668 ;
  assign n16670 = ~n16667 & n16669 ;
  assign n16671 = n16670 ^ n7432 ^ 1'b0 ;
  assign n16672 = n15226 & n16671 ;
  assign n16673 = n8822 & n16672 ;
  assign n16674 = n5914 ^ n3626 ^ 1'b0 ;
  assign n16675 = n4899 & n16674 ;
  assign n16676 = n16675 ^ n5773 ^ n5533 ;
  assign n16677 = n16676 ^ n16082 ^ n6078 ;
  assign n16678 = n16677 ^ n8262 ^ n5404 ;
  assign n16680 = ( n2380 & n4754 ) | ( n2380 & ~n13500 ) | ( n4754 & ~n13500 ) ;
  assign n16679 = n10700 ^ n3380 ^ 1'b0 ;
  assign n16681 = n16680 ^ n16679 ^ n2943 ;
  assign n16682 = n16681 ^ n3230 ^ n3190 ;
  assign n16685 = n1648 | n6265 ;
  assign n16686 = n6265 & ~n16685 ;
  assign n16687 = n2192 | n3562 ;
  assign n16688 = n2192 & ~n16687 ;
  assign n16689 = n5121 | n16688 ;
  assign n16690 = n16686 & ~n16689 ;
  assign n16691 = n662 & ~n3530 ;
  assign n16692 = ( n4348 & n16690 ) | ( n4348 & ~n16691 ) | ( n16690 & ~n16691 ) ;
  assign n16683 = ~n1581 & n13519 ;
  assign n16684 = ~n6384 & n16683 ;
  assign n16693 = n16692 ^ n16684 ^ n7774 ;
  assign n16694 = ( ~n2375 & n4147 ) | ( ~n2375 & n9365 ) | ( n4147 & n9365 ) ;
  assign n16695 = n16694 ^ n13906 ^ n2553 ;
  assign n16696 = n7633 ^ n4899 ^ n1813 ;
  assign n16697 = n1725 & ~n16696 ;
  assign n16698 = n9949 ^ n6106 ^ n436 ;
  assign n16699 = ~n7493 & n11784 ;
  assign n16701 = n6297 ^ n4747 ^ 1'b0 ;
  assign n16702 = ( x15 & n10911 ) | ( x15 & n16701 ) | ( n10911 & n16701 ) ;
  assign n16703 = n807 & n16702 ;
  assign n16704 = n14542 ^ n9448 ^ 1'b0 ;
  assign n16705 = n8634 & n16704 ;
  assign n16706 = n16705 ^ n12302 ^ x30 ;
  assign n16707 = ( n6780 & n16703 ) | ( n6780 & ~n16706 ) | ( n16703 & ~n16706 ) ;
  assign n16700 = n15433 | n15669 ;
  assign n16708 = n16707 ^ n16700 ^ 1'b0 ;
  assign n16709 = n868 ^ x72 ^ 1'b0 ;
  assign n16710 = ~n14552 & n16709 ;
  assign n16711 = n3796 & n9026 ;
  assign n16712 = n4848 & n16711 ;
  assign n16713 = n7815 & ~n16712 ;
  assign n16714 = ( ~n2351 & n2899 ) | ( ~n2351 & n15984 ) | ( n2899 & n15984 ) ;
  assign n16715 = ( n525 & ~n5890 ) | ( n525 & n16714 ) | ( ~n5890 & n16714 ) ;
  assign n16716 = n16713 | n16715 ;
  assign n16717 = ( n3344 & n9489 ) | ( n3344 & n10095 ) | ( n9489 & n10095 ) ;
  assign n16718 = n15550 ^ n10472 ^ 1'b0 ;
  assign n16719 = ~n16717 & n16718 ;
  assign n16720 = n4804 ^ n4052 ^ 1'b0 ;
  assign n16721 = ( n7117 & n13132 ) | ( n7117 & ~n16720 ) | ( n13132 & ~n16720 ) ;
  assign n16722 = ( n2313 & n5352 ) | ( n2313 & ~n10828 ) | ( n5352 & ~n10828 ) ;
  assign n16723 = n16722 ^ n13886 ^ n1773 ;
  assign n16724 = ( n9969 & ~n10677 ) | ( n9969 & n11848 ) | ( ~n10677 & n11848 ) ;
  assign n16725 = n16724 ^ n13992 ^ n5589 ;
  assign n16726 = n15040 ^ n3948 ^ 1'b0 ;
  assign n16727 = ( ~n2057 & n16725 ) | ( ~n2057 & n16726 ) | ( n16725 & n16726 ) ;
  assign n16728 = ~n598 & n1113 ;
  assign n16729 = n16728 ^ n697 ^ 1'b0 ;
  assign n16730 = ( ~n7705 & n12740 ) | ( ~n7705 & n16729 ) | ( n12740 & n16729 ) ;
  assign n16731 = n16730 ^ n13788 ^ n4365 ;
  assign n16732 = x51 & n6633 ;
  assign n16733 = n3537 & n11077 ;
  assign n16734 = n16733 ^ x126 ^ 1'b0 ;
  assign n16735 = n16732 | n16734 ;
  assign n16736 = n16735 ^ n5665 ^ 1'b0 ;
  assign n16737 = ( n3025 & n3522 ) | ( n3025 & n3799 ) | ( n3522 & n3799 ) ;
  assign n16738 = ~n16736 & n16737 ;
  assign n16739 = ( x208 & ~n4662 ) | ( x208 & n16738 ) | ( ~n4662 & n16738 ) ;
  assign n16745 = ( n1575 & ~n3254 ) | ( n1575 & n7014 ) | ( ~n3254 & n7014 ) ;
  assign n16743 = n11511 ^ n7518 ^ n4144 ;
  assign n16741 = n9448 ^ n4141 ^ n2070 ;
  assign n16740 = n6104 | n8719 ;
  assign n16742 = n16741 ^ n16740 ^ 1'b0 ;
  assign n16744 = n16743 ^ n16742 ^ n7919 ;
  assign n16746 = n16745 ^ n16744 ^ n8813 ;
  assign n16747 = n1637 & ~n1676 ;
  assign n16748 = ~n16746 & n16747 ;
  assign n16749 = n16145 ^ n5302 ^ n4822 ;
  assign n16750 = n8748 | n11554 ;
  assign n16751 = n13045 ^ n8134 ^ n3668 ;
  assign n16752 = n12563 ^ n5978 ^ n3085 ;
  assign n16753 = n16752 ^ n7791 ^ n2450 ;
  assign n16754 = ( n3259 & n10052 ) | ( n3259 & n10308 ) | ( n10052 & n10308 ) ;
  assign n16755 = ( n7126 & ~n10881 ) | ( n7126 & n13061 ) | ( ~n10881 & n13061 ) ;
  assign n16756 = ( n16753 & n16754 ) | ( n16753 & n16755 ) | ( n16754 & n16755 ) ;
  assign n16757 = n10212 ^ n6143 ^ n1158 ;
  assign n16759 = n16496 ^ n6743 ^ n3644 ;
  assign n16758 = n2681 | n13103 ;
  assign n16760 = n16759 ^ n16758 ^ 1'b0 ;
  assign n16761 = n1809 | n16760 ;
  assign n16762 = n10679 ^ n9121 ^ n4532 ;
  assign n16763 = n16762 ^ n1039 ^ 1'b0 ;
  assign n16764 = n6873 ^ n5204 ^ n1315 ;
  assign n16765 = n8785 ^ n1906 ^ 1'b0 ;
  assign n16766 = n16764 & n16765 ;
  assign n16767 = n16766 ^ n10337 ^ 1'b0 ;
  assign n16768 = n13801 & ~n16767 ;
  assign n16769 = ( n12278 & ~n16763 ) | ( n12278 & n16768 ) | ( ~n16763 & n16768 ) ;
  assign n16770 = n13709 ^ n355 ^ 1'b0 ;
  assign n16771 = ~n1293 & n16770 ;
  assign n16772 = n16771 ^ n9947 ^ 1'b0 ;
  assign n16773 = ( n625 & n3167 ) | ( n625 & n8465 ) | ( n3167 & n8465 ) ;
  assign n16774 = n2127 | n4454 ;
  assign n16775 = n16773 | n16774 ;
  assign n16776 = n11079 & n16775 ;
  assign n16777 = n16776 ^ n11670 ^ x81 ;
  assign n16778 = n15363 ^ n10052 ^ n1960 ;
  assign n16779 = n429 | n3358 ;
  assign n16780 = ~n5839 & n11686 ;
  assign n16781 = ~n439 & n16780 ;
  assign n16789 = n14381 ^ n1718 ^ 1'b0 ;
  assign n16790 = ~n1425 & n16789 ;
  assign n16783 = n791 & ~n5102 ;
  assign n16784 = n1333 & n16783 ;
  assign n16782 = n3887 & ~n5013 ;
  assign n16785 = n16784 ^ n16782 ^ 1'b0 ;
  assign n16786 = ~n1676 & n3365 ;
  assign n16787 = n16786 ^ n10042 ^ 1'b0 ;
  assign n16788 = n16785 & n16787 ;
  assign n16791 = n16790 ^ n16788 ^ 1'b0 ;
  assign n16792 = ~n16781 & n16791 ;
  assign n16793 = n16792 ^ n10446 ^ 1'b0 ;
  assign n16794 = n1069 & n4106 ;
  assign n16795 = ( n2173 & ~n3314 ) | ( n2173 & n5387 ) | ( ~n3314 & n5387 ) ;
  assign n16796 = n3331 ^ n2859 ^ n2010 ;
  assign n16797 = n16795 & n16796 ;
  assign n16798 = n6531 & ~n10138 ;
  assign n16799 = n16798 ^ n14593 ^ x37 ;
  assign n16800 = ( ~n5135 & n8898 ) | ( ~n5135 & n16333 ) | ( n8898 & n16333 ) ;
  assign n16801 = n2065 & n14449 ;
  assign n16802 = n12122 & n16801 ;
  assign n16803 = x192 & n13432 ;
  assign n16804 = n2904 & ~n11952 ;
  assign n16805 = n5362 ^ n5361 ^ 1'b0 ;
  assign n16806 = ( ~n4493 & n11171 ) | ( ~n4493 & n15702 ) | ( n11171 & n15702 ) ;
  assign n16807 = n11195 ^ n3132 ^ 1'b0 ;
  assign n16808 = ( n1003 & n8923 ) | ( n1003 & ~n12979 ) | ( n8923 & ~n12979 ) ;
  assign n16809 = n7880 ^ n6756 ^ n1315 ;
  assign n16810 = n7369 ^ n3368 ^ 1'b0 ;
  assign n16811 = ( n615 & ~n5385 ) | ( n615 & n10946 ) | ( ~n5385 & n10946 ) ;
  assign n16812 = n16811 ^ n4046 ^ 1'b0 ;
  assign n16813 = n5553 ^ n4696 ^ 1'b0 ;
  assign n16814 = n16762 ^ n12515 ^ 1'b0 ;
  assign n16815 = ~n898 & n16814 ;
  assign n16816 = ( n9142 & n16813 ) | ( n9142 & n16815 ) | ( n16813 & n16815 ) ;
  assign n16817 = n16238 ^ n13617 ^ n3814 ;
  assign n16818 = n6094 ^ n3221 ^ 1'b0 ;
  assign n16819 = n9570 & n16818 ;
  assign n16820 = ( ~n3124 & n8503 ) | ( ~n3124 & n9489 ) | ( n8503 & n9489 ) ;
  assign n16821 = n16820 ^ n16213 ^ n6006 ;
  assign n16822 = n10996 ^ x55 ^ 1'b0 ;
  assign n16823 = ~n11529 & n16822 ;
  assign n16824 = ( n3293 & n4585 ) | ( n3293 & ~n12060 ) | ( n4585 & ~n12060 ) ;
  assign n16825 = n16824 ^ n9325 ^ n946 ;
  assign n16826 = ( ~n662 & n13486 ) | ( ~n662 & n15157 ) | ( n13486 & n15157 ) ;
  assign n16827 = n6076 | n6503 ;
  assign n16828 = n16827 ^ n9043 ^ 1'b0 ;
  assign n16829 = n6035 ^ n4804 ^ 1'b0 ;
  assign n16830 = n16829 ^ n6992 ^ n2790 ;
  assign n16832 = n3237 | n3768 ;
  assign n16831 = ( ~n6294 & n8567 ) | ( ~n6294 & n10205 ) | ( n8567 & n10205 ) ;
  assign n16833 = n16832 ^ n16831 ^ 1'b0 ;
  assign n16834 = ~n16830 & n16833 ;
  assign n16835 = n10057 & ~n13929 ;
  assign n16836 = n16835 ^ n3174 ^ 1'b0 ;
  assign n16837 = n6706 & ~n7565 ;
  assign n16838 = n6162 ^ n1602 ^ n1308 ;
  assign n16839 = n4562 ^ n2779 ^ 1'b0 ;
  assign n16840 = ( n10494 & n16838 ) | ( n10494 & n16839 ) | ( n16838 & n16839 ) ;
  assign n16841 = ( n541 & ~n16837 ) | ( n541 & n16840 ) | ( ~n16837 & n16840 ) ;
  assign n16842 = ( n2940 & ~n3503 ) | ( n2940 & n3861 ) | ( ~n3503 & n3861 ) ;
  assign n16843 = n16842 ^ n1277 ^ 1'b0 ;
  assign n16844 = n15884 & n16843 ;
  assign n16845 = n16844 ^ n8506 ^ 1'b0 ;
  assign n16846 = n6828 & ~n16845 ;
  assign n16847 = ( n2638 & ~n4182 ) | ( n2638 & n8659 ) | ( ~n4182 & n8659 ) ;
  assign n16848 = ( n16841 & n16846 ) | ( n16841 & n16847 ) | ( n16846 & n16847 ) ;
  assign n16849 = ( x109 & ~n2490 ) | ( x109 & n3753 ) | ( ~n2490 & n3753 ) ;
  assign n16850 = n16849 ^ n9914 ^ n2121 ;
  assign n16851 = n3579 & ~n14620 ;
  assign n16852 = ~n16546 & n16851 ;
  assign n16853 = n12486 ^ n7434 ^ n3794 ;
  assign n16854 = n16853 ^ n14172 ^ n12889 ;
  assign n16855 = ~n7203 & n10067 ;
  assign n16856 = n11917 ^ n8527 ^ x12 ;
  assign n16857 = n16856 ^ n7654 ^ n4090 ;
  assign n16858 = ~n2589 & n4571 ;
  assign n16859 = n16857 | n16858 ;
  assign n16860 = n16859 ^ n10468 ^ 1'b0 ;
  assign n16861 = n4334 & n10379 ;
  assign n16862 = n4824 ^ n2619 ^ 1'b0 ;
  assign n16863 = ~n10054 & n12573 ;
  assign n16864 = n16863 ^ n5464 ^ 1'b0 ;
  assign n16865 = n5693 & n16864 ;
  assign n16866 = ~x188 & n1220 ;
  assign n16867 = ~n3083 & n12089 ;
  assign n16868 = n16867 ^ n6806 ^ 1'b0 ;
  assign n16869 = n8607 ^ n4245 ^ 1'b0 ;
  assign n16870 = n8250 & n16869 ;
  assign n16871 = n16870 ^ n8094 ^ 1'b0 ;
  assign n16872 = ( n16866 & ~n16868 ) | ( n16866 & n16871 ) | ( ~n16868 & n16871 ) ;
  assign n16876 = ~n784 & n6477 ;
  assign n16877 = n16876 ^ n260 ^ 1'b0 ;
  assign n16873 = n5410 ^ n4923 ^ 1'b0 ;
  assign n16874 = n16873 ^ n16670 ^ 1'b0 ;
  assign n16875 = n16874 ^ n9671 ^ n6428 ;
  assign n16878 = n16877 ^ n16875 ^ n2104 ;
  assign n16879 = ( ~n2191 & n7147 ) | ( ~n2191 & n11349 ) | ( n7147 & n11349 ) ;
  assign n16880 = ( n6773 & ~n15640 ) | ( n6773 & n16879 ) | ( ~n15640 & n16879 ) ;
  assign n16882 = n16597 ^ n10836 ^ n1538 ;
  assign n16881 = n5662 & ~n5921 ;
  assign n16883 = n16882 ^ n16881 ^ 1'b0 ;
  assign n16884 = ( n9418 & n15941 ) | ( n9418 & n16883 ) | ( n15941 & n16883 ) ;
  assign n16885 = n3715 ^ n3492 ^ 1'b0 ;
  assign n16886 = n16885 ^ n3775 ^ 1'b0 ;
  assign n16887 = n15681 ^ n1634 ^ 1'b0 ;
  assign n16888 = n16887 ^ n679 ^ 1'b0 ;
  assign n16889 = ( n2928 & n16886 ) | ( n2928 & n16888 ) | ( n16886 & n16888 ) ;
  assign n16890 = ( n4332 & n5683 ) | ( n4332 & n7675 ) | ( n5683 & n7675 ) ;
  assign n16891 = n15104 ^ n4063 ^ 1'b0 ;
  assign n16892 = n287 & n16891 ;
  assign n16893 = ( n16813 & ~n16890 ) | ( n16813 & n16892 ) | ( ~n16890 & n16892 ) ;
  assign n16899 = n10019 ^ n6581 ^ 1'b0 ;
  assign n16900 = n6758 & n16899 ;
  assign n16894 = n6543 ^ n6427 ^ 1'b0 ;
  assign n16895 = n12865 ^ n4236 ^ n3042 ;
  assign n16896 = n16894 | n16895 ;
  assign n16897 = n16896 ^ n6393 ^ 1'b0 ;
  assign n16898 = n3630 & ~n16897 ;
  assign n16901 = n16900 ^ n16898 ^ 1'b0 ;
  assign n16902 = n5752 & n16901 ;
  assign n16903 = ( n6091 & n6162 ) | ( n6091 & n10475 ) | ( n6162 & n10475 ) ;
  assign n16904 = ~n2707 & n16903 ;
  assign n16906 = x131 & ~n12460 ;
  assign n16907 = n3204 & n16906 ;
  assign n16905 = n14019 ^ n10710 ^ n10009 ;
  assign n16908 = n16907 ^ n16905 ^ 1'b0 ;
  assign n16909 = n16904 & ~n16908 ;
  assign n16911 = n2214 | n4384 ;
  assign n16910 = n15575 ^ n7900 ^ 1'b0 ;
  assign n16912 = n16911 ^ n16910 ^ 1'b0 ;
  assign n16913 = n16909 & ~n16912 ;
  assign n16914 = ~n6822 & n12114 ;
  assign n16915 = n16913 & n16914 ;
  assign n16916 = n1922 & ~n11190 ;
  assign n16917 = n3648 & n16916 ;
  assign n16918 = ( ~n5373 & n5857 ) | ( ~n5373 & n16917 ) | ( n5857 & n16917 ) ;
  assign n16919 = ( n8623 & n13190 ) | ( n8623 & ~n16918 ) | ( n13190 & ~n16918 ) ;
  assign n16925 = n1934 ^ n988 ^ n778 ;
  assign n16926 = n16925 ^ n3527 ^ 1'b0 ;
  assign n16927 = n13557 & ~n16926 ;
  assign n16928 = n16927 ^ n3383 ^ 1'b0 ;
  assign n16920 = ~n4344 & n14784 ;
  assign n16921 = n13658 ^ n955 ^ x240 ;
  assign n16922 = n4192 & ~n16921 ;
  assign n16923 = n4443 & n10958 ;
  assign n16924 = ( n16920 & n16922 ) | ( n16920 & n16923 ) | ( n16922 & n16923 ) ;
  assign n16929 = n16928 ^ n16924 ^ n5895 ;
  assign n16930 = n3025 & n10834 ;
  assign n16931 = ~n2686 & n15436 ;
  assign n16932 = ~n16930 & n16931 ;
  assign n16933 = ~n16929 & n16932 ;
  assign n16934 = n2173 & ~n8979 ;
  assign n16935 = n16934 ^ n3406 ^ 1'b0 ;
  assign n16936 = ( n11545 & n12605 ) | ( n11545 & n16935 ) | ( n12605 & n16935 ) ;
  assign n16937 = n1890 | n16936 ;
  assign n16938 = n16937 ^ n8750 ^ 1'b0 ;
  assign n16939 = n16938 ^ n10895 ^ 1'b0 ;
  assign n16940 = ~n6799 & n9204 ;
  assign n16941 = n2776 ^ n1494 ^ 1'b0 ;
  assign n16942 = n15929 | n16941 ;
  assign n16943 = n16942 ^ n2609 ^ n2456 ;
  assign n16944 = n16943 ^ n14186 ^ n7940 ;
  assign n16945 = n8684 | n16944 ;
  assign n16946 = n14892 & ~n16945 ;
  assign n16950 = ( ~n3140 & n10042 ) | ( ~n3140 & n11927 ) | ( n10042 & n11927 ) ;
  assign n16947 = n1745 & ~n11995 ;
  assign n16948 = ~n9247 & n16947 ;
  assign n16949 = n15488 | n16948 ;
  assign n16951 = n16950 ^ n16949 ^ 1'b0 ;
  assign n16952 = n16951 ^ n401 ^ 1'b0 ;
  assign n16953 = n16946 | n16952 ;
  assign n16954 = n10740 ^ n4422 ^ 1'b0 ;
  assign n16955 = n16954 ^ n15909 ^ n9059 ;
  assign n16956 = n16955 ^ n2215 ^ 1'b0 ;
  assign n16957 = ~n12408 & n16956 ;
  assign n16958 = n10118 & n16957 ;
  assign n16959 = n16958 ^ n8926 ^ 1'b0 ;
  assign n16960 = ~n5180 & n16959 ;
  assign n16962 = n6359 & n10039 ;
  assign n16963 = n2199 & ~n16962 ;
  assign n16964 = n16963 ^ n4295 ^ 1'b0 ;
  assign n16961 = n2315 & ~n4594 ;
  assign n16965 = n16964 ^ n16961 ^ 1'b0 ;
  assign n16966 = n3056 | n9206 ;
  assign n16967 = n16966 ^ n12887 ^ 1'b0 ;
  assign n16968 = n7636 ^ n2959 ^ n1034 ;
  assign n16969 = n3749 & n16968 ;
  assign n16970 = ( n7325 & n16967 ) | ( n7325 & ~n16969 ) | ( n16967 & ~n16969 ) ;
  assign n16971 = ~n3922 & n9022 ;
  assign n16972 = ( n3103 & n16970 ) | ( n3103 & ~n16971 ) | ( n16970 & ~n16971 ) ;
  assign n16973 = ( n12415 & n12443 ) | ( n12415 & ~n16972 ) | ( n12443 & ~n16972 ) ;
  assign n16974 = n1152 & ~n13559 ;
  assign n16975 = n16974 ^ n8751 ^ n7867 ;
  assign n16976 = n3407 ^ n997 ^ 1'b0 ;
  assign n16977 = n13112 & n16976 ;
  assign n16978 = n2220 & n16977 ;
  assign n16979 = n6955 & n16978 ;
  assign n16980 = ( ~n1562 & n3624 ) | ( ~n1562 & n10385 ) | ( n3624 & n10385 ) ;
  assign n16981 = ( n15201 & ~n15863 ) | ( n15201 & n16980 ) | ( ~n15863 & n16980 ) ;
  assign n16982 = ( n7723 & n16979 ) | ( n7723 & n16981 ) | ( n16979 & n16981 ) ;
  assign n16983 = n15813 ^ n7812 ^ n4095 ;
  assign n16984 = n8841 | n16983 ;
  assign n16985 = n16984 ^ n3929 ^ 1'b0 ;
  assign n16986 = n16985 ^ n14939 ^ 1'b0 ;
  assign n16987 = n6410 & n16986 ;
  assign n16988 = n16249 ^ n12420 ^ n513 ;
  assign n16989 = ~n12269 & n16988 ;
  assign n16990 = n1510 & ~n16989 ;
  assign n16994 = n1031 | n7083 ;
  assign n16995 = n16994 ^ n7395 ^ 1'b0 ;
  assign n16992 = n3228 ^ n2074 ^ 1'b0 ;
  assign n16993 = ~n11992 & n16992 ;
  assign n16991 = x89 & n268 ;
  assign n16996 = n16995 ^ n16993 ^ n16991 ;
  assign n16997 = n16759 ^ n7323 ^ n7108 ;
  assign n16998 = n16997 ^ n16829 ^ n12930 ;
  assign n16999 = n14730 ^ n14583 ^ n11868 ;
  assign n17000 = ~n7230 & n14083 ;
  assign n17001 = ~n16999 & n17000 ;
  assign n17002 = n7581 ^ n808 ^ 1'b0 ;
  assign n17003 = n2521 & n17002 ;
  assign n17004 = ( n7223 & ~n8094 ) | ( n7223 & n12618 ) | ( ~n8094 & n12618 ) ;
  assign n17005 = n17004 ^ n1354 ^ 1'b0 ;
  assign n17007 = ~n6053 & n11073 ;
  assign n17008 = ~n6045 & n17007 ;
  assign n17006 = n2553 & ~n6648 ;
  assign n17009 = n17008 ^ n17006 ^ 1'b0 ;
  assign n17010 = n10361 & n13594 ;
  assign n17011 = n7177 & n16604 ;
  assign n17012 = n17011 ^ x161 ^ 1'b0 ;
  assign n17013 = n17012 ^ n14210 ^ n13209 ;
  assign n17014 = n17010 & ~n17013 ;
  assign n17015 = ( n627 & n815 ) | ( n627 & ~n14507 ) | ( n815 & ~n14507 ) ;
  assign n17016 = n7903 | n17015 ;
  assign n17017 = n6962 | n17016 ;
  assign n17020 = ~n270 & n7704 ;
  assign n17021 = n8330 & n17020 ;
  assign n17022 = n17021 ^ n7150 ^ 1'b0 ;
  assign n17023 = n4924 & ~n17022 ;
  assign n17024 = n17023 ^ n10327 ^ n9584 ;
  assign n17018 = ( ~n3215 & n7101 ) | ( ~n3215 & n10792 ) | ( n7101 & n10792 ) ;
  assign n17019 = n17018 ^ n3055 ^ 1'b0 ;
  assign n17025 = n17024 ^ n17019 ^ 1'b0 ;
  assign n17026 = n17017 & ~n17025 ;
  assign n17027 = n17026 ^ n1952 ^ 1'b0 ;
  assign n17028 = n5868 & n17027 ;
  assign n17029 = x167 & ~n1489 ;
  assign n17030 = n8551 & n17029 ;
  assign n17031 = n11848 | n17030 ;
  assign n17032 = ( n11661 & n13977 ) | ( n11661 & ~n17031 ) | ( n13977 & ~n17031 ) ;
  assign n17033 = ( n2680 & n2686 ) | ( n2680 & ~n5618 ) | ( n2686 & ~n5618 ) ;
  assign n17034 = ( n5676 & n14392 ) | ( n5676 & n17033 ) | ( n14392 & n17033 ) ;
  assign n17035 = n8857 ^ n4458 ^ n1528 ;
  assign n17036 = n15114 ^ n11590 ^ n9952 ;
  assign n17037 = n935 & n7640 ;
  assign n17038 = n17037 ^ n2838 ^ 1'b0 ;
  assign n17039 = n17038 ^ n8527 ^ 1'b0 ;
  assign n17040 = n17036 | n17039 ;
  assign n17045 = ~n4750 & n9535 ;
  assign n17046 = n17045 ^ n3375 ^ 1'b0 ;
  assign n17043 = ( n517 & ~n628 ) | ( n517 & n763 ) | ( ~n628 & n763 ) ;
  assign n17044 = n4404 | n17043 ;
  assign n17041 = ( n3865 & n5737 ) | ( n3865 & ~n14452 ) | ( n5737 & ~n14452 ) ;
  assign n17042 = ( n2662 & ~n6100 ) | ( n2662 & n17041 ) | ( ~n6100 & n17041 ) ;
  assign n17047 = n17046 ^ n17044 ^ n17042 ;
  assign n17048 = ( n14172 & ~n14416 ) | ( n14172 & n17047 ) | ( ~n14416 & n17047 ) ;
  assign n17049 = n17048 ^ n4346 ^ 1'b0 ;
  assign n17050 = n17049 ^ n13900 ^ n6829 ;
  assign n17051 = n2790 & ~n6269 ;
  assign n17052 = n17051 ^ n15232 ^ 1'b0 ;
  assign n17053 = n12989 ^ n2796 ^ n1508 ;
  assign n17054 = ( ~n8822 & n13430 ) | ( ~n8822 & n17053 ) | ( n13430 & n17053 ) ;
  assign n17055 = n17054 ^ n7448 ^ 1'b0 ;
  assign n17056 = n4753 | n17055 ;
  assign n17057 = ~n2950 & n6622 ;
  assign n17058 = n6270 & ~n17057 ;
  assign n17059 = n14112 ^ n12475 ^ n3655 ;
  assign n17060 = ~n17058 & n17059 ;
  assign n17061 = n14633 ^ n9257 ^ 1'b0 ;
  assign n17062 = n9182 & ~n17061 ;
  assign n17063 = n13879 & ~n17062 ;
  assign n17064 = n10647 ^ n6319 ^ 1'b0 ;
  assign n17065 = ~n2838 & n17064 ;
  assign n17066 = n7597 | n13149 ;
  assign n17067 = n17065 | n17066 ;
  assign n17068 = n17067 ^ n14967 ^ n5935 ;
  assign n17069 = n7557 ^ n2947 ^ n1359 ;
  assign n17070 = n10151 | n17069 ;
  assign n17071 = n17070 ^ n16419 ^ 1'b0 ;
  assign n17072 = n7129 ^ n4294 ^ 1'b0 ;
  assign n17073 = n3679 | n17072 ;
  assign n17074 = ( n9154 & n13915 ) | ( n9154 & n17073 ) | ( n13915 & n17073 ) ;
  assign n17079 = n423 | n539 ;
  assign n17080 = n8964 ^ n1723 ^ 1'b0 ;
  assign n17081 = n17079 & ~n17080 ;
  assign n17077 = n6159 ^ n4309 ^ n3209 ;
  assign n17078 = ~n8282 & n17077 ;
  assign n17082 = n17081 ^ n17078 ^ n14385 ;
  assign n17075 = ( n2023 & ~n4118 ) | ( n2023 & n15423 ) | ( ~n4118 & n15423 ) ;
  assign n17076 = n17075 ^ n14656 ^ n13042 ;
  assign n17083 = n17082 ^ n17076 ^ n11218 ;
  assign n17084 = n6615 ^ x150 ^ 1'b0 ;
  assign n17085 = n6913 | n17084 ;
  assign n17086 = n8689 ^ n6464 ^ n2693 ;
  assign n17087 = n16257 ^ n3303 ^ n2117 ;
  assign n17088 = n11074 | n17087 ;
  assign n17089 = n17086 & ~n17088 ;
  assign n17091 = n9324 ^ n6558 ^ n3430 ;
  assign n17090 = ~n4883 & n13319 ;
  assign n17092 = n17091 ^ n17090 ^ 1'b0 ;
  assign n17093 = n4642 ^ n4577 ^ n2390 ;
  assign n17094 = ( n7178 & n12660 ) | ( n7178 & n17093 ) | ( n12660 & n17093 ) ;
  assign n17095 = n10564 ^ n8212 ^ n3787 ;
  assign n17096 = ( n10641 & ~n11003 ) | ( n10641 & n13167 ) | ( ~n11003 & n13167 ) ;
  assign n17097 = n6956 ^ n745 ^ 1'b0 ;
  assign n17098 = ( ~n3911 & n4240 ) | ( ~n3911 & n8755 ) | ( n4240 & n8755 ) ;
  assign n17099 = ~n17097 & n17098 ;
  assign n17100 = n9997 ^ n884 ^ 1'b0 ;
  assign n17101 = n8847 & ~n17100 ;
  assign n17102 = ~n7946 & n16259 ;
  assign n17104 = n11387 ^ n3671 ^ n1077 ;
  assign n17103 = n1740 | n6702 ;
  assign n17105 = n17104 ^ n17103 ^ 1'b0 ;
  assign n17106 = ~n3608 & n4350 ;
  assign n17107 = ~n12300 & n17106 ;
  assign n17108 = n7164 ^ n861 ^ 1'b0 ;
  assign n17109 = n1494 & ~n10811 ;
  assign n17110 = ( ~n2184 & n6368 ) | ( ~n2184 & n9736 ) | ( n6368 & n9736 ) ;
  assign n17111 = n17110 ^ n11513 ^ 1'b0 ;
  assign n17112 = ( ~n6442 & n10587 ) | ( ~n6442 & n10904 ) | ( n10587 & n10904 ) ;
  assign n17113 = n12240 | n17112 ;
  assign n17128 = n10372 | n11837 ;
  assign n17129 = n463 | n17128 ;
  assign n17121 = n3922 | n7749 ;
  assign n17122 = n17121 ^ n2446 ^ 1'b0 ;
  assign n17114 = n8911 ^ n536 ^ 1'b0 ;
  assign n17115 = ( n6992 & n9119 ) | ( n6992 & ~n17114 ) | ( n9119 & ~n17114 ) ;
  assign n17116 = n7859 ^ n360 ^ 1'b0 ;
  assign n17117 = n8135 & n17116 ;
  assign n17118 = n17117 ^ n16287 ^ 1'b0 ;
  assign n17119 = ~n17115 & n17118 ;
  assign n17120 = n16567 & n17119 ;
  assign n17123 = n17122 ^ n17120 ^ x238 ;
  assign n17124 = ~n2841 & n4760 ;
  assign n17125 = n17124 ^ n13082 ^ 1'b0 ;
  assign n17126 = ~n15014 & n17125 ;
  assign n17127 = n17123 & n17126 ;
  assign n17130 = n17129 ^ n17127 ^ n8446 ;
  assign n17131 = n6832 ^ n4035 ^ 1'b0 ;
  assign n17132 = n534 | n17131 ;
  assign n17133 = n17132 ^ n3430 ^ 1'b0 ;
  assign n17134 = n12804 ^ n8514 ^ 1'b0 ;
  assign n17135 = n14583 & ~n17134 ;
  assign n17136 = n4414 & ~n17135 ;
  assign n17137 = ~n1550 & n17136 ;
  assign n17138 = n7409 & n17137 ;
  assign n17139 = n6989 ^ n6131 ^ n5724 ;
  assign n17140 = ( n2401 & n15783 ) | ( n2401 & n17139 ) | ( n15783 & n17139 ) ;
  assign n17141 = n17140 ^ n16616 ^ 1'b0 ;
  assign n17142 = n17141 ^ n4623 ^ n3646 ;
  assign n17143 = n15207 ^ n14534 ^ n5839 ;
  assign n17148 = ( n2503 & n4266 ) | ( n2503 & ~n9397 ) | ( n4266 & ~n9397 ) ;
  assign n17144 = n3577 & n7709 ;
  assign n17145 = n5926 & ~n17144 ;
  assign n17146 = n17145 ^ n8599 ^ 1'b0 ;
  assign n17147 = n17146 ^ x3 ^ 1'b0 ;
  assign n17149 = n17148 ^ n17147 ^ n2962 ;
  assign n17150 = n13153 ^ n10817 ^ n6493 ;
  assign n17151 = ( ~n753 & n4285 ) | ( ~n753 & n6379 ) | ( n4285 & n6379 ) ;
  assign n17152 = ( n7082 & ~n16245 ) | ( n7082 & n17151 ) | ( ~n16245 & n17151 ) ;
  assign n17153 = ~n17150 & n17152 ;
  assign n17154 = n13658 ^ n3210 ^ 1'b0 ;
  assign n17155 = n17154 ^ n7747 ^ n5715 ;
  assign n17156 = n13099 ^ n4674 ^ n1282 ;
  assign n17157 = n17156 ^ n4486 ^ 1'b0 ;
  assign n17158 = n17155 & n17157 ;
  assign n17160 = ( ~n6873 & n7824 ) | ( ~n6873 & n10345 ) | ( n7824 & n10345 ) ;
  assign n17159 = n8134 ^ n3454 ^ 1'b0 ;
  assign n17161 = n17160 ^ n17159 ^ n9162 ;
  assign n17166 = n13135 ^ n6168 ^ n1851 ;
  assign n17162 = n4090 & n11392 ;
  assign n17163 = ~n11379 & n17162 ;
  assign n17164 = n17163 ^ n12661 ^ 1'b0 ;
  assign n17165 = n5738 & ~n17164 ;
  assign n17167 = n17166 ^ n17165 ^ 1'b0 ;
  assign n17172 = n4972 ^ n4821 ^ 1'b0 ;
  assign n17168 = n8565 ^ n6622 ^ 1'b0 ;
  assign n17169 = n12161 & ~n17168 ;
  assign n17170 = n15792 ^ n9217 ^ x112 ;
  assign n17171 = ( n3630 & ~n17169 ) | ( n3630 & n17170 ) | ( ~n17169 & n17170 ) ;
  assign n17173 = n17172 ^ n17171 ^ n3155 ;
  assign n17174 = n4932 & n9702 ;
  assign n17175 = n407 & n17174 ;
  assign n17176 = n14158 & n16037 ;
  assign n17181 = n11089 ^ n8587 ^ n1972 ;
  assign n17177 = ~n704 & n8048 ;
  assign n17178 = n17177 ^ n10712 ^ 1'b0 ;
  assign n17179 = n17178 ^ n10302 ^ 1'b0 ;
  assign n17180 = n17179 ^ n13958 ^ n9976 ;
  assign n17182 = n17181 ^ n17180 ^ n1311 ;
  assign n17186 = n6928 ^ n5865 ^ n632 ;
  assign n17183 = n14431 ^ n5139 ^ 1'b0 ;
  assign n17184 = ( n1141 & n7292 ) | ( n1141 & n17183 ) | ( n7292 & n17183 ) ;
  assign n17185 = ( n811 & n2486 ) | ( n811 & n17184 ) | ( n2486 & n17184 ) ;
  assign n17187 = n17186 ^ n17185 ^ n670 ;
  assign n17191 = ( n941 & ~n6591 ) | ( n941 & n13390 ) | ( ~n6591 & n13390 ) ;
  assign n17190 = ( n6773 & n9606 ) | ( n6773 & n15678 ) | ( n9606 & n15678 ) ;
  assign n17188 = ( n9167 & n15159 ) | ( n9167 & n16244 ) | ( n15159 & n16244 ) ;
  assign n17189 = ( n4179 & ~n13027 ) | ( n4179 & n17188 ) | ( ~n13027 & n17188 ) ;
  assign n17192 = n17191 ^ n17190 ^ n17189 ;
  assign n17196 = n4581 ^ n3026 ^ 1'b0 ;
  assign n17197 = n14501 ^ n9208 ^ 1'b0 ;
  assign n17198 = n17196 | n17197 ;
  assign n17199 = n17198 ^ n8965 ^ 1'b0 ;
  assign n17193 = ( n949 & n8574 ) | ( n949 & n12457 ) | ( n8574 & n12457 ) ;
  assign n17194 = n15079 ^ n7565 ^ 1'b0 ;
  assign n17195 = n17193 | n17194 ;
  assign n17200 = n17199 ^ n17195 ^ n5501 ;
  assign n17201 = ( n1280 & ~n4604 ) | ( n1280 & n16775 ) | ( ~n4604 & n16775 ) ;
  assign n17202 = n17201 ^ n2735 ^ 1'b0 ;
  assign n17205 = n2580 | n15422 ;
  assign n17204 = n2692 ^ n1644 ^ n912 ;
  assign n17206 = n17205 ^ n17204 ^ n9211 ;
  assign n17207 = ( ~n2210 & n4676 ) | ( ~n2210 & n17206 ) | ( n4676 & n17206 ) ;
  assign n17203 = n3417 ^ n1988 ^ 1'b0 ;
  assign n17208 = n17207 ^ n17203 ^ 1'b0 ;
  assign n17209 = n17202 & ~n17208 ;
  assign n17210 = n5828 & n10808 ;
  assign n17213 = n6907 ^ n3233 ^ x222 ;
  assign n17211 = n2242 | n2602 ;
  assign n17212 = ~n4367 & n17211 ;
  assign n17214 = n17213 ^ n17212 ^ 1'b0 ;
  assign n17215 = ( ~n3625 & n15641 ) | ( ~n3625 & n17214 ) | ( n15641 & n17214 ) ;
  assign n17216 = n6561 & ~n16159 ;
  assign n17217 = ( n1124 & n6987 ) | ( n1124 & ~n17216 ) | ( n6987 & ~n17216 ) ;
  assign n17219 = n17058 ^ n12875 ^ n7756 ;
  assign n17218 = n9848 ^ n8133 ^ n1445 ;
  assign n17220 = n17219 ^ n17218 ^ n5383 ;
  assign n17221 = n9231 ^ n6204 ^ n2350 ;
  assign n17224 = n14873 ^ n9053 ^ 1'b0 ;
  assign n17225 = n6944 | n8689 ;
  assign n17226 = n4191 & ~n17225 ;
  assign n17227 = ~n14129 & n17226 ;
  assign n17228 = ~n17224 & n17227 ;
  assign n17229 = n15470 | n17228 ;
  assign n17230 = n17229 ^ x222 ^ 1'b0 ;
  assign n17222 = n10514 ^ n9678 ^ n4056 ;
  assign n17223 = n5421 & n17222 ;
  assign n17231 = n17230 ^ n17223 ^ 1'b0 ;
  assign n17232 = n4248 & ~n7567 ;
  assign n17233 = n17232 ^ n3166 ^ 1'b0 ;
  assign n17234 = n10913 & n17233 ;
  assign n17235 = n15694 ^ n8512 ^ 1'b0 ;
  assign n17236 = ~n5701 & n5798 ;
  assign n17237 = ~n1479 & n17236 ;
  assign n17238 = n17237 ^ n13580 ^ 1'b0 ;
  assign n17239 = n2176 & ~n5711 ;
  assign n17240 = ( n3833 & ~n17238 ) | ( n3833 & n17239 ) | ( ~n17238 & n17239 ) ;
  assign n17241 = ( n15856 & n17235 ) | ( n15856 & ~n17240 ) | ( n17235 & ~n17240 ) ;
  assign n17242 = ~n5860 & n10094 ;
  assign n17243 = n13117 & n17242 ;
  assign n17244 = n9637 ^ n2111 ^ n754 ;
  assign n17245 = ( n3605 & n17243 ) | ( n3605 & n17244 ) | ( n17243 & n17244 ) ;
  assign n17246 = n17245 ^ n2600 ^ n1230 ;
  assign n17247 = n17246 ^ n7900 ^ 1'b0 ;
  assign n17248 = n326 & n5665 ;
  assign n17249 = n4320 & n17248 ;
  assign n17250 = n17249 ^ n6207 ^ 1'b0 ;
  assign n17251 = n3503 | n3540 ;
  assign n17252 = n17251 ^ n8835 ^ 1'b0 ;
  assign n17253 = ~n6236 & n17252 ;
  assign n17254 = ~n2493 & n17253 ;
  assign n17255 = ( n4950 & n8260 ) | ( n4950 & n13164 ) | ( n8260 & n13164 ) ;
  assign n17256 = ( n6307 & n6728 ) | ( n6307 & ~n17255 ) | ( n6728 & ~n17255 ) ;
  assign n17257 = n7663 ^ n2195 ^ 1'b0 ;
  assign n17258 = n4744 & n17257 ;
  assign n17259 = n5641 & n8355 ;
  assign n17260 = ~n17258 & n17259 ;
  assign n17261 = n17260 ^ n4941 ^ 1'b0 ;
  assign n17264 = n14279 ^ n9170 ^ n266 ;
  assign n17265 = n17264 ^ n5486 ^ n4157 ;
  assign n17266 = n17265 ^ n9142 ^ n487 ;
  assign n17267 = x208 & n3984 ;
  assign n17268 = n17266 & n17267 ;
  assign n17262 = n9295 ^ n8200 ^ n5302 ;
  assign n17263 = n17262 ^ n13664 ^ 1'b0 ;
  assign n17269 = n17268 ^ n17263 ^ 1'b0 ;
  assign n17270 = n9084 ^ n5236 ^ x83 ;
  assign n17271 = n17270 ^ n12703 ^ n4153 ;
  assign n17272 = ( n4770 & ~n5189 ) | ( n4770 & n6214 ) | ( ~n5189 & n6214 ) ;
  assign n17273 = ( ~n879 & n1960 ) | ( ~n879 & n17272 ) | ( n1960 & n17272 ) ;
  assign n17274 = n4807 & ~n6452 ;
  assign n17275 = ( n7811 & n8949 ) | ( n7811 & ~n17274 ) | ( n8949 & ~n17274 ) ;
  assign n17276 = ( n10765 & n17273 ) | ( n10765 & n17275 ) | ( n17273 & n17275 ) ;
  assign n17277 = n5580 ^ n4129 ^ 1'b0 ;
  assign n17278 = n1610 & n17277 ;
  assign n17279 = n17278 ^ n3678 ^ n1718 ;
  assign n17280 = n10928 ^ n3545 ^ 1'b0 ;
  assign n17281 = ~n17279 & n17280 ;
  assign n17282 = n16487 ^ n13158 ^ 1'b0 ;
  assign n17283 = ( ~n8904 & n9994 ) | ( ~n8904 & n14723 ) | ( n9994 & n14723 ) ;
  assign n17284 = ( n5348 & n7070 ) | ( n5348 & n12176 ) | ( n7070 & n12176 ) ;
  assign n17285 = n10069 | n17284 ;
  assign n17286 = n13052 & n13678 ;
  assign n17287 = ~n10681 & n16050 ;
  assign n17288 = ~n4726 & n17287 ;
  assign n17289 = ( ~n17285 & n17286 ) | ( ~n17285 & n17288 ) | ( n17286 & n17288 ) ;
  assign n17290 = ( ~n14946 & n17283 ) | ( ~n14946 & n17289 ) | ( n17283 & n17289 ) ;
  assign n17291 = n9892 ^ n811 ^ 1'b0 ;
  assign n17292 = n14380 & n17291 ;
  assign n17293 = n9017 ^ n539 ^ 1'b0 ;
  assign n17294 = n17292 & n17293 ;
  assign n17295 = n3433 ^ n3049 ^ 1'b0 ;
  assign n17296 = ( n6948 & ~n17294 ) | ( n6948 & n17295 ) | ( ~n17294 & n17295 ) ;
  assign n17297 = n10974 ^ n10804 ^ n6463 ;
  assign n17298 = n17297 ^ n4370 ^ 1'b0 ;
  assign n17299 = n13052 & n17298 ;
  assign n17300 = n17299 ^ n12037 ^ n2858 ;
  assign n17301 = n438 & n9928 ;
  assign n17302 = n17301 ^ n16483 ^ 1'b0 ;
  assign n17303 = ~n924 & n15046 ;
  assign n17304 = n3555 & n17303 ;
  assign n17305 = n4802 & ~n12497 ;
  assign n17306 = n17305 ^ n1792 ^ 1'b0 ;
  assign n17307 = n17306 ^ n14387 ^ n5791 ;
  assign n17308 = ~n5840 & n9291 ;
  assign n17309 = ( ~n5990 & n17307 ) | ( ~n5990 & n17308 ) | ( n17307 & n17308 ) ;
  assign n17310 = ~n9280 & n17309 ;
  assign n17311 = n6314 ^ n5015 ^ n3826 ;
  assign n17312 = n17311 ^ n4902 ^ 1'b0 ;
  assign n17313 = n5517 ^ n4092 ^ n2083 ;
  assign n17314 = n17313 ^ n6967 ^ 1'b0 ;
  assign n17315 = x90 & ~n17314 ;
  assign n17316 = n16583 ^ n2362 ^ 1'b0 ;
  assign n17317 = ( ~n13354 & n17315 ) | ( ~n13354 & n17316 ) | ( n17315 & n17316 ) ;
  assign n17327 = n4571 ^ n2521 ^ 1'b0 ;
  assign n17318 = ( ~n3485 & n5099 ) | ( ~n3485 & n13123 ) | ( n5099 & n13123 ) ;
  assign n17322 = n10304 ^ n4171 ^ n2149 ;
  assign n17321 = n12675 ^ n3803 ^ n1358 ;
  assign n17323 = n17322 ^ n17321 ^ 1'b0 ;
  assign n17324 = n13195 | n17323 ;
  assign n17319 = n1014 | n5715 ;
  assign n17320 = n17319 ^ n8813 ^ 1'b0 ;
  assign n17325 = n17324 ^ n17320 ^ 1'b0 ;
  assign n17326 = n17318 | n17325 ;
  assign n17328 = n17327 ^ n17326 ^ n7238 ;
  assign n17329 = n2300 | n15029 ;
  assign n17330 = x248 | n17329 ;
  assign n17331 = ( n5564 & n12875 ) | ( n5564 & ~n13489 ) | ( n12875 & ~n13489 ) ;
  assign n17332 = ( n5543 & n17330 ) | ( n5543 & ~n17331 ) | ( n17330 & ~n17331 ) ;
  assign n17333 = n9455 ^ n8526 ^ n4204 ;
  assign n17334 = ( ~n7779 & n8880 ) | ( ~n7779 & n17333 ) | ( n8880 & n17333 ) ;
  assign n17340 = ( n3538 & n11737 ) | ( n3538 & ~n11866 ) | ( n11737 & ~n11866 ) ;
  assign n17335 = n3348 & ~n6635 ;
  assign n17336 = ~n2954 & n17335 ;
  assign n17337 = n17336 ^ n10280 ^ 1'b0 ;
  assign n17338 = n15785 | n17337 ;
  assign n17339 = n10538 | n17338 ;
  assign n17341 = n17340 ^ n17339 ^ 1'b0 ;
  assign n17344 = n6111 ^ n3428 ^ x221 ;
  assign n17345 = n11489 | n17344 ;
  assign n17346 = n1948 & ~n17345 ;
  assign n17342 = ~n6787 & n10468 ;
  assign n17343 = n17342 ^ n1078 ^ 1'b0 ;
  assign n17347 = n17346 ^ n17343 ^ 1'b0 ;
  assign n17348 = ( n399 & n4738 ) | ( n399 & n17056 ) | ( n4738 & n17056 ) ;
  assign n17350 = x100 & n2853 ;
  assign n17351 = n4333 & n17350 ;
  assign n17349 = n6785 & ~n14539 ;
  assign n17352 = n17351 ^ n17349 ^ 1'b0 ;
  assign n17353 = ~n14840 & n17352 ;
  assign n17354 = ~n483 & n17353 ;
  assign n17355 = n1506 | n17354 ;
  assign n17356 = n4763 & ~n17355 ;
  assign n17357 = n11301 | n17356 ;
  assign n17359 = n1192 & ~n10613 ;
  assign n17360 = n1124 & n17359 ;
  assign n17361 = n4644 | n17360 ;
  assign n17358 = ( ~n2374 & n7710 ) | ( ~n2374 & n16388 ) | ( n7710 & n16388 ) ;
  assign n17362 = n17361 ^ n17358 ^ x110 ;
  assign n17363 = n11632 ^ n5314 ^ n5298 ;
  assign n17364 = n539 | n8649 ;
  assign n17365 = n17363 & ~n17364 ;
  assign n17366 = ( ~n7314 & n7365 ) | ( ~n7314 & n7899 ) | ( n7365 & n7899 ) ;
  assign n17367 = n5328 ^ n1506 ^ 1'b0 ;
  assign n17368 = n2246 | n17367 ;
  assign n17369 = n3924 & n7736 ;
  assign n17370 = ( n1500 & n6997 ) | ( n1500 & ~n7125 ) | ( n6997 & ~n7125 ) ;
  assign n17371 = n628 & n9055 ;
  assign n17372 = ~n17370 & n17371 ;
  assign n17373 = n17369 & ~n17372 ;
  assign n17374 = n16019 & n17373 ;
  assign n17375 = ( n8447 & ~n17368 ) | ( n8447 & n17374 ) | ( ~n17368 & n17374 ) ;
  assign n17377 = ( ~n1375 & n6291 ) | ( ~n1375 & n9905 ) | ( n6291 & n9905 ) ;
  assign n17376 = ( n642 & n650 ) | ( n642 & ~n10370 ) | ( n650 & ~n10370 ) ;
  assign n17378 = n17377 ^ n17376 ^ n4765 ;
  assign n17379 = ( n279 & n6246 ) | ( n279 & ~n16422 ) | ( n6246 & ~n16422 ) ;
  assign n17380 = n15439 & n17379 ;
  assign n17381 = n589 | n5458 ;
  assign n17382 = ~n9785 & n11195 ;
  assign n17383 = n17381 & n17382 ;
  assign n17384 = n4696 & n5576 ;
  assign n17385 = n17384 ^ n3786 ^ 1'b0 ;
  assign n17386 = ( ~n1440 & n9180 ) | ( ~n1440 & n11084 ) | ( n9180 & n11084 ) ;
  assign n17387 = n17386 ^ n472 ^ 1'b0 ;
  assign n17388 = n17385 & ~n17387 ;
  assign n17389 = ( ~n5787 & n10483 ) | ( ~n5787 & n14164 ) | ( n10483 & n14164 ) ;
  assign n17390 = n17389 ^ n5702 ^ n4004 ;
  assign n17391 = n11635 ^ n3472 ^ n947 ;
  assign n17392 = n17391 ^ n5726 ^ n1262 ;
  assign n17396 = n9560 ^ n4332 ^ 1'b0 ;
  assign n17397 = n17396 ^ n7265 ^ 1'b0 ;
  assign n17393 = ( n3129 & n3588 ) | ( n3129 & ~n14295 ) | ( n3588 & ~n14295 ) ;
  assign n17394 = ~n980 & n10377 ;
  assign n17395 = ( n16049 & n17393 ) | ( n16049 & ~n17394 ) | ( n17393 & ~n17394 ) ;
  assign n17398 = n17397 ^ n17395 ^ 1'b0 ;
  assign n17399 = n16272 & ~n17398 ;
  assign n17400 = ( n803 & n7255 ) | ( n803 & ~n7485 ) | ( n7255 & ~n7485 ) ;
  assign n17401 = n6132 & ~n17400 ;
  assign n17405 = n10671 ^ n10359 ^ 1'b0 ;
  assign n17406 = n17405 ^ n8638 ^ 1'b0 ;
  assign n17402 = n1003 & ~n11203 ;
  assign n17403 = n17402 ^ n15799 ^ 1'b0 ;
  assign n17404 = n17403 ^ n9264 ^ n6983 ;
  assign n17407 = n17406 ^ n17404 ^ n2891 ;
  assign n17408 = n13822 ^ n8403 ^ 1'b0 ;
  assign n17409 = n8159 & ~n17408 ;
  assign n17411 = n10115 & n11010 ;
  assign n17412 = n17411 ^ x166 ^ 1'b0 ;
  assign n17413 = n17412 ^ n1699 ^ 1'b0 ;
  assign n17414 = ( n675 & n9506 ) | ( n675 & n16317 ) | ( n9506 & n16317 ) ;
  assign n17415 = ( n4499 & ~n7743 ) | ( n4499 & n14020 ) | ( ~n7743 & n14020 ) ;
  assign n17416 = ( n17413 & n17414 ) | ( n17413 & n17415 ) | ( n17414 & n17415 ) ;
  assign n17410 = n9629 ^ n3462 ^ 1'b0 ;
  assign n17417 = n17416 ^ n17410 ^ n901 ;
  assign n17418 = ( n2935 & n10840 ) | ( n2935 & ~n17379 ) | ( n10840 & ~n17379 ) ;
  assign n17419 = x108 & n15912 ;
  assign n17420 = ~n11868 & n17419 ;
  assign n17426 = n7766 ^ n6357 ^ n2915 ;
  assign n17427 = ( n1841 & n8313 ) | ( n1841 & n17426 ) | ( n8313 & n17426 ) ;
  assign n17421 = ( n2813 & n6727 ) | ( n2813 & ~n10769 ) | ( n6727 & ~n10769 ) ;
  assign n17422 = ( x59 & n7598 ) | ( x59 & ~n17421 ) | ( n7598 & ~n17421 ) ;
  assign n17423 = n17422 ^ n1671 ^ 1'b0 ;
  assign n17424 = n450 | n17423 ;
  assign n17425 = ( n7461 & n14978 ) | ( n7461 & ~n17424 ) | ( n14978 & ~n17424 ) ;
  assign n17428 = n17427 ^ n17425 ^ n3248 ;
  assign n17429 = n13860 | n15109 ;
  assign n17430 = n1906 | n7384 ;
  assign n17431 = n17430 ^ n12641 ^ n938 ;
  assign n17432 = ~n7549 & n17431 ;
  assign n17433 = ( n5121 & ~n5378 ) | ( n5121 & n17432 ) | ( ~n5378 & n17432 ) ;
  assign n17434 = ( n1609 & n3864 ) | ( n1609 & ~n13372 ) | ( n3864 & ~n13372 ) ;
  assign n17435 = n17434 ^ n15460 ^ n7642 ;
  assign n17436 = ( n2410 & n2583 ) | ( n2410 & n17435 ) | ( n2583 & n17435 ) ;
  assign n17437 = ~n17433 & n17436 ;
  assign n17438 = n3677 ^ n624 ^ 1'b0 ;
  assign n17439 = n7264 & n17438 ;
  assign n17440 = ~n4363 & n17439 ;
  assign n17441 = n3066 & ~n17440 ;
  assign n17442 = x152 & n6954 ;
  assign n17443 = ~n11271 & n17442 ;
  assign n17444 = ( n5354 & ~n11266 ) | ( n5354 & n17443 ) | ( ~n11266 & n17443 ) ;
  assign n17445 = n8985 ^ n7596 ^ n2865 ;
  assign n17446 = ( ~n8122 & n10537 ) | ( ~n8122 & n17445 ) | ( n10537 & n17445 ) ;
  assign n17447 = n17372 | n17446 ;
  assign n17448 = n17444 & ~n17447 ;
  assign n17449 = n17448 ^ n5515 ^ n3179 ;
  assign n17450 = x208 & ~n15593 ;
  assign n17451 = n3831 & n17450 ;
  assign n17452 = n17449 | n17451 ;
  assign n17456 = n7423 ^ n7253 ^ 1'b0 ;
  assign n17457 = n2915 & n17456 ;
  assign n17453 = ( ~n7139 & n7856 ) | ( ~n7139 & n10558 ) | ( n7856 & n10558 ) ;
  assign n17454 = n13557 & ~n17453 ;
  assign n17455 = n17454 ^ n8836 ^ 1'b0 ;
  assign n17458 = n17457 ^ n17455 ^ n2150 ;
  assign n17459 = n15781 ^ n6871 ^ n2748 ;
  assign n17460 = ~n9688 & n10278 ;
  assign n17461 = ( n4794 & n6678 ) | ( n4794 & n12912 ) | ( n6678 & n12912 ) ;
  assign n17462 = ( n8903 & n17460 ) | ( n8903 & ~n17461 ) | ( n17460 & ~n17461 ) ;
  assign n17463 = n17462 ^ n8636 ^ n2754 ;
  assign n17464 = ( n7994 & ~n14928 ) | ( n7994 & n17463 ) | ( ~n14928 & n17463 ) ;
  assign n17466 = n4638 ^ n3420 ^ 1'b0 ;
  assign n17465 = n12510 ^ n3453 ^ 1'b0 ;
  assign n17467 = n17466 ^ n17465 ^ n14565 ;
  assign n17468 = ( x64 & n2051 ) | ( x64 & n10281 ) | ( n2051 & n10281 ) ;
  assign n17469 = ( n2140 & n6250 ) | ( n2140 & n17468 ) | ( n6250 & n17468 ) ;
  assign n17470 = n17469 ^ n5310 ^ 1'b0 ;
  assign n17471 = n4488 & ~n17470 ;
  assign n17472 = ~n751 & n17471 ;
  assign n17473 = n2727 & n7300 ;
  assign n17474 = ~n17472 & n17473 ;
  assign n17481 = n2332 & n8693 ;
  assign n17482 = n17481 ^ n13692 ^ 1'b0 ;
  assign n17475 = ( x234 & ~n1587 ) | ( x234 & n3462 ) | ( ~n1587 & n3462 ) ;
  assign n17476 = n17475 ^ n5165 ^ n4645 ;
  assign n17477 = ( n3789 & n5128 ) | ( n3789 & n17476 ) | ( n5128 & n17476 ) ;
  assign n17478 = ~n2769 & n17477 ;
  assign n17479 = n4479 & n17478 ;
  assign n17480 = n17479 ^ n16546 ^ n13159 ;
  assign n17483 = n17482 ^ n17480 ^ n2064 ;
  assign n17484 = ( n2480 & ~n17474 ) | ( n2480 & n17483 ) | ( ~n17474 & n17483 ) ;
  assign n17485 = n5321 & ~n9126 ;
  assign n17486 = ~n6891 & n17485 ;
  assign n17487 = n893 | n2950 ;
  assign n17488 = n17487 ^ n6562 ^ 1'b0 ;
  assign n17489 = ( n4362 & n9918 ) | ( n4362 & ~n17488 ) | ( n9918 & ~n17488 ) ;
  assign n17490 = n17489 ^ n8937 ^ n3538 ;
  assign n17491 = ( ~n16710 & n17486 ) | ( ~n16710 & n17490 ) | ( n17486 & n17490 ) ;
  assign n17494 = ( n1748 & n4023 ) | ( n1748 & n5293 ) | ( n4023 & n5293 ) ;
  assign n17492 = n4319 & n5393 ;
  assign n17493 = n9535 & ~n17492 ;
  assign n17495 = n17494 ^ n17493 ^ 1'b0 ;
  assign n17496 = ( n2314 & ~n3705 ) | ( n2314 & n9092 ) | ( ~n3705 & n9092 ) ;
  assign n17497 = ~n5781 & n17496 ;
  assign n17498 = n17497 ^ n7698 ^ n2102 ;
  assign n17499 = n10936 | n14446 ;
  assign n17500 = n17498 | n17499 ;
  assign n17501 = ( n3516 & ~n6557 ) | ( n3516 & n17500 ) | ( ~n6557 & n17500 ) ;
  assign n17502 = ( n3169 & n3392 ) | ( n3169 & n4798 ) | ( n3392 & n4798 ) ;
  assign n17503 = n17502 ^ n12144 ^ n3081 ;
  assign n17504 = n10386 | n17503 ;
  assign n17505 = n2684 & n6981 ;
  assign n17506 = n11242 & ~n12014 ;
  assign n17507 = ~x94 & n17506 ;
  assign n17508 = n17507 ^ n2397 ^ 1'b0 ;
  assign n17509 = ~n10151 & n10875 ;
  assign n17510 = n17509 ^ n17174 ^ 1'b0 ;
  assign n17512 = n8239 ^ n3125 ^ 1'b0 ;
  assign n17513 = n2547 & ~n17512 ;
  assign n17514 = n17513 ^ n3293 ^ 1'b0 ;
  assign n17511 = n8722 ^ n4198 ^ n3598 ;
  assign n17515 = n17514 ^ n17511 ^ 1'b0 ;
  assign n17516 = n17515 ^ n11869 ^ n7268 ;
  assign n17517 = ( n17309 & n17510 ) | ( n17309 & ~n17516 ) | ( n17510 & ~n17516 ) ;
  assign n17519 = n2089 & ~n4491 ;
  assign n17520 = n17519 ^ n5272 ^ 1'b0 ;
  assign n17518 = ~n6889 & n14230 ;
  assign n17521 = n17520 ^ n17518 ^ 1'b0 ;
  assign n17523 = ( ~n5223 & n6548 ) | ( ~n5223 & n10490 ) | ( n6548 & n10490 ) ;
  assign n17522 = ~n13529 & n16474 ;
  assign n17524 = n17523 ^ n17522 ^ 1'b0 ;
  assign n17525 = n2474 ^ n872 ^ 1'b0 ;
  assign n17526 = n6396 & ~n17525 ;
  assign n17527 = n5882 & n17526 ;
  assign n17531 = n6010 ^ n5166 ^ 1'b0 ;
  assign n17532 = ~n9922 & n17531 ;
  assign n17528 = n1887 ^ x180 ^ x22 ;
  assign n17529 = n17528 ^ x192 ^ 1'b0 ;
  assign n17530 = n5659 | n17529 ;
  assign n17533 = n17532 ^ n17530 ^ n10693 ;
  assign n17534 = ( n1669 & ~n2367 ) | ( n1669 & n7657 ) | ( ~n2367 & n7657 ) ;
  assign n17535 = ~n399 & n17534 ;
  assign n17536 = ( n11073 & n15518 ) | ( n11073 & ~n17535 ) | ( n15518 & ~n17535 ) ;
  assign n17537 = n7014 & ~n11246 ;
  assign n17548 = ( n2192 & ~n7200 ) | ( n2192 & n8235 ) | ( ~n7200 & n8235 ) ;
  assign n17549 = n17548 ^ n4286 ^ 1'b0 ;
  assign n17538 = x5 & n3094 ;
  assign n17539 = ~n8903 & n17538 ;
  assign n17540 = n10412 ^ n8601 ^ n952 ;
  assign n17541 = ( ~n6726 & n6758 ) | ( ~n6726 & n17540 ) | ( n6758 & n17540 ) ;
  assign n17542 = ~n17539 & n17541 ;
  assign n17543 = n17542 ^ n456 ^ 1'b0 ;
  assign n17544 = ~n4484 & n5960 ;
  assign n17545 = ~n4681 & n6885 ;
  assign n17546 = ( ~n12362 & n17544 ) | ( ~n12362 & n17545 ) | ( n17544 & n17545 ) ;
  assign n17547 = ( ~n4319 & n17543 ) | ( ~n4319 & n17546 ) | ( n17543 & n17546 ) ;
  assign n17550 = n17549 ^ n17547 ^ n7595 ;
  assign n17551 = ( n267 & n7097 ) | ( n267 & ~n15510 ) | ( n7097 & ~n15510 ) ;
  assign n17552 = n2425 ^ x41 ^ 1'b0 ;
  assign n17553 = n5363 & n17552 ;
  assign n17554 = n17553 ^ n6300 ^ 1'b0 ;
  assign n17555 = n9635 ^ n6887 ^ 1'b0 ;
  assign n17556 = n17555 ^ n12086 ^ n3951 ;
  assign n17557 = ( ~n15776 & n17554 ) | ( ~n15776 & n17556 ) | ( n17554 & n17556 ) ;
  assign n17558 = ~n11796 & n17557 ;
  assign n17559 = n17558 ^ n6022 ^ 1'b0 ;
  assign n17560 = n13006 ^ n8117 ^ 1'b0 ;
  assign n17561 = x122 & ~n4707 ;
  assign n17562 = n17561 ^ n9593 ^ 1'b0 ;
  assign n17563 = ( ~n3921 & n13212 ) | ( ~n3921 & n17562 ) | ( n13212 & n17562 ) ;
  assign n17564 = n6601 ^ n1796 ^ 1'b0 ;
  assign n17565 = n17564 ^ n11538 ^ n3290 ;
  assign n17566 = n9390 | n12326 ;
  assign n17567 = n4827 & ~n17566 ;
  assign n17574 = n8027 & ~n8926 ;
  assign n17568 = n7072 | n12804 ;
  assign n17569 = n17568 ^ n2878 ^ 1'b0 ;
  assign n17570 = n992 & ~n17569 ;
  assign n17571 = n17570 ^ n5583 ^ n2184 ;
  assign n17572 = n17571 ^ x97 ^ 1'b0 ;
  assign n17573 = ~n1098 & n17572 ;
  assign n17575 = n17574 ^ n17573 ^ n12757 ;
  assign n17576 = n11967 ^ n10552 ^ x48 ;
  assign n17577 = n11984 ^ n550 ^ 1'b0 ;
  assign n17578 = ~n3254 & n17577 ;
  assign n17579 = ~n16317 & n17578 ;
  assign n17580 = ( n696 & n17576 ) | ( n696 & ~n17579 ) | ( n17576 & ~n17579 ) ;
  assign n17581 = n4593 & ~n5342 ;
  assign n17582 = n17581 ^ n912 ^ 1'b0 ;
  assign n17583 = ~n5722 & n17582 ;
  assign n17584 = n4673 & n17583 ;
  assign n17585 = ~n3999 & n10127 ;
  assign n17586 = n17585 ^ n3188 ^ 1'b0 ;
  assign n17587 = ~n17584 & n17586 ;
  assign n17588 = n4713 & ~n9799 ;
  assign n17589 = ( n4076 & n4412 ) | ( n4076 & n9909 ) | ( n4412 & n9909 ) ;
  assign n17590 = n470 & n2370 ;
  assign n17591 = ( n4939 & n14194 ) | ( n4939 & ~n17590 ) | ( n14194 & ~n17590 ) ;
  assign n17592 = x237 & n1863 ;
  assign n17593 = n17592 ^ n12338 ^ 1'b0 ;
  assign n17594 = ( ~n2875 & n7450 ) | ( ~n2875 & n17593 ) | ( n7450 & n17593 ) ;
  assign n17595 = n17594 ^ n13332 ^ n4834 ;
  assign n17596 = n11691 & ~n16376 ;
  assign n17597 = ~n17595 & n17596 ;
  assign n17598 = n1340 ^ n1294 ^ 1'b0 ;
  assign n17599 = n17598 ^ n5511 ^ n428 ;
  assign n17600 = n17599 ^ n10317 ^ n2898 ;
  assign n17601 = ~n1708 & n17600 ;
  assign n17602 = n15498 & n17601 ;
  assign n17603 = ( ~n5128 & n6807 ) | ( ~n5128 & n17151 ) | ( n6807 & n17151 ) ;
  assign n17604 = n6660 ^ n5172 ^ 1'b0 ;
  assign n17605 = n17604 ^ n10733 ^ 1'b0 ;
  assign n17606 = n7474 ^ n6664 ^ 1'b0 ;
  assign n17613 = n5839 & n8508 ;
  assign n17607 = ( n488 & ~n3956 ) | ( n488 & n9643 ) | ( ~n3956 & n9643 ) ;
  assign n17608 = n3846 ^ n2347 ^ 1'b0 ;
  assign n17609 = n17607 | n17608 ;
  assign n17610 = ( n1803 & n5076 ) | ( n1803 & ~n17609 ) | ( n5076 & ~n17609 ) ;
  assign n17611 = n17610 ^ n2045 ^ 1'b0 ;
  assign n17612 = n17611 ^ n10765 ^ 1'b0 ;
  assign n17614 = n17613 ^ n17612 ^ n546 ;
  assign n17615 = n9218 | n16236 ;
  assign n17616 = n11121 ^ n5171 ^ 1'b0 ;
  assign n17617 = ~n17615 & n17616 ;
  assign n17618 = n12143 ^ n6998 ^ 1'b0 ;
  assign n17619 = n17617 & ~n17618 ;
  assign n17620 = ( ~n1691 & n17614 ) | ( ~n1691 & n17619 ) | ( n17614 & n17619 ) ;
  assign n17622 = n11798 ^ n3647 ^ 1'b0 ;
  assign n17621 = n10380 ^ n9308 ^ n4874 ;
  assign n17623 = n17622 ^ n17621 ^ n13904 ;
  assign n17624 = n11887 ^ n5053 ^ 1'b0 ;
  assign n17625 = n14109 & n17624 ;
  assign n17626 = ( n5405 & n7446 ) | ( n5405 & ~n8616 ) | ( n7446 & ~n8616 ) ;
  assign n17627 = n15945 ^ x134 ^ 1'b0 ;
  assign n17628 = n17627 ^ n12080 ^ 1'b0 ;
  assign n17629 = n15794 & n17628 ;
  assign n17630 = n17626 & ~n17629 ;
  assign n17631 = n9938 & ~n11149 ;
  assign n17632 = n17631 ^ n4153 ^ 1'b0 ;
  assign n17633 = ( n1109 & ~n10577 ) | ( n1109 & n17632 ) | ( ~n10577 & n17632 ) ;
  assign n17634 = ~n1010 & n5281 ;
  assign n17635 = n17634 ^ n7124 ^ 1'b0 ;
  assign n17637 = n3851 ^ n3375 ^ x230 ;
  assign n17636 = n5733 | n5800 ;
  assign n17638 = n17637 ^ n17636 ^ n2748 ;
  assign n17639 = n517 & n17638 ;
  assign n17640 = ( n2937 & ~n6206 ) | ( n2937 & n17639 ) | ( ~n6206 & n17639 ) ;
  assign n17641 = n17640 ^ n9357 ^ 1'b0 ;
  assign n17642 = n17635 & n17641 ;
  assign n17643 = n17642 ^ n12339 ^ n5092 ;
  assign n17644 = n17412 ^ n5373 ^ n4674 ;
  assign n17645 = ~n2791 & n17644 ;
  assign n17646 = ~n3592 & n17645 ;
  assign n17647 = ( x144 & n12763 ) | ( x144 & ~n15071 ) | ( n12763 & ~n15071 ) ;
  assign n17648 = n17026 ^ n12447 ^ 1'b0 ;
  assign n17649 = n13176 ^ x81 ^ 1'b0 ;
  assign n17650 = n17590 ^ n12249 ^ 1'b0 ;
  assign n17651 = n17650 ^ n11891 ^ n5539 ;
  assign n17652 = n8863 ^ n792 ^ 1'b0 ;
  assign n17653 = ~n10843 & n17652 ;
  assign n17654 = n17653 ^ n14797 ^ n7795 ;
  assign n17655 = n5924 & n6500 ;
  assign n17656 = ~n5924 & n17655 ;
  assign n17657 = ( n4405 & n5702 ) | ( n4405 & n5891 ) | ( n5702 & n5891 ) ;
  assign n17658 = n6367 & n8340 ;
  assign n17659 = n17657 & ~n17658 ;
  assign n17660 = n17656 & n17659 ;
  assign n17661 = n4812 ^ n2628 ^ 1'b0 ;
  assign n17662 = n672 | n17661 ;
  assign n17663 = n12595 | n17662 ;
  assign n17664 = ( n6188 & n15390 ) | ( n6188 & ~n17663 ) | ( n15390 & ~n17663 ) ;
  assign n17665 = n14645 ^ n7520 ^ 1'b0 ;
  assign n17666 = ~n9478 & n17665 ;
  assign n17667 = n7117 & n17666 ;
  assign n17668 = n10029 ^ n5232 ^ n1343 ;
  assign n17669 = ( n6531 & n10467 ) | ( n6531 & n17668 ) | ( n10467 & n17668 ) ;
  assign n17670 = ( n1544 & n1599 ) | ( n1544 & n6076 ) | ( n1599 & n6076 ) ;
  assign n17671 = ( n5006 & n13122 ) | ( n5006 & ~n17670 ) | ( n13122 & ~n17670 ) ;
  assign n17672 = ( ~n2364 & n17669 ) | ( ~n2364 & n17671 ) | ( n17669 & n17671 ) ;
  assign n17674 = n17082 ^ n555 ^ 1'b0 ;
  assign n17675 = n3891 | n17674 ;
  assign n17673 = ( n8545 & n14697 ) | ( n8545 & ~n15491 ) | ( n14697 & ~n15491 ) ;
  assign n17676 = n17675 ^ n17673 ^ n5251 ;
  assign n17677 = ( ~n8215 & n10175 ) | ( ~n8215 & n14181 ) | ( n10175 & n14181 ) ;
  assign n17680 = n4815 ^ n2498 ^ 1'b0 ;
  assign n17678 = n10611 ^ x36 ^ 1'b0 ;
  assign n17679 = ~n7596 & n17678 ;
  assign n17681 = n17680 ^ n17679 ^ 1'b0 ;
  assign n17682 = n4266 & n17681 ;
  assign n17683 = n4866 & n17682 ;
  assign n17684 = n7027 | n11057 ;
  assign n17685 = n16164 ^ n11460 ^ 1'b0 ;
  assign n17686 = n13689 | n14186 ;
  assign n17687 = n17686 ^ n13926 ^ 1'b0 ;
  assign n17688 = n14614 & ~n17687 ;
  assign n17689 = ~n10333 & n17688 ;
  assign n17690 = n13803 ^ n3130 ^ 1'b0 ;
  assign n17691 = n1815 | n2365 ;
  assign n17693 = n3381 & ~n11679 ;
  assign n17692 = ( ~n1929 & n4139 ) | ( ~n1929 & n16762 ) | ( n4139 & n16762 ) ;
  assign n17694 = n17693 ^ n17692 ^ 1'b0 ;
  assign n17696 = n13728 ^ n1430 ^ 1'b0 ;
  assign n17697 = n14787 & ~n17696 ;
  assign n17698 = n7900 & n17697 ;
  assign n17699 = ( n2355 & n7601 ) | ( n2355 & ~n17698 ) | ( n7601 & ~n17698 ) ;
  assign n17695 = ( ~n2904 & n3582 ) | ( ~n2904 & n4873 ) | ( n3582 & n4873 ) ;
  assign n17700 = n17699 ^ n17695 ^ n4664 ;
  assign n17701 = n11350 ^ n1003 ^ 1'b0 ;
  assign n17702 = n17700 & ~n17701 ;
  assign n17703 = n459 & ~n15657 ;
  assign n17704 = n17703 ^ n12339 ^ 1'b0 ;
  assign n17705 = n5566 & ~n12633 ;
  assign n17706 = n17705 ^ n7753 ^ 1'b0 ;
  assign n17707 = ( n5806 & n12544 ) | ( n5806 & n17706 ) | ( n12544 & n17706 ) ;
  assign n17708 = ~n6887 & n17707 ;
  assign n17710 = ( n838 & n2055 ) | ( n838 & n9094 ) | ( n2055 & n9094 ) ;
  assign n17709 = n13041 | n14716 ;
  assign n17711 = n17710 ^ n17709 ^ 1'b0 ;
  assign n17712 = ~n5121 & n8635 ;
  assign n17713 = ~n8184 & n9193 ;
  assign n17714 = n17388 & ~n17713 ;
  assign n17715 = n17712 & n17714 ;
  assign n17716 = ~n5097 & n13211 ;
  assign n17717 = n6083 & ~n6101 ;
  assign n17718 = ( n5875 & n6934 ) | ( n5875 & n17308 ) | ( n6934 & n17308 ) ;
  assign n17719 = ~n4263 & n10834 ;
  assign n17720 = n17719 ^ n9670 ^ 1'b0 ;
  assign n17721 = n17720 ^ n6275 ^ n2766 ;
  assign n17727 = n3625 ^ n542 ^ 1'b0 ;
  assign n17723 = n8026 ^ n1609 ^ 1'b0 ;
  assign n17724 = n8157 & n17723 ;
  assign n17722 = n5367 & n15673 ;
  assign n17725 = n17724 ^ n17722 ^ 1'b0 ;
  assign n17726 = n13008 | n17725 ;
  assign n17728 = n17727 ^ n17726 ^ 1'b0 ;
  assign n17729 = n17728 ^ n13035 ^ n7370 ;
  assign n17730 = ~n466 & n6539 ;
  assign n17731 = ~n3350 & n17730 ;
  assign n17732 = n4201 | n7582 ;
  assign n17733 = ( n1831 & ~n9814 ) | ( n1831 & n17732 ) | ( ~n9814 & n17732 ) ;
  assign n17734 = ( ~n9611 & n17731 ) | ( ~n9611 & n17733 ) | ( n17731 & n17733 ) ;
  assign n17735 = n17500 ^ n11884 ^ n10376 ;
  assign n17736 = n16047 | n17735 ;
  assign n17737 = n6923 | n10116 ;
  assign n17738 = n5980 & n9534 ;
  assign n17739 = ~n8136 & n17738 ;
  assign n17740 = n17739 ^ n8619 ^ n1428 ;
  assign n17741 = ( n5918 & n17737 ) | ( n5918 & n17740 ) | ( n17737 & n17740 ) ;
  assign n17742 = n3493 & n11329 ;
  assign n17743 = ~n1351 & n17742 ;
  assign n17744 = n13648 & ~n17743 ;
  assign n17745 = n17744 ^ n12471 ^ 1'b0 ;
  assign n17746 = x198 & n10548 ;
  assign n17747 = ~n6185 & n17746 ;
  assign n17748 = ( ~n755 & n1046 ) | ( ~n755 & n4009 ) | ( n1046 & n4009 ) ;
  assign n17752 = n8558 ^ n7277 ^ n4198 ;
  assign n17749 = n6044 ^ n425 ^ 1'b0 ;
  assign n17750 = n3397 & n17749 ;
  assign n17751 = ~n10306 & n17750 ;
  assign n17753 = n17752 ^ n17751 ^ 1'b0 ;
  assign n17754 = ( n3380 & ~n17748 ) | ( n3380 & n17753 ) | ( ~n17748 & n17753 ) ;
  assign n17755 = n329 ^ x22 ^ 1'b0 ;
  assign n17756 = n4339 ^ n1603 ^ 1'b0 ;
  assign n17757 = n12199 & n17756 ;
  assign n17758 = ( ~n1358 & n17755 ) | ( ~n1358 & n17757 ) | ( n17755 & n17757 ) ;
  assign n17759 = n15359 ^ n12398 ^ n8544 ;
  assign n17760 = n9461 | n9620 ;
  assign n17761 = n12751 | n17760 ;
  assign n17762 = ( n4926 & n15259 ) | ( n4926 & n17761 ) | ( n15259 & n17761 ) ;
  assign n17763 = n7800 & n17762 ;
  assign n17764 = n6755 & n17763 ;
  assign n17765 = ~n1260 & n7799 ;
  assign n17766 = ~n6574 & n17765 ;
  assign n17768 = n10424 ^ n4044 ^ 1'b0 ;
  assign n17769 = ~n14516 & n17768 ;
  assign n17767 = ( n933 & n2417 ) | ( n933 & n14648 ) | ( n2417 & n14648 ) ;
  assign n17770 = n17769 ^ n17767 ^ n2610 ;
  assign n17771 = n17770 ^ n12887 ^ 1'b0 ;
  assign n17772 = ~n17021 & n17771 ;
  assign n17773 = ( n3561 & n10799 ) | ( n3561 & ~n17379 ) | ( n10799 & ~n17379 ) ;
  assign n17774 = ~n5753 & n17773 ;
  assign n17775 = n1104 & n2404 ;
  assign n17776 = ( n3972 & n11529 ) | ( n3972 & ~n17775 ) | ( n11529 & ~n17775 ) ;
  assign n17777 = ( n602 & n6168 ) | ( n602 & n14525 ) | ( n6168 & n14525 ) ;
  assign n17778 = n16530 ^ n2183 ^ 1'b0 ;
  assign n17779 = ~n6657 & n17778 ;
  assign n17780 = n17779 ^ n10373 ^ n1228 ;
  assign n17783 = n11800 ^ n10149 ^ n7641 ;
  assign n17784 = ( n14332 & ~n14811 ) | ( n14332 & n17783 ) | ( ~n14811 & n17783 ) ;
  assign n17781 = ( ~n1815 & n2878 ) | ( ~n1815 & n4334 ) | ( n2878 & n4334 ) ;
  assign n17782 = n13142 | n17781 ;
  assign n17785 = n17784 ^ n17782 ^ 1'b0 ;
  assign n17790 = ( ~n4434 & n10825 ) | ( ~n4434 & n13724 ) | ( n10825 & n13724 ) ;
  assign n17786 = n5784 & ~n7162 ;
  assign n17787 = n2923 & n17786 ;
  assign n17788 = ( n2092 & n13090 ) | ( n2092 & n17787 ) | ( n13090 & n17787 ) ;
  assign n17789 = ( n4343 & ~n8515 ) | ( n4343 & n17788 ) | ( ~n8515 & n17788 ) ;
  assign n17791 = n17790 ^ n17789 ^ n17132 ;
  assign n17792 = n17791 ^ n7004 ^ 1'b0 ;
  assign n17793 = n8402 ^ n2799 ^ 1'b0 ;
  assign n17794 = n8743 & n17793 ;
  assign n17795 = n15596 ^ n5032 ^ n2495 ;
  assign n17796 = n703 | n17795 ;
  assign n17797 = n10629 & ~n17796 ;
  assign n17798 = n9505 & ~n17797 ;
  assign n17799 = n7085 & n7894 ;
  assign n17800 = n3388 & ~n17799 ;
  assign n17801 = n16217 | n17800 ;
  assign n17802 = n17798 | n17801 ;
  assign n17803 = n7640 ^ n1691 ^ 1'b0 ;
  assign n17804 = n17803 ^ n2407 ^ 1'b0 ;
  assign n17805 = n5831 | n17804 ;
  assign n17806 = n6240 | n17805 ;
  assign n17807 = n10203 ^ n459 ^ 1'b0 ;
  assign n17808 = ( n959 & n7660 ) | ( n959 & ~n17807 ) | ( n7660 & ~n17807 ) ;
  assign n17809 = n17808 ^ n9887 ^ 1'b0 ;
  assign n17810 = n5963 ^ n2913 ^ 1'b0 ;
  assign n17811 = n2140 & n16267 ;
  assign n17812 = n7216 ^ n4747 ^ 1'b0 ;
  assign n17813 = n12097 ^ n9087 ^ 1'b0 ;
  assign n17814 = n14337 & n17813 ;
  assign n17815 = ( n6918 & ~n17812 ) | ( n6918 & n17814 ) | ( ~n17812 & n17814 ) ;
  assign n17816 = ( n14798 & n17811 ) | ( n14798 & ~n17815 ) | ( n17811 & ~n17815 ) ;
  assign n17817 = ( n5228 & ~n6981 ) | ( n5228 & n17816 ) | ( ~n6981 & n17816 ) ;
  assign n17818 = ( n4128 & n4995 ) | ( n4128 & ~n17817 ) | ( n4995 & ~n17817 ) ;
  assign n17819 = n6326 ^ n5092 ^ 1'b0 ;
  assign n17820 = ~n4927 & n17819 ;
  assign n17821 = n6930 & n17820 ;
  assign n17822 = n15906 & ~n17821 ;
  assign n17823 = ( n7490 & n17528 ) | ( n7490 & ~n17822 ) | ( n17528 & ~n17822 ) ;
  assign n17824 = ( ~n286 & n2169 ) | ( ~n286 & n3213 ) | ( n2169 & n3213 ) ;
  assign n17825 = n12249 ^ n2620 ^ 1'b0 ;
  assign n17826 = n17824 & n17825 ;
  assign n17827 = ( ~n5269 & n13290 ) | ( ~n5269 & n17826 ) | ( n13290 & n17826 ) ;
  assign n17830 = ~n2778 & n8813 ;
  assign n17831 = n4134 & n17830 ;
  assign n17832 = n7901 & ~n17831 ;
  assign n17833 = n4227 & n17832 ;
  assign n17829 = n12050 & n17017 ;
  assign n17834 = n17833 ^ n17829 ^ n4017 ;
  assign n17828 = n3407 & n16504 ;
  assign n17835 = n17834 ^ n17828 ^ 1'b0 ;
  assign n17836 = n9879 ^ n3212 ^ 1'b0 ;
  assign n17837 = n9925 & ~n17836 ;
  assign n17838 = n17837 ^ n15383 ^ 1'b0 ;
  assign n17839 = n17625 & n17838 ;
  assign n17840 = n13543 ^ n3943 ^ x3 ;
  assign n17841 = n17840 ^ n17067 ^ 1'b0 ;
  assign n17842 = n1763 | n9279 ;
  assign n17843 = n17842 ^ n7618 ^ 1'b0 ;
  assign n17844 = ( ~n9063 & n11887 ) | ( ~n9063 & n17843 ) | ( n11887 & n17843 ) ;
  assign n17845 = n9218 | n17844 ;
  assign n17846 = n7198 ^ n4434 ^ 1'b0 ;
  assign n17847 = ~n3354 & n17539 ;
  assign n17848 = n1446 | n17847 ;
  assign n17849 = n2964 & ~n17848 ;
  assign n17851 = ( n1317 & ~n6510 ) | ( n1317 & n11704 ) | ( ~n6510 & n11704 ) ;
  assign n17852 = ~n7258 & n17851 ;
  assign n17850 = n8496 & n10678 ;
  assign n17853 = n17852 ^ n17850 ^ n16054 ;
  assign n17854 = ( n3259 & n7468 ) | ( n3259 & n17853 ) | ( n7468 & n17853 ) ;
  assign n17855 = n14292 ^ n1918 ^ n314 ;
  assign n17856 = n7843 ^ n7137 ^ 1'b0 ;
  assign n17857 = ~n17855 & n17856 ;
  assign n17858 = ( n3906 & ~n7144 ) | ( n3906 & n15260 ) | ( ~n7144 & n15260 ) ;
  assign n17859 = n14917 ^ n9623 ^ n4958 ;
  assign n17860 = n6981 & n8168 ;
  assign n17861 = ~n923 & n17860 ;
  assign n17862 = n17859 & n17861 ;
  assign n17863 = n3065 & ~n17862 ;
  assign n17864 = ( n5669 & ~n17858 ) | ( n5669 & n17863 ) | ( ~n17858 & n17863 ) ;
  assign n17865 = ( n9036 & n10259 ) | ( n9036 & n17622 ) | ( n10259 & n17622 ) ;
  assign n17866 = n1073 | n7009 ;
  assign n17867 = n16548 ^ n6976 ^ 1'b0 ;
  assign n17868 = ( ~n8388 & n17866 ) | ( ~n8388 & n17867 ) | ( n17866 & n17867 ) ;
  assign n17869 = n9013 | n9961 ;
  assign n17870 = ( n5478 & n11298 ) | ( n5478 & ~n15458 ) | ( n11298 & ~n15458 ) ;
  assign n17871 = n17870 ^ n5938 ^ n628 ;
  assign n17872 = n3753 & n6042 ;
  assign n17873 = n9875 | n17872 ;
  assign n17874 = n4512 ^ n2942 ^ 1'b0 ;
  assign n17875 = n2472 & n17874 ;
  assign n17876 = n431 | n7747 ;
  assign n17877 = n14603 | n17876 ;
  assign n17878 = x2 & ~n1776 ;
  assign n17879 = n6509 & n17878 ;
  assign n17880 = n17879 ^ n10449 ^ n4853 ;
  assign n17881 = n17880 ^ n3290 ^ 1'b0 ;
  assign n17882 = n16046 ^ n10163 ^ n504 ;
  assign n17883 = n14651 & ~n17882 ;
  assign n17884 = n308 & n17883 ;
  assign n17885 = x196 & ~n17884 ;
  assign n17886 = ~n17881 & n17885 ;
  assign n17891 = n17075 ^ n8849 ^ n7957 ;
  assign n17892 = x72 & ~n1083 ;
  assign n17893 = n17891 & n17892 ;
  assign n17888 = n4275 ^ n3870 ^ n3738 ;
  assign n17887 = n813 & ~n8779 ;
  assign n17889 = n17888 ^ n17887 ^ 1'b0 ;
  assign n17890 = n10887 | n17889 ;
  assign n17894 = n17893 ^ n17890 ^ 1'b0 ;
  assign n17895 = ~n6540 & n6915 ;
  assign n17896 = n17895 ^ n16146 ^ n8524 ;
  assign n17897 = n15562 ^ n14085 ^ 1'b0 ;
  assign n17898 = n13483 & n17897 ;
  assign n17899 = n3751 & ~n13622 ;
  assign n17900 = n17899 ^ n3948 ^ 1'b0 ;
  assign n17901 = ( ~n9671 & n17898 ) | ( ~n9671 & n17900 ) | ( n17898 & n17900 ) ;
  assign n17902 = n5276 & n9185 ;
  assign n17903 = n17902 ^ n12202 ^ 1'b0 ;
  assign n17904 = n3119 | n8270 ;
  assign n17905 = n17904 ^ n7133 ^ 1'b0 ;
  assign n17906 = n17905 ^ n5231 ^ n2209 ;
  assign n17909 = ( n679 & n2066 ) | ( n679 & ~n2343 ) | ( n2066 & ~n2343 ) ;
  assign n17907 = ~n5111 & n5267 ;
  assign n17908 = n2256 & n17907 ;
  assign n17910 = n17909 ^ n17908 ^ n2474 ;
  assign n17911 = n14324 ^ n6903 ^ 1'b0 ;
  assign n17912 = ~n17910 & n17911 ;
  assign n17913 = ~n17906 & n17912 ;
  assign n17914 = n17913 ^ n11139 ^ 1'b0 ;
  assign n17915 = n10222 & ~n15334 ;
  assign n17916 = n17915 ^ n17135 ^ 1'b0 ;
  assign n17917 = ( n13161 & n17914 ) | ( n13161 & n17916 ) | ( n17914 & n17916 ) ;
  assign n17918 = n5958 ^ n5461 ^ 1'b0 ;
  assign n17919 = n1492 | n17918 ;
  assign n17920 = n9017 & ~n17919 ;
  assign n17921 = n13011 ^ n5223 ^ 1'b0 ;
  assign n17922 = ~n13261 & n17921 ;
  assign n17923 = n9220 ^ n4517 ^ 1'b0 ;
  assign n17924 = n1187 | n17923 ;
  assign n17925 = n4831 | n17924 ;
  assign n17926 = n4041 & ~n17925 ;
  assign n17927 = n17926 ^ n3156 ^ n1047 ;
  assign n17928 = ( n1879 & n2869 ) | ( n1879 & ~n17927 ) | ( n2869 & ~n17927 ) ;
  assign n17929 = n17922 & n17928 ;
  assign n17930 = n10473 ^ n5611 ^ n1614 ;
  assign n17931 = n3213 & ~n7698 ;
  assign n17932 = n17931 ^ n12441 ^ 1'b0 ;
  assign n17933 = n17932 ^ n13390 ^ 1'b0 ;
  assign n17934 = ( n7914 & n8349 ) | ( n7914 & ~n13175 ) | ( n8349 & ~n13175 ) ;
  assign n17935 = ( n5521 & ~n16266 ) | ( n5521 & n17343 ) | ( ~n16266 & n17343 ) ;
  assign n17936 = n287 | n4753 ;
  assign n17937 = n16811 ^ n2165 ^ n445 ;
  assign n17938 = n2039 | n2424 ;
  assign n17939 = n843 | n17938 ;
  assign n17940 = n17939 ^ n17264 ^ n2954 ;
  assign n17941 = ( ~n14387 & n17937 ) | ( ~n14387 & n17940 ) | ( n17937 & n17940 ) ;
  assign n17942 = ( n8049 & ~n17936 ) | ( n8049 & n17941 ) | ( ~n17936 & n17941 ) ;
  assign n17952 = ( n2985 & ~n8234 ) | ( n2985 & n14571 ) | ( ~n8234 & n14571 ) ;
  assign n17949 = n7988 ^ n7389 ^ n717 ;
  assign n17950 = n17949 ^ n6329 ^ 1'b0 ;
  assign n17943 = n16393 ^ n6689 ^ 1'b0 ;
  assign n17944 = n17943 ^ n13563 ^ n10363 ;
  assign n17945 = ~n286 & n1122 ;
  assign n17946 = n17945 ^ x136 ^ 1'b0 ;
  assign n17947 = n17946 ^ n15445 ^ 1'b0 ;
  assign n17948 = ~n17944 & n17947 ;
  assign n17951 = n17950 ^ n17948 ^ 1'b0 ;
  assign n17953 = n17952 ^ n17951 ^ 1'b0 ;
  assign n17958 = n5101 | n17787 ;
  assign n17959 = n3789 & ~n17958 ;
  assign n17954 = n14818 ^ n11430 ^ 1'b0 ;
  assign n17955 = n15986 ^ n10104 ^ n4619 ;
  assign n17956 = n17954 & ~n17955 ;
  assign n17957 = n17956 ^ n9128 ^ 1'b0 ;
  assign n17960 = n17959 ^ n17957 ^ n8983 ;
  assign n17961 = n10507 | n17960 ;
  assign n17962 = n1064 & n14962 ;
  assign n17963 = n17962 ^ n12602 ^ 1'b0 ;
  assign n17964 = ( ~n13722 & n15079 ) | ( ~n13722 & n17963 ) | ( n15079 & n17963 ) ;
  assign n17969 = n2715 | n12654 ;
  assign n17965 = ~n4152 & n5616 ;
  assign n17966 = ~n2676 & n17965 ;
  assign n17967 = n6486 & ~n8644 ;
  assign n17968 = n17966 | n17967 ;
  assign n17970 = n17969 ^ n17968 ^ n2632 ;
  assign n17980 = ~n7754 & n12835 ;
  assign n17979 = ( x95 & ~n4687 ) | ( x95 & n6615 ) | ( ~n4687 & n6615 ) ;
  assign n17971 = n16060 ^ n5063 ^ n3573 ;
  assign n17972 = ~n4868 & n5764 ;
  assign n17973 = ~n17971 & n17972 ;
  assign n17974 = ( n610 & ~n1487 ) | ( n610 & n9238 ) | ( ~n1487 & n9238 ) ;
  assign n17975 = n17974 ^ n1768 ^ n1574 ;
  assign n17976 = ~n17973 & n17975 ;
  assign n17977 = ~n3151 & n3875 ;
  assign n17978 = ~n17976 & n17977 ;
  assign n17981 = n17980 ^ n17979 ^ n17978 ;
  assign n17982 = ~n2810 & n3295 ;
  assign n17983 = n17982 ^ n7851 ^ n1813 ;
  assign n17984 = ( n5095 & ~n7973 ) | ( n5095 & n17983 ) | ( ~n7973 & n17983 ) ;
  assign n17985 = ( n1138 & n3412 ) | ( n1138 & ~n8320 ) | ( n3412 & ~n8320 ) ;
  assign n17986 = n2357 | n17985 ;
  assign n17987 = n17986 ^ n6857 ^ 1'b0 ;
  assign n17988 = n17987 ^ n16419 ^ 1'b0 ;
  assign n17989 = n15474 & n17988 ;
  assign n17990 = n7504 & ~n10334 ;
  assign n17991 = n12288 ^ n5025 ^ 1'b0 ;
  assign n17992 = ~n17990 & n17991 ;
  assign n17993 = x227 & n10243 ;
  assign n17994 = ~n2162 & n17993 ;
  assign n17995 = n17994 ^ n6711 ^ 1'b0 ;
  assign n17996 = n15016 | n15929 ;
  assign n17997 = n13780 & ~n17996 ;
  assign n17998 = n9622 ^ n5923 ^ n1910 ;
  assign n17999 = ~n14006 & n17998 ;
  assign n18000 = n17999 ^ n3257 ^ 1'b0 ;
  assign n18001 = n18000 ^ n7677 ^ 1'b0 ;
  assign n18002 = n18001 ^ n12766 ^ n4709 ;
  assign n18015 = n6430 | n12974 ;
  assign n18011 = ~n876 & n3571 ;
  assign n18012 = n1129 | n18011 ;
  assign n18013 = n18012 ^ n991 ^ 1'b0 ;
  assign n18008 = n17696 ^ n13875 ^ n3545 ;
  assign n18009 = n18008 ^ n13618 ^ 1'b0 ;
  assign n18010 = n9358 & ~n18009 ;
  assign n18014 = n18013 ^ n18010 ^ 1'b0 ;
  assign n18003 = n1864 & ~n16935 ;
  assign n18004 = n4371 & n18003 ;
  assign n18005 = n10124 ^ n4592 ^ 1'b0 ;
  assign n18006 = n7085 & ~n18005 ;
  assign n18007 = ~n18004 & n18006 ;
  assign n18016 = n18015 ^ n18014 ^ n18007 ;
  assign n18017 = x120 & ~n16752 ;
  assign n18018 = n18017 ^ n13922 ^ 1'b0 ;
  assign n18019 = ~n10832 & n13630 ;
  assign n18020 = n18019 ^ n1373 ^ 1'b0 ;
  assign n18021 = ~n18018 & n18020 ;
  assign n18022 = n18021 ^ n8927 ^ 1'b0 ;
  assign n18023 = n7811 & ~n18022 ;
  assign n18024 = n16868 & n18023 ;
  assign n18025 = n11190 ^ n9511 ^ n4345 ;
  assign n18026 = n8782 ^ n3143 ^ 1'b0 ;
  assign n18027 = n18025 | n18026 ;
  assign n18028 = n12919 ^ n10012 ^ 1'b0 ;
  assign n18031 = ( n2620 & n3684 ) | ( n2620 & n8667 ) | ( n3684 & n8667 ) ;
  assign n18029 = n8706 & ~n11158 ;
  assign n18030 = n18029 ^ n12692 ^ 1'b0 ;
  assign n18032 = n18031 ^ n18030 ^ n10669 ;
  assign n18033 = n15035 ^ n12199 ^ n6267 ;
  assign n18034 = ( n10054 & ~n12489 ) | ( n10054 & n18033 ) | ( ~n12489 & n18033 ) ;
  assign n18035 = n13042 ^ n7905 ^ n4290 ;
  assign n18036 = ( n5814 & n12679 ) | ( n5814 & n18035 ) | ( n12679 & n18035 ) ;
  assign n18038 = n6005 & ~n6630 ;
  assign n18039 = n3040 & n18038 ;
  assign n18040 = ( ~n589 & n7475 ) | ( ~n589 & n18039 ) | ( n7475 & n18039 ) ;
  assign n18037 = n16151 ^ n3896 ^ n3224 ;
  assign n18041 = n18040 ^ n18037 ^ n11727 ;
  assign n18042 = n18041 ^ n384 ^ 1'b0 ;
  assign n18043 = n3290 | n18042 ;
  assign n18044 = n18043 ^ n10732 ^ 1'b0 ;
  assign n18045 = n18036 | n18044 ;
  assign n18046 = n1138 & ~n3309 ;
  assign n18047 = n18046 ^ n2288 ^ 1'b0 ;
  assign n18048 = n18047 ^ n8877 ^ n1184 ;
  assign n18049 = n16131 ^ n11715 ^ n1960 ;
  assign n18050 = ~n5241 & n15216 ;
  assign n18051 = n8764 & n18050 ;
  assign n18052 = n5617 & ~n16428 ;
  assign n18053 = n9122 & n18052 ;
  assign n18054 = n17154 & n18053 ;
  assign n18055 = n3750 ^ n1436 ^ 1'b0 ;
  assign n18056 = ~n427 & n18055 ;
  assign n18057 = n17555 ^ n14883 ^ 1'b0 ;
  assign n18058 = ( n1734 & n6404 ) | ( n1734 & ~n18057 ) | ( n6404 & ~n18057 ) ;
  assign n18059 = n18058 ^ n9025 ^ 1'b0 ;
  assign n18060 = n18056 & ~n18059 ;
  assign n18061 = n10008 ^ n3467 ^ 1'b0 ;
  assign n18062 = n18061 ^ n10068 ^ 1'b0 ;
  assign n18063 = n18062 ^ n15513 ^ n8527 ;
  assign n18064 = n11680 ^ n4782 ^ 1'b0 ;
  assign n18065 = n14503 | n16109 ;
  assign n18066 = n18065 ^ n7934 ^ 1'b0 ;
  assign n18067 = n18066 ^ n5882 ^ 1'b0 ;
  assign n18068 = n18064 | n18067 ;
  assign n18072 = n6981 ^ n3813 ^ n306 ;
  assign n18071 = n7097 ^ n1578 ^ n280 ;
  assign n18073 = n18072 ^ n18071 ^ n8217 ;
  assign n18074 = ( n2702 & n12770 ) | ( n2702 & n18073 ) | ( n12770 & n18073 ) ;
  assign n18075 = n18074 ^ n6379 ^ n4917 ;
  assign n18076 = n7543 & n18075 ;
  assign n18077 = ~n17949 & n18076 ;
  assign n18069 = n8699 ^ n6904 ^ n5604 ;
  assign n18070 = n18069 ^ n6682 ^ n2688 ;
  assign n18078 = n18077 ^ n18070 ^ 1'b0 ;
  assign n18093 = n739 | n6180 ;
  assign n18079 = n6649 & n7283 ;
  assign n18080 = n2314 & n18079 ;
  assign n18081 = n2597 | n18080 ;
  assign n18082 = n3730 & ~n18081 ;
  assign n18083 = ( n2110 & n3837 ) | ( n2110 & n18082 ) | ( n3837 & n18082 ) ;
  assign n18084 = ( n1751 & n4259 ) | ( n1751 & n5427 ) | ( n4259 & n5427 ) ;
  assign n18085 = n18084 ^ n12833 ^ 1'b0 ;
  assign n18086 = n2759 & n8431 ;
  assign n18087 = n18086 ^ n3226 ^ 1'b0 ;
  assign n18088 = ~n8686 & n18087 ;
  assign n18089 = n12487 ^ n3616 ^ 1'b0 ;
  assign n18090 = n18088 | n18089 ;
  assign n18091 = ~n18085 & n18090 ;
  assign n18092 = n18083 & ~n18091 ;
  assign n18094 = n18093 ^ n18092 ^ 1'b0 ;
  assign n18095 = n4416 & n15182 ;
  assign n18096 = n18095 ^ n5310 ^ 1'b0 ;
  assign n18097 = n13053 & n18096 ;
  assign n18098 = n18097 ^ n7752 ^ 1'b0 ;
  assign n18099 = n5860 ^ n3921 ^ 1'b0 ;
  assign n18100 = ~n2787 & n18099 ;
  assign n18101 = ~n1670 & n8900 ;
  assign n18102 = n18100 & n18101 ;
  assign n18103 = n14641 ^ n10659 ^ n10261 ;
  assign n18104 = n8427 ^ x174 ^ 1'b0 ;
  assign n18105 = n3991 & n18104 ;
  assign n18106 = n3335 & n18105 ;
  assign n18107 = n18106 ^ n3439 ^ 1'b0 ;
  assign n18108 = ( n848 & n9023 ) | ( n848 & n15191 ) | ( n9023 & n15191 ) ;
  assign n18109 = n18108 ^ n15659 ^ n5084 ;
  assign n18111 = ( n498 & ~n7832 ) | ( n498 & n10832 ) | ( ~n7832 & n10832 ) ;
  assign n18112 = n4295 & n18111 ;
  assign n18110 = ~n10681 & n17143 ;
  assign n18113 = n18112 ^ n18110 ^ 1'b0 ;
  assign n18114 = n17873 ^ n17460 ^ 1'b0 ;
  assign n18115 = ~n2114 & n2187 ;
  assign n18116 = ~n6525 & n18115 ;
  assign n18117 = n16625 ^ n13377 ^ n3790 ;
  assign n18118 = ( n9546 & ~n18116 ) | ( n9546 & n18117 ) | ( ~n18116 & n18117 ) ;
  assign n18119 = ~n7335 & n18118 ;
  assign n18120 = n7221 ^ x203 ^ 1'b0 ;
  assign n18121 = n18120 ^ n9823 ^ n2819 ;
  assign n18122 = x24 & ~n1780 ;
  assign n18123 = ~n12854 & n18122 ;
  assign n18124 = n18123 ^ n5593 ^ 1'b0 ;
  assign n18125 = ~n11139 & n18124 ;
  assign n18126 = n1139 & ~n2819 ;
  assign n18127 = ( ~n835 & n18125 ) | ( ~n835 & n18126 ) | ( n18125 & n18126 ) ;
  assign n18128 = n3115 & ~n11285 ;
  assign n18132 = ( n2412 & n9618 ) | ( n2412 & ~n13075 ) | ( n9618 & ~n13075 ) ;
  assign n18129 = n1356 ^ n1105 ^ 1'b0 ;
  assign n18130 = n18129 ^ n9652 ^ 1'b0 ;
  assign n18131 = ( n8461 & n16161 ) | ( n8461 & n18130 ) | ( n16161 & n18130 ) ;
  assign n18133 = n18132 ^ n18131 ^ n15109 ;
  assign n18134 = n14471 ^ n594 ^ 1'b0 ;
  assign n18135 = n18133 & ~n18134 ;
  assign n18136 = n12872 ^ n3211 ^ n3004 ;
  assign n18137 = n13153 ^ n9957 ^ n2469 ;
  assign n18138 = n18136 | n18137 ;
  assign n18139 = ( x41 & n9791 ) | ( x41 & n18138 ) | ( n9791 & n18138 ) ;
  assign n18140 = ( n510 & n3431 ) | ( n510 & n15169 ) | ( n3431 & n15169 ) ;
  assign n18141 = n18140 ^ n9380 ^ n399 ;
  assign n18142 = n5787 ^ x179 ^ 1'b0 ;
  assign n18143 = n9548 & n18142 ;
  assign n18144 = n4842 | n18143 ;
  assign n18145 = n18144 ^ n12236 ^ n8085 ;
  assign n18146 = n6202 & ~n9404 ;
  assign n18147 = n18146 ^ n5671 ^ 1'b0 ;
  assign n18148 = n18147 ^ n8378 ^ 1'b0 ;
  assign n18149 = ~n6838 & n14837 ;
  assign n18150 = n11173 & n18149 ;
  assign n18151 = x38 | n4978 ;
  assign n18152 = ~n6433 & n6893 ;
  assign n18153 = n8492 & n18152 ;
  assign n18154 = ( n1131 & n18151 ) | ( n1131 & ~n18153 ) | ( n18151 & ~n18153 ) ;
  assign n18155 = ( n17501 & n18150 ) | ( n17501 & n18154 ) | ( n18150 & n18154 ) ;
  assign n18156 = n6237 | n13394 ;
  assign n18157 = ~n1098 & n18156 ;
  assign n18158 = ~n6613 & n18157 ;
  assign n18160 = n7588 ^ n6362 ^ n3178 ;
  assign n18159 = n13115 ^ n3682 ^ n2106 ;
  assign n18161 = n18160 ^ n18159 ^ n5878 ;
  assign n18162 = n18161 ^ n14781 ^ n11992 ;
  assign n18163 = ( n7514 & ~n7851 ) | ( n7514 & n10009 ) | ( ~n7851 & n10009 ) ;
  assign n18164 = n18163 ^ n10173 ^ n6966 ;
  assign n18165 = n15649 & ~n15963 ;
  assign n18166 = n18165 ^ n4340 ^ 1'b0 ;
  assign n18167 = ( n8876 & n14803 ) | ( n8876 & n15575 ) | ( n14803 & n15575 ) ;
  assign n18168 = n8915 & ~n9814 ;
  assign n18169 = ~n18167 & n18168 ;
  assign n18170 = n589 | n18169 ;
  assign n18171 = n18166 | n18170 ;
  assign n18174 = n7571 | n8178 ;
  assign n18172 = ~n6053 & n12230 ;
  assign n18173 = n2064 & n18172 ;
  assign n18175 = n18174 ^ n18173 ^ 1'b0 ;
  assign n18176 = n5707 & ~n18175 ;
  assign n18177 = n18176 ^ n13103 ^ n6522 ;
  assign n18178 = n3720 | n18177 ;
  assign n18180 = n13615 ^ n3912 ^ n2623 ;
  assign n18179 = ( n10692 & n10998 ) | ( n10692 & n11360 ) | ( n10998 & n11360 ) ;
  assign n18181 = n18180 ^ n18179 ^ 1'b0 ;
  assign n18182 = ~n1771 & n1773 ;
  assign n18183 = n1988 & n9338 ;
  assign n18184 = ~n15959 & n18183 ;
  assign n18185 = ( n8428 & ~n18182 ) | ( n8428 & n18184 ) | ( ~n18182 & n18184 ) ;
  assign n18186 = n6337 & n7494 ;
  assign n18187 = ~n8883 & n18186 ;
  assign n18188 = n14514 ^ n7563 ^ n331 ;
  assign n18189 = n18187 & n18188 ;
  assign n18193 = ( n3790 & n3994 ) | ( n3790 & n12206 ) | ( n3994 & n12206 ) ;
  assign n18194 = ( ~n5106 & n11046 ) | ( ~n5106 & n18193 ) | ( n11046 & n18193 ) ;
  assign n18192 = n5707 ^ n4228 ^ n1840 ;
  assign n18190 = n15454 ^ n7342 ^ 1'b0 ;
  assign n18191 = n2801 & ~n18190 ;
  assign n18195 = n18194 ^ n18192 ^ n18191 ;
  assign n18196 = n11112 & ~n18195 ;
  assign n18197 = n11261 ^ n6195 ^ n2306 ;
  assign n18198 = n18197 ^ n3101 ^ n2121 ;
  assign n18199 = n4288 | n18198 ;
  assign n18200 = n7708 | n18199 ;
  assign n18201 = n7031 | n18200 ;
  assign n18202 = ( n3918 & n9582 ) | ( n3918 & n18201 ) | ( n9582 & n18201 ) ;
  assign n18203 = ( ~n5487 & n15757 ) | ( ~n5487 & n17687 ) | ( n15757 & n17687 ) ;
  assign n18205 = n4180 & n8723 ;
  assign n18206 = n18205 ^ n4678 ^ 1'b0 ;
  assign n18204 = n7106 ^ n1448 ^ 1'b0 ;
  assign n18207 = n18206 ^ n18204 ^ 1'b0 ;
  assign n18208 = n18207 ^ n7989 ^ n5126 ;
  assign n18209 = n1611 & ~n7732 ;
  assign n18210 = n18209 ^ n10753 ^ n9187 ;
  assign n18211 = n3448 | n9724 ;
  assign n18212 = n14685 & ~n18211 ;
  assign n18213 = n5217 ^ n3678 ^ 1'b0 ;
  assign n18214 = ( n3646 & ~n4990 ) | ( n3646 & n18213 ) | ( ~n4990 & n18213 ) ;
  assign n18215 = n3826 ^ n540 ^ 1'b0 ;
  assign n18216 = ~n9471 & n18215 ;
  assign n18217 = ~n13160 & n18216 ;
  assign n18218 = n18217 ^ n9852 ^ 1'b0 ;
  assign n18219 = n2327 & ~n18218 ;
  assign n18220 = n16322 ^ n14670 ^ n8456 ;
  assign n18221 = ~n4224 & n12565 ;
  assign n18222 = n8558 & ~n18221 ;
  assign n18223 = n15071 ^ n13273 ^ 1'b0 ;
  assign n18224 = n16369 & n18223 ;
  assign n18232 = n12884 ^ n12239 ^ 1'b0 ;
  assign n18233 = n6981 & n18232 ;
  assign n18225 = n2991 | n3368 ;
  assign n18226 = n18225 ^ n5902 ^ 1'b0 ;
  assign n18227 = x126 & n1319 ;
  assign n18228 = n9485 & n18227 ;
  assign n18229 = ( n4053 & ~n18226 ) | ( n4053 & n18228 ) | ( ~n18226 & n18228 ) ;
  assign n18230 = n18229 ^ n14350 ^ 1'b0 ;
  assign n18231 = n9539 | n18230 ;
  assign n18234 = n18233 ^ n18231 ^ 1'b0 ;
  assign n18235 = n5981 ^ n5908 ^ 1'b0 ;
  assign n18236 = n18235 ^ n9552 ^ 1'b0 ;
  assign n18237 = n14155 & ~n18236 ;
  assign n18238 = ( n2886 & ~n7578 ) | ( n2886 & n18237 ) | ( ~n7578 & n18237 ) ;
  assign n18242 = ( ~n3586 & n3931 ) | ( ~n3586 & n5128 ) | ( n3931 & n5128 ) ;
  assign n18243 = n18242 ^ n10485 ^ 1'b0 ;
  assign n18239 = ( n2188 & n12222 ) | ( n2188 & n12285 ) | ( n12222 & n12285 ) ;
  assign n18240 = n11673 ^ n4946 ^ n4724 ;
  assign n18241 = ( n9122 & ~n18239 ) | ( n9122 & n18240 ) | ( ~n18239 & n18240 ) ;
  assign n18244 = n18243 ^ n18241 ^ n5303 ;
  assign n18245 = n7139 ^ n1422 ^ 1'b0 ;
  assign n18246 = n12976 | n18245 ;
  assign n18247 = ( n1491 & n5110 ) | ( n1491 & n18246 ) | ( n5110 & n18246 ) ;
  assign n18248 = n18046 ^ n3037 ^ 1'b0 ;
  assign n18249 = n15305 ^ n2495 ^ 1'b0 ;
  assign n18250 = ~n18248 & n18249 ;
  assign n18251 = n18250 ^ n4166 ^ 1'b0 ;
  assign n18252 = n13671 & ~n15750 ;
  assign n18253 = n12243 ^ n7504 ^ 1'b0 ;
  assign n18254 = n1372 | n18253 ;
  assign n18255 = ( n9796 & n12082 ) | ( n9796 & ~n18254 ) | ( n12082 & ~n18254 ) ;
  assign n18256 = n6640 | n17985 ;
  assign n18257 = n18256 ^ n7878 ^ 1'b0 ;
  assign n18258 = ( n3187 & n6650 ) | ( n3187 & n18257 ) | ( n6650 & n18257 ) ;
  assign n18259 = ~n18255 & n18258 ;
  assign n18260 = n18259 ^ n15637 ^ 1'b0 ;
  assign n18261 = ~n16159 & n18260 ;
  assign n18262 = ~n11354 & n15184 ;
  assign n18263 = ~n9140 & n18262 ;
  assign n18264 = n10845 ^ n4644 ^ 1'b0 ;
  assign n18265 = n2587 & n16225 ;
  assign n18266 = n14577 & n18265 ;
  assign n18267 = n3298 & ~n14788 ;
  assign n18268 = n18267 ^ n6592 ^ x199 ;
  assign n18269 = ( n2310 & ~n18266 ) | ( n2310 & n18268 ) | ( ~n18266 & n18268 ) ;
  assign n18270 = ~n18264 & n18269 ;
  assign n18271 = n12936 & n13884 ;
  assign n18272 = ~n7295 & n13126 ;
  assign n18273 = ( n11748 & n17882 ) | ( n11748 & ~n18272 ) | ( n17882 & ~n18272 ) ;
  assign n18274 = n6249 ^ n4209 ^ 1'b0 ;
  assign n18275 = n614 & ~n18274 ;
  assign n18276 = ( n7147 & n8665 ) | ( n7147 & n18275 ) | ( n8665 & n18275 ) ;
  assign n18279 = n6219 ^ n3220 ^ 1'b0 ;
  assign n18280 = n18279 ^ x121 ^ 1'b0 ;
  assign n18281 = n18280 ^ n4536 ^ 1'b0 ;
  assign n18277 = n9161 ^ n5307 ^ 1'b0 ;
  assign n18278 = ( n6070 & n6498 ) | ( n6070 & ~n18277 ) | ( n6498 & ~n18277 ) ;
  assign n18282 = n18281 ^ n18278 ^ 1'b0 ;
  assign n18283 = n18276 & n18282 ;
  assign n18284 = n11674 ^ n2572 ^ n1320 ;
  assign n18285 = n339 & ~n18284 ;
  assign n18286 = n1602 | n18285 ;
  assign n18287 = n9730 ^ n5803 ^ 1'b0 ;
  assign n18288 = n4216 | n18287 ;
  assign n18289 = n18288 ^ n11873 ^ 1'b0 ;
  assign n18290 = ~n7815 & n8611 ;
  assign n18291 = n3970 & n18290 ;
  assign n18292 = ~n4085 & n14889 ;
  assign n18293 = n7906 ^ n6643 ^ 1'b0 ;
  assign n18294 = n8768 ^ n4504 ^ n1993 ;
  assign n18295 = n18294 ^ n15434 ^ 1'b0 ;
  assign n18296 = ~n18293 & n18295 ;
  assign n18297 = ( n7827 & n9940 ) | ( n7827 & n15833 ) | ( n9940 & n15833 ) ;
  assign n18298 = ( n346 & n3360 ) | ( n346 & n10887 ) | ( n3360 & n10887 ) ;
  assign n18299 = n3064 | n4653 ;
  assign n18300 = n18298 & ~n18299 ;
  assign n18301 = n18297 & n18300 ;
  assign n18302 = n11717 ^ n7210 ^ 1'b0 ;
  assign n18303 = n18301 & n18302 ;
  assign n18304 = n8827 ^ n5782 ^ 1'b0 ;
  assign n18305 = ( n13580 & ~n16724 ) | ( n13580 & n18304 ) | ( ~n16724 & n18304 ) ;
  assign n18306 = n13063 ^ n5836 ^ n5624 ;
  assign n18310 = n3329 ^ x9 ^ 1'b0 ;
  assign n18307 = n14912 ^ n7795 ^ 1'b0 ;
  assign n18308 = n14789 | n18307 ;
  assign n18309 = n18308 ^ n14428 ^ 1'b0 ;
  assign n18311 = n18310 ^ n18309 ^ n14568 ;
  assign n18312 = ( n1961 & ~n6000 ) | ( n1961 & n16885 ) | ( ~n6000 & n16885 ) ;
  assign n18313 = n18312 ^ n7551 ^ 1'b0 ;
  assign n18314 = n18311 & ~n18313 ;
  assign n18315 = ~n18306 & n18314 ;
  assign n18316 = ~n1941 & n18315 ;
  assign n18317 = n12834 ^ n2585 ^ 1'b0 ;
  assign n18318 = n14778 ^ n4017 ^ n901 ;
  assign n18319 = n18318 ^ n492 ^ x142 ;
  assign n18323 = ~n13929 & n16580 ;
  assign n18321 = n11294 ^ n5449 ^ x252 ;
  assign n18320 = ~n1201 & n10889 ;
  assign n18322 = n18321 ^ n18320 ^ n5728 ;
  assign n18324 = n18323 ^ n18322 ^ n7463 ;
  assign n18329 = ( n6223 & n11045 ) | ( n6223 & ~n16896 ) | ( n11045 & ~n16896 ) ;
  assign n18330 = n18329 ^ n4405 ^ n1222 ;
  assign n18325 = ( x160 & n1653 ) | ( x160 & ~n4492 ) | ( n1653 & ~n4492 ) ;
  assign n18326 = n5500 & ~n18325 ;
  assign n18327 = n11056 ^ n6310 ^ 1'b0 ;
  assign n18328 = n18326 & ~n18327 ;
  assign n18331 = n18330 ^ n18328 ^ 1'b0 ;
  assign n18332 = n1356 & n5454 ;
  assign n18333 = ~n6170 & n18332 ;
  assign n18334 = ( ~n5731 & n6976 ) | ( ~n5731 & n7395 ) | ( n6976 & n7395 ) ;
  assign n18335 = n18334 ^ n9775 ^ 1'b0 ;
  assign n18336 = n18333 | n18335 ;
  assign n18337 = n6039 ^ n4224 ^ 1'b0 ;
  assign n18338 = n18337 ^ n6382 ^ x94 ;
  assign n18339 = n862 ^ n470 ^ 1'b0 ;
  assign n18340 = ( n818 & ~n12072 ) | ( n818 & n16237 ) | ( ~n12072 & n16237 ) ;
  assign n18341 = n8042 ^ n1087 ^ 1'b0 ;
  assign n18342 = n9751 & n18341 ;
  assign n18343 = ~n18248 & n18342 ;
  assign n18344 = n18343 ^ x48 ^ 1'b0 ;
  assign n18345 = n11772 ^ n3046 ^ 1'b0 ;
  assign n18346 = n12778 ^ n1246 ^ 1'b0 ;
  assign n18347 = ~n18345 & n18346 ;
  assign n18348 = ( n5589 & n6681 ) | ( n5589 & n17924 ) | ( n6681 & n17924 ) ;
  assign n18349 = ~n2965 & n9435 ;
  assign n18350 = n18349 ^ n1249 ^ 1'b0 ;
  assign n18351 = ( n4652 & n18348 ) | ( n4652 & n18350 ) | ( n18348 & n18350 ) ;
  assign n18352 = n10401 ^ n2131 ^ n362 ;
  assign n18353 = n18352 ^ n17867 ^ n1733 ;
  assign n18354 = n5681 | n6354 ;
  assign n18355 = n18354 ^ n14293 ^ n8584 ;
  assign n18356 = n2672 & n18355 ;
  assign n18357 = ~n18353 & n18356 ;
  assign n18358 = n4454 ^ n914 ^ x21 ;
  assign n18359 = n18358 ^ n4085 ^ 1'b0 ;
  assign n18360 = ( n5517 & n15017 ) | ( n5517 & n18359 ) | ( n15017 & n18359 ) ;
  assign n18361 = n5687 & ~n7174 ;
  assign n18362 = ( n6442 & n10887 ) | ( n6442 & n18361 ) | ( n10887 & n18361 ) ;
  assign n18363 = n5179 ^ n2706 ^ 1'b0 ;
  assign n18364 = n18363 ^ n16943 ^ 1'b0 ;
  assign n18365 = n16557 ^ n16143 ^ n3629 ;
  assign n18366 = n1638 & ~n2813 ;
  assign n18367 = ~n2316 & n18366 ;
  assign n18368 = n18367 ^ n1422 ^ 1'b0 ;
  assign n18369 = n9247 & ~n18368 ;
  assign n18370 = ( n1543 & ~n2172 ) | ( n1543 & n5931 ) | ( ~n2172 & n5931 ) ;
  assign n18371 = ~n11607 & n18370 ;
  assign n18372 = n18371 ^ n9282 ^ 1'b0 ;
  assign n18373 = ( n2204 & n10658 ) | ( n2204 & ~n18372 ) | ( n10658 & ~n18372 ) ;
  assign n18375 = ~n5731 & n7345 ;
  assign n18374 = n12116 ^ n8212 ^ 1'b0 ;
  assign n18376 = n18375 ^ n18374 ^ n9471 ;
  assign n18377 = n18376 ^ n8595 ^ n4811 ;
  assign n18386 = ~n1969 & n7283 ;
  assign n18385 = n10681 ^ n2440 ^ 1'b0 ;
  assign n18378 = n4990 ^ n647 ^ 1'b0 ;
  assign n18379 = n9385 & n18378 ;
  assign n18380 = n11767 & ~n18379 ;
  assign n18381 = n4833 ^ n2052 ^ 1'b0 ;
  assign n18382 = n2070 & n18381 ;
  assign n18383 = n18382 ^ n13929 ^ 1'b0 ;
  assign n18384 = n18380 & ~n18383 ;
  assign n18387 = n18386 ^ n18385 ^ n18384 ;
  assign n18388 = ( n1423 & n1624 ) | ( n1423 & ~n8538 ) | ( n1624 & ~n8538 ) ;
  assign n18389 = ( ~x222 & n2242 ) | ( ~x222 & n5482 ) | ( n2242 & n5482 ) ;
  assign n18390 = n18388 | n18389 ;
  assign n18394 = n14860 ^ n9025 ^ n332 ;
  assign n18391 = ~n3773 & n6396 ;
  assign n18392 = n4686 & n18391 ;
  assign n18393 = n18392 ^ n7079 ^ n4334 ;
  assign n18395 = n18394 ^ n18393 ^ n4788 ;
  assign n18396 = n6469 | n10784 ;
  assign n18397 = n14868 ^ n1932 ^ 1'b0 ;
  assign n18398 = ( n2260 & n12897 ) | ( n2260 & ~n14168 ) | ( n12897 & ~n14168 ) ;
  assign n18399 = ( n3518 & n16066 ) | ( n3518 & n18398 ) | ( n16066 & n18398 ) ;
  assign n18400 = n15357 ^ n14245 ^ n12230 ;
  assign n18401 = n5043 ^ n2240 ^ n1880 ;
  assign n18402 = ( n3741 & n13780 ) | ( n3741 & ~n14730 ) | ( n13780 & ~n14730 ) ;
  assign n18403 = ( n13292 & ~n18401 ) | ( n13292 & n18402 ) | ( ~n18401 & n18402 ) ;
  assign n18404 = n13759 ^ n13358 ^ n1504 ;
  assign n18405 = ~n15521 & n18404 ;
  assign n18406 = n18403 & n18405 ;
  assign n18407 = n11634 & ~n13980 ;
  assign n18408 = ~n14169 & n18407 ;
  assign n18409 = ( n4727 & n16660 ) | ( n4727 & n16918 ) | ( n16660 & n16918 ) ;
  assign n18410 = n2095 & n6987 ;
  assign n18411 = n18410 ^ n14741 ^ n2418 ;
  assign n18412 = n11682 ^ n3854 ^ 1'b0 ;
  assign n18413 = n3994 & n18412 ;
  assign n18414 = n18413 ^ n16054 ^ 1'b0 ;
  assign n18415 = n2426 | n18414 ;
  assign n18416 = x138 & n13741 ;
  assign n18417 = n11350 & n18416 ;
  assign n18418 = ( ~n1505 & n6229 ) | ( ~n1505 & n10724 ) | ( n6229 & n10724 ) ;
  assign n18419 = n18418 ^ n7664 ^ n1233 ;
  assign n18420 = n13841 ^ n7072 ^ n3721 ;
  assign n18421 = n1046 & ~n3753 ;
  assign n18422 = n2185 | n18421 ;
  assign n18423 = n18422 ^ n10488 ^ 1'b0 ;
  assign n18424 = n18423 ^ n13726 ^ n7013 ;
  assign n18425 = n10302 | n18424 ;
  assign n18426 = n1078 | n18425 ;
  assign n18428 = n2039 | n2992 ;
  assign n18429 = n18428 ^ n7150 ^ n3111 ;
  assign n18430 = n18429 ^ n15642 ^ n10972 ;
  assign n18427 = n3320 | n4814 ;
  assign n18431 = n18430 ^ n18427 ^ 1'b0 ;
  assign n18432 = n1266 | n2185 ;
  assign n18433 = n18432 ^ n16231 ^ 1'b0 ;
  assign n18436 = ( x78 & n3577 ) | ( x78 & ~n9425 ) | ( n3577 & ~n9425 ) ;
  assign n18434 = n17174 ^ n7388 ^ n4310 ;
  assign n18435 = ( n6051 & n6695 ) | ( n6051 & n18434 ) | ( n6695 & n18434 ) ;
  assign n18437 = n18436 ^ n18435 ^ n8946 ;
  assign n18438 = n12262 & ~n15521 ;
  assign n18441 = n11310 ^ n8235 ^ 1'b0 ;
  assign n18440 = x230 & ~n4605 ;
  assign n18442 = n18441 ^ n18440 ^ 1'b0 ;
  assign n18439 = n10443 ^ n7602 ^ n1257 ;
  assign n18443 = n18442 ^ n18439 ^ n5353 ;
  assign n18444 = n18443 ^ n5541 ^ 1'b0 ;
  assign n18445 = ( n1751 & ~n3891 ) | ( n1751 & n3955 ) | ( ~n3891 & n3955 ) ;
  assign n18446 = n18445 ^ n15575 ^ n2192 ;
  assign n18447 = n10196 ^ x88 ^ 1'b0 ;
  assign n18448 = ( n4171 & n9053 ) | ( n4171 & n18447 ) | ( n9053 & n18447 ) ;
  assign n18449 = n5316 ^ n3013 ^ n988 ;
  assign n18450 = n17638 ^ n6805 ^ 1'b0 ;
  assign n18451 = ( n1463 & ~n8422 ) | ( n1463 & n18450 ) | ( ~n8422 & n18450 ) ;
  assign n18452 = n7470 ^ n448 ^ x151 ;
  assign n18453 = n11122 & n18452 ;
  assign n18454 = n18453 ^ n2194 ^ 1'b0 ;
  assign n18455 = ( x128 & ~n6867 ) | ( x128 & n18454 ) | ( ~n6867 & n18454 ) ;
  assign n18456 = ( ~n465 & n8757 ) | ( ~n465 & n11320 ) | ( n8757 & n11320 ) ;
  assign n18457 = n18456 ^ n1062 ^ 1'b0 ;
  assign n18458 = ~n18455 & n18457 ;
  assign n18459 = ~n13024 & n18458 ;
  assign n18460 = ( n2001 & n6626 ) | ( n2001 & ~n6670 ) | ( n6626 & ~n6670 ) ;
  assign n18461 = n10270 & ~n18460 ;
  assign n18462 = ( n12841 & ~n16993 ) | ( n12841 & n18461 ) | ( ~n16993 & n18461 ) ;
  assign n18475 = n3061 & ~n13430 ;
  assign n18476 = ~n4302 & n18475 ;
  assign n18469 = ( n277 & n5648 ) | ( n277 & n7098 ) | ( n5648 & n7098 ) ;
  assign n18470 = ~n922 & n1865 ;
  assign n18471 = ~n14279 & n18470 ;
  assign n18472 = n8334 | n18471 ;
  assign n18473 = n18469 | n18472 ;
  assign n18474 = n6386 & n18473 ;
  assign n18477 = n18476 ^ n18474 ^ 1'b0 ;
  assign n18478 = n18477 ^ n5598 ^ 1'b0 ;
  assign n18464 = ( n2021 & ~n5688 ) | ( n2021 & n5949 ) | ( ~n5688 & n5949 ) ;
  assign n18465 = ~n5353 & n18215 ;
  assign n18466 = n18464 & n18465 ;
  assign n18467 = n6289 | n18466 ;
  assign n18468 = n18467 ^ n8794 ^ 1'b0 ;
  assign n18463 = n13408 ^ n6369 ^ n810 ;
  assign n18479 = n18478 ^ n18468 ^ n18463 ;
  assign n18480 = ( n5585 & ~n6596 ) | ( n5585 & n18479 ) | ( ~n6596 & n18479 ) ;
  assign n18481 = n11375 ^ n1629 ^ n331 ;
  assign n18482 = ( x202 & ~n6774 ) | ( x202 & n18481 ) | ( ~n6774 & n18481 ) ;
  assign n18488 = n12570 ^ n10014 ^ n2867 ;
  assign n18485 = n6023 ^ n4161 ^ n3942 ;
  assign n18486 = n1685 | n2696 ;
  assign n18487 = ( n5064 & ~n18485 ) | ( n5064 & n18486 ) | ( ~n18485 & n18486 ) ;
  assign n18483 = n7279 ^ n1293 ^ 1'b0 ;
  assign n18484 = n18483 ^ n13338 ^ 1'b0 ;
  assign n18489 = n18488 ^ n18487 ^ n18484 ;
  assign n18491 = ( n1046 & ~n5368 ) | ( n1046 & n10453 ) | ( ~n5368 & n10453 ) ;
  assign n18490 = n2978 | n11274 ;
  assign n18492 = n18491 ^ n18490 ^ 1'b0 ;
  assign n18494 = n2527 ^ n1759 ^ 1'b0 ;
  assign n18493 = n1411 & ~n10314 ;
  assign n18495 = n18494 ^ n18493 ^ 1'b0 ;
  assign n18496 = ( n3076 & ~n4914 ) | ( n3076 & n18495 ) | ( ~n4914 & n18495 ) ;
  assign n18497 = ( n8337 & n10609 ) | ( n8337 & ~n18496 ) | ( n10609 & ~n18496 ) ;
  assign n18501 = n721 & ~n9356 ;
  assign n18502 = n18501 ^ n2337 ^ 1'b0 ;
  assign n18498 = ( n13814 & n14995 ) | ( n13814 & ~n15840 ) | ( n14995 & ~n15840 ) ;
  assign n18499 = n3950 | n7684 ;
  assign n18500 = n18498 & ~n18499 ;
  assign n18503 = n18502 ^ n18500 ^ n1560 ;
  assign n18504 = ( n710 & ~n857 ) | ( n710 & n2177 ) | ( ~n857 & n2177 ) ;
  assign n18505 = n8247 ^ n6550 ^ 1'b0 ;
  assign n18506 = n8505 & ~n18505 ;
  assign n18507 = ( ~n13694 & n18504 ) | ( ~n13694 & n18506 ) | ( n18504 & n18506 ) ;
  assign n18508 = n11229 ^ n6559 ^ n1399 ;
  assign n18509 = ( n1353 & n2004 ) | ( n1353 & n18508 ) | ( n2004 & n18508 ) ;
  assign n18510 = n18509 ^ n11937 ^ n4966 ;
  assign n18511 = ~n15687 & n18510 ;
  assign n18512 = n10854 & n12775 ;
  assign n18513 = n8037 ^ n5963 ^ n3349 ;
  assign n18514 = x130 & n759 ;
  assign n18515 = x206 & ~n14105 ;
  assign n18516 = ~n2029 & n18515 ;
  assign n18517 = n6298 | n18516 ;
  assign n18518 = n18517 ^ n5041 ^ 1'b0 ;
  assign n18519 = ( ~n1854 & n6155 ) | ( ~n1854 & n18518 ) | ( n6155 & n18518 ) ;
  assign n18520 = n18519 ^ n15221 ^ n4673 ;
  assign n18521 = ( ~n18513 & n18514 ) | ( ~n18513 & n18520 ) | ( n18514 & n18520 ) ;
  assign n18522 = ( n12129 & n17567 ) | ( n12129 & ~n18521 ) | ( n17567 & ~n18521 ) ;
  assign n18523 = x182 & ~n3420 ;
  assign n18524 = n18523 ^ n8731 ^ 1'b0 ;
  assign n18525 = n18524 ^ n1162 ^ x156 ;
  assign n18526 = n18525 ^ n10546 ^ n3220 ;
  assign n18527 = n2649 & n5676 ;
  assign n18528 = n16989 ^ n4084 ^ 1'b0 ;
  assign n18529 = n18527 & ~n18528 ;
  assign n18530 = n9172 ^ n7776 ^ 1'b0 ;
  assign n18531 = n12972 & ~n18530 ;
  assign n18532 = ~n1372 & n10395 ;
  assign n18533 = n6001 ^ n3754 ^ 1'b0 ;
  assign n18534 = ( n1713 & ~n18532 ) | ( n1713 & n18533 ) | ( ~n18532 & n18533 ) ;
  assign n18535 = n18534 ^ n17955 ^ n14170 ;
  assign n18536 = n2596 ^ n2139 ^ n628 ;
  assign n18537 = n9418 ^ n2704 ^ 1'b0 ;
  assign n18538 = ( n10335 & ~n18536 ) | ( n10335 & n18537 ) | ( ~n18536 & n18537 ) ;
  assign n18539 = n3646 & n12001 ;
  assign n18544 = n1469 | n16230 ;
  assign n18545 = n18544 ^ n6998 ^ n643 ;
  assign n18543 = n5342 & n10921 ;
  assign n18540 = ( n8256 & ~n9844 ) | ( n8256 & n16887 ) | ( ~n9844 & n16887 ) ;
  assign n18541 = n6916 | n18540 ;
  assign n18542 = n4247 | n18541 ;
  assign n18546 = n18545 ^ n18543 ^ n18542 ;
  assign n18547 = n8545 | n16741 ;
  assign n18548 = n13864 | n18547 ;
  assign n18549 = n439 & n5913 ;
  assign n18550 = n18549 ^ n11197 ^ n5079 ;
  assign n18551 = n1743 | n18550 ;
  assign n18552 = n5558 ^ n1724 ^ n448 ;
  assign n18553 = n9074 & ~n18552 ;
  assign n18554 = ~n4483 & n18553 ;
  assign n18555 = n12354 ^ n6455 ^ 1'b0 ;
  assign n18556 = n18555 ^ n12388 ^ n7021 ;
  assign n18557 = ( x51 & n10453 ) | ( x51 & ~n13250 ) | ( n10453 & ~n13250 ) ;
  assign n18558 = x245 | n7116 ;
  assign n18559 = n8917 ^ n1682 ^ 1'b0 ;
  assign n18560 = n8867 | n18559 ;
  assign n18561 = n18558 & ~n18560 ;
  assign n18562 = n18561 ^ n11696 ^ 1'b0 ;
  assign n18563 = n9340 ^ n7903 ^ n2549 ;
  assign n18564 = n4972 & ~n13158 ;
  assign n18565 = n18564 ^ n9409 ^ 1'b0 ;
  assign n18566 = ( n11009 & n18563 ) | ( n11009 & n18565 ) | ( n18563 & n18565 ) ;
  assign n18570 = ( n2845 & n6611 ) | ( n2845 & n7150 ) | ( n6611 & n7150 ) ;
  assign n18571 = ( ~n13109 & n13670 ) | ( ~n13109 & n18570 ) | ( n13670 & n18570 ) ;
  assign n18567 = n1197 & n5717 ;
  assign n18568 = n18567 ^ n343 ^ 1'b0 ;
  assign n18569 = x209 & ~n18568 ;
  assign n18572 = n18571 ^ n18569 ^ x84 ;
  assign n18573 = n14677 ^ n10140 ^ 1'b0 ;
  assign n18574 = n1821 & ~n18573 ;
  assign n18575 = n18574 ^ n16737 ^ n4877 ;
  assign n18576 = n6355 ^ n2858 ^ n2419 ;
  assign n18577 = ~n3033 & n5213 ;
  assign n18578 = n18577 ^ n8937 ^ 1'b0 ;
  assign n18579 = n8462 ^ n2545 ^ n317 ;
  assign n18580 = ( n18576 & n18578 ) | ( n18576 & ~n18579 ) | ( n18578 & ~n18579 ) ;
  assign n18581 = n18580 ^ n17821 ^ n3125 ;
  assign n18582 = n4680 & n18581 ;
  assign n18583 = ~n18575 & n18582 ;
  assign n18584 = n17712 ^ n16775 ^ n10854 ;
  assign n18585 = ( n587 & n4767 ) | ( n587 & n18584 ) | ( n4767 & n18584 ) ;
  assign n18586 = n2711 ^ x253 ^ 1'b0 ;
  assign n18587 = n12291 | n13673 ;
  assign n18589 = ( n4221 & n6645 ) | ( n4221 & ~n7087 ) | ( n6645 & ~n7087 ) ;
  assign n18590 = n18589 ^ n7472 ^ 1'b0 ;
  assign n18588 = ( n5901 & n8095 ) | ( n5901 & n9310 ) | ( n8095 & n9310 ) ;
  assign n18591 = n18590 ^ n18588 ^ 1'b0 ;
  assign n18592 = x11 & ~n18591 ;
  assign n18593 = n18592 ^ n11429 ^ n5637 ;
  assign n18594 = n18587 & n18593 ;
  assign n18595 = ( n10429 & n18586 ) | ( n10429 & n18594 ) | ( n18586 & n18594 ) ;
  assign n18596 = x29 & n12148 ;
  assign n18597 = n17770 ^ n15798 ^ 1'b0 ;
  assign n18598 = n12435 & ~n18597 ;
  assign n18599 = n18598 ^ n12511 ^ 1'b0 ;
  assign n18601 = n18584 ^ n10544 ^ n2711 ;
  assign n18600 = n5991 | n10619 ;
  assign n18602 = n18601 ^ n18600 ^ n13705 ;
  assign n18603 = n6417 ^ n4737 ^ 1'b0 ;
  assign n18604 = n4109 & ~n18603 ;
  assign n18605 = ~n8880 & n18604 ;
  assign n18606 = n356 & n18605 ;
  assign n18607 = ~n17803 & n18606 ;
  assign n18608 = ~n4491 & n7923 ;
  assign n18609 = n18608 ^ n10732 ^ 1'b0 ;
  assign n18610 = n2022 | n3560 ;
  assign n18611 = n13608 & ~n18610 ;
  assign n18612 = ( n14446 & n18442 ) | ( n14446 & ~n18611 ) | ( n18442 & ~n18611 ) ;
  assign n18613 = n18609 & n18612 ;
  assign n18614 = n18613 ^ n18064 ^ n14501 ;
  assign n18616 = ( ~n1289 & n3430 ) | ( ~n1289 & n12591 ) | ( n3430 & n12591 ) ;
  assign n18617 = ( ~n971 & n6187 ) | ( ~n971 & n18616 ) | ( n6187 & n18616 ) ;
  assign n18615 = n11010 ^ n10885 ^ n2822 ;
  assign n18618 = n18617 ^ n18615 ^ 1'b0 ;
  assign n18619 = ( n5938 & n7708 ) | ( n5938 & ~n11008 ) | ( n7708 & ~n11008 ) ;
  assign n18620 = ( n6178 & n11692 ) | ( n6178 & ~n18619 ) | ( n11692 & ~n18619 ) ;
  assign n18621 = n18620 ^ n14745 ^ 1'b0 ;
  assign n18622 = n447 | n11415 ;
  assign n18623 = n9257 & ~n18622 ;
  assign n18624 = n1469 | n18623 ;
  assign n18625 = n2398 & ~n18624 ;
  assign n18626 = n6007 ^ n4404 ^ 1'b0 ;
  assign n18627 = ~n1828 & n18626 ;
  assign n18628 = ( ~n1879 & n13190 ) | ( ~n1879 & n18627 ) | ( n13190 & n18627 ) ;
  assign n18629 = ~n7563 & n12919 ;
  assign n18630 = n3480 & n18629 ;
  assign n18631 = n15877 ^ n11357 ^ n6431 ;
  assign n18632 = ~n18630 & n18631 ;
  assign n18633 = ( ~n4507 & n15244 ) | ( ~n4507 & n18632 ) | ( n15244 & n18632 ) ;
  assign n18634 = n18628 & ~n18633 ;
  assign n18635 = n18634 ^ n10611 ^ 1'b0 ;
  assign n18636 = n18635 ^ n8726 ^ n2463 ;
  assign n18637 = ~n356 & n6028 ;
  assign n18638 = n15767 | n18637 ;
  assign n18639 = n11655 | n18638 ;
  assign n18640 = n18639 ^ n9924 ^ 1'b0 ;
  assign n18641 = n17582 ^ n4415 ^ 1'b0 ;
  assign n18642 = n6562 | n18641 ;
  assign n18645 = n7700 | n8750 ;
  assign n18643 = n7611 ^ n5907 ^ 1'b0 ;
  assign n18644 = n977 & ~n18643 ;
  assign n18646 = n18645 ^ n18644 ^ 1'b0 ;
  assign n18647 = n1449 | n18646 ;
  assign n18648 = n12802 & n12805 ;
  assign n18649 = n18648 ^ n11647 ^ 1'b0 ;
  assign n18650 = ( n2724 & n4624 ) | ( n2724 & n7376 ) | ( n4624 & n7376 ) ;
  assign n18651 = n18650 ^ n4175 ^ n1461 ;
  assign n18652 = n7870 & ~n18651 ;
  assign n18653 = ( n1237 & n4158 ) | ( n1237 & n6810 ) | ( n4158 & n6810 ) ;
  assign n18654 = ( n3600 & n8558 ) | ( n3600 & ~n11321 ) | ( n8558 & ~n11321 ) ;
  assign n18655 = n18654 ^ n11638 ^ 1'b0 ;
  assign n18656 = ( n11529 & n18653 ) | ( n11529 & n18655 ) | ( n18653 & n18655 ) ;
  assign n18657 = n12351 ^ n5980 ^ 1'b0 ;
  assign n18658 = ~n433 & n1829 ;
  assign n18659 = n18658 ^ n18519 ^ 1'b0 ;
  assign n18660 = n12249 & ~n18659 ;
  assign n18661 = n10364 ^ n5714 ^ n4084 ;
  assign n18662 = n10546 ^ n10530 ^ 1'b0 ;
  assign n18663 = ~n1916 & n18662 ;
  assign n18664 = ( n8770 & ~n18661 ) | ( n8770 & n18663 ) | ( ~n18661 & n18663 ) ;
  assign n18665 = ( n1784 & ~n7633 ) | ( n1784 & n13934 ) | ( ~n7633 & n13934 ) ;
  assign n18666 = n4055 | n18665 ;
  assign n18667 = n18666 ^ n4598 ^ 1'b0 ;
  assign n18668 = n18667 ^ n12850 ^ 1'b0 ;
  assign n18669 = n11504 & n16481 ;
  assign n18670 = n2666 & ~n12461 ;
  assign n18671 = n4770 ^ n2793 ^ 1'b0 ;
  assign n18672 = n7045 & ~n18671 ;
  assign n18673 = ( n11226 & n18670 ) | ( n11226 & n18672 ) | ( n18670 & n18672 ) ;
  assign n18675 = ( n645 & n9476 ) | ( n645 & ~n9909 ) | ( n9476 & ~n9909 ) ;
  assign n18676 = ( ~n4782 & n9482 ) | ( ~n4782 & n18675 ) | ( n9482 & n18675 ) ;
  assign n18674 = n8455 | n13742 ;
  assign n18677 = n18676 ^ n18674 ^ 1'b0 ;
  assign n18678 = n11018 ^ n7706 ^ n6753 ;
  assign n18679 = n18678 ^ n12923 ^ n7200 ;
  assign n18680 = n3897 & n18679 ;
  assign n18681 = n18677 & n18680 ;
  assign n18682 = n14821 ^ n7663 ^ 1'b0 ;
  assign n18683 = ~n18681 & n18682 ;
  assign n18686 = n6712 ^ n4167 ^ x42 ;
  assign n18687 = n7783 & ~n18686 ;
  assign n18684 = ~n3853 & n6466 ;
  assign n18685 = n9720 & ~n18684 ;
  assign n18688 = n18687 ^ n18685 ^ n10353 ;
  assign n18689 = n18688 ^ n11932 ^ n6471 ;
  assign n18690 = n10685 ^ n1445 ^ 1'b0 ;
  assign n18691 = n7792 & ~n18690 ;
  assign n18692 = n9433 & ~n14799 ;
  assign n18693 = n511 & ~n1690 ;
  assign n18694 = x84 & ~n14540 ;
  assign n18695 = n3156 & n18694 ;
  assign n18696 = n18695 ^ n10152 ^ n7486 ;
  assign n18697 = n18693 | n18696 ;
  assign n18698 = ( n7743 & ~n14507 ) | ( n7743 & n18697 ) | ( ~n14507 & n18697 ) ;
  assign n18699 = n18513 ^ n469 ^ 1'b0 ;
  assign n18700 = n18698 & ~n18699 ;
  assign n18701 = n9667 ^ n5984 ^ 1'b0 ;
  assign n18702 = n718 | n13120 ;
  assign n18703 = n3870 & ~n18702 ;
  assign n18704 = ( ~n1786 & n16356 ) | ( ~n1786 & n18703 ) | ( n16356 & n18703 ) ;
  assign n18705 = n18704 ^ n6959 ^ n2838 ;
  assign n18706 = n18091 ^ n4896 ^ 1'b0 ;
  assign n18707 = n11149 & ~n18418 ;
  assign n18708 = n18707 ^ n17699 ^ 1'b0 ;
  assign n18709 = ( n1953 & n8076 ) | ( n1953 & ~n14547 ) | ( n8076 & ~n14547 ) ;
  assign n18710 = n3161 | n4752 ;
  assign n18711 = n18710 ^ n9217 ^ 1'b0 ;
  assign n18712 = n10819 & ~n18711 ;
  assign n18713 = n18712 ^ n15895 ^ 1'b0 ;
  assign n18714 = n18713 ^ n1062 ^ 1'b0 ;
  assign n18715 = n6731 ^ n3417 ^ n2553 ;
  assign n18716 = n18715 ^ n9935 ^ n1730 ;
  assign n18717 = n16511 & n18716 ;
  assign n18718 = n13312 ^ n273 ^ 1'b0 ;
  assign n18719 = n4032 & ~n18718 ;
  assign n18722 = n8811 ^ n8570 ^ n3776 ;
  assign n18720 = n13201 ^ n518 ^ 1'b0 ;
  assign n18721 = n436 | n18720 ;
  assign n18723 = n18722 ^ n18721 ^ n914 ;
  assign n18724 = n14820 ^ n1180 ^ 1'b0 ;
  assign n18725 = n1846 & ~n18724 ;
  assign n18732 = n1121 & n3144 ;
  assign n18733 = n3324 & ~n13063 ;
  assign n18734 = n18732 & n18733 ;
  assign n18726 = x252 & n819 ;
  assign n18727 = n18726 ^ x111 ^ 1'b0 ;
  assign n18728 = ( x232 & ~n10019 ) | ( x232 & n18727 ) | ( ~n10019 & n18727 ) ;
  assign n18729 = n18728 ^ n12215 ^ 1'b0 ;
  assign n18730 = n8072 & n18729 ;
  assign n18731 = n8357 & n18730 ;
  assign n18735 = n18734 ^ n18731 ^ 1'b0 ;
  assign n18737 = ( n1319 & n8937 ) | ( n1319 & n9696 ) | ( n8937 & n9696 ) ;
  assign n18736 = n1034 ^ n767 ^ 1'b0 ;
  assign n18738 = n18737 ^ n18736 ^ n6776 ;
  assign n18739 = n3898 ^ n3885 ^ 1'b0 ;
  assign n18740 = n12917 ^ n3648 ^ 1'b0 ;
  assign n18741 = ~n12035 & n18740 ;
  assign n18742 = x88 & ~n18715 ;
  assign n18743 = n12486 ^ n1122 ^ 1'b0 ;
  assign n18746 = ( n885 & ~n4554 ) | ( n885 & n5902 ) | ( ~n4554 & n5902 ) ;
  assign n18747 = n18746 ^ n6877 ^ n2588 ;
  assign n18744 = n14468 ^ n12624 ^ n627 ;
  assign n18745 = n18744 ^ n5732 ^ n4000 ;
  assign n18748 = n18747 ^ n18745 ^ n16140 ;
  assign n18749 = ( n1032 & ~n13878 ) | ( n1032 & n17560 ) | ( ~n13878 & n17560 ) ;
  assign n18750 = n16428 ^ n7641 ^ n5048 ;
  assign n18751 = n853 | n11824 ;
  assign n18752 = ( n508 & n4245 ) | ( n508 & ~n14054 ) | ( n4245 & ~n14054 ) ;
  assign n18753 = ( n6370 & n18751 ) | ( n6370 & n18752 ) | ( n18751 & n18752 ) ;
  assign n18754 = ( n776 & n7314 ) | ( n776 & ~n18753 ) | ( n7314 & ~n18753 ) ;
  assign n18755 = n1221 & n10070 ;
  assign n18756 = n18755 ^ n12390 ^ n785 ;
  assign n18757 = n18756 ^ n1282 ^ 1'b0 ;
  assign n18758 = n18754 & ~n18757 ;
  assign n18759 = ( n2232 & n14116 ) | ( n2232 & n18648 ) | ( n14116 & n18648 ) ;
  assign n18760 = ( n3671 & ~n3889 ) | ( n3671 & n8446 ) | ( ~n3889 & n8446 ) ;
  assign n18761 = n10784 & n18760 ;
  assign n18762 = n17939 ^ n9632 ^ n592 ;
  assign n18763 = n16749 & ~n18762 ;
  assign n18764 = n10827 ^ x193 ^ 1'b0 ;
  assign n18766 = n1893 | n3166 ;
  assign n18767 = n18766 ^ n5472 ^ 1'b0 ;
  assign n18768 = n8301 & ~n18767 ;
  assign n18769 = x144 & n18768 ;
  assign n18765 = ( n3081 & n4584 ) | ( n3081 & ~n4721 ) | ( n4584 & ~n4721 ) ;
  assign n18770 = n18769 ^ n18765 ^ n15812 ;
  assign n18775 = n7834 ^ n2148 ^ 1'b0 ;
  assign n18776 = ( ~n2160 & n17725 ) | ( ~n2160 & n18775 ) | ( n17725 & n18775 ) ;
  assign n18777 = n10162 | n18776 ;
  assign n18778 = n18777 ^ n9599 ^ 1'b0 ;
  assign n18772 = n17611 ^ n16490 ^ n12495 ;
  assign n18773 = n18772 ^ n12222 ^ n5060 ;
  assign n18774 = ~n8692 & n18773 ;
  assign n18779 = n18778 ^ n18774 ^ 1'b0 ;
  assign n18780 = n18779 ^ n5150 ^ n2097 ;
  assign n18771 = n14856 ^ n9052 ^ 1'b0 ;
  assign n18781 = n18780 ^ n18771 ^ n5222 ;
  assign n18782 = n7697 | n9566 ;
  assign n18783 = n18782 ^ n15180 ^ n736 ;
  assign n18784 = ( n1989 & n15423 ) | ( n1989 & n18783 ) | ( n15423 & n18783 ) ;
  assign n18785 = n18784 ^ n4236 ^ 1'b0 ;
  assign n18786 = n10525 & ~n18785 ;
  assign n18787 = n18786 ^ n16089 ^ 1'b0 ;
  assign n18788 = n5939 | n10390 ;
  assign n18789 = n8389 ^ n5881 ^ 1'b0 ;
  assign n18790 = n18789 ^ n13552 ^ 1'b0 ;
  assign n18791 = n5053 | n18790 ;
  assign n18792 = ( n701 & n3633 ) | ( n701 & n4255 ) | ( n3633 & n4255 ) ;
  assign n18793 = ( n8465 & ~n18068 ) | ( n8465 & n18792 ) | ( ~n18068 & n18792 ) ;
  assign n18794 = n9413 & n16559 ;
  assign n18795 = n12874 & n18794 ;
  assign n18796 = n18795 ^ n13482 ^ n10420 ;
  assign n18797 = n10400 ^ n1700 ^ 1'b0 ;
  assign n18798 = n18797 ^ n13760 ^ n4872 ;
  assign n18799 = n7600 & ~n8762 ;
  assign n18800 = n18799 ^ n12959 ^ 1'b0 ;
  assign n18801 = n12537 ^ n11083 ^ n3439 ;
  assign n18802 = n9678 | n17943 ;
  assign n18803 = n18801 & n18802 ;
  assign n18804 = n18800 & ~n18803 ;
  assign n18805 = n18804 ^ n17800 ^ 1'b0 ;
  assign n18806 = x190 & ~n18805 ;
  assign n18811 = n17819 ^ n5976 ^ n1780 ;
  assign n18812 = n3428 & ~n7827 ;
  assign n18813 = ~n18811 & n18812 ;
  assign n18807 = ( n2693 & ~n9063 ) | ( n2693 & n16744 ) | ( ~n9063 & n16744 ) ;
  assign n18808 = n584 & n18807 ;
  assign n18809 = ~n13837 & n18808 ;
  assign n18810 = ( ~n5681 & n13305 ) | ( ~n5681 & n18809 ) | ( n13305 & n18809 ) ;
  assign n18814 = n18813 ^ n18810 ^ 1'b0 ;
  assign n18815 = n11122 ^ n3456 ^ n511 ;
  assign n18816 = n2933 & n18815 ;
  assign n18817 = ~n260 & n10835 ;
  assign n18819 = n12460 ^ n6061 ^ n3431 ;
  assign n18818 = ( n1657 & n7961 ) | ( n1657 & n9369 ) | ( n7961 & n9369 ) ;
  assign n18820 = n18819 ^ n18818 ^ 1'b0 ;
  assign n18821 = n17814 ^ n8168 ^ 1'b0 ;
  assign n18822 = ( n7889 & n8864 ) | ( n7889 & n18821 ) | ( n8864 & n18821 ) ;
  assign n18823 = n11413 ^ n5595 ^ n2957 ;
  assign n18824 = n18823 ^ n16664 ^ n12179 ;
  assign n18825 = n3834 & n18663 ;
  assign n18827 = ( n2970 & n4822 ) | ( n2970 & n7906 ) | ( n4822 & n7906 ) ;
  assign n18826 = n4381 & ~n13314 ;
  assign n18828 = n18827 ^ n18826 ^ n18588 ;
  assign n18829 = n11366 ^ x37 ^ 1'b0 ;
  assign n18830 = n15422 ^ n15182 ^ n10696 ;
  assign n18831 = n16125 & n18830 ;
  assign n18832 = n14744 & n18831 ;
  assign n18833 = n18829 | n18832 ;
  assign n18834 = n1408 & ~n18833 ;
  assign n18835 = n12868 ^ n3911 ^ 1'b0 ;
  assign n18836 = n5074 ^ n577 ^ 1'b0 ;
  assign n18837 = n10859 ^ n1030 ^ 1'b0 ;
  assign n18838 = n18836 & n18837 ;
  assign n18839 = ( n7011 & n18835 ) | ( n7011 & n18838 ) | ( n18835 & n18838 ) ;
  assign n18840 = ( n1274 & n6833 ) | ( n1274 & n18839 ) | ( n6833 & n18839 ) ;
  assign n18841 = ( ~n376 & n7928 ) | ( ~n376 & n14123 ) | ( n7928 & n14123 ) ;
  assign n18844 = n6424 ^ n3793 ^ n1569 ;
  assign n18842 = n14288 ^ n13300 ^ n12725 ;
  assign n18843 = n18842 ^ n10797 ^ n7636 ;
  assign n18845 = n18844 ^ n18843 ^ 1'b0 ;
  assign n18846 = ~n3206 & n18845 ;
  assign n18847 = n3255 & n18846 ;
  assign n18848 = ~n18841 & n18847 ;
  assign n18849 = n11725 ^ n10742 ^ 1'b0 ;
  assign n18850 = n5987 & ~n18849 ;
  assign n18851 = n14246 ^ n11432 ^ 1'b0 ;
  assign n18852 = n6439 | n18851 ;
  assign n18853 = n18850 | n18852 ;
  assign n18860 = n10505 & n11354 ;
  assign n18854 = n776 & n1164 ;
  assign n18855 = n1609 & n18854 ;
  assign n18856 = n18855 ^ n7665 ^ n432 ;
  assign n18857 = n862 & ~n9580 ;
  assign n18858 = n18857 ^ n787 ^ 1'b0 ;
  assign n18859 = n18856 & ~n18858 ;
  assign n18861 = n18860 ^ n18859 ^ 1'b0 ;
  assign n18862 = n7779 & ~n18861 ;
  assign n18863 = n6214 & n18862 ;
  assign n18864 = ( n2948 & n18853 ) | ( n2948 & ~n18863 ) | ( n18853 & ~n18863 ) ;
  assign n18865 = ( n1162 & ~n9746 ) | ( n1162 & n16364 ) | ( ~n9746 & n16364 ) ;
  assign n18866 = n18865 ^ n18772 ^ 1'b0 ;
  assign n18867 = ~n2482 & n18866 ;
  assign n18868 = ( ~n2176 & n11937 ) | ( ~n2176 & n18867 ) | ( n11937 & n18867 ) ;
  assign n18869 = ( n7301 & ~n11229 ) | ( n7301 & n18868 ) | ( ~n11229 & n18868 ) ;
  assign n18874 = n5769 ^ n3658 ^ n2522 ;
  assign n18875 = n18874 ^ n1680 ^ n317 ;
  assign n18870 = n8130 ^ n3125 ^ n2776 ;
  assign n18871 = n3828 & n6933 ;
  assign n18872 = ~n8891 & n18871 ;
  assign n18873 = n18870 & ~n18872 ;
  assign n18876 = n18875 ^ n18873 ^ 1'b0 ;
  assign n18880 = n17613 ^ n15126 ^ n14665 ;
  assign n18881 = n18880 ^ n5322 ^ 1'b0 ;
  assign n18877 = ( n3379 & ~n5431 ) | ( n3379 & n9131 ) | ( ~n5431 & n9131 ) ;
  assign n18878 = n18877 ^ n15887 ^ n378 ;
  assign n18879 = ~n5645 & n18878 ;
  assign n18882 = n18881 ^ n18879 ^ 1'b0 ;
  assign n18883 = n1922 | n8063 ;
  assign n18884 = n18496 & n18883 ;
  assign n18885 = ~n8435 & n18884 ;
  assign n18886 = n18885 ^ n17777 ^ 1'b0 ;
  assign n18887 = ( ~n946 & n3140 ) | ( ~n946 & n3839 ) | ( n3140 & n3839 ) ;
  assign n18888 = n12863 & ~n18887 ;
  assign n18893 = n11727 & ~n17905 ;
  assign n18894 = n7663 | n18893 ;
  assign n18895 = n18894 ^ n1768 ^ 1'b0 ;
  assign n18896 = n550 | n18895 ;
  assign n18889 = ( ~n4807 & n14374 ) | ( ~n4807 & n14964 ) | ( n14374 & n14964 ) ;
  assign n18890 = n8126 & n18889 ;
  assign n18891 = n18890 ^ n2375 ^ 1'b0 ;
  assign n18892 = n5237 & ~n18891 ;
  assign n18897 = n18896 ^ n18892 ^ n5426 ;
  assign n18898 = n17580 ^ n8302 ^ 1'b0 ;
  assign n18899 = n4922 & ~n15586 ;
  assign n18900 = ~n4922 & n18899 ;
  assign n18901 = ( n4880 & ~n14135 ) | ( n4880 & n18900 ) | ( ~n14135 & n18900 ) ;
  assign n18902 = n9626 ^ n4136 ^ 1'b0 ;
  assign n18903 = n14946 & n16745 ;
  assign n18904 = n18902 & n18903 ;
  assign n18905 = n13552 ^ n10909 ^ n3922 ;
  assign n18906 = n18221 | n18905 ;
  assign n18907 = ( ~n3226 & n4808 ) | ( ~n3226 & n8503 ) | ( n4808 & n8503 ) ;
  assign n18908 = n291 & n3155 ;
  assign n18909 = n18908 ^ n8327 ^ 1'b0 ;
  assign n18910 = ( ~n6218 & n18907 ) | ( ~n6218 & n18909 ) | ( n18907 & n18909 ) ;
  assign n18911 = ( ~n8693 & n12478 ) | ( ~n8693 & n18550 ) | ( n12478 & n18550 ) ;
  assign n18912 = n14860 ^ n12052 ^ n2956 ;
  assign n18913 = n18912 ^ n2424 ^ 1'b0 ;
  assign n18914 = n1087 & ~n18913 ;
  assign n18915 = ~n3838 & n18914 ;
  assign n18916 = n18911 & n18915 ;
  assign n18917 = n4451 & ~n18916 ;
  assign n18918 = n6681 ^ n2196 ^ 1'b0 ;
  assign n18919 = n10846 & n18918 ;
  assign n18920 = n2551 & n11836 ;
  assign n18923 = n16625 ^ n4846 ^ n4819 ;
  assign n18921 = n6681 | n8848 ;
  assign n18922 = n9482 | n18921 ;
  assign n18924 = n18923 ^ n18922 ^ n18000 ;
  assign n18925 = ( n4866 & ~n8777 ) | ( n4866 & n18924 ) | ( ~n8777 & n18924 ) ;
  assign n18926 = ( n8774 & n10761 ) | ( n8774 & n18925 ) | ( n10761 & n18925 ) ;
  assign n18927 = n12958 ^ n4633 ^ n3268 ;
  assign n18928 = ~n978 & n1494 ;
  assign n18929 = n18928 ^ n12015 ^ 1'b0 ;
  assign n18930 = n18929 ^ n2912 ^ 1'b0 ;
  assign n18931 = n7329 & n18930 ;
  assign n18937 = n5551 & n8611 ;
  assign n18932 = n10040 ^ n5786 ^ x32 ;
  assign n18934 = n11617 ^ n557 ^ 1'b0 ;
  assign n18933 = ~n3320 & n13277 ;
  assign n18935 = n18934 ^ n18933 ^ x27 ;
  assign n18936 = ( n15498 & n18932 ) | ( n15498 & ~n18935 ) | ( n18932 & ~n18935 ) ;
  assign n18938 = n18937 ^ n18936 ^ 1'b0 ;
  assign n18939 = ~n268 & n18938 ;
  assign n18940 = ( n11319 & ~n12243 ) | ( n11319 & n18939 ) | ( ~n12243 & n18939 ) ;
  assign n18941 = n1073 & n8276 ;
  assign n18942 = n17764 & n18941 ;
  assign n18943 = n10089 & ~n18942 ;
  assign n18945 = n10206 ^ n2048 ^ 1'b0 ;
  assign n18944 = n9751 ^ n7812 ^ n1208 ;
  assign n18946 = n18945 ^ n18944 ^ n4804 ;
  assign n18947 = n3218 ^ n1103 ^ 1'b0 ;
  assign n18949 = ( n626 & n6520 ) | ( n626 & ~n9338 ) | ( n6520 & ~n9338 ) ;
  assign n18950 = ( n3037 & n14106 ) | ( n3037 & ~n18949 ) | ( n14106 & ~n18949 ) ;
  assign n18948 = n540 & ~n9943 ;
  assign n18951 = n18950 ^ n18948 ^ 1'b0 ;
  assign n18952 = n18951 ^ n12550 ^ n12244 ;
  assign n18953 = n4222 & ~n15752 ;
  assign n18954 = ~n18952 & n18953 ;
  assign n18955 = ( ~n1779 & n12998 ) | ( ~n1779 & n15641 ) | ( n12998 & n15641 ) ;
  assign n18956 = n1078 ^ x26 ^ 1'b0 ;
  assign n18957 = ~n1304 & n18956 ;
  assign n18958 = n7031 | n14454 ;
  assign n18959 = n18958 ^ n17234 ^ 1'b0 ;
  assign n18960 = n18516 | n18959 ;
  assign n18961 = n13165 ^ n5657 ^ 1'b0 ;
  assign n18962 = ( ~n15979 & n18477 ) | ( ~n15979 & n18961 ) | ( n18477 & n18961 ) ;
  assign n18963 = n18962 ^ n11463 ^ n11451 ;
  assign n18964 = n1427 & ~n3653 ;
  assign n18965 = ~n2309 & n7255 ;
  assign n18966 = ( n8306 & ~n18964 ) | ( n8306 & n18965 ) | ( ~n18964 & n18965 ) ;
  assign n18967 = n6076 | n18519 ;
  assign n18968 = n18967 ^ n1776 ^ 1'b0 ;
  assign n18981 = n8407 ^ n4797 ^ n3530 ;
  assign n18982 = n18981 ^ n3273 ^ n1042 ;
  assign n18979 = n7007 ^ n4249 ^ 1'b0 ;
  assign n18975 = n5891 ^ n5657 ^ n2060 ;
  assign n18976 = ~n11521 & n18975 ;
  assign n18977 = ~n7477 & n18976 ;
  assign n18978 = n11858 & ~n18977 ;
  assign n18980 = n18979 ^ n18978 ^ 1'b0 ;
  assign n18972 = n13465 ^ n10410 ^ 1'b0 ;
  assign n18973 = n3752 | n18972 ;
  assign n18970 = ( n6378 & n10043 ) | ( n6378 & ~n10664 ) | ( n10043 & ~n10664 ) ;
  assign n18971 = n18970 ^ n18293 ^ n14022 ;
  assign n18969 = n13991 ^ n6274 ^ 1'b0 ;
  assign n18974 = n18973 ^ n18971 ^ n18969 ;
  assign n18983 = n18982 ^ n18980 ^ n18974 ;
  assign n18984 = ~n720 & n2547 ;
  assign n18985 = n1943 & ~n3427 ;
  assign n18986 = n18985 ^ n6039 ^ 1'b0 ;
  assign n18987 = ~n9360 & n18986 ;
  assign n18988 = n11322 ^ n8139 ^ 1'b0 ;
  assign n18989 = ( n4741 & n5650 ) | ( n4741 & n13047 ) | ( n5650 & n13047 ) ;
  assign n18990 = n4625 & n7386 ;
  assign n18991 = n18990 ^ n16597 ^ 1'b0 ;
  assign n18992 = ( n3583 & n6182 ) | ( n3583 & n7277 ) | ( n6182 & n7277 ) ;
  assign n18993 = ( n7719 & n18991 ) | ( n7719 & n18992 ) | ( n18991 & n18992 ) ;
  assign n18994 = n6193 ^ n5927 ^ 1'b0 ;
  assign n18995 = ~n2191 & n4848 ;
  assign n18998 = n10920 ^ n4075 ^ 1'b0 ;
  assign n18996 = n2899 ^ n2523 ^ 1'b0 ;
  assign n18997 = n12970 & n18996 ;
  assign n18999 = n18998 ^ n18997 ^ 1'b0 ;
  assign n19001 = n9365 & n16548 ;
  assign n19000 = n5726 | n16989 ;
  assign n19002 = n19001 ^ n19000 ^ 1'b0 ;
  assign n19005 = x142 & n8169 ;
  assign n19006 = ~n10483 & n19005 ;
  assign n19003 = n14481 ^ n8801 ^ n7771 ;
  assign n19004 = n18192 & n19003 ;
  assign n19007 = n19006 ^ n19004 ^ n17245 ;
  assign n19008 = n8287 | n15644 ;
  assign n19009 = ( n1165 & n2106 ) | ( n1165 & ~n5232 ) | ( n2106 & ~n5232 ) ;
  assign n19010 = n4556 & ~n19009 ;
  assign n19011 = ~n7511 & n10738 ;
  assign n19012 = n19011 ^ n15716 ^ 1'b0 ;
  assign n19013 = ( n19008 & n19010 ) | ( n19008 & n19012 ) | ( n19010 & n19012 ) ;
  assign n19017 = ( n2157 & ~n2374 ) | ( n2157 & n2752 ) | ( ~n2374 & n2752 ) ;
  assign n19014 = n7989 ^ n6430 ^ 1'b0 ;
  assign n19015 = n9160 & n19014 ;
  assign n19016 = n19015 ^ n854 ^ 1'b0 ;
  assign n19018 = n19017 ^ n19016 ^ n18398 ;
  assign n19021 = n13460 ^ n2763 ^ 1'b0 ;
  assign n19019 = ( n670 & n2682 ) | ( n670 & n3706 ) | ( n2682 & n3706 ) ;
  assign n19020 = n9269 | n19019 ;
  assign n19022 = n19021 ^ n19020 ^ 1'b0 ;
  assign n19023 = ( n1600 & n11322 ) | ( n1600 & ~n14294 ) | ( n11322 & ~n14294 ) ;
  assign n19024 = n19023 ^ n16909 ^ n2355 ;
  assign n19025 = ( n6171 & n19022 ) | ( n6171 & ~n19024 ) | ( n19022 & ~n19024 ) ;
  assign n19026 = n9765 & ~n13352 ;
  assign n19027 = n13481 | n19026 ;
  assign n19028 = ( ~n7374 & n11269 ) | ( ~n7374 & n18679 ) | ( n11269 & n18679 ) ;
  assign n19029 = n19028 ^ n10592 ^ 1'b0 ;
  assign n19030 = n3043 & n19029 ;
  assign n19031 = n18916 & n19030 ;
  assign n19032 = n15290 ^ n11918 ^ n1686 ;
  assign n19033 = ~n4076 & n8744 ;
  assign n19035 = n12739 ^ n5649 ^ n3662 ;
  assign n19036 = n19035 ^ n13096 ^ n12975 ;
  assign n19037 = n19036 ^ n620 ^ 1'b0 ;
  assign n19038 = n19037 ^ n9916 ^ n8401 ;
  assign n19034 = n4128 | n4846 ;
  assign n19039 = n19038 ^ n19034 ^ 1'b0 ;
  assign n19040 = ( n10062 & ~n19033 ) | ( n10062 & n19039 ) | ( ~n19033 & n19039 ) ;
  assign n19041 = ~n3253 & n17554 ;
  assign n19042 = n17351 & n19041 ;
  assign n19044 = n2932 ^ n2409 ^ 1'b0 ;
  assign n19043 = n17799 ^ n4227 ^ n1566 ;
  assign n19045 = n19044 ^ n19043 ^ n9681 ;
  assign n19046 = n19045 ^ n718 ^ 1'b0 ;
  assign n19047 = n19042 | n19046 ;
  assign n19048 = n18682 ^ n14685 ^ n2217 ;
  assign n19049 = ( n1525 & ~n7525 ) | ( n1525 & n7722 ) | ( ~n7525 & n7722 ) ;
  assign n19050 = ~n1626 & n3493 ;
  assign n19051 = n3420 & n19050 ;
  assign n19052 = n19051 ^ n10302 ^ n5928 ;
  assign n19053 = ( ~n11801 & n19049 ) | ( ~n11801 & n19052 ) | ( n19049 & n19052 ) ;
  assign n19054 = n19053 ^ n14009 ^ n9314 ;
  assign n19057 = n5883 & ~n18695 ;
  assign n19058 = n13282 & n19057 ;
  assign n19055 = n3109 & ~n10776 ;
  assign n19056 = n4422 & n19055 ;
  assign n19059 = n19058 ^ n19056 ^ 1'b0 ;
  assign n19060 = ~n1993 & n5760 ;
  assign n19061 = ( n707 & n12015 ) | ( n707 & ~n12265 ) | ( n12015 & ~n12265 ) ;
  assign n19062 = n19061 ^ n432 ^ 1'b0 ;
  assign n19063 = ~n18973 & n19062 ;
  assign n19071 = n13271 ^ n3810 ^ x226 ;
  assign n19069 = n16405 ^ n4354 ^ 1'b0 ;
  assign n19070 = n9717 & n19069 ;
  assign n19072 = n19071 ^ n19070 ^ 1'b0 ;
  assign n19073 = ~n11759 & n19072 ;
  assign n19074 = n19073 ^ n18072 ^ n10516 ;
  assign n19066 = n6601 & n7771 ;
  assign n19067 = n2461 & n19066 ;
  assign n19064 = n7799 ^ n5537 ^ n286 ;
  assign n19065 = n19064 ^ n1100 ^ n721 ;
  assign n19068 = n19067 ^ n19065 ^ 1'b0 ;
  assign n19075 = n19074 ^ n19068 ^ n8723 ;
  assign n19076 = n7707 & n8386 ;
  assign n19077 = ~n701 & n19076 ;
  assign n19078 = ~n8664 & n19077 ;
  assign n19079 = n721 & n16603 ;
  assign n19080 = n5773 ^ n542 ^ 1'b0 ;
  assign n19081 = n19080 ^ n15827 ^ 1'b0 ;
  assign n19082 = n19079 & ~n19081 ;
  assign n19084 = n1766 | n5793 ;
  assign n19083 = n4119 ^ n1295 ^ 1'b0 ;
  assign n19085 = n19084 ^ n19083 ^ 1'b0 ;
  assign n19088 = n3701 ^ n3179 ^ n2121 ;
  assign n19086 = n3841 ^ n3309 ^ n2051 ;
  assign n19087 = ( n6240 & ~n7223 ) | ( n6240 & n19086 ) | ( ~n7223 & n19086 ) ;
  assign n19089 = n19088 ^ n19087 ^ n16281 ;
  assign n19090 = n15169 ^ n7407 ^ n2917 ;
  assign n19091 = n3374 & n16729 ;
  assign n19092 = n6541 & n19091 ;
  assign n19093 = ( n8634 & n17872 ) | ( n8634 & n19092 ) | ( n17872 & n19092 ) ;
  assign n19098 = n18424 ^ n12974 ^ 1'b0 ;
  assign n19094 = n13720 ^ n388 ^ 1'b0 ;
  assign n19095 = n3530 & n19094 ;
  assign n19096 = n19095 ^ n14394 ^ n8640 ;
  assign n19097 = ( n5129 & n13820 ) | ( n5129 & n19096 ) | ( n13820 & n19096 ) ;
  assign n19099 = n19098 ^ n19097 ^ 1'b0 ;
  assign n19100 = n17279 ^ x141 ^ 1'b0 ;
  assign n19101 = n8452 | n19100 ;
  assign n19102 = n1264 & n9341 ;
  assign n19103 = n19101 & n19102 ;
  assign n19104 = n19103 ^ n4593 ^ 1'b0 ;
  assign n19105 = x161 & n4875 ;
  assign n19106 = n7311 ^ n3339 ^ 1'b0 ;
  assign n19107 = n19106 ^ n8994 ^ n8915 ;
  assign n19108 = n12155 ^ n6756 ^ 1'b0 ;
  assign n19109 = n19107 & n19108 ;
  assign n19110 = n577 & n15838 ;
  assign n19111 = n10672 ^ n3437 ^ 1'b0 ;
  assign n19112 = ~n15745 & n19111 ;
  assign n19113 = n15384 | n19112 ;
  assign n19114 = n12419 & ~n19113 ;
  assign n19115 = ~n12073 & n19114 ;
  assign n19116 = n10981 ^ n969 ^ 1'b0 ;
  assign n19117 = n13558 | n19116 ;
  assign n19118 = n18337 | n19117 ;
  assign n19119 = n12586 | n19118 ;
  assign n19120 = n19119 ^ n6874 ^ 1'b0 ;
  assign n19121 = n6509 ^ n541 ^ n360 ;
  assign n19122 = n19121 ^ n18630 ^ n17079 ;
  assign n19123 = ( n9464 & n10123 ) | ( n9464 & n10961 ) | ( n10123 & n10961 ) ;
  assign n19124 = n19123 ^ n15298 ^ 1'b0 ;
  assign n19125 = n19122 | n19124 ;
  assign n19126 = n19125 ^ n12640 ^ n9058 ;
  assign n19130 = n10263 ^ n1667 ^ 1'b0 ;
  assign n19131 = n6907 & ~n19130 ;
  assign n19127 = n10294 ^ n9416 ^ n2979 ;
  assign n19128 = n15540 ^ n5556 ^ 1'b0 ;
  assign n19129 = ( n12000 & n19127 ) | ( n12000 & ~n19128 ) | ( n19127 & ~n19128 ) ;
  assign n19132 = n19131 ^ n19129 ^ 1'b0 ;
  assign n19137 = ( n5935 & n8163 ) | ( n5935 & ~n18784 ) | ( n8163 & ~n18784 ) ;
  assign n19133 = n8548 | n8680 ;
  assign n19134 = ~n6059 & n12746 ;
  assign n19135 = ~n19133 & n19134 ;
  assign n19136 = n13441 | n19135 ;
  assign n19138 = n19137 ^ n19136 ^ 1'b0 ;
  assign n19139 = n4315 ^ n627 ^ 1'b0 ;
  assign n19140 = n3653 & ~n19139 ;
  assign n19141 = n19140 ^ n1666 ^ 1'b0 ;
  assign n19142 = n9503 ^ n5561 ^ 1'b0 ;
  assign n19143 = n19142 ^ n4085 ^ 1'b0 ;
  assign n19144 = n1678 & n19143 ;
  assign n19145 = n19144 ^ n18779 ^ n10492 ;
  assign n19146 = ~n3163 & n19145 ;
  assign n19147 = ~n19141 & n19146 ;
  assign n19148 = ~n2148 & n11817 ;
  assign n19149 = ~n6878 & n19148 ;
  assign n19150 = n19149 ^ n17664 ^ n3811 ;
  assign n19157 = n11848 ^ n2800 ^ 1'b0 ;
  assign n19158 = ( n2201 & n15021 ) | ( n2201 & n19157 ) | ( n15021 & n19157 ) ;
  assign n19151 = n16585 ^ n16449 ^ n3059 ;
  assign n19152 = n19151 ^ n16045 ^ 1'b0 ;
  assign n19153 = n3832 ^ n3042 ^ 1'b0 ;
  assign n19154 = n1589 & n19153 ;
  assign n19155 = ( ~n5277 & n19152 ) | ( ~n5277 & n19154 ) | ( n19152 & n19154 ) ;
  assign n19156 = ~n4494 & n19155 ;
  assign n19159 = n19158 ^ n19156 ^ 1'b0 ;
  assign n19160 = n14781 ^ n5787 ^ 1'b0 ;
  assign n19161 = n15062 & ~n19160 ;
  assign n19162 = ( n9613 & n19159 ) | ( n9613 & ~n19161 ) | ( n19159 & ~n19161 ) ;
  assign n19166 = n3005 & ~n7683 ;
  assign n19167 = ~n8693 & n19166 ;
  assign n19168 = n19167 ^ n6135 ^ 1'b0 ;
  assign n19163 = ( n2271 & n7722 ) | ( n2271 & n14998 ) | ( n7722 & n14998 ) ;
  assign n19164 = n19163 ^ n18695 ^ n9320 ;
  assign n19165 = n9066 & n19164 ;
  assign n19169 = n19168 ^ n19165 ^ 1'b0 ;
  assign n19171 = n11010 ^ n4210 ^ n2006 ;
  assign n19170 = n14178 ^ n3571 ^ 1'b0 ;
  assign n19172 = n19171 ^ n19170 ^ 1'b0 ;
  assign n19173 = n1900 | n11407 ;
  assign n19174 = n19173 ^ n7697 ^ 1'b0 ;
  assign n19175 = ( n7670 & n8006 ) | ( n7670 & n19174 ) | ( n8006 & n19174 ) ;
  assign n19176 = n16316 | n19175 ;
  assign n19177 = n3028 | n17807 ;
  assign n19178 = n4981 & ~n19177 ;
  assign n19179 = n19178 ^ n10980 ^ n5111 ;
  assign n19180 = n7327 & ~n10790 ;
  assign n19181 = n19180 ^ n9226 ^ 1'b0 ;
  assign n19182 = n18024 ^ n16668 ^ 1'b0 ;
  assign n19183 = n14032 ^ n9461 ^ n8840 ;
  assign n19184 = n7722 & ~n19183 ;
  assign n19185 = n19184 ^ n13475 ^ 1'b0 ;
  assign n19186 = n4932 & ~n14795 ;
  assign n19187 = ~n8106 & n19186 ;
  assign n19188 = ~n2191 & n11389 ;
  assign n19189 = n19188 ^ n9409 ^ 1'b0 ;
  assign n19190 = n9597 ^ n4642 ^ n2238 ;
  assign n19191 = ( ~n19187 & n19189 ) | ( ~n19187 & n19190 ) | ( n19189 & n19190 ) ;
  assign n19192 = n19191 ^ n4773 ^ 1'b0 ;
  assign n19193 = n17273 & n19192 ;
  assign n19194 = n19193 ^ n16416 ^ n9447 ;
  assign n19195 = n10639 ^ n5126 ^ n3184 ;
  assign n19196 = ~n10412 & n18215 ;
  assign n19197 = ~n19195 & n19196 ;
  assign n19198 = n19197 ^ n16057 ^ n12086 ;
  assign n19200 = ( ~n8136 & n8807 ) | ( ~n8136 & n9232 ) | ( n8807 & n9232 ) ;
  assign n19199 = n12441 & n13695 ;
  assign n19201 = n19200 ^ n19199 ^ 1'b0 ;
  assign n19202 = ( n660 & n9073 ) | ( n660 & ~n13682 ) | ( n9073 & ~n13682 ) ;
  assign n19203 = n11274 | n19202 ;
  assign n19204 = n19201 | n19203 ;
  assign n19205 = n9297 ^ n7887 ^ n3738 ;
  assign n19206 = n19205 ^ n15985 ^ n9728 ;
  assign n19207 = n16595 ^ n10352 ^ 1'b0 ;
  assign n19209 = ~n9444 & n18684 ;
  assign n19208 = n13586 ^ n2829 ^ 1'b0 ;
  assign n19210 = n19209 ^ n19208 ^ 1'b0 ;
  assign n19211 = n12717 | n19210 ;
  assign n19212 = n6955 | n11851 ;
  assign n19213 = n19212 ^ n11420 ^ n893 ;
  assign n19214 = n19213 ^ n2464 ^ n688 ;
  assign n19215 = n8359 ^ n7023 ^ n291 ;
  assign n19216 = ( n1394 & ~n13794 ) | ( n1394 & n19215 ) | ( ~n13794 & n19215 ) ;
  assign n19217 = n19214 | n19216 ;
  assign n19218 = n19211 & ~n19217 ;
  assign n19219 = ~n517 & n10261 ;
  assign n19220 = ~n5589 & n19219 ;
  assign n19221 = n11590 & ~n19220 ;
  assign n19222 = n8803 & n19221 ;
  assign n19223 = ( n4416 & n13247 ) | ( n4416 & ~n19222 ) | ( n13247 & ~n19222 ) ;
  assign n19224 = n19223 ^ n9678 ^ n7334 ;
  assign n19225 = ~n2633 & n19224 ;
  assign n19226 = ( n1352 & n12697 ) | ( n1352 & n18545 ) | ( n12697 & n18545 ) ;
  assign n19227 = n8966 ^ n6292 ^ 1'b0 ;
  assign n19228 = n11045 | n19227 ;
  assign n19229 = n8180 ^ n2248 ^ 1'b0 ;
  assign n19230 = n19229 ^ n18929 ^ x122 ;
  assign n19231 = n9921 ^ n1032 ^ n539 ;
  assign n19232 = n9160 & n19231 ;
  assign n19233 = x72 | x108 ;
  assign n19234 = ~n6622 & n19233 ;
  assign n19235 = n19234 ^ n9252 ^ 1'b0 ;
  assign n19236 = n4017 ^ n2405 ^ 1'b0 ;
  assign n19237 = ~n19235 & n19236 ;
  assign n19238 = ( n7164 & n10915 ) | ( n7164 & ~n12623 ) | ( n10915 & ~n12623 ) ;
  assign n19239 = ~n17905 & n19238 ;
  assign n19240 = n19239 ^ n18037 ^ 1'b0 ;
  assign n19241 = ( ~n7292 & n19237 ) | ( ~n7292 & n19240 ) | ( n19237 & n19240 ) ;
  assign n19242 = n2273 ^ n947 ^ 1'b0 ;
  assign n19243 = n3266 ^ n2152 ^ 1'b0 ;
  assign n19244 = n19242 & n19243 ;
  assign n19245 = x230 | n2763 ;
  assign n19246 = ( n11683 & n13103 ) | ( n11683 & n19245 ) | ( n13103 & n19245 ) ;
  assign n19247 = ~n1679 & n19246 ;
  assign n19248 = ( n4786 & n10068 ) | ( n4786 & n19247 ) | ( n10068 & n19247 ) ;
  assign n19249 = ( n12578 & ~n19244 ) | ( n12578 & n19248 ) | ( ~n19244 & n19248 ) ;
  assign n19250 = n15164 ^ n14234 ^ n5908 ;
  assign n19254 = n2675 & n6301 ;
  assign n19251 = n4569 ^ n2629 ^ 1'b0 ;
  assign n19252 = n9370 ^ n8122 ^ 1'b0 ;
  assign n19253 = ( ~n7661 & n19251 ) | ( ~n7661 & n19252 ) | ( n19251 & n19252 ) ;
  assign n19255 = n19254 ^ n19253 ^ 1'b0 ;
  assign n19256 = n19250 & n19255 ;
  assign n19257 = n11402 ^ n5132 ^ n2887 ;
  assign n19258 = n11251 ^ n10551 ^ 1'b0 ;
  assign n19259 = ( n1352 & n7490 ) | ( n1352 & ~n11717 ) | ( n7490 & ~n11717 ) ;
  assign n19260 = ( n19257 & n19258 ) | ( n19257 & ~n19259 ) | ( n19258 & ~n19259 ) ;
  assign n19261 = n19260 ^ n6565 ^ n3814 ;
  assign n19262 = n2367 | n12250 ;
  assign n19263 = n15703 ^ n14024 ^ n8205 ;
  assign n19264 = ~n1651 & n8403 ;
  assign n19265 = ~n2610 & n10098 ;
  assign n19266 = n19264 & ~n19265 ;
  assign n19267 = ~n2433 & n19266 ;
  assign n19268 = n7814 ^ n7780 ^ n7696 ;
  assign n19269 = n8291 | n19268 ;
  assign n19270 = n19269 ^ n9180 ^ 1'b0 ;
  assign n19271 = n5193 | n19270 ;
  assign n19272 = ~n11173 & n19271 ;
  assign n19274 = n6967 & ~n12261 ;
  assign n19275 = n19274 ^ n7685 ^ 1'b0 ;
  assign n19273 = n3704 & ~n16715 ;
  assign n19276 = n19275 ^ n19273 ^ 1'b0 ;
  assign n19277 = n19276 ^ n1666 ^ 1'b0 ;
  assign n19278 = n19272 & ~n19277 ;
  assign n19279 = ~n5619 & n9205 ;
  assign n19280 = n19279 ^ n11303 ^ n5108 ;
  assign n19281 = n3603 | n5761 ;
  assign n19282 = n19281 ^ n17239 ^ 1'b0 ;
  assign n19283 = n19280 & ~n19282 ;
  assign n19284 = ( ~n3364 & n11354 ) | ( ~n3364 & n12460 ) | ( n11354 & n12460 ) ;
  assign n19285 = n1271 | n19284 ;
  assign n19286 = n19285 ^ n1669 ^ x7 ;
  assign n19287 = ( n6562 & n12097 ) | ( n6562 & ~n19209 ) | ( n12097 & ~n19209 ) ;
  assign n19288 = n13361 ^ n11756 ^ n6263 ;
  assign n19289 = n14931 ^ n10544 ^ n4018 ;
  assign n19290 = n6400 ^ n4559 ^ n686 ;
  assign n19291 = ( n1673 & ~n2472 ) | ( n1673 & n19290 ) | ( ~n2472 & n19290 ) ;
  assign n19292 = ( n13247 & n19289 ) | ( n13247 & ~n19291 ) | ( n19289 & ~n19291 ) ;
  assign n19293 = ( ~n10788 & n14790 ) | ( ~n10788 & n16779 ) | ( n14790 & n16779 ) ;
  assign n19294 = n15044 ^ n13216 ^ n7429 ;
  assign n19295 = n15974 ^ n6327 ^ n3729 ;
  assign n19296 = ( x234 & n5953 ) | ( x234 & ~n19295 ) | ( n5953 & ~n19295 ) ;
  assign n19297 = ~n2546 & n19296 ;
  assign n19298 = n2861 & n19297 ;
  assign n19299 = n4507 | n19298 ;
  assign n19300 = n13722 ^ n6797 ^ 1'b0 ;
  assign n19301 = n19299 & ~n19300 ;
  assign n19302 = ~n6266 & n8550 ;
  assign n19303 = n19302 ^ n3446 ^ 1'b0 ;
  assign n19304 = n17769 | n19303 ;
  assign n19305 = n19304 ^ n707 ^ 1'b0 ;
  assign n19306 = ( ~n1385 & n2998 ) | ( ~n1385 & n16200 ) | ( n2998 & n16200 ) ;
  assign n19307 = n19306 ^ n4209 ^ n1876 ;
  assign n19308 = n3081 & ~n4904 ;
  assign n19309 = ~n6320 & n19308 ;
  assign n19310 = ( n3620 & n7405 ) | ( n3620 & ~n19309 ) | ( n7405 & ~n19309 ) ;
  assign n19311 = n2609 & n5254 ;
  assign n19312 = n19311 ^ n14202 ^ 1'b0 ;
  assign n19313 = ~n19310 & n19312 ;
  assign n19314 = n3582 & n10854 ;
  assign n19315 = ( n2935 & ~n8342 ) | ( n2935 & n19314 ) | ( ~n8342 & n19314 ) ;
  assign n19316 = ( ~n1275 & n12415 ) | ( ~n1275 & n19315 ) | ( n12415 & n19315 ) ;
  assign n19317 = ~n1736 & n2118 ;
  assign n19318 = n19316 & n19317 ;
  assign n19319 = n17132 ^ n2372 ^ n1570 ;
  assign n19320 = n19319 ^ n13755 ^ n11448 ;
  assign n19321 = n9980 ^ n8561 ^ n5972 ;
  assign n19322 = n7281 ^ n6987 ^ n5645 ;
  assign n19323 = n10081 & ~n19322 ;
  assign n19324 = n11935 ^ n9266 ^ 1'b0 ;
  assign n19325 = n4938 & n19324 ;
  assign n19326 = n19323 & n19325 ;
  assign n19327 = n6300 & ~n10151 ;
  assign n19328 = n18160 & n19327 ;
  assign n19329 = ( n836 & n13422 ) | ( n836 & ~n19328 ) | ( n13422 & ~n19328 ) ;
  assign n19330 = n5509 & n19329 ;
  assign n19331 = n11651 & n19330 ;
  assign n19332 = n721 & ~n16877 ;
  assign n19333 = n19331 & n19332 ;
  assign n19334 = n19333 ^ n2947 ^ n2787 ;
  assign n19335 = n10056 ^ n1254 ^ n541 ;
  assign n19336 = ( n2954 & n9434 ) | ( n2954 & n14219 ) | ( n9434 & n14219 ) ;
  assign n19337 = n1705 & ~n2605 ;
  assign n19338 = ~n19336 & n19337 ;
  assign n19339 = ( n1632 & ~n2095 ) | ( n1632 & n3101 ) | ( ~n2095 & n3101 ) ;
  assign n19340 = n19339 ^ n9013 ^ n8621 ;
  assign n19341 = n12193 ^ n10815 ^ n6150 ;
  assign n19342 = ( n2690 & n4990 ) | ( n2690 & ~n5723 ) | ( n4990 & ~n5723 ) ;
  assign n19343 = ~n3385 & n19342 ;
  assign n19344 = n19341 & n19343 ;
  assign n19345 = n5663 & ~n19344 ;
  assign n19346 = ( ~n5147 & n8266 ) | ( ~n5147 & n8972 ) | ( n8266 & n8972 ) ;
  assign n19347 = x144 & n14191 ;
  assign n19349 = n10815 ^ n5519 ^ 1'b0 ;
  assign n19350 = n2493 & n19349 ;
  assign n19351 = n19350 ^ n2055 ^ 1'b0 ;
  assign n19352 = n591 & ~n19351 ;
  assign n19348 = ( n1034 & ~n12252 ) | ( n1034 & n14459 ) | ( ~n12252 & n14459 ) ;
  assign n19353 = n19352 ^ n19348 ^ n4831 ;
  assign n19354 = ( n19346 & ~n19347 ) | ( n19346 & n19353 ) | ( ~n19347 & n19353 ) ;
  assign n19355 = n19354 ^ n14776 ^ 1'b0 ;
  assign n19356 = ( n19340 & n19345 ) | ( n19340 & ~n19355 ) | ( n19345 & ~n19355 ) ;
  assign n19357 = n10546 ^ n2201 ^ x218 ;
  assign n19360 = n2062 & n7150 ;
  assign n19358 = n9121 ^ n3715 ^ n3579 ;
  assign n19359 = n19358 ^ n8848 ^ 1'b0 ;
  assign n19361 = n19360 ^ n19359 ^ n5693 ;
  assign n19362 = ( ~n18409 & n19357 ) | ( ~n18409 & n19361 ) | ( n19357 & n19361 ) ;
  assign n19363 = n10137 ^ n3151 ^ 1'b0 ;
  assign n19364 = n1122 & ~n19363 ;
  assign n19365 = n14958 & n19364 ;
  assign n19366 = ( n8446 & ~n8536 ) | ( n8446 & n15693 ) | ( ~n8536 & n15693 ) ;
  assign n19367 = n8048 ^ n5176 ^ 1'b0 ;
  assign n19370 = n14476 ^ n1583 ^ n817 ;
  assign n19371 = n19370 ^ n5509 ^ n701 ;
  assign n19368 = n11630 ^ n9232 ^ n8229 ;
  assign n19369 = n19368 ^ n6460 ^ 1'b0 ;
  assign n19372 = n19371 ^ n19369 ^ 1'b0 ;
  assign n19373 = n11073 ^ n8007 ^ n2829 ;
  assign n19374 = n19373 ^ n15235 ^ x211 ;
  assign n19375 = n9177 | n19374 ;
  assign n19376 = n6015 ^ n2204 ^ 1'b0 ;
  assign n19377 = ~n15015 & n19376 ;
  assign n19378 = ~n4138 & n19377 ;
  assign n19379 = n19378 ^ n10450 ^ n2705 ;
  assign n19380 = n19379 ^ n14747 ^ n6058 ;
  assign n19383 = n8111 ^ n4764 ^ n459 ;
  assign n19381 = n11554 ^ n3762 ^ 1'b0 ;
  assign n19382 = n14369 & ~n19381 ;
  assign n19384 = n19383 ^ n19382 ^ 1'b0 ;
  assign n19385 = ~n17219 & n19384 ;
  assign n19386 = n18633 ^ n7139 ^ 1'b0 ;
  assign n19387 = n7129 & n19386 ;
  assign n19388 = n4167 & ~n4697 ;
  assign n19389 = n8699 & n19388 ;
  assign n19390 = n19389 ^ n15529 ^ n394 ;
  assign n19391 = ( n1198 & n4375 ) | ( n1198 & n16603 ) | ( n4375 & n16603 ) ;
  assign n19392 = ( n13974 & ~n18441 ) | ( n13974 & n19391 ) | ( ~n18441 & n19391 ) ;
  assign n19393 = ( n7297 & n12940 ) | ( n7297 & n19392 ) | ( n12940 & n19392 ) ;
  assign n19394 = n19393 ^ n12493 ^ n2405 ;
  assign n19395 = n10077 ^ n5335 ^ n3405 ;
  assign n19396 = n19395 ^ n11312 ^ 1'b0 ;
  assign n19402 = n15426 ^ n13670 ^ n11721 ;
  assign n19397 = n5524 & ~n17180 ;
  assign n19398 = n8651 & n19397 ;
  assign n19399 = x47 & ~n9322 ;
  assign n19400 = n19398 & n19399 ;
  assign n19401 = n11880 | n19400 ;
  assign n19403 = n19402 ^ n19401 ^ 1'b0 ;
  assign n19404 = n19403 ^ n11633 ^ n7627 ;
  assign n19405 = ( n834 & ~n1672 ) | ( n834 & n18537 ) | ( ~n1672 & n18537 ) ;
  assign n19406 = n19404 | n19405 ;
  assign n19407 = n19406 ^ n6815 ^ 1'b0 ;
  assign n19413 = n5268 & ~n16482 ;
  assign n19408 = ( n7926 & n8812 ) | ( n7926 & ~n10116 ) | ( n8812 & ~n10116 ) ;
  assign n19409 = ( n6462 & n14471 ) | ( n6462 & n19408 ) | ( n14471 & n19408 ) ;
  assign n19410 = n11393 & n18569 ;
  assign n19411 = n19410 ^ n4153 ^ 1'b0 ;
  assign n19412 = ( n2096 & n19409 ) | ( n2096 & ~n19411 ) | ( n19409 & ~n19411 ) ;
  assign n19414 = n19413 ^ n19412 ^ n8867 ;
  assign n19415 = ~n8703 & n14106 ;
  assign n19416 = n19415 ^ n16334 ^ 1'b0 ;
  assign n19417 = ~n5231 & n17556 ;
  assign n19418 = n19417 ^ n16330 ^ 1'b0 ;
  assign n19419 = ~n7169 & n19242 ;
  assign n19420 = n1286 & n19419 ;
  assign n19421 = n19420 ^ n4420 ^ 1'b0 ;
  assign n19423 = n5548 ^ n5260 ^ n3946 ;
  assign n19424 = n9275 & ~n10020 ;
  assign n19425 = n2791 | n2979 ;
  assign n19426 = n19424 & n19425 ;
  assign n19427 = ~n19423 & n19426 ;
  assign n19422 = ~n8599 & n14194 ;
  assign n19428 = n19427 ^ n19422 ^ 1'b0 ;
  assign n19429 = ( n2556 & ~n2991 ) | ( n2556 & n19428 ) | ( ~n2991 & n19428 ) ;
  assign n19430 = ( n1703 & ~n7042 ) | ( n1703 & n8606 ) | ( ~n7042 & n8606 ) ;
  assign n19431 = n19430 ^ n7471 ^ 1'b0 ;
  assign n19432 = n6293 & ~n11650 ;
  assign n19433 = n19432 ^ n7766 ^ 1'b0 ;
  assign n19434 = ~n14776 & n19433 ;
  assign n19435 = n19434 ^ n13543 ^ 1'b0 ;
  assign n19436 = n14046 | n19435 ;
  assign n19437 = ( n2517 & n3566 ) | ( n2517 & ~n19436 ) | ( n3566 & ~n19436 ) ;
  assign n19439 = n362 | n3626 ;
  assign n19438 = n3779 | n7262 ;
  assign n19440 = n19439 ^ n19438 ^ 1'b0 ;
  assign n19441 = x116 | n6659 ;
  assign n19442 = ( n2070 & n6892 ) | ( n2070 & ~n7721 ) | ( n6892 & ~n7721 ) ;
  assign n19443 = n11890 | n19442 ;
  assign n19444 = n9418 | n19443 ;
  assign n19445 = n12021 | n19328 ;
  assign n19446 = n3433 & ~n19445 ;
  assign n19447 = n6509 | n19446 ;
  assign n19448 = x174 & ~n18214 ;
  assign n19449 = n19448 ^ n16155 ^ 1'b0 ;
  assign n19450 = n17809 & n19038 ;
  assign n19451 = n7403 ^ n3543 ^ 1'b0 ;
  assign n19452 = n5555 & n19451 ;
  assign n19453 = n2570 | n4520 ;
  assign n19454 = n13502 | n19453 ;
  assign n19455 = ( n11389 & n12799 ) | ( n11389 & ~n19454 ) | ( n12799 & ~n19454 ) ;
  assign n19456 = n19455 ^ n16334 ^ 1'b0 ;
  assign n19457 = n19284 | n19456 ;
  assign n19460 = n18194 ^ n7236 ^ n2064 ;
  assign n19461 = n19460 ^ n8892 ^ 1'b0 ;
  assign n19459 = n6341 ^ n836 ^ 1'b0 ;
  assign n19458 = n12824 ^ n10226 ^ n5921 ;
  assign n19462 = n19461 ^ n19459 ^ n19458 ;
  assign n19463 = n7877 ^ n5866 ^ 1'b0 ;
  assign n19464 = n9096 ^ n2453 ^ 1'b0 ;
  assign n19465 = n19464 ^ n8638 ^ 1'b0 ;
  assign n19466 = n19463 & n19465 ;
  assign n19467 = n13747 ^ n2842 ^ 1'b0 ;
  assign n19468 = ( n3516 & n19466 ) | ( n3516 & ~n19467 ) | ( n19466 & ~n19467 ) ;
  assign n19469 = ( n2572 & ~n7611 ) | ( n2572 & n13035 ) | ( ~n7611 & n13035 ) ;
  assign n19470 = n9664 & ~n19469 ;
  assign n19471 = n19470 ^ n4580 ^ 1'b0 ;
  assign n19472 = ~n5696 & n19471 ;
  assign n19473 = n19472 ^ n18789 ^ n7664 ;
  assign n19474 = ( ~n5818 & n8737 ) | ( ~n5818 & n16417 ) | ( n8737 & n16417 ) ;
  assign n19475 = n19474 ^ n18107 ^ n6147 ;
  assign n19476 = n11028 ^ n773 ^ 1'b0 ;
  assign n19477 = n7229 ^ n4402 ^ 1'b0 ;
  assign n19478 = n16308 ^ x185 ^ 1'b0 ;
  assign n19479 = n2540 & ~n19478 ;
  assign n19480 = ~n19477 & n19479 ;
  assign n19481 = n9281 & n19480 ;
  assign n19482 = n12993 ^ n1572 ^ 1'b0 ;
  assign n19483 = n1524 & n7439 ;
  assign n19484 = ( ~n10376 & n14322 ) | ( ~n10376 & n17811 ) | ( n14322 & n17811 ) ;
  assign n19485 = n2285 & ~n11426 ;
  assign n19486 = n19485 ^ n16369 ^ 1'b0 ;
  assign n19487 = n19486 ^ n2829 ^ 1'b0 ;
  assign n19488 = n7182 & n19487 ;
  assign n19489 = ~n1468 & n11728 ;
  assign n19490 = ( n13591 & n15118 ) | ( n13591 & n19489 ) | ( n15118 & n19489 ) ;
  assign n19493 = ( ~n2046 & n6497 ) | ( ~n2046 & n16844 ) | ( n6497 & n16844 ) ;
  assign n19491 = n10226 ^ n9648 ^ 1'b0 ;
  assign n19492 = ~n9329 & n19491 ;
  assign n19494 = n19493 ^ n19492 ^ 1'b0 ;
  assign n19495 = n18704 ^ n12643 ^ 1'b0 ;
  assign n19503 = ~n1484 & n7098 ;
  assign n19496 = ( n5110 & ~n7119 ) | ( n5110 & n9922 ) | ( ~n7119 & n9922 ) ;
  assign n19497 = n6698 ^ n1642 ^ n387 ;
  assign n19498 = n852 | n19497 ;
  assign n19499 = n3987 & ~n19498 ;
  assign n19500 = n19499 ^ n16776 ^ 1'b0 ;
  assign n19501 = n6649 & n19500 ;
  assign n19502 = ( n13616 & n19496 ) | ( n13616 & n19501 ) | ( n19496 & n19501 ) ;
  assign n19504 = n19503 ^ n19502 ^ 1'b0 ;
  assign n19505 = n3198 & ~n16850 ;
  assign n19506 = n19505 ^ n10907 ^ 1'b0 ;
  assign n19507 = n5581 | n16117 ;
  assign n19508 = n3476 & ~n19507 ;
  assign n19509 = ~n2463 & n19508 ;
  assign n19510 = n4582 | n9552 ;
  assign n19511 = n19510 ^ n5217 ^ 1'b0 ;
  assign n19512 = n19511 ^ n15681 ^ n1282 ;
  assign n19513 = ~n2791 & n13318 ;
  assign n19514 = n4811 ^ n4454 ^ 1'b0 ;
  assign n19515 = ~n2300 & n19514 ;
  assign n19516 = n5257 ^ n2617 ^ 1'b0 ;
  assign n19517 = n19515 & ~n19516 ;
  assign n19518 = n19517 ^ n3145 ^ n2006 ;
  assign n19519 = n16948 ^ n16923 ^ 1'b0 ;
  assign n19520 = n6068 & n16273 ;
  assign n19521 = ( n19518 & n19519 ) | ( n19518 & n19520 ) | ( n19519 & n19520 ) ;
  assign n19522 = n9464 & ~n19521 ;
  assign n19523 = ( n1839 & n11406 ) | ( n1839 & n15276 ) | ( n11406 & n15276 ) ;
  assign n19524 = ~n2146 & n16405 ;
  assign n19525 = n1108 ^ n761 ^ 1'b0 ;
  assign n19526 = ( n7096 & n19524 ) | ( n7096 & n19525 ) | ( n19524 & n19525 ) ;
  assign n19527 = n19526 ^ n12653 ^ n890 ;
  assign n19528 = x108 & ~n19044 ;
  assign n19529 = ( n6934 & ~n16734 ) | ( n6934 & n17344 ) | ( ~n16734 & n17344 ) ;
  assign n19530 = n19528 & n19529 ;
  assign n19531 = ( n19523 & n19527 ) | ( n19523 & ~n19530 ) | ( n19527 & ~n19530 ) ;
  assign n19533 = ( x179 & ~n7103 ) | ( x179 & n7723 ) | ( ~n7103 & n7723 ) ;
  assign n19532 = n8233 & ~n18277 ;
  assign n19534 = n19533 ^ n19532 ^ 1'b0 ;
  assign n19535 = n17983 ^ n5643 ^ 1'b0 ;
  assign n19536 = n7435 & n19535 ;
  assign n19537 = n19536 ^ n5526 ^ 1'b0 ;
  assign n19538 = n721 & ~n6033 ;
  assign n19539 = n9103 & n19538 ;
  assign n19540 = n19539 ^ n10858 ^ n2131 ;
  assign n19541 = n10345 ^ n4605 ^ n1640 ;
  assign n19542 = n1122 & n19541 ;
  assign n19543 = n4772 ^ n4227 ^ n3068 ;
  assign n19544 = n17024 ^ n6275 ^ 1'b0 ;
  assign n19545 = ~n19543 & n19544 ;
  assign n19546 = ( x75 & n19542 ) | ( x75 & n19545 ) | ( n19542 & n19545 ) ;
  assign n19547 = x174 & n19546 ;
  assign n19548 = ~n19540 & n19547 ;
  assign n19549 = ( ~n2417 & n12647 ) | ( ~n2417 & n18940 ) | ( n12647 & n18940 ) ;
  assign n19550 = n6124 ^ n3813 ^ n3482 ;
  assign n19551 = n3441 ^ n2087 ^ 1'b0 ;
  assign n19552 = n8873 | n19551 ;
  assign n19553 = n19552 ^ n6211 ^ 1'b0 ;
  assign n19554 = n12764 & ~n15703 ;
  assign n19555 = n19176 & n19554 ;
  assign n19561 = n1109 | n9672 ;
  assign n19556 = x158 & ~n293 ;
  assign n19557 = n19556 ^ n7853 ^ 1'b0 ;
  assign n19558 = n19557 ^ n12409 ^ n4603 ;
  assign n19559 = n19558 ^ n7065 ^ n5642 ;
  assign n19560 = n19559 ^ n892 ^ 1'b0 ;
  assign n19562 = n19561 ^ n19560 ^ n19441 ;
  assign n19570 = n1723 & n8723 ;
  assign n19567 = ~n871 & n6005 ;
  assign n19568 = n4889 & n19567 ;
  assign n19569 = ~n16244 & n19568 ;
  assign n19571 = n19570 ^ n19569 ^ n11121 ;
  assign n19563 = n2864 & ~n12739 ;
  assign n19564 = n19563 ^ n5791 ^ 1'b0 ;
  assign n19565 = ( ~n1401 & n13589 ) | ( ~n1401 & n19564 ) | ( n13589 & n19564 ) ;
  assign n19566 = n19565 ^ n17073 ^ n526 ;
  assign n19572 = n19571 ^ n19566 ^ n6987 ;
  assign n19573 = n1850 | n4773 ;
  assign n19574 = n19573 ^ n15491 ^ 1'b0 ;
  assign n19575 = n10242 ^ n3329 ^ 1'b0 ;
  assign n19576 = ~n8407 & n19575 ;
  assign n19577 = n17937 ^ n6797 ^ 1'b0 ;
  assign n19578 = n19577 ^ n5535 ^ n1366 ;
  assign n19585 = n17585 ^ n7871 ^ n793 ;
  assign n19584 = n18505 ^ n7625 ^ 1'b0 ;
  assign n19579 = n11978 ^ n9199 ^ 1'b0 ;
  assign n19580 = n7982 & ~n19579 ;
  assign n19581 = ( ~n4858 & n7434 ) | ( ~n4858 & n17998 ) | ( n7434 & n17998 ) ;
  assign n19582 = n19580 & n19581 ;
  assign n19583 = ~n4257 & n19582 ;
  assign n19586 = n19585 ^ n19584 ^ n19583 ;
  assign n19587 = n2362 & n19586 ;
  assign n19588 = n8454 ^ n2850 ^ 1'b0 ;
  assign n19589 = ( ~n1022 & n13460 ) | ( ~n1022 & n14139 ) | ( n13460 & n14139 ) ;
  assign n19590 = n19589 ^ n5546 ^ n3303 ;
  assign n19591 = ~n19588 & n19590 ;
  assign n19592 = n1709 & n12970 ;
  assign n19593 = ~n12970 & n19592 ;
  assign n19594 = ( ~n955 & n6307 ) | ( ~n955 & n19593 ) | ( n6307 & n19593 ) ;
  assign n19595 = n16376 ^ n1064 ^ 1'b0 ;
  assign n19596 = n11166 | n19595 ;
  assign n19597 = n4478 | n19596 ;
  assign n19598 = n6776 & n16811 ;
  assign n19599 = x65 & ~n7674 ;
  assign n19600 = n17154 | n19599 ;
  assign n19601 = n11951 ^ n3174 ^ 1'b0 ;
  assign n19602 = n19601 ^ n5328 ^ n4685 ;
  assign n19603 = n2140 | n14987 ;
  assign n19604 = n19603 ^ n803 ^ 1'b0 ;
  assign n19605 = n19604 ^ n495 ^ 1'b0 ;
  assign n19606 = ( n690 & ~n3481 ) | ( n690 & n19341 ) | ( ~n3481 & n19341 ) ;
  assign n19607 = n19606 ^ n5967 ^ 1'b0 ;
  assign n19608 = ( n19602 & ~n19605 ) | ( n19602 & n19607 ) | ( ~n19605 & n19607 ) ;
  assign n19609 = n18041 ^ n17680 ^ 1'b0 ;
  assign n19616 = n15615 ^ n3034 ^ 1'b0 ;
  assign n19617 = ~n11925 & n19616 ;
  assign n19613 = n4559 ^ n401 ^ 1'b0 ;
  assign n19614 = ~n13031 & n19613 ;
  assign n19610 = n8124 ^ n7384 ^ 1'b0 ;
  assign n19611 = ( x132 & n2579 ) | ( x132 & n19610 ) | ( n2579 & n19610 ) ;
  assign n19612 = n6065 & ~n19611 ;
  assign n19615 = n19614 ^ n19612 ^ 1'b0 ;
  assign n19618 = n19617 ^ n19615 ^ n7347 ;
  assign n19619 = n9437 & n9455 ;
  assign n19620 = n19619 ^ n9238 ^ 1'b0 ;
  assign n19621 = ( n12213 & n14683 ) | ( n12213 & ~n19620 ) | ( n14683 & ~n19620 ) ;
  assign n19622 = ( n14744 & n14849 ) | ( n14744 & n19621 ) | ( n14849 & n19621 ) ;
  assign n19623 = n18048 ^ n10372 ^ n10350 ;
  assign n19625 = n10781 | n15144 ;
  assign n19626 = n16422 & ~n19625 ;
  assign n19624 = ~n3220 & n12468 ;
  assign n19627 = n19626 ^ n19624 ^ n18728 ;
  assign n19641 = ~n4311 & n7829 ;
  assign n19642 = n7749 & n19641 ;
  assign n19643 = ( n2102 & n6940 ) | ( n2102 & ~n19642 ) | ( n6940 & ~n19642 ) ;
  assign n19628 = ( ~n1093 & n1993 ) | ( ~n1093 & n5905 ) | ( n1993 & n5905 ) ;
  assign n19629 = n3462 & n6188 ;
  assign n19630 = n19629 ^ n15946 ^ n10642 ;
  assign n19638 = ( n1255 & n4371 ) | ( n1255 & n8431 ) | ( n4371 & n8431 ) ;
  assign n19633 = n447 | n10215 ;
  assign n19634 = n19633 ^ n5732 ^ 1'b0 ;
  assign n19632 = n3255 & ~n5867 ;
  assign n19635 = n19634 ^ n19632 ^ 1'b0 ;
  assign n19636 = n7175 & n9351 ;
  assign n19637 = n19635 & n19636 ;
  assign n19631 = ( n2978 & ~n9143 ) | ( n2978 & n13581 ) | ( ~n9143 & n13581 ) ;
  assign n19639 = n19638 ^ n19637 ^ n19631 ;
  assign n19640 = ( n19628 & ~n19630 ) | ( n19628 & n19639 ) | ( ~n19630 & n19639 ) ;
  assign n19644 = n19643 ^ n19640 ^ n2472 ;
  assign n19645 = x253 & ~n9332 ;
  assign n19646 = n5217 | n19645 ;
  assign n19647 = n10292 & n19646 ;
  assign n19648 = ( n13388 & n13794 ) | ( n13388 & ~n15615 ) | ( n13794 & ~n15615 ) ;
  assign n19649 = ~n834 & n19648 ;
  assign n19650 = ~n19647 & n19649 ;
  assign n19651 = ~n2343 & n17392 ;
  assign n19652 = ( n1219 & n2716 ) | ( n1219 & ~n6334 ) | ( n2716 & ~n6334 ) ;
  assign n19653 = n19652 ^ n8066 ^ 1'b0 ;
  assign n19654 = n14536 | n19653 ;
  assign n19656 = ( n538 & n9383 ) | ( n538 & ~n18611 ) | ( n9383 & ~n18611 ) ;
  assign n19655 = n18478 ^ n7661 ^ 1'b0 ;
  assign n19657 = n19656 ^ n19655 ^ n12422 ;
  assign n19658 = ~n7018 & n10633 ;
  assign n19659 = ( n779 & ~n5896 ) | ( n779 & n19658 ) | ( ~n5896 & n19658 ) ;
  assign n19660 = n9155 ^ x184 ^ 1'b0 ;
  assign n19661 = ~n5253 & n19660 ;
  assign n19662 = ( ~n17765 & n19659 ) | ( ~n17765 & n19661 ) | ( n19659 & n19661 ) ;
  assign n19663 = ( ~n2996 & n4137 ) | ( ~n2996 & n11170 ) | ( n4137 & n11170 ) ;
  assign n19664 = n5623 | n9648 ;
  assign n19665 = n19664 ^ n9336 ^ 1'b0 ;
  assign n19666 = n5116 | n19665 ;
  assign n19667 = n19663 & ~n19666 ;
  assign n19668 = ( n18004 & n19451 ) | ( n18004 & n19667 ) | ( n19451 & n19667 ) ;
  assign n19670 = ( x149 & n1047 ) | ( x149 & n5638 ) | ( n1047 & n5638 ) ;
  assign n19671 = ~n4974 & n7548 ;
  assign n19672 = ~n19670 & n19671 ;
  assign n19669 = ~n3133 & n14444 ;
  assign n19673 = n19672 ^ n19669 ^ 1'b0 ;
  assign n19674 = n9487 ^ n868 ^ 1'b0 ;
  assign n19675 = n19674 ^ n12500 ^ 1'b0 ;
  assign n19676 = n19675 ^ n13021 ^ n10544 ;
  assign n19677 = n12527 ^ x50 ^ 1'b0 ;
  assign n19678 = ( x191 & n1276 ) | ( x191 & ~n7450 ) | ( n1276 & ~n7450 ) ;
  assign n19679 = n5628 & n19678 ;
  assign n19680 = n5838 & n19679 ;
  assign n19681 = n19680 ^ n2937 ^ 1'b0 ;
  assign n19682 = ~n9444 & n16092 ;
  assign n19683 = n19682 ^ n6037 ^ 1'b0 ;
  assign n19684 = ~n14261 & n15021 ;
  assign n19685 = x143 & n13977 ;
  assign n19686 = ( n5947 & ~n7606 ) | ( n5947 & n19685 ) | ( ~n7606 & n19685 ) ;
  assign n19687 = n7663 | n14330 ;
  assign n19688 = n5542 & n19687 ;
  assign n19689 = ~n2293 & n19688 ;
  assign n19690 = n19689 ^ n5803 ^ 1'b0 ;
  assign n19691 = ~n322 & n8534 ;
  assign n19692 = ~n3981 & n19691 ;
  assign n19693 = n19692 ^ n5613 ^ 1'b0 ;
  assign n19694 = n2918 & ~n19693 ;
  assign n19695 = n10426 ^ n5758 ^ 1'b0 ;
  assign n19696 = n1419 & n19695 ;
  assign n19698 = n13027 ^ n655 ^ n391 ;
  assign n19697 = n10538 & ~n13090 ;
  assign n19699 = n19698 ^ n19697 ^ 1'b0 ;
  assign n19700 = ( n1333 & n5919 ) | ( n1333 & ~n8043 ) | ( n5919 & ~n8043 ) ;
  assign n19702 = n14740 ^ n10400 ^ 1'b0 ;
  assign n19703 = ~n4976 & n19702 ;
  assign n19701 = ~n2634 & n10967 ;
  assign n19704 = n19703 ^ n19701 ^ 1'b0 ;
  assign n19705 = n471 & ~n6297 ;
  assign n19706 = n8028 ^ n7224 ^ n853 ;
  assign n19707 = ~n3831 & n19706 ;
  assign n19708 = ~n19705 & n19707 ;
  assign n19709 = ( n261 & n6209 ) | ( n261 & ~n13918 ) | ( n6209 & ~n13918 ) ;
  assign n19710 = n19709 ^ n10472 ^ n3863 ;
  assign n19711 = n19710 ^ n7541 ^ 1'b0 ;
  assign n19713 = ~n1400 & n9387 ;
  assign n19712 = n8962 & ~n15502 ;
  assign n19714 = n19713 ^ n19712 ^ n1714 ;
  assign n19715 = ( n16725 & ~n19711 ) | ( n16725 & n19714 ) | ( ~n19711 & n19714 ) ;
  assign n19717 = ( n8006 & n18310 ) | ( n8006 & n18518 ) | ( n18310 & n18518 ) ;
  assign n19716 = n9386 & ~n15998 ;
  assign n19718 = n19717 ^ n19716 ^ 1'b0 ;
  assign n19719 = n13018 & n18602 ;
  assign n19720 = ~n12085 & n19719 ;
  assign n19721 = n5978 & ~n14029 ;
  assign n19722 = n8859 & n19721 ;
  assign n19723 = n19722 ^ n13084 ^ 1'b0 ;
  assign n19724 = n11312 & n19723 ;
  assign n19725 = n15820 ^ n1731 ^ 1'b0 ;
  assign n19726 = ( n5919 & n13813 ) | ( n5919 & ~n17182 ) | ( n13813 & ~n17182 ) ;
  assign n19727 = n5792 | n8566 ;
  assign n19728 = n7228 & n19727 ;
  assign n19729 = n19728 ^ n16435 ^ 1'b0 ;
  assign n19742 = n4033 & ~n16891 ;
  assign n19739 = ( n3746 & ~n5006 ) | ( n3746 & n9435 ) | ( ~n5006 & n9435 ) ;
  assign n19736 = n7072 ^ n4460 ^ 1'b0 ;
  assign n19737 = n13328 & n19736 ;
  assign n19738 = n19737 ^ n2956 ^ 1'b0 ;
  assign n19740 = n19739 ^ n19738 ^ n1286 ;
  assign n19730 = ( n4067 & ~n11844 ) | ( n4067 & n17012 ) | ( ~n11844 & n17012 ) ;
  assign n19731 = n1666 & n2634 ;
  assign n19732 = n19731 ^ n8138 ^ 1'b0 ;
  assign n19733 = n11933 | n19732 ;
  assign n19734 = n12321 | n19733 ;
  assign n19735 = ~n19730 & n19734 ;
  assign n19741 = n19740 ^ n19735 ^ n5378 ;
  assign n19743 = n19742 ^ n19741 ^ 1'b0 ;
  assign n19744 = n18584 ^ n884 ^ 1'b0 ;
  assign n19745 = n19744 ^ n8375 ^ n5026 ;
  assign n19746 = n11406 ^ n4265 ^ n4083 ;
  assign n19747 = n19746 ^ n16101 ^ n2641 ;
  assign n19749 = n2940 & ~n6141 ;
  assign n19748 = n3353 ^ n407 ^ 1'b0 ;
  assign n19750 = n19749 ^ n19748 ^ n539 ;
  assign n19754 = n18830 ^ n13846 ^ n9151 ;
  assign n19751 = n7457 ^ n4099 ^ n2486 ;
  assign n19752 = n19751 ^ n12550 ^ 1'b0 ;
  assign n19753 = n6025 & n19752 ;
  assign n19755 = n19754 ^ n19753 ^ 1'b0 ;
  assign n19756 = n19750 | n19755 ;
  assign n19757 = ( n5303 & n8282 ) | ( n5303 & ~n8659 ) | ( n8282 & ~n8659 ) ;
  assign n19758 = ( n1494 & n18087 ) | ( n1494 & ~n19757 ) | ( n18087 & ~n19757 ) ;
  assign n19759 = n17520 ^ n12411 ^ n9938 ;
  assign n19760 = n3067 & ~n13215 ;
  assign n19761 = n3272 & ~n4892 ;
  assign n19762 = ~n2884 & n19761 ;
  assign n19763 = n19762 ^ n7077 ^ n573 ;
  assign n19764 = n19763 ^ n7774 ^ 1'b0 ;
  assign n19765 = n19760 & ~n19764 ;
  assign n19766 = n15719 ^ n5106 ^ 1'b0 ;
  assign n19767 = n11800 ^ n4337 ^ 1'b0 ;
  assign n19768 = n19766 & ~n19767 ;
  assign n19769 = ~n6334 & n19768 ;
  assign n19770 = ~n7262 & n19769 ;
  assign n19771 = ( n1884 & n5809 ) | ( n1884 & ~n15211 ) | ( n5809 & ~n15211 ) ;
  assign n19772 = n11286 ^ n1916 ^ 1'b0 ;
  assign n19773 = ~n3615 & n19772 ;
  assign n19774 = n446 & ~n5780 ;
  assign n19775 = n8984 | n9135 ;
  assign n19776 = n3349 | n19775 ;
  assign n19777 = ( n1673 & ~n3010 ) | ( n1673 & n19776 ) | ( ~n3010 & n19776 ) ;
  assign n19778 = n19774 | n19777 ;
  assign n19779 = n8455 ^ n7520 ^ n639 ;
  assign n19780 = ~n12104 & n19779 ;
  assign n19781 = n19780 ^ n2272 ^ n1755 ;
  assign n19782 = ( n3112 & n7531 ) | ( n3112 & n13020 ) | ( n7531 & n13020 ) ;
  assign n19783 = n19782 ^ n13766 ^ n8536 ;
  assign n19784 = n9420 | n15823 ;
  assign n19785 = n19784 ^ n1200 ^ 1'b0 ;
  assign n19786 = ( ~n663 & n2970 ) | ( ~n663 & n10086 ) | ( n2970 & n10086 ) ;
  assign n19787 = n19786 ^ n7014 ^ n2856 ;
  assign n19788 = n1595 & ~n6488 ;
  assign n19789 = ~n19787 & n19788 ;
  assign n19790 = n13521 ^ n7721 ^ 1'b0 ;
  assign n19791 = n10849 ^ n5500 ^ 1'b0 ;
  assign n19792 = ( ~n401 & n18385 ) | ( ~n401 & n19791 ) | ( n18385 & n19791 ) ;
  assign n19793 = ( n9652 & n12099 ) | ( n9652 & n19792 ) | ( n12099 & n19792 ) ;
  assign n19796 = n15121 ^ n14485 ^ n3494 ;
  assign n19794 = n15781 ^ n11087 ^ 1'b0 ;
  assign n19795 = n5244 | n19794 ;
  assign n19797 = n19796 ^ n19795 ^ 1'b0 ;
  assign n19798 = n8051 ^ n4297 ^ 1'b0 ;
  assign n19799 = n2386 | n19798 ;
  assign n19800 = ~n2679 & n19799 ;
  assign n19801 = n2183 & n3097 ;
  assign n19802 = ( n3142 & n8755 ) | ( n3142 & ~n19801 ) | ( n8755 & ~n19801 ) ;
  assign n19803 = n2123 & n3081 ;
  assign n19804 = n19803 ^ n3658 ^ 1'b0 ;
  assign n19805 = x138 & ~n1010 ;
  assign n19806 = n19805 ^ n1262 ^ 1'b0 ;
  assign n19807 = n1763 & ~n19806 ;
  assign n19808 = n19807 ^ n7479 ^ n7057 ;
  assign n19809 = ( n16559 & ~n19804 ) | ( n16559 & n19808 ) | ( ~n19804 & n19808 ) ;
  assign n19810 = ( ~n3589 & n19802 ) | ( ~n3589 & n19809 ) | ( n19802 & n19809 ) ;
  assign n19811 = ( n1156 & n4204 ) | ( n1156 & n4619 ) | ( n4204 & n4619 ) ;
  assign n19812 = n19811 ^ n2195 ^ n1829 ;
  assign n19813 = ( n974 & n3900 ) | ( n974 & ~n19812 ) | ( n3900 & ~n19812 ) ;
  assign n19814 = n4652 & n9144 ;
  assign n19815 = n19814 ^ n4750 ^ 1'b0 ;
  assign n19816 = n18952 & ~n19815 ;
  assign n19817 = n14292 & n19776 ;
  assign n19818 = n2446 & n19817 ;
  assign n19819 = n12511 & ~n19818 ;
  assign n19820 = n19819 ^ n2705 ^ 1'b0 ;
  assign n19821 = n389 & n19820 ;
  assign n19822 = n19821 ^ n9121 ^ 1'b0 ;
  assign n19823 = ( n1853 & ~n2932 ) | ( n1853 & n3236 ) | ( ~n2932 & n3236 ) ;
  assign n19824 = n19823 ^ n12544 ^ 1'b0 ;
  assign n19825 = n19824 ^ n7706 ^ 1'b0 ;
  assign n19826 = n18653 ^ n3200 ^ 1'b0 ;
  assign n19827 = n19825 & ~n19826 ;
  assign n19834 = n7035 ^ n5983 ^ 1'b0 ;
  assign n19835 = n7009 & n19834 ;
  assign n19828 = n8752 ^ n3911 ^ 1'b0 ;
  assign n19829 = ~n18686 & n19828 ;
  assign n19830 = ( n589 & n10277 ) | ( n589 & ~n19829 ) | ( n10277 & ~n19829 ) ;
  assign n19831 = n4553 & ~n19830 ;
  assign n19832 = ( ~n10756 & n11824 ) | ( ~n10756 & n12701 ) | ( n11824 & n12701 ) ;
  assign n19833 = ( ~n9405 & n19831 ) | ( ~n9405 & n19832 ) | ( n19831 & n19832 ) ;
  assign n19836 = n19835 ^ n19833 ^ 1'b0 ;
  assign n19837 = n13969 ^ n5929 ^ 1'b0 ;
  assign n19838 = x198 & ~n19837 ;
  assign n19839 = ~n2520 & n9385 ;
  assign n19840 = n19839 ^ n7316 ^ 1'b0 ;
  assign n19841 = n19838 & ~n19840 ;
  assign n19842 = n19841 ^ n1358 ^ 1'b0 ;
  assign n19843 = ( ~n1997 & n8689 ) | ( ~n1997 & n19842 ) | ( n8689 & n19842 ) ;
  assign n19844 = n11310 ^ n6652 ^ n2764 ;
  assign n19845 = n19844 ^ n19342 ^ n9317 ;
  assign n19846 = n5024 | n8482 ;
  assign n19847 = n1130 & ~n5158 ;
  assign n19848 = ~n2354 & n19847 ;
  assign n19849 = ( n3208 & n7631 ) | ( n3208 & ~n19848 ) | ( n7631 & ~n19848 ) ;
  assign n19850 = ( n15240 & n19846 ) | ( n15240 & n19849 ) | ( n19846 & n19849 ) ;
  assign n19851 = n3007 & ~n10375 ;
  assign n19852 = n293 & n19851 ;
  assign n19853 = n10920 & ~n19852 ;
  assign n19854 = n5513 & n19853 ;
  assign n19855 = n16306 ^ n1659 ^ 1'b0 ;
  assign n19856 = n19855 ^ n1733 ^ 1'b0 ;
  assign n19857 = n19854 | n19856 ;
  assign n19858 = n8883 & ~n15745 ;
  assign n19859 = n12750 ^ n7551 ^ n6815 ;
  assign n19860 = ( n7747 & n19154 ) | ( n7747 & n19859 ) | ( n19154 & n19859 ) ;
  assign n19861 = ( n2149 & n3598 ) | ( n2149 & n18153 ) | ( n3598 & n18153 ) ;
  assign n19862 = n8609 & ~n10055 ;
  assign n19863 = ~n16988 & n19862 ;
  assign n19864 = n17258 ^ n6391 ^ n3611 ;
  assign n19867 = n4904 | n17530 ;
  assign n19868 = n7023 & ~n19867 ;
  assign n19869 = n15121 & ~n19868 ;
  assign n19870 = n19869 ^ n8862 ^ 1'b0 ;
  assign n19865 = n15258 ^ n8380 ^ n6390 ;
  assign n19866 = n6176 & ~n19865 ;
  assign n19871 = n19870 ^ n19866 ^ 1'b0 ;
  assign n19872 = n13956 ^ n8149 ^ 1'b0 ;
  assign n19873 = n6203 ^ n2433 ^ 1'b0 ;
  assign n19874 = n19873 ^ n14191 ^ 1'b0 ;
  assign n19875 = ~n706 & n19874 ;
  assign n19876 = n19875 ^ n15009 ^ n6457 ;
  assign n19877 = ( ~n5359 & n11609 ) | ( ~n5359 & n18008 ) | ( n11609 & n18008 ) ;
  assign n19878 = ( n16306 & n18054 ) | ( n16306 & n19877 ) | ( n18054 & n19877 ) ;
  assign n19879 = n3710 | n3987 ;
  assign n19880 = ~n15024 & n19879 ;
  assign n19881 = n5412 ^ n1088 ^ 1'b0 ;
  assign n19882 = n14665 & n19881 ;
  assign n19883 = n19882 ^ n13557 ^ 1'b0 ;
  assign n19885 = ( n870 & n3809 ) | ( n870 & ~n6226 ) | ( n3809 & ~n6226 ) ;
  assign n19886 = n19885 ^ n13797 ^ n10794 ;
  assign n19884 = ~n1439 & n7220 ;
  assign n19887 = n19886 ^ n19884 ^ 1'b0 ;
  assign n19888 = n5328 ^ n1461 ^ 1'b0 ;
  assign n19889 = n19888 ^ n19390 ^ n15278 ;
  assign n19895 = n15422 ^ n2137 ^ 1'b0 ;
  assign n19890 = n4841 ^ n2255 ^ 1'b0 ;
  assign n19891 = n4937 & n19890 ;
  assign n19892 = n11638 & ~n19891 ;
  assign n19893 = n7293 & n11386 ;
  assign n19894 = n19892 & n19893 ;
  assign n19896 = n19895 ^ n19894 ^ 1'b0 ;
  assign n19897 = n7946 & n19896 ;
  assign n19898 = n17421 ^ n1813 ^ 1'b0 ;
  assign n19899 = n11143 ^ n10267 ^ n1468 ;
  assign n19900 = n2500 | n10397 ;
  assign n19901 = n9275 | n19900 ;
  assign n19902 = n2090 & n19901 ;
  assign n19903 = n17879 ^ x19 ^ 1'b0 ;
  assign n19904 = n3297 ^ n2631 ^ n1346 ;
  assign n19905 = n8350 & n19904 ;
  assign n19906 = n19905 ^ n18784 ^ n15751 ;
  assign n19907 = n11065 ^ n8038 ^ n5544 ;
  assign n19908 = n19312 ^ n15927 ^ n11697 ;
  assign n19909 = ~n7874 & n11305 ;
  assign n19910 = n19909 ^ n10795 ^ 1'b0 ;
  assign n19911 = ( n19907 & ~n19908 ) | ( n19907 & n19910 ) | ( ~n19908 & n19910 ) ;
  assign n19912 = ( ~n391 & n19906 ) | ( ~n391 & n19911 ) | ( n19906 & n19911 ) ;
  assign n19913 = n17528 ^ n1616 ^ 1'b0 ;
  assign n19914 = n19913 ^ n18542 ^ n2205 ;
  assign n19915 = n16274 ^ n11451 ^ n6319 ;
  assign n19916 = ( n10337 & ~n14358 ) | ( n10337 & n19915 ) | ( ~n14358 & n19915 ) ;
  assign n19917 = n3504 ^ n3313 ^ 1'b0 ;
  assign n19918 = n13581 | n19917 ;
  assign n19919 = n17281 & ~n19918 ;
  assign n19920 = n18685 ^ n3838 ^ 1'b0 ;
  assign n19921 = n16925 ^ n16266 ^ n7672 ;
  assign n19922 = n19920 | n19921 ;
  assign n19923 = n19922 ^ n6915 ^ 1'b0 ;
  assign n19924 = ( n2671 & ~n15790 ) | ( n2671 & n19923 ) | ( ~n15790 & n19923 ) ;
  assign n19925 = n4277 | n6324 ;
  assign n19926 = n19925 ^ n9134 ^ 1'b0 ;
  assign n19927 = n19926 ^ n4753 ^ n499 ;
  assign n19928 = n12725 ^ n9670 ^ n2139 ;
  assign n19929 = n5263 & ~n19732 ;
  assign n19930 = n19928 & n19929 ;
  assign n19934 = n9013 ^ n2120 ^ 1'b0 ;
  assign n19931 = ~n3148 & n3699 ;
  assign n19932 = n5970 ^ n3886 ^ n3057 ;
  assign n19933 = ( ~n3948 & n19931 ) | ( ~n3948 & n19932 ) | ( n19931 & n19932 ) ;
  assign n19935 = n19934 ^ n19933 ^ n1914 ;
  assign n19936 = n17361 ^ n8615 ^ n6735 ;
  assign n19937 = n14303 ^ n6631 ^ n4733 ;
  assign n19938 = n4676 ^ n4255 ^ 1'b0 ;
  assign n19939 = ~n4594 & n19938 ;
  assign n19940 = ( n15337 & n19937 ) | ( n15337 & ~n19939 ) | ( n19937 & ~n19939 ) ;
  assign n19941 = n16187 ^ n13716 ^ 1'b0 ;
  assign n19942 = ( n14134 & n15989 ) | ( n14134 & n19941 ) | ( n15989 & n19941 ) ;
  assign n19947 = x29 & n5180 ;
  assign n19948 = n19947 ^ n7809 ^ 1'b0 ;
  assign n19949 = n19948 ^ n14381 ^ n2512 ;
  assign n19944 = ( ~n885 & n1203 ) | ( ~n885 & n4598 ) | ( n1203 & n4598 ) ;
  assign n19945 = n19944 ^ n6099 ^ n5616 ;
  assign n19946 = n19945 ^ n8929 ^ 1'b0 ;
  assign n19943 = ~n5126 & n19400 ;
  assign n19950 = n19949 ^ n19946 ^ n19943 ;
  assign n19955 = n7007 ^ n3677 ^ 1'b0 ;
  assign n19954 = n7318 & n13736 ;
  assign n19951 = n12017 ^ n6735 ^ 1'b0 ;
  assign n19952 = n16604 & n19951 ;
  assign n19953 = n19952 ^ n5628 ^ n4549 ;
  assign n19956 = n19955 ^ n19954 ^ n19953 ;
  assign n19957 = ( n2574 & ~n6332 ) | ( n2574 & n7213 ) | ( ~n6332 & n7213 ) ;
  assign n19958 = n5601 ^ n3111 ^ 1'b0 ;
  assign n19959 = n11937 ^ n5968 ^ 1'b0 ;
  assign n19960 = n15027 | n19959 ;
  assign n19961 = n9869 ^ n1422 ^ 1'b0 ;
  assign n19962 = ( n12487 & ~n14934 ) | ( n12487 & n19961 ) | ( ~n14934 & n19961 ) ;
  assign n19965 = n971 & n9023 ;
  assign n19966 = ~n3351 & n19965 ;
  assign n19963 = n1638 & ~n10259 ;
  assign n19964 = n19963 ^ n7211 ^ 1'b0 ;
  assign n19967 = n19966 ^ n19964 ^ 1'b0 ;
  assign n19969 = n16393 ^ n502 ^ 1'b0 ;
  assign n19968 = n2540 & n12511 ;
  assign n19970 = n19969 ^ n19968 ^ 1'b0 ;
  assign n19971 = n19970 ^ n18237 ^ n14250 ;
  assign n19972 = n13534 ^ n5738 ^ 1'b0 ;
  assign n19973 = n19972 ^ n11192 ^ n4089 ;
  assign n19974 = n19849 & ~n19973 ;
  assign n19975 = n18195 & n19974 ;
  assign n19976 = ( ~n3487 & n12239 ) | ( ~n3487 & n18382 ) | ( n12239 & n18382 ) ;
  assign n19977 = n1733 & ~n13388 ;
  assign n19978 = ~n19976 & n19977 ;
  assign n19979 = n10785 & ~n15562 ;
  assign n19980 = n16494 ^ n12147 ^ n4617 ;
  assign n19981 = n19980 ^ n8138 ^ 1'b0 ;
  assign n19982 = n5855 & n19981 ;
  assign n19983 = n19982 ^ n3155 ^ 1'b0 ;
  assign n19984 = ( n435 & ~n2130 ) | ( n435 & n5939 ) | ( ~n2130 & n5939 ) ;
  assign n19985 = ~n1184 & n19984 ;
  assign n19986 = n7022 & n19985 ;
  assign n19987 = n2733 | n19986 ;
  assign n19988 = n17051 ^ n16815 ^ 1'b0 ;
  assign n19989 = n11885 | n19988 ;
  assign n19990 = n19989 ^ n4960 ^ 1'b0 ;
  assign n19991 = ( ~n7234 & n8538 ) | ( ~n7234 & n18964 ) | ( n8538 & n18964 ) ;
  assign n19992 = n19991 ^ n3793 ^ 1'b0 ;
  assign n19994 = n7184 | n17043 ;
  assign n19995 = n19994 ^ n10550 ^ 1'b0 ;
  assign n19993 = ~n4393 & n7625 ;
  assign n19996 = n19995 ^ n19993 ^ 1'b0 ;
  assign n19997 = ~n19992 & n19996 ;
  assign n19999 = n10553 | n18775 ;
  assign n20000 = n19999 ^ n13087 ^ 1'b0 ;
  assign n20001 = n20000 ^ n910 ^ 1'b0 ;
  assign n19998 = ~n6095 & n11559 ;
  assign n20002 = n20001 ^ n19998 ^ 1'b0 ;
  assign n20003 = n5029 & n7418 ;
  assign n20004 = n15486 | n20003 ;
  assign n20005 = ( ~n13837 & n18048 ) | ( ~n13837 & n18442 ) | ( n18048 & n18442 ) ;
  assign n20006 = n13292 & ~n14272 ;
  assign n20007 = n20006 ^ n10505 ^ 1'b0 ;
  assign n20017 = n2304 & ~n3983 ;
  assign n20018 = n1612 & ~n20017 ;
  assign n20019 = n1173 & n20018 ;
  assign n20015 = n8349 ^ n2012 ^ 1'b0 ;
  assign n20012 = n491 | n10579 ;
  assign n20013 = n20012 ^ n6032 ^ 1'b0 ;
  assign n20014 = n20013 ^ n15495 ^ n3057 ;
  assign n20016 = n20015 ^ n20014 ^ n8574 ;
  assign n20020 = n20019 ^ n20016 ^ 1'b0 ;
  assign n20021 = n10577 & n20020 ;
  assign n20008 = n6448 & n11023 ;
  assign n20009 = n2183 & ~n20008 ;
  assign n20010 = n6143 & n20009 ;
  assign n20011 = x159 & ~n20010 ;
  assign n20022 = n20021 ^ n20011 ^ 1'b0 ;
  assign n20023 = n19796 ^ n4621 ^ 1'b0 ;
  assign n20024 = ( n2183 & ~n3885 ) | ( n2183 & n6249 ) | ( ~n3885 & n6249 ) ;
  assign n20025 = n18093 ^ n1969 ^ 1'b0 ;
  assign n20026 = n7592 & n20025 ;
  assign n20027 = n20026 ^ n13154 ^ n1886 ;
  assign n20028 = n20024 & ~n20027 ;
  assign n20030 = ~n1588 & n5134 ;
  assign n20031 = ~n7763 & n20030 ;
  assign n20032 = n2051 & n9606 ;
  assign n20033 = n20031 & n20032 ;
  assign n20034 = ~n3776 & n20033 ;
  assign n20029 = n5638 & ~n6846 ;
  assign n20035 = n20034 ^ n20029 ^ n12529 ;
  assign n20036 = n20035 ^ n19035 ^ n14509 ;
  assign n20037 = n19815 ^ n13580 ^ 1'b0 ;
  assign n20038 = ~n5300 & n20037 ;
  assign n20039 = n20038 ^ n11380 ^ 1'b0 ;
  assign n20040 = n7144 ^ n5615 ^ 1'b0 ;
  assign n20041 = n20040 ^ n8856 ^ n8063 ;
  assign n20042 = n20039 | n20041 ;
  assign n20043 = n20042 ^ n793 ^ 1'b0 ;
  assign n20044 = n11174 & n20043 ;
  assign n20045 = n20044 ^ n3725 ^ 1'b0 ;
  assign n20046 = n20045 ^ n17018 ^ n6215 ;
  assign n20047 = n5896 ^ n3146 ^ 1'b0 ;
  assign n20048 = ~n6998 & n20047 ;
  assign n20049 = n4974 & n20048 ;
  assign n20050 = n8216 & n9655 ;
  assign n20051 = n7213 ^ n6364 ^ n4585 ;
  assign n20052 = ( n792 & n1965 ) | ( n792 & n8607 ) | ( n1965 & n8607 ) ;
  assign n20053 = ( ~n291 & n20051 ) | ( ~n291 & n20052 ) | ( n20051 & n20052 ) ;
  assign n20054 = n16918 ^ n9456 ^ n2009 ;
  assign n20056 = x80 & ~n2579 ;
  assign n20055 = n17879 ^ n10465 ^ n858 ;
  assign n20057 = n20056 ^ n20055 ^ n9952 ;
  assign n20058 = n20057 ^ n10146 ^ n9505 ;
  assign n20059 = ( n20053 & ~n20054 ) | ( n20053 & n20058 ) | ( ~n20054 & n20058 ) ;
  assign n20060 = n13393 ^ n5475 ^ n3858 ;
  assign n20062 = ( n3633 & n5518 ) | ( n3633 & n5688 ) | ( n5518 & n5688 ) ;
  assign n20061 = n14118 ^ n13726 ^ n898 ;
  assign n20063 = n20062 ^ n20061 ^ n1597 ;
  assign n20064 = n20063 ^ n19980 ^ 1'b0 ;
  assign n20068 = n891 & ~n16234 ;
  assign n20069 = n7690 & n20068 ;
  assign n20066 = ( n393 & ~n1865 ) | ( n393 & n4875 ) | ( ~n1865 & n4875 ) ;
  assign n20065 = n14844 | n18409 ;
  assign n20067 = n20066 ^ n20065 ^ 1'b0 ;
  assign n20070 = n20069 ^ n20067 ^ n15490 ;
  assign n20071 = ( ~n544 & n2538 ) | ( ~n544 & n20070 ) | ( n2538 & n20070 ) ;
  assign n20072 = n4234 & ~n11987 ;
  assign n20073 = ( n2549 & n3294 ) | ( n2549 & ~n5497 ) | ( n3294 & ~n5497 ) ;
  assign n20074 = n20073 ^ n9614 ^ n5359 ;
  assign n20077 = n3325 ^ n1330 ^ 1'b0 ;
  assign n20075 = n7927 | n15668 ;
  assign n20076 = n20075 ^ n12005 ^ 1'b0 ;
  assign n20078 = n20077 ^ n20076 ^ n6800 ;
  assign n20079 = n16364 ^ n9267 ^ n7425 ;
  assign n20080 = ( ~n5158 & n7678 ) | ( ~n5158 & n20079 ) | ( n7678 & n20079 ) ;
  assign n20081 = ( ~n5193 & n13988 ) | ( ~n5193 & n20080 ) | ( n13988 & n20080 ) ;
  assign n20082 = n20081 ^ x14 ^ 1'b0 ;
  assign n20083 = n20082 ^ n17446 ^ 1'b0 ;
  assign n20084 = n14279 ^ n8198 ^ 1'b0 ;
  assign n20085 = x218 & ~n20084 ;
  assign n20087 = ( n1394 & n5464 ) | ( n1394 & n11884 ) | ( n5464 & n11884 ) ;
  assign n20086 = n19322 ^ n5622 ^ 1'b0 ;
  assign n20088 = n20087 ^ n20086 ^ n13797 ;
  assign n20089 = n20085 & n20088 ;
  assign n20090 = n3187 & n20089 ;
  assign n20091 = ~n2770 & n6113 ;
  assign n20092 = ( ~n1034 & n2514 ) | ( ~n1034 & n12551 ) | ( n2514 & n12551 ) ;
  assign n20093 = n20091 & n20092 ;
  assign n20094 = n2456 & n20093 ;
  assign n20096 = n18033 ^ n11158 ^ 1'b0 ;
  assign n20097 = ~n3801 & n20096 ;
  assign n20098 = n20097 ^ n12510 ^ 1'b0 ;
  assign n20095 = ~n1063 & n16255 ;
  assign n20099 = n20098 ^ n20095 ^ n15117 ;
  assign n20100 = n1865 & ~n3254 ;
  assign n20101 = ( n11275 & ~n12830 ) | ( n11275 & n15767 ) | ( ~n12830 & n15767 ) ;
  assign n20102 = ( n7182 & ~n15742 ) | ( n7182 & n20101 ) | ( ~n15742 & n20101 ) ;
  assign n20103 = n9773 | n20102 ;
  assign n20104 = n20103 ^ n3329 ^ 1'b0 ;
  assign n20106 = ( n466 & n7439 ) | ( n466 & ~n10802 ) | ( n7439 & ~n10802 ) ;
  assign n20105 = n1802 ^ n1164 ^ 1'b0 ;
  assign n20107 = n20106 ^ n20105 ^ n3595 ;
  assign n20108 = n16287 ^ n8168 ^ n1506 ;
  assign n20109 = n20108 ^ n9118 ^ n3983 ;
  assign n20110 = n15466 ^ n10848 ^ n1934 ;
  assign n20111 = n655 | n10300 ;
  assign n20112 = n20111 ^ n18693 ^ 1'b0 ;
  assign n20113 = ~n5561 & n18428 ;
  assign n20114 = ( ~n5587 & n20112 ) | ( ~n5587 & n20113 ) | ( n20112 & n20113 ) ;
  assign n20115 = n3364 | n5310 ;
  assign n20116 = n7463 | n20115 ;
  assign n20117 = ( n1786 & n7094 ) | ( n1786 & ~n10454 ) | ( n7094 & ~n10454 ) ;
  assign n20119 = n4850 ^ n688 ^ 1'b0 ;
  assign n20118 = ~n2127 & n3722 ;
  assign n20120 = n20119 ^ n20118 ^ 1'b0 ;
  assign n20121 = n5836 | n12053 ;
  assign n20122 = n20121 ^ n14374 ^ 1'b0 ;
  assign n20123 = n3255 ^ n1071 ^ x130 ;
  assign n20124 = ( n4583 & ~n15429 ) | ( n4583 & n20123 ) | ( ~n15429 & n20123 ) ;
  assign n20125 = n20124 ^ n1175 ^ n779 ;
  assign n20130 = ~n5815 & n12065 ;
  assign n20126 = n17414 ^ n3097 ^ 1'b0 ;
  assign n20127 = n20126 ^ n9295 ^ n6721 ;
  assign n20128 = n1308 & n13962 ;
  assign n20129 = ~n20127 & n20128 ;
  assign n20131 = n20130 ^ n20129 ^ 1'b0 ;
  assign n20132 = ~n2951 & n12679 ;
  assign n20135 = ( ~n3974 & n5820 ) | ( ~n3974 & n9949 ) | ( n5820 & n9949 ) ;
  assign n20134 = n12701 ^ n11470 ^ n9558 ;
  assign n20136 = n20135 ^ n20134 ^ 1'b0 ;
  assign n20133 = n3359 & ~n11210 ;
  assign n20137 = n20136 ^ n20133 ^ 1'b0 ;
  assign n20142 = n3147 ^ x78 ^ 1'b0 ;
  assign n20143 = n6188 & n20142 ;
  assign n20144 = ( ~n1610 & n12735 ) | ( ~n1610 & n20143 ) | ( n12735 & n20143 ) ;
  assign n20145 = n20144 ^ n8990 ^ 1'b0 ;
  assign n20146 = n5833 & ~n20145 ;
  assign n20147 = n1166 & n9531 ;
  assign n20148 = n8920 | n20147 ;
  assign n20149 = n20146 | n20148 ;
  assign n20140 = n3087 ^ n547 ^ 1'b0 ;
  assign n20141 = n11694 | n20140 ;
  assign n20138 = ( n660 & n1899 ) | ( n660 & n7536 ) | ( n1899 & n7536 ) ;
  assign n20139 = ( n6789 & n8409 ) | ( n6789 & ~n20138 ) | ( n8409 & ~n20138 ) ;
  assign n20150 = n20149 ^ n20141 ^ n20139 ;
  assign n20151 = n13531 ^ n11910 ^ n8251 ;
  assign n20152 = ( n5121 & ~n7266 ) | ( n5121 & n20151 ) | ( ~n7266 & n20151 ) ;
  assign n20153 = n4280 | n20152 ;
  assign n20154 = n20153 ^ n4998 ^ 1'b0 ;
  assign n20155 = ( x94 & n13574 ) | ( x94 & ~n20154 ) | ( n13574 & ~n20154 ) ;
  assign n20156 = n5720 ^ n883 ^ 1'b0 ;
  assign n20157 = x55 & n12422 ;
  assign n20158 = n7160 & n20157 ;
  assign n20159 = n20158 ^ n13427 ^ 1'b0 ;
  assign n20160 = n20156 & ~n20159 ;
  assign n20161 = n10569 ^ n3256 ^ 1'b0 ;
  assign n20162 = n9609 ^ n7968 ^ 1'b0 ;
  assign n20163 = ( n13859 & n14007 ) | ( n13859 & n20162 ) | ( n14007 & n20162 ) ;
  assign n20164 = n12626 & ~n20163 ;
  assign n20165 = n6887 & n20164 ;
  assign n20166 = n5492 | n6802 ;
  assign n20167 = n3871 & ~n20166 ;
  assign n20168 = ( n2475 & ~n6581 ) | ( n2475 & n20167 ) | ( ~n6581 & n20167 ) ;
  assign n20169 = n20168 ^ n7102 ^ 1'b0 ;
  assign n20170 = n20165 | n20169 ;
  assign n20171 = n7896 | n20170 ;
  assign n20172 = ~n270 & n3347 ;
  assign n20173 = n20172 ^ n922 ^ n518 ;
  assign n20178 = ( n13056 & n15154 ) | ( n13056 & n20135 ) | ( n15154 & n20135 ) ;
  assign n20174 = n15612 ^ n6239 ^ n541 ;
  assign n20175 = n19358 ^ n8968 ^ n2158 ;
  assign n20176 = ( n5409 & n9567 ) | ( n5409 & n20175 ) | ( n9567 & n20175 ) ;
  assign n20177 = ( n10207 & n20174 ) | ( n10207 & ~n20176 ) | ( n20174 & ~n20176 ) ;
  assign n20179 = n20178 ^ n20177 ^ 1'b0 ;
  assign n20180 = n11976 ^ n9319 ^ 1'b0 ;
  assign n20181 = n1363 & ~n4356 ;
  assign n20182 = ~n20180 & n20181 ;
  assign n20183 = ( n3955 & ~n7079 ) | ( n3955 & n7168 ) | ( ~n7079 & n7168 ) ;
  assign n20184 = ~n7722 & n15795 ;
  assign n20185 = ~n2978 & n16839 ;
  assign n20186 = n20185 ^ n11370 ^ 1'b0 ;
  assign n20187 = ( n11851 & n19608 ) | ( n11851 & ~n20186 ) | ( n19608 & ~n20186 ) ;
  assign n20188 = n1980 | n6074 ;
  assign n20189 = n20188 ^ n7133 ^ 1'b0 ;
  assign n20190 = n18229 ^ n2544 ^ 1'b0 ;
  assign n20191 = n19125 | n20190 ;
  assign n20192 = n20189 & ~n20191 ;
  assign n20193 = ( n2400 & n4055 ) | ( n2400 & n4475 ) | ( n4055 & n4475 ) ;
  assign n20194 = ( n7598 & ~n9686 ) | ( n7598 & n15438 ) | ( ~n9686 & n15438 ) ;
  assign n20195 = n2729 & ~n3786 ;
  assign n20196 = n17018 & n20195 ;
  assign n20197 = n17461 ^ n7618 ^ n2172 ;
  assign n20198 = n4305 & ~n19982 ;
  assign n20199 = ~n8354 & n9742 ;
  assign n20200 = n852 & n20199 ;
  assign n20201 = x154 & n14889 ;
  assign n20202 = n20201 ^ n6102 ^ 1'b0 ;
  assign n20203 = n4857 ^ n2009 ^ 1'b0 ;
  assign n20204 = n15895 ^ n11514 ^ 1'b0 ;
  assign n20205 = n20203 | n20204 ;
  assign n20206 = n10286 ^ n5933 ^ n2702 ;
  assign n20207 = ~n8937 & n20206 ;
  assign n20208 = n20207 ^ n1680 ^ 1'b0 ;
  assign n20209 = n14684 & ~n20208 ;
  assign n20210 = ( ~n7049 & n20205 ) | ( ~n7049 & n20209 ) | ( n20205 & n20209 ) ;
  assign n20211 = n20210 ^ n15282 ^ 1'b0 ;
  assign n20212 = ( n5723 & n6119 ) | ( n5723 & n15402 ) | ( n6119 & n15402 ) ;
  assign n20216 = n20112 ^ n12654 ^ n10971 ;
  assign n20213 = n15953 | n17033 ;
  assign n20214 = ( n13152 & n19257 ) | ( n13152 & ~n20213 ) | ( n19257 & ~n20213 ) ;
  assign n20215 = n20214 ^ n7396 ^ n2375 ;
  assign n20217 = n20216 ^ n20215 ^ n19949 ;
  assign n20218 = n15115 ^ n14697 ^ n5971 ;
  assign n20220 = n5269 & n6129 ;
  assign n20221 = n20220 ^ n422 ^ 1'b0 ;
  assign n20219 = n1557 & ~n1786 ;
  assign n20222 = n20221 ^ n20219 ^ 1'b0 ;
  assign n20223 = n4375 | n15692 ;
  assign n20224 = n15468 & ~n20223 ;
  assign n20225 = ~n8055 & n19569 ;
  assign n20226 = ( n19539 & n20224 ) | ( n19539 & ~n20225 ) | ( n20224 & ~n20225 ) ;
  assign n20227 = ( n8294 & n20222 ) | ( n8294 & ~n20226 ) | ( n20222 & ~n20226 ) ;
  assign n20228 = n7962 | n20227 ;
  assign n20229 = ~n14748 & n15419 ;
  assign n20230 = n20229 ^ n11861 ^ 1'b0 ;
  assign n20231 = n18821 & n20230 ;
  assign n20232 = ( n2947 & n3540 ) | ( n2947 & n7470 ) | ( n3540 & n7470 ) ;
  assign n20233 = n12140 & ~n12680 ;
  assign n20234 = n20233 ^ n10732 ^ 1'b0 ;
  assign n20235 = n20234 ^ n19163 ^ n7806 ;
  assign n20236 = n1351 & ~n20235 ;
  assign n20239 = n2107 ^ x42 ^ 1'b0 ;
  assign n20240 = ~n2657 & n20239 ;
  assign n20237 = n14233 ^ n9247 ^ n2555 ;
  assign n20238 = ( n4445 & n11104 ) | ( n4445 & ~n20237 ) | ( n11104 & ~n20237 ) ;
  assign n20241 = n20240 ^ n20238 ^ n5209 ;
  assign n20242 = ( n20232 & n20236 ) | ( n20232 & ~n20241 ) | ( n20236 & ~n20241 ) ;
  assign n20243 = ( ~n13426 & n13587 ) | ( ~n13426 & n15234 ) | ( n13587 & n15234 ) ;
  assign n20244 = n877 | n4346 ;
  assign n20245 = n20244 ^ n4220 ^ 1'b0 ;
  assign n20246 = n20245 ^ n3585 ^ x163 ;
  assign n20247 = ( n6318 & n20243 ) | ( n6318 & n20246 ) | ( n20243 & n20246 ) ;
  assign n20248 = ~n5520 & n20247 ;
  assign n20249 = n20248 ^ n7316 ^ 1'b0 ;
  assign n20250 = n20249 ^ n7384 ^ n3017 ;
  assign n20251 = n15584 ^ n7022 ^ n440 ;
  assign n20252 = n10981 | n13247 ;
  assign n20253 = n2021 & ~n20252 ;
  assign n20254 = n10886 ^ n2086 ^ 1'b0 ;
  assign n20255 = n5926 & ~n20254 ;
  assign n20256 = n14845 & n20255 ;
  assign n20257 = ~n8794 & n20256 ;
  assign n20258 = ( n975 & ~n6843 ) | ( n975 & n20257 ) | ( ~n6843 & n20257 ) ;
  assign n20259 = ( x30 & ~n3889 ) | ( x30 & n17154 ) | ( ~n3889 & n17154 ) ;
  assign n20260 = ( n11845 & n20258 ) | ( n11845 & n20259 ) | ( n20258 & n20259 ) ;
  assign n20261 = n20253 | n20260 ;
  assign n20262 = n15573 | n20261 ;
  assign n20272 = n10735 & ~n12409 ;
  assign n20263 = n18093 ^ n14980 ^ x204 ;
  assign n20264 = n2415 & n20263 ;
  assign n20265 = ~n1478 & n20264 ;
  assign n20266 = x20 & ~n7553 ;
  assign n20267 = n20266 ^ n7553 ^ 1'b0 ;
  assign n20268 = n20267 ^ n6403 ^ 1'b0 ;
  assign n20269 = ~n20265 & n20268 ;
  assign n20270 = n20269 ^ x148 ^ 1'b0 ;
  assign n20271 = ~n533 & n20270 ;
  assign n20273 = n20272 ^ n20271 ^ n8766 ;
  assign n20274 = ~n3450 & n14942 ;
  assign n20275 = n3916 & n20274 ;
  assign n20276 = ( ~n3864 & n20273 ) | ( ~n3864 & n20275 ) | ( n20273 & n20275 ) ;
  assign n20277 = n13519 ^ n4857 ^ x149 ;
  assign n20278 = n1966 ^ n1800 ^ 1'b0 ;
  assign n20279 = ~n20277 & n20278 ;
  assign n20280 = n19718 & n20279 ;
  assign n20281 = n6456 & ~n8684 ;
  assign n20282 = ( n4478 & ~n6483 ) | ( n4478 & n10222 ) | ( ~n6483 & n10222 ) ;
  assign n20283 = n1062 | n20282 ;
  assign n20284 = ( n734 & n20281 ) | ( n734 & ~n20283 ) | ( n20281 & ~n20283 ) ;
  assign n20285 = n20284 ^ n6795 ^ n3435 ;
  assign n20286 = ~n539 & n9128 ;
  assign n20287 = ~n1007 & n15845 ;
  assign n20288 = n275 & n20287 ;
  assign n20289 = n20288 ^ n13974 ^ n5357 ;
  assign n20290 = ( n11803 & n14867 ) | ( n11803 & ~n20289 ) | ( n14867 & ~n20289 ) ;
  assign n20291 = n1824 | n17446 ;
  assign n20292 = ( x225 & n4977 ) | ( x225 & ~n8386 ) | ( n4977 & ~n8386 ) ;
  assign n20295 = ~n2666 & n16647 ;
  assign n20296 = n4492 & ~n20295 ;
  assign n20297 = n9363 & n20296 ;
  assign n20293 = n1043 | n4137 ;
  assign n20294 = ~n20114 & n20293 ;
  assign n20298 = n20297 ^ n20294 ^ 1'b0 ;
  assign n20299 = n5351 | n8871 ;
  assign n20300 = n1305 & ~n20299 ;
  assign n20301 = ( n633 & ~n2065 ) | ( n633 & n3049 ) | ( ~n2065 & n3049 ) ;
  assign n20302 = ~n10395 & n20301 ;
  assign n20303 = ( n10873 & n20300 ) | ( n10873 & ~n20302 ) | ( n20300 & ~n20302 ) ;
  assign n20304 = ( x36 & n5354 ) | ( x36 & n8597 ) | ( n5354 & n8597 ) ;
  assign n20305 = ( ~n6251 & n12659 ) | ( ~n6251 & n14950 ) | ( n12659 & n14950 ) ;
  assign n20306 = ( n11819 & ~n13426 ) | ( n11819 & n20305 ) | ( ~n13426 & n20305 ) ;
  assign n20307 = n20304 & ~n20306 ;
  assign n20308 = ( n4596 & ~n6091 ) | ( n4596 & n7680 ) | ( ~n6091 & n7680 ) ;
  assign n20309 = ~n2952 & n20308 ;
  assign n20310 = n20309 ^ n10014 ^ 1'b0 ;
  assign n20311 = ~n8251 & n20310 ;
  assign n20312 = n1896 & ~n5076 ;
  assign n20313 = n20312 ^ n11625 ^ 1'b0 ;
  assign n20314 = n7253 ^ n4010 ^ 1'b0 ;
  assign n20315 = x221 & ~n20314 ;
  assign n20316 = n17244 & n20315 ;
  assign n20317 = n20316 ^ n10310 ^ 1'b0 ;
  assign n20318 = n17909 ^ n1192 ^ n1036 ;
  assign n20319 = n6850 ^ n1374 ^ 1'b0 ;
  assign n20320 = n15914 & n20319 ;
  assign n20321 = ( n18279 & ~n20318 ) | ( n18279 & n20320 ) | ( ~n20318 & n20320 ) ;
  assign n20322 = ~n20317 & n20321 ;
  assign n20323 = ~n20313 & n20322 ;
  assign n20324 = n20311 & ~n20323 ;
  assign n20325 = n20324 ^ n13773 ^ 1'b0 ;
  assign n20326 = n12148 & n20325 ;
  assign n20328 = n1887 & ~n6622 ;
  assign n20329 = n20328 ^ n8177 ^ 1'b0 ;
  assign n20330 = n20329 ^ n2987 ^ 1'b0 ;
  assign n20327 = ~n3562 & n6587 ;
  assign n20331 = n20330 ^ n20327 ^ 1'b0 ;
  assign n20332 = n8614 & n18586 ;
  assign n20333 = ( n6534 & n20331 ) | ( n6534 & ~n20332 ) | ( n20331 & ~n20332 ) ;
  assign n20334 = ( ~n763 & n924 ) | ( ~n763 & n11767 ) | ( n924 & n11767 ) ;
  assign n20335 = n7014 ^ n6574 ^ n3772 ;
  assign n20336 = n20335 ^ n2596 ^ n701 ;
  assign n20337 = ( n7603 & n12623 ) | ( n7603 & ~n20336 ) | ( n12623 & ~n20336 ) ;
  assign n20338 = ( x94 & ~n2707 ) | ( x94 & n3552 ) | ( ~n2707 & n3552 ) ;
  assign n20339 = ( n1542 & ~n9041 ) | ( n1542 & n20338 ) | ( ~n9041 & n20338 ) ;
  assign n20340 = n20339 ^ n9125 ^ 1'b0 ;
  assign n20341 = ( n20334 & ~n20337 ) | ( n20334 & n20340 ) | ( ~n20337 & n20340 ) ;
  assign n20342 = n20341 ^ n15651 ^ n11082 ;
  assign n20343 = ( n493 & n5643 ) | ( n493 & ~n16943 ) | ( n5643 & ~n16943 ) ;
  assign n20344 = n20343 ^ n12032 ^ n2976 ;
  assign n20345 = ( ~n10817 & n15175 ) | ( ~n10817 & n20344 ) | ( n15175 & n20344 ) ;
  assign n20346 = ( n1036 & n9028 ) | ( n1036 & n13058 ) | ( n9028 & n13058 ) ;
  assign n20347 = n8481 ^ n7913 ^ 1'b0 ;
  assign n20348 = ~n20346 & n20347 ;
  assign n20349 = n20348 ^ n953 ^ 1'b0 ;
  assign n20350 = n3467 & ~n12623 ;
  assign n20351 = n20349 & n20350 ;
  assign n20352 = ( n9556 & n13344 ) | ( n9556 & ~n15485 ) | ( n13344 & ~n15485 ) ;
  assign n20353 = ( n1532 & n9538 ) | ( n1532 & n20352 ) | ( n9538 & n20352 ) ;
  assign n20354 = n7588 ^ n6945 ^ n6727 ;
  assign n20355 = ( n4074 & ~n19945 ) | ( n4074 & n20354 ) | ( ~n19945 & n20354 ) ;
  assign n20356 = n9865 | n20355 ;
  assign n20357 = n15008 & ~n20356 ;
  assign n20358 = n20357 ^ n18197 ^ n17671 ;
  assign n20359 = ~n7126 & n12852 ;
  assign n20360 = n4884 & n20359 ;
  assign n20361 = n20360 ^ n8922 ^ n1139 ;
  assign n20362 = n7224 ^ n6783 ^ n1567 ;
  assign n20363 = n6611 ^ n943 ^ 1'b0 ;
  assign n20364 = ~n13976 & n20363 ;
  assign n20365 = n20364 ^ n19952 ^ 1'b0 ;
  assign n20366 = ( n1428 & n3535 ) | ( n1428 & ~n6181 ) | ( n3535 & ~n6181 ) ;
  assign n20367 = ~n15498 & n20366 ;
  assign n20368 = n20367 ^ n12742 ^ 1'b0 ;
  assign n20369 = ( n2073 & ~n7448 ) | ( n2073 & n19049 ) | ( ~n7448 & n19049 ) ;
  assign n20370 = n18101 ^ n7184 ^ 1'b0 ;
  assign n20371 = ~n14788 & n20370 ;
  assign n20372 = ( n6863 & ~n20369 ) | ( n6863 & n20371 ) | ( ~n20369 & n20371 ) ;
  assign n20375 = n10610 ^ n2899 ^ 1'b0 ;
  assign n20376 = n7262 & n20375 ;
  assign n20373 = n12269 ^ n4430 ^ 1'b0 ;
  assign n20374 = n20373 ^ n17331 ^ n10697 ;
  assign n20377 = n20376 ^ n20374 ^ n9909 ;
  assign n20378 = ( x62 & n8393 ) | ( x62 & ~n10913 ) | ( n8393 & ~n10913 ) ;
  assign n20379 = ( n4118 & ~n16552 ) | ( n4118 & n20378 ) | ( ~n16552 & n20378 ) ;
  assign n20380 = n20379 ^ n3909 ^ 1'b0 ;
  assign n20381 = n7947 ^ n1257 ^ 1'b0 ;
  assign n20382 = n8984 ^ n7175 ^ n3760 ;
  assign n20383 = n7726 | n14079 ;
  assign n20384 = n20382 & ~n20383 ;
  assign n20385 = n20384 ^ n10015 ^ 1'b0 ;
  assign n20386 = n16442 ^ n8130 ^ 1'b0 ;
  assign n20387 = ~n10669 & n20386 ;
  assign n20388 = ( ~n1175 & n20385 ) | ( ~n1175 & n20387 ) | ( n20385 & n20387 ) ;
  assign n20389 = ( n11458 & ~n13322 ) | ( n11458 & n16679 ) | ( ~n13322 & n16679 ) ;
  assign n20390 = n20389 ^ n3214 ^ 1'b0 ;
  assign n20391 = n18670 ^ n10732 ^ n3420 ;
  assign n20392 = n20391 ^ n10874 ^ 1'b0 ;
  assign n20395 = ( ~n3791 & n4555 ) | ( ~n3791 & n11190 ) | ( n4555 & n11190 ) ;
  assign n20396 = ( n4094 & n7819 ) | ( n4094 & ~n20395 ) | ( n7819 & ~n20395 ) ;
  assign n20393 = ( n2634 & ~n4283 ) | ( n2634 & n6753 ) | ( ~n4283 & n6753 ) ;
  assign n20394 = ~n17910 & n20393 ;
  assign n20397 = n20396 ^ n20394 ^ n14245 ;
  assign n20399 = n17696 ^ n3358 ^ 1'b0 ;
  assign n20398 = ( n1411 & ~n6036 ) | ( n1411 & n10439 ) | ( ~n6036 & n10439 ) ;
  assign n20400 = n20399 ^ n20398 ^ n11527 ;
  assign n20402 = n2471 ^ x118 ^ 1'b0 ;
  assign n20403 = n3545 & n20402 ;
  assign n20404 = n935 & n7997 ;
  assign n20405 = ( ~n15425 & n20403 ) | ( ~n15425 & n20404 ) | ( n20403 & n20404 ) ;
  assign n20401 = ( n4010 & n6483 ) | ( n4010 & n12047 ) | ( n6483 & n12047 ) ;
  assign n20406 = n20405 ^ n20401 ^ n11105 ;
  assign n20407 = ( ~n2769 & n9349 ) | ( ~n2769 & n15844 ) | ( n9349 & n15844 ) ;
  assign n20408 = n2993 ^ n1470 ^ 1'b0 ;
  assign n20409 = n20408 ^ n2490 ^ 1'b0 ;
  assign n20410 = ~n2076 & n20409 ;
  assign n20411 = ~n10343 & n20410 ;
  assign n20412 = n14840 & n15577 ;
  assign n20413 = n20377 ^ n17443 ^ n14132 ;
  assign n20414 = n3460 & ~n13513 ;
  assign n20415 = ( n1457 & n3354 ) | ( n1457 & ~n20414 ) | ( n3354 & ~n20414 ) ;
  assign n20416 = n20415 ^ n6860 ^ n4302 ;
  assign n20421 = n724 & ~n5864 ;
  assign n20419 = n11803 ^ n6301 ^ n5884 ;
  assign n20420 = n19685 & ~n20419 ;
  assign n20422 = n20421 ^ n20420 ^ 1'b0 ;
  assign n20418 = n3710 & ~n13899 ;
  assign n20423 = n20422 ^ n20418 ^ 1'b0 ;
  assign n20417 = n3559 | n13899 ;
  assign n20424 = n20423 ^ n20417 ^ n2585 ;
  assign n20425 = n19796 ^ n17692 ^ 1'b0 ;
  assign n20426 = n6119 ^ n3164 ^ 1'b0 ;
  assign n20427 = n20426 ^ n9512 ^ 1'b0 ;
  assign n20428 = ~n1575 & n3785 ;
  assign n20429 = n7591 & n20428 ;
  assign n20430 = n10270 ^ n1370 ^ 1'b0 ;
  assign n20431 = n5505 & ~n20430 ;
  assign n20432 = ~n5312 & n9552 ;
  assign n20433 = n9114 & n20432 ;
  assign n20434 = ( n14086 & ~n20431 ) | ( n14086 & n20433 ) | ( ~n20431 & n20433 ) ;
  assign n20435 = ( n5146 & ~n9784 ) | ( n5146 & n20434 ) | ( ~n9784 & n20434 ) ;
  assign n20436 = n3666 ^ n2726 ^ 1'b0 ;
  assign n20437 = n13006 | n14219 ;
  assign n20438 = n1977 & ~n20437 ;
  assign n20439 = ( ~n5346 & n16993 ) | ( ~n5346 & n17076 ) | ( n16993 & n17076 ) ;
  assign n20440 = n20000 ^ n19803 ^ 1'b0 ;
  assign n20441 = ( ~n3243 & n4442 ) | ( ~n3243 & n12249 ) | ( n4442 & n12249 ) ;
  assign n20442 = n960 | n20441 ;
  assign n20443 = ( n2208 & n15131 ) | ( n2208 & n20442 ) | ( n15131 & n20442 ) ;
  assign n20450 = ( n800 & n1848 ) | ( n800 & n6062 ) | ( n1848 & n6062 ) ;
  assign n20448 = n7198 ^ n2317 ^ n1743 ;
  assign n20449 = ( n4374 & n5789 ) | ( n4374 & ~n20448 ) | ( n5789 & ~n20448 ) ;
  assign n20446 = n15692 ^ n1994 ^ 1'b0 ;
  assign n20444 = n12432 ^ n3420 ^ n516 ;
  assign n20445 = n20444 ^ n1475 ^ 1'b0 ;
  assign n20447 = n20446 ^ n20445 ^ 1'b0 ;
  assign n20451 = n20450 ^ n20449 ^ n20447 ;
  assign n20452 = n11344 ^ x164 ^ 1'b0 ;
  assign n20453 = n5446 & ~n20452 ;
  assign n20454 = ( n3672 & ~n4649 ) | ( n3672 & n9720 ) | ( ~n4649 & n9720 ) ;
  assign n20455 = n10933 | n14433 ;
  assign n20456 = n2666 & ~n20455 ;
  assign n20457 = n20454 & n20456 ;
  assign n20458 = n20457 ^ n10491 ^ n2549 ;
  assign n20459 = n20458 ^ n4791 ^ 1'b0 ;
  assign n20460 = ~n1580 & n18894 ;
  assign n20461 = n20460 ^ n17712 ^ n11186 ;
  assign n20462 = n6338 ^ n4686 ^ 1'b0 ;
  assign n20466 = ( n1028 & n2851 ) | ( n1028 & n12392 ) | ( n2851 & n12392 ) ;
  assign n20467 = n1957 | n20466 ;
  assign n20468 = n20467 ^ n5539 ^ 1'b0 ;
  assign n20469 = n18704 | n20468 ;
  assign n20463 = n15035 ^ n8179 ^ 1'b0 ;
  assign n20464 = x163 & ~n20463 ;
  assign n20465 = n20464 ^ n19741 ^ n1449 ;
  assign n20470 = n20469 ^ n20465 ^ n11655 ;
  assign n20471 = n10386 ^ n4209 ^ 1'b0 ;
  assign n20472 = ~n5214 & n14622 ;
  assign n20473 = n20471 & n20472 ;
  assign n20474 = n20473 ^ n14800 ^ 1'b0 ;
  assign n20475 = n1659 & ~n20474 ;
  assign n20476 = n4766 & n12158 ;
  assign n20477 = ( n12916 & n17824 ) | ( n12916 & n20476 ) | ( n17824 & n20476 ) ;
  assign n20478 = ( n9248 & n12463 ) | ( n9248 & n17549 ) | ( n12463 & n17549 ) ;
  assign n20479 = n19477 ^ n12799 ^ x189 ;
  assign n20480 = n4498 | n7087 ;
  assign n20481 = n387 & ~n12141 ;
  assign n20482 = n3487 ^ n3109 ^ 1'b0 ;
  assign n20483 = n2059 | n20482 ;
  assign n20484 = n7341 & ~n15495 ;
  assign n20485 = ~n20483 & n20484 ;
  assign n20487 = n15013 ^ n8403 ^ n3036 ;
  assign n20486 = n1532 & n18844 ;
  assign n20488 = n20487 ^ n20486 ^ n17274 ;
  assign n20489 = n7207 & ~n19247 ;
  assign n20490 = n7870 ^ n7639 ^ n5369 ;
  assign n20491 = n19803 & n20490 ;
  assign n20492 = ( n3263 & n5459 ) | ( n3263 & n20491 ) | ( n5459 & n20491 ) ;
  assign n20494 = n3154 & n4996 ;
  assign n20493 = n15334 ^ n8155 ^ n355 ;
  assign n20495 = n20494 ^ n20493 ^ n3172 ;
  assign n20496 = n3283 | n5667 ;
  assign n20497 = n6705 & ~n20496 ;
  assign n20498 = n10499 | n20497 ;
  assign n20499 = n9551 | n20498 ;
  assign n20500 = ~n20495 & n20499 ;
  assign n20501 = n20500 ^ n14909 ^ n6867 ;
  assign n20502 = ( n2591 & n14479 ) | ( n2591 & n20501 ) | ( n14479 & n20501 ) ;
  assign n20503 = ( ~n13997 & n14090 ) | ( ~n13997 & n17699 ) | ( n14090 & n17699 ) ;
  assign n20504 = ( n1250 & n9694 ) | ( n1250 & ~n14029 ) | ( n9694 & ~n14029 ) ;
  assign n20505 = n5921 & n20504 ;
  assign n20506 = n12881 & n20505 ;
  assign n20507 = ( ~n2036 & n4010 ) | ( ~n2036 & n20506 ) | ( n4010 & n20506 ) ;
  assign n20508 = ~n4634 & n10732 ;
  assign n20509 = n15347 ^ n286 ^ 1'b0 ;
  assign n20510 = n12729 ^ n12607 ^ n5803 ;
  assign n20511 = ~n16011 & n20510 ;
  assign n20512 = ( n20508 & n20509 ) | ( n20508 & ~n20511 ) | ( n20509 & ~n20511 ) ;
  assign n20513 = n1708 | n20512 ;
  assign n20514 = n20513 ^ n5241 ^ 1'b0 ;
  assign n20515 = n18980 ^ n3636 ^ 1'b0 ;
  assign n20516 = n13324 & n20515 ;
  assign n20517 = n15353 & n20516 ;
  assign n20518 = n17644 ^ n12292 ^ n6250 ;
  assign n20519 = n6330 ^ n989 ^ 1'b0 ;
  assign n20520 = ( n1722 & n2556 ) | ( n1722 & ~n8534 ) | ( n2556 & ~n8534 ) ;
  assign n20521 = n7794 | n20520 ;
  assign n20522 = n4804 ^ n3732 ^ 1'b0 ;
  assign n20523 = ( ~n304 & n1020 ) | ( ~n304 & n20522 ) | ( n1020 & n20522 ) ;
  assign n20524 = n20523 ^ n7626 ^ n7311 ;
  assign n20525 = n9362 ^ n6558 ^ 1'b0 ;
  assign n20526 = n18692 & n20525 ;
  assign n20528 = n5165 & n8311 ;
  assign n20527 = n1289 | n9974 ;
  assign n20529 = n20528 ^ n20527 ^ 1'b0 ;
  assign n20530 = n20529 ^ n19663 ^ n1982 ;
  assign n20535 = n10743 ^ n6573 ^ 1'b0 ;
  assign n20536 = x144 | n20535 ;
  assign n20537 = n7399 | n20536 ;
  assign n20531 = ( n663 & n2751 ) | ( n663 & n3441 ) | ( n2751 & n3441 ) ;
  assign n20532 = n20531 ^ n9362 ^ 1'b0 ;
  assign n20533 = n15346 & n20532 ;
  assign n20534 = ~n15147 & n20533 ;
  assign n20538 = n20537 ^ n20534 ^ 1'b0 ;
  assign n20539 = ( n11062 & n15245 ) | ( n11062 & n20538 ) | ( n15245 & n20538 ) ;
  assign n20540 = ( x111 & ~n17023 ) | ( x111 & n18394 ) | ( ~n17023 & n18394 ) ;
  assign n20541 = n9281 & n18907 ;
  assign n20542 = n20541 ^ n15649 ^ 1'b0 ;
  assign n20543 = ( ~n5456 & n20540 ) | ( ~n5456 & n20542 ) | ( n20540 & n20542 ) ;
  assign n20544 = n2889 | n11719 ;
  assign n20545 = ( n3897 & ~n9212 ) | ( n3897 & n12243 ) | ( ~n9212 & n12243 ) ;
  assign n20546 = n8103 ^ n3527 ^ n2107 ;
  assign n20547 = ~n19139 & n20546 ;
  assign n20548 = n1792 & n20547 ;
  assign n20549 = n20033 ^ n8303 ^ 1'b0 ;
  assign n20550 = n4229 ^ n1067 ^ 1'b0 ;
  assign n20551 = n5688 | n20550 ;
  assign n20552 = n1507 ^ n1246 ^ 1'b0 ;
  assign n20553 = ( n10680 & ~n20551 ) | ( n10680 & n20552 ) | ( ~n20551 & n20552 ) ;
  assign n20554 = n20549 & n20553 ;
  assign n20556 = n18934 ^ n11314 ^ n10631 ;
  assign n20555 = n1157 | n8603 ;
  assign n20557 = n20556 ^ n20555 ^ 1'b0 ;
  assign n20558 = n3404 & ~n4333 ;
  assign n20559 = ~n2100 & n20558 ;
  assign n20560 = n19679 & ~n20559 ;
  assign n20561 = n6904 & ~n10996 ;
  assign n20562 = n20561 ^ n1858 ^ 1'b0 ;
  assign n20563 = ( n9527 & n10597 ) | ( n9527 & ~n20562 ) | ( n10597 & ~n20562 ) ;
  assign n20565 = ( n1081 & ~n7795 ) | ( n1081 & n15256 ) | ( ~n7795 & n15256 ) ;
  assign n20564 = n14413 ^ n10520 ^ n8440 ;
  assign n20566 = n20565 ^ n20564 ^ n20207 ;
  assign n20567 = ( x155 & n10739 ) | ( x155 & n12647 ) | ( n10739 & n12647 ) ;
  assign n20568 = n984 & n20567 ;
  assign n20569 = n20566 & n20568 ;
  assign n20570 = ( n5905 & ~n10840 ) | ( n5905 & n11649 ) | ( ~n10840 & n11649 ) ;
  assign n20571 = n16256 ^ n14370 ^ n7833 ;
  assign n20572 = n7323 & ~n20571 ;
  assign n20573 = n3906 & n20572 ;
  assign n20574 = ~n20531 & n20573 ;
  assign n20575 = n1124 & ~n20574 ;
  assign n20576 = n16391 ^ n6061 ^ 1'b0 ;
  assign n20577 = n16209 & n20576 ;
  assign n20578 = n14800 ^ n7453 ^ 1'b0 ;
  assign n20579 = n12780 ^ n12715 ^ n10531 ;
  assign n20580 = n20579 ^ n7819 ^ 1'b0 ;
  assign n20581 = n15319 ^ n3931 ^ 1'b0 ;
  assign n20582 = ( n1790 & n19112 ) | ( n1790 & n20581 ) | ( n19112 & n20581 ) ;
  assign n20583 = n20582 ^ n16784 ^ n986 ;
  assign n20584 = n6300 & n20583 ;
  assign n20585 = n6720 ^ n4104 ^ n1096 ;
  assign n20586 = n8027 & ~n20585 ;
  assign n20587 = n20586 ^ n7419 ^ 1'b0 ;
  assign n20588 = n20587 ^ n17539 ^ n5541 ;
  assign n20589 = ~n10410 & n20588 ;
  assign n20590 = ~n12062 & n20589 ;
  assign n20591 = n8296 ^ n5362 ^ 1'b0 ;
  assign n20592 = n9503 & n20591 ;
  assign n20593 = ( n603 & n14195 ) | ( n603 & n20592 ) | ( n14195 & n20592 ) ;
  assign n20594 = n6301 ^ n5643 ^ 1'b0 ;
  assign n20595 = n20594 ^ n8407 ^ 1'b0 ;
  assign n20596 = n1026 & n20595 ;
  assign n20597 = n20596 ^ n15524 ^ n8425 ;
  assign n20599 = n3403 ^ n2318 ^ n2265 ;
  assign n20600 = n20599 ^ n6649 ^ 1'b0 ;
  assign n20601 = n19873 & n20600 ;
  assign n20598 = n7272 ^ n6317 ^ x64 ;
  assign n20602 = n20601 ^ n20598 ^ n15258 ;
  assign n20603 = ( n562 & n20597 ) | ( n562 & n20602 ) | ( n20597 & n20602 ) ;
  assign n20604 = n8822 ^ n914 ^ 1'b0 ;
  assign n20605 = n7504 | n20604 ;
  assign n20606 = n7618 & ~n20605 ;
  assign n20607 = n4495 & ~n18389 ;
  assign n20608 = n20607 ^ n13969 ^ 1'b0 ;
  assign n20611 = n1624 ^ x206 ^ 1'b0 ;
  assign n20609 = n2445 & n16655 ;
  assign n20610 = n4398 & n20609 ;
  assign n20612 = n20611 ^ n20610 ^ n9218 ;
  assign n20613 = ( n6122 & n6507 ) | ( n6122 & n17330 ) | ( n6507 & n17330 ) ;
  assign n20614 = n20613 ^ n7658 ^ n1388 ;
  assign n20615 = n3861 | n3918 ;
  assign n20616 = n18752 ^ n6326 ^ 1'b0 ;
  assign n20617 = n6418 & ~n20616 ;
  assign n20618 = n20617 ^ n20553 ^ n10269 ;
  assign n20619 = n3916 & ~n9881 ;
  assign n20620 = n4857 & n8233 ;
  assign n20621 = n1378 & n20620 ;
  assign n20622 = ( ~n600 & n5854 ) | ( ~n600 & n13989 ) | ( n5854 & n13989 ) ;
  assign n20623 = n15876 ^ n4621 ^ n3123 ;
  assign n20624 = ~n17940 & n20623 ;
  assign n20625 = ~n20622 & n20624 ;
  assign n20626 = n20621 | n20625 ;
  assign n20627 = n20626 ^ n4609 ^ 1'b0 ;
  assign n20628 = ~n20619 & n20627 ;
  assign n20629 = n14583 ^ n9867 ^ n4539 ;
  assign n20631 = n4477 ^ n2188 ^ 1'b0 ;
  assign n20632 = n5314 & n20631 ;
  assign n20630 = x193 & n4046 ;
  assign n20633 = n20632 ^ n20630 ^ 1'b0 ;
  assign n20634 = ( ~n3914 & n4862 ) | ( ~n3914 & n6464 ) | ( n4862 & n6464 ) ;
  assign n20635 = ( n2776 & n20633 ) | ( n2776 & n20634 ) | ( n20633 & n20634 ) ;
  assign n20636 = n15571 ^ n13722 ^ 1'b0 ;
  assign n20637 = n5600 & n20636 ;
  assign n20638 = n13985 & n16329 ;
  assign n20639 = n20638 ^ n10921 ^ 1'b0 ;
  assign n20640 = ~n991 & n20639 ;
  assign n20641 = n12064 ^ n10765 ^ 1'b0 ;
  assign n20642 = x13 & ~n20641 ;
  assign n20643 = n20642 ^ n16729 ^ 1'b0 ;
  assign n20644 = n20643 ^ n16164 ^ n8914 ;
  assign n20645 = n7651 ^ n343 ^ 1'b0 ;
  assign n20646 = n20645 ^ n20224 ^ n6504 ;
  assign n20647 = n15505 ^ n6600 ^ n3191 ;
  assign n20650 = n5095 ^ n2726 ^ n660 ;
  assign n20648 = n3569 | n8563 ;
  assign n20649 = n12382 | n20648 ;
  assign n20651 = n20650 ^ n20649 ^ 1'b0 ;
  assign n20652 = n8168 ^ n4089 ^ 1'b0 ;
  assign n20653 = n20652 ^ n1390 ^ 1'b0 ;
  assign n20654 = ( x195 & ~n8413 ) | ( x195 & n10272 ) | ( ~n8413 & n10272 ) ;
  assign n20655 = n5574 & ~n10319 ;
  assign n20656 = ( n4547 & n20654 ) | ( n4547 & ~n20655 ) | ( n20654 & ~n20655 ) ;
  assign n20657 = ~n20653 & n20656 ;
  assign n20658 = n20657 ^ n15926 ^ 1'b0 ;
  assign n20659 = n16911 ^ n325 ^ 1'b0 ;
  assign n20660 = n12513 & ~n20659 ;
  assign n20661 = n4049 | n20660 ;
  assign n20662 = n10724 ^ n7234 ^ n2111 ;
  assign n20663 = ( ~n4998 & n8531 ) | ( ~n4998 & n13513 ) | ( n8531 & n13513 ) ;
  assign n20664 = n20663 ^ n1087 ^ 1'b0 ;
  assign n20665 = ~n18101 & n20664 ;
  assign n20666 = ( n3054 & ~n20662 ) | ( n3054 & n20665 ) | ( ~n20662 & n20665 ) ;
  assign n20667 = ( n8445 & ~n11094 ) | ( n8445 & n20625 ) | ( ~n11094 & n20625 ) ;
  assign n20670 = ( ~n1632 & n3018 ) | ( ~n1632 & n3749 ) | ( n3018 & n3749 ) ;
  assign n20668 = ~n3892 & n5363 ;
  assign n20669 = n20668 ^ n2633 ^ 1'b0 ;
  assign n20671 = n20670 ^ n20669 ^ n2744 ;
  assign n20672 = n9001 & n20671 ;
  assign n20673 = ~n4623 & n20672 ;
  assign n20674 = n11572 & ~n20673 ;
  assign n20675 = n20674 ^ n6265 ^ 1'b0 ;
  assign n20676 = ( n13919 & n18377 ) | ( n13919 & ~n19895 ) | ( n18377 & ~n19895 ) ;
  assign n20677 = ( n4775 & ~n4794 ) | ( n4775 & n8206 ) | ( ~n4794 & n8206 ) ;
  assign n20678 = n14294 & ~n20677 ;
  assign n20679 = n20678 ^ n11525 ^ 1'b0 ;
  assign n20680 = n13022 ^ n4789 ^ 1'b0 ;
  assign n20681 = n20679 & n20680 ;
  assign n20682 = ( n2099 & ~n11784 ) | ( n2099 & n14022 ) | ( ~n11784 & n14022 ) ;
  assign n20683 = ( ~n2247 & n7606 ) | ( ~n2247 & n7640 ) | ( n7606 & n7640 ) ;
  assign n20684 = n20683 ^ n19137 ^ 1'b0 ;
  assign n20685 = ~n6174 & n20684 ;
  assign n20686 = n3548 | n13985 ;
  assign n20687 = n20686 ^ n13764 ^ n13589 ;
  assign n20689 = n1562 & ~n5245 ;
  assign n20690 = n4106 & n20689 ;
  assign n20688 = n16859 ^ n10123 ^ n525 ;
  assign n20691 = n20690 ^ n20688 ^ 1'b0 ;
  assign n20692 = ( ~n20279 & n20687 ) | ( ~n20279 & n20691 ) | ( n20687 & n20691 ) ;
  assign n20693 = n20685 & n20692 ;
  assign n20695 = n8742 ^ n2320 ^ 1'b0 ;
  assign n20696 = ( n7139 & n8139 ) | ( n7139 & ~n20695 ) | ( n8139 & ~n20695 ) ;
  assign n20694 = n6559 | n9230 ;
  assign n20697 = n20696 ^ n20694 ^ 1'b0 ;
  assign n20698 = n2256 | n20697 ;
  assign n20699 = n8750 ^ n3492 ^ 1'b0 ;
  assign n20700 = n8847 & n20699 ;
  assign n20701 = ~n13271 & n20700 ;
  assign n20702 = ( ~n11702 & n20698 ) | ( ~n11702 & n20701 ) | ( n20698 & n20701 ) ;
  assign n20703 = n5387 ^ n1257 ^ n511 ;
  assign n20704 = n9741 ^ n7409 ^ n6022 ;
  assign n20705 = n20703 | n20704 ;
  assign n20706 = n20705 ^ n17422 ^ n15013 ;
  assign n20707 = n9410 & n20144 ;
  assign n20708 = n6005 & n20707 ;
  assign n20709 = ( n10942 & n11777 ) | ( n10942 & n14188 ) | ( n11777 & n14188 ) ;
  assign n20710 = ~n1469 & n5957 ;
  assign n20711 = n2062 & n20710 ;
  assign n20712 = ( n3568 & n3832 ) | ( n3568 & ~n13587 ) | ( n3832 & ~n13587 ) ;
  assign n20713 = ~n20711 & n20712 ;
  assign n20714 = ~n20709 & n20713 ;
  assign n20715 = ( n1676 & n8211 ) | ( n1676 & n14489 ) | ( n8211 & n14489 ) ;
  assign n20716 = ~n9148 & n20715 ;
  assign n20717 = n20716 ^ n3408 ^ 1'b0 ;
  assign n20718 = n6076 | n20717 ;
  assign n20723 = n14789 ^ n8583 ^ 1'b0 ;
  assign n20724 = n15835 | n20723 ;
  assign n20719 = n2372 | n8894 ;
  assign n20720 = n9067 | n20719 ;
  assign n20721 = n19648 & ~n19868 ;
  assign n20722 = ~n20720 & n20721 ;
  assign n20725 = n20724 ^ n20722 ^ n13198 ;
  assign n20727 = n15885 ^ n11538 ^ n7753 ;
  assign n20728 = ( n8060 & n11893 ) | ( n8060 & n20727 ) | ( n11893 & n20727 ) ;
  assign n20726 = n8466 ^ n6326 ^ n3335 ;
  assign n20729 = n20728 ^ n20726 ^ n13231 ;
  assign n20730 = n10770 & ~n20729 ;
  assign n20733 = ~n3143 & n19762 ;
  assign n20734 = ( x53 & n7516 ) | ( x53 & n20733 ) | ( n7516 & n20733 ) ;
  assign n20731 = ~n11153 & n13819 ;
  assign n20732 = n20731 ^ n493 ^ 1'b0 ;
  assign n20735 = n20734 ^ n20732 ^ n8551 ;
  assign n20739 = ( n1666 & ~n3303 ) | ( n1666 & n19891 ) | ( ~n3303 & n19891 ) ;
  assign n20740 = n1705 & ~n16649 ;
  assign n20741 = n7778 & n20740 ;
  assign n20742 = n20741 ^ n16392 ^ 1'b0 ;
  assign n20743 = n20739 & n20742 ;
  assign n20744 = n12777 | n20743 ;
  assign n20736 = x187 & n8962 ;
  assign n20737 = n8132 & n20736 ;
  assign n20738 = n6577 | n20737 ;
  assign n20745 = n20744 ^ n20738 ^ 1'b0 ;
  assign n20747 = n20237 ^ n6166 ^ 1'b0 ;
  assign n20746 = ( ~n1828 & n9013 ) | ( ~n1828 & n9794 ) | ( n9013 & n9794 ) ;
  assign n20748 = n20747 ^ n20746 ^ n12290 ;
  assign n20749 = n3415 | n12737 ;
  assign n20750 = n11956 & ~n20749 ;
  assign n20751 = n3142 & n3536 ;
  assign n20752 = n20751 ^ n7692 ^ 1'b0 ;
  assign n20753 = n20752 ^ n18819 ^ 1'b0 ;
  assign n20754 = ~n7037 & n20753 ;
  assign n20755 = ( n1892 & ~n4208 ) | ( n1892 & n4475 ) | ( ~n4208 & n4475 ) ;
  assign n20756 = n20755 ^ n11823 ^ 1'b0 ;
  assign n20757 = n9182 ^ n838 ^ 1'b0 ;
  assign n20758 = n11773 | n20744 ;
  assign n20763 = ( ~n857 & n6214 ) | ( ~n857 & n11257 ) | ( n6214 & n11257 ) ;
  assign n20764 = n20763 ^ n13222 ^ n8228 ;
  assign n20765 = n6969 & n15202 ;
  assign n20766 = n20764 & n20765 ;
  assign n20767 = n20766 ^ n8276 ^ n1370 ;
  assign n20759 = n7309 | n7681 ;
  assign n20760 = n3402 | n17410 ;
  assign n20761 = n20759 | n20760 ;
  assign n20762 = n20761 ^ n8119 ^ 1'b0 ;
  assign n20768 = n20767 ^ n20762 ^ n8218 ;
  assign n20769 = ( n1466 & n6768 ) | ( n1466 & ~n20768 ) | ( n6768 & ~n20768 ) ;
  assign n20770 = n20769 ^ n13815 ^ n9984 ;
  assign n20771 = ( ~n1331 & n12408 ) | ( ~n1331 & n20533 ) | ( n12408 & n20533 ) ;
  assign n20776 = n1330 ^ n1087 ^ 1'b0 ;
  assign n20772 = n2445 ^ n2178 ^ 1'b0 ;
  assign n20773 = n20772 ^ n2356 ^ 1'b0 ;
  assign n20774 = n20773 ^ n1020 ^ n533 ;
  assign n20775 = n11231 & n20774 ;
  assign n20777 = n20776 ^ n20775 ^ 1'b0 ;
  assign n20782 = ( n547 & ~n5946 ) | ( n547 & n16039 ) | ( ~n5946 & n16039 ) ;
  assign n20783 = n16373 & ~n20782 ;
  assign n20784 = n20783 ^ n9616 ^ 1'b0 ;
  assign n20778 = n4516 ^ x92 ^ 1'b0 ;
  assign n20779 = n7664 ^ n4032 ^ n2856 ;
  assign n20780 = ( n8990 & n17482 ) | ( n8990 & n20779 ) | ( n17482 & n20779 ) ;
  assign n20781 = n20778 | n20780 ;
  assign n20785 = n20784 ^ n20781 ^ n12062 ;
  assign n20786 = ( n3994 & ~n6926 ) | ( n3994 & n8807 ) | ( ~n6926 & n8807 ) ;
  assign n20787 = ( ~x54 & n14067 ) | ( ~x54 & n20786 ) | ( n14067 & n20786 ) ;
  assign n20788 = n7688 | n20109 ;
  assign n20789 = n9589 | n20788 ;
  assign n20790 = n12887 & ~n15568 ;
  assign n20791 = n20790 ^ n14303 ^ 1'b0 ;
  assign n20794 = n9772 ^ n9167 ^ n1340 ;
  assign n20793 = ~n2233 & n9973 ;
  assign n20792 = n4941 | n7458 ;
  assign n20795 = n20794 ^ n20793 ^ n20792 ;
  assign n20796 = n2589 & n6739 ;
  assign n20797 = n4297 ^ n2906 ^ x26 ;
  assign n20798 = ( n1680 & n1746 ) | ( n1680 & ~n20797 ) | ( n1746 & ~n20797 ) ;
  assign n20799 = n12931 ^ n6975 ^ n1831 ;
  assign n20800 = n13134 & ~n20799 ;
  assign n20801 = n930 & n17211 ;
  assign n20802 = n7651 & n20801 ;
  assign n20803 = n20802 ^ n18504 ^ 1'b0 ;
  assign n20804 = n13277 ^ n7322 ^ n533 ;
  assign n20805 = n20804 ^ n8648 ^ n1403 ;
  assign n20806 = n6634 & n17851 ;
  assign n20807 = ~n10336 & n20806 ;
  assign n20808 = n20807 ^ n11811 ^ 1'b0 ;
  assign n20809 = n5414 | n6020 ;
  assign n20810 = n20808 | n20809 ;
  assign n20811 = ( n556 & n8415 ) | ( n556 & n9071 ) | ( n8415 & n9071 ) ;
  assign n20812 = x101 & n20811 ;
  assign n20813 = n813 & n13175 ;
  assign n20814 = ( ~n7233 & n11205 ) | ( ~n7233 & n16640 ) | ( n11205 & n16640 ) ;
  assign n20815 = n20813 & n20814 ;
  assign n20816 = n16684 & n20815 ;
  assign n20817 = n19995 & ~n20816 ;
  assign n20818 = ( n1886 & ~n10649 ) | ( n1886 & n15282 ) | ( ~n10649 & n15282 ) ;
  assign n20819 = n687 | n20818 ;
  assign n20820 = x182 & ~n3256 ;
  assign n20821 = n20820 ^ n6527 ^ 1'b0 ;
  assign n20822 = n20821 ^ n17795 ^ n7736 ;
  assign n20824 = n10915 ^ n6693 ^ 1'b0 ;
  assign n20823 = n18627 ^ n6061 ^ n1951 ;
  assign n20825 = n20824 ^ n20823 ^ 1'b0 ;
  assign n20826 = ~n8676 & n20825 ;
  assign n20827 = n20826 ^ n9616 ^ 1'b0 ;
  assign n20828 = n959 & ~n8906 ;
  assign n20829 = n20828 ^ n11809 ^ 1'b0 ;
  assign n20830 = ~n13290 & n20829 ;
  assign n20831 = n19322 & n20830 ;
  assign n20832 = n16789 ^ n12882 ^ 1'b0 ;
  assign n20833 = ~x187 & n2381 ;
  assign n20834 = ~n4960 & n19648 ;
  assign n20835 = n20834 ^ n5818 ^ 1'b0 ;
  assign n20837 = x28 & n663 ;
  assign n20836 = n882 & ~n7932 ;
  assign n20838 = n20837 ^ n20836 ^ 1'b0 ;
  assign n20839 = n1404 & ~n2598 ;
  assign n20840 = n20839 ^ n16742 ^ 1'b0 ;
  assign n20841 = n13534 ^ n7377 ^ n1336 ;
  assign n20842 = ( ~n10316 & n11976 ) | ( ~n10316 & n20841 ) | ( n11976 & n20841 ) ;
  assign n20843 = ( n16701 & n20840 ) | ( n16701 & ~n20842 ) | ( n20840 & ~n20842 ) ;
  assign n20844 = n16498 ^ n7987 ^ n7940 ;
  assign n20845 = n8749 ^ n6917 ^ n2759 ;
  assign n20846 = n6424 & n20845 ;
  assign n20847 = n12977 ^ n9201 ^ 1'b0 ;
  assign n20848 = ( n603 & ~n20846 ) | ( n603 & n20847 ) | ( ~n20846 & n20847 ) ;
  assign n20849 = n770 | n2031 ;
  assign n20850 = ( n11570 & n15063 ) | ( n11570 & ~n20849 ) | ( n15063 & ~n20849 ) ;
  assign n20851 = ( n6883 & n7579 ) | ( n6883 & n7640 ) | ( n7579 & n7640 ) ;
  assign n20852 = n20851 ^ n8728 ^ n812 ;
  assign n20853 = ~n8649 & n12557 ;
  assign n20854 = n20853 ^ n6817 ^ 1'b0 ;
  assign n20855 = ~n3252 & n20854 ;
  assign n20856 = n20855 ^ n4346 ^ 1'b0 ;
  assign n20857 = ~n6418 & n20856 ;
  assign n20858 = n19284 ^ n16078 ^ 1'b0 ;
  assign n20859 = n9644 | n20858 ;
  assign n20860 = n4575 ^ n1206 ^ n960 ;
  assign n20861 = n13767 & n20860 ;
  assign n20862 = n5816 | n7113 ;
  assign n20863 = n20862 ^ n1465 ^ 1'b0 ;
  assign n20864 = ~n17866 & n20863 ;
  assign n20865 = n2393 & ~n4042 ;
  assign n20866 = ( n3274 & n14657 ) | ( n3274 & ~n20865 ) | ( n14657 & ~n20865 ) ;
  assign n20867 = n20866 ^ n8372 ^ 1'b0 ;
  assign n20868 = n5912 | n20867 ;
  assign n20869 = n20868 ^ n7627 ^ 1'b0 ;
  assign n20871 = n724 & n2552 ;
  assign n20872 = n20871 ^ n7175 ^ 1'b0 ;
  assign n20870 = n4475 | n8911 ;
  assign n20873 = n20872 ^ n20870 ^ 1'b0 ;
  assign n20874 = ( n533 & n17461 ) | ( n533 & ~n20873 ) | ( n17461 & ~n20873 ) ;
  assign n20875 = n4859 ^ n2372 ^ 1'b0 ;
  assign n20876 = ( n5941 & ~n16738 ) | ( n5941 & n20875 ) | ( ~n16738 & n20875 ) ;
  assign n20878 = n5213 & ~n8902 ;
  assign n20879 = n20878 ^ n13767 ^ 1'b0 ;
  assign n20880 = n5369 ^ n4932 ^ 1'b0 ;
  assign n20881 = n20879 & n20880 ;
  assign n20877 = n12059 & n12915 ;
  assign n20882 = n20881 ^ n20877 ^ 1'b0 ;
  assign n20883 = ( n3546 & n11339 ) | ( n3546 & n20882 ) | ( n11339 & n20882 ) ;
  assign n20890 = n3550 & n11527 ;
  assign n20891 = n11378 | n20890 ;
  assign n20892 = n20891 ^ n20639 ^ 1'b0 ;
  assign n20884 = ~n7200 & n10173 ;
  assign n20885 = n20884 ^ n539 ^ 1'b0 ;
  assign n20886 = ~n773 & n20885 ;
  assign n20887 = ( n2168 & ~n16107 ) | ( n2168 & n20886 ) | ( ~n16107 & n20886 ) ;
  assign n20888 = n20887 ^ n311 ^ 1'b0 ;
  assign n20889 = n3627 & n20888 ;
  assign n20893 = n20892 ^ n20889 ^ n2071 ;
  assign n20894 = n20893 ^ n8784 ^ 1'b0 ;
  assign n20895 = ( n5587 & ~n5836 ) | ( n5587 & n14788 ) | ( ~n5836 & n14788 ) ;
  assign n20896 = n1396 | n9471 ;
  assign n20897 = n20895 & ~n20896 ;
  assign n20898 = n6953 ^ n3352 ^ n2270 ;
  assign n20899 = ~n10104 & n20898 ;
  assign n20900 = n20899 ^ n4725 ^ 1'b0 ;
  assign n20901 = ~n742 & n20900 ;
  assign n20902 = n20901 ^ n6444 ^ 1'b0 ;
  assign n20903 = ~n20897 & n20902 ;
  assign n20904 = n14432 ^ n13156 ^ 1'b0 ;
  assign n20905 = n12089 & ~n20904 ;
  assign n20906 = n20905 ^ n15989 ^ 1'b0 ;
  assign n20914 = n1004 & ~n3156 ;
  assign n20915 = n18488 & n20914 ;
  assign n20911 = ( n3370 & ~n4623 ) | ( n3370 & n5027 ) | ( ~n4623 & n5027 ) ;
  assign n20912 = n20911 ^ n12891 ^ 1'b0 ;
  assign n20913 = ~n6888 & n20912 ;
  assign n20908 = n7670 ^ n1510 ^ 1'b0 ;
  assign n20909 = ~n3565 & n20908 ;
  assign n20907 = n17021 | n17110 ;
  assign n20910 = n20909 ^ n20907 ^ 1'b0 ;
  assign n20916 = n20915 ^ n20913 ^ n20910 ;
  assign n20917 = n10825 ^ n8726 ^ n1777 ;
  assign n20921 = n631 | n2114 ;
  assign n20922 = ( ~n13943 & n14673 ) | ( ~n13943 & n20921 ) | ( n14673 & n20921 ) ;
  assign n20918 = ( n2148 & ~n4902 ) | ( n2148 & n9108 ) | ( ~n4902 & n9108 ) ;
  assign n20919 = n2169 | n20918 ;
  assign n20920 = n20919 ^ n1722 ^ 1'b0 ;
  assign n20923 = n20922 ^ n20920 ^ 1'b0 ;
  assign n20924 = n6099 & ~n20923 ;
  assign n20925 = n15783 ^ n2911 ^ n1425 ;
  assign n20926 = ( n8451 & n13167 ) | ( n8451 & n20925 ) | ( n13167 & n20925 ) ;
  assign n20927 = n19049 & ~n20926 ;
  assign n20928 = n20927 ^ n2709 ^ 1'b0 ;
  assign n20932 = ( n6328 & ~n8270 ) | ( n6328 & n9727 ) | ( ~n8270 & n9727 ) ;
  assign n20931 = n14588 ^ n4027 ^ 1'b0 ;
  assign n20929 = n16491 ^ n3892 ^ 1'b0 ;
  assign n20930 = n7313 & ~n20929 ;
  assign n20933 = n20932 ^ n20931 ^ n20930 ;
  assign n20934 = n13670 ^ n4818 ^ n1367 ;
  assign n20935 = n20934 ^ n12471 ^ n4927 ;
  assign n20936 = ~n9689 & n20935 ;
  assign n20939 = n3929 | n9885 ;
  assign n20937 = ( n2722 & n4152 ) | ( n2722 & ~n5159 ) | ( n4152 & ~n5159 ) ;
  assign n20938 = n20937 ^ n3024 ^ 1'b0 ;
  assign n20940 = n20939 ^ n20938 ^ n475 ;
  assign n20943 = n2682 | n3255 ;
  assign n20944 = n20943 ^ n6743 ^ 1'b0 ;
  assign n20941 = n13505 ^ n5738 ^ 1'b0 ;
  assign n20942 = ~n16032 & n20941 ;
  assign n20945 = n20944 ^ n20942 ^ n8461 ;
  assign n20946 = n20945 ^ n11231 ^ n7238 ;
  assign n20947 = n15829 ^ n13534 ^ 1'b0 ;
  assign n20948 = n7374 | n20947 ;
  assign n20949 = ( n12157 & n20066 ) | ( n12157 & ~n20948 ) | ( n20066 & ~n20948 ) ;
  assign n20950 = n2217 & ~n5239 ;
  assign n20951 = n517 & n20950 ;
  assign n20952 = n317 & ~n17086 ;
  assign n20953 = n20952 ^ n2105 ^ 1'b0 ;
  assign n20954 = n1647 | n20953 ;
  assign n20955 = n20954 ^ n14750 ^ 1'b0 ;
  assign n20956 = ( ~n8160 & n12607 ) | ( ~n8160 & n14973 ) | ( n12607 & n14973 ) ;
  assign n20957 = n20956 ^ n2837 ^ 1'b0 ;
  assign n20958 = n20957 ^ n4483 ^ n648 ;
  assign n20959 = ~n1081 & n4809 ;
  assign n20960 = n19618 ^ n8945 ^ 1'b0 ;
  assign n20961 = n1786 | n20960 ;
  assign n20962 = n10800 ^ n10576 ^ n1198 ;
  assign n20963 = n13599 | n14061 ;
  assign n20964 = n20962 & ~n20963 ;
  assign n20965 = n10304 ^ n9709 ^ 1'b0 ;
  assign n20966 = n5026 ^ n1761 ^ 1'b0 ;
  assign n20967 = n10607 | n12674 ;
  assign n20968 = n20966 & ~n20967 ;
  assign n20969 = ( ~n13093 & n20965 ) | ( ~n13093 & n20968 ) | ( n20965 & n20968 ) ;
  assign n20970 = n3107 & ~n20969 ;
  assign n20971 = n4240 ^ n1637 ^ 1'b0 ;
  assign n20972 = n12859 & n20971 ;
  assign n20973 = ( ~n18893 & n20461 ) | ( ~n18893 & n20972 ) | ( n20461 & n20972 ) ;
  assign n20974 = n17595 ^ n1140 ^ 1'b0 ;
  assign n20975 = n9973 & n20974 ;
  assign n20976 = n13961 ^ n6020 ^ n1578 ;
  assign n20977 = ( n5343 & n13837 ) | ( n5343 & ~n20976 ) | ( n13837 & ~n20976 ) ;
  assign n20978 = n20977 ^ n19016 ^ n7174 ;
  assign n20979 = n19868 | n20978 ;
  assign n20980 = n20979 ^ n16794 ^ 1'b0 ;
  assign n20981 = n4340 ^ n716 ^ 1'b0 ;
  assign n20982 = n9685 & n20981 ;
  assign n20983 = n17843 ^ n3028 ^ 1'b0 ;
  assign n20988 = n3466 & ~n7013 ;
  assign n20989 = ~n4228 & n20988 ;
  assign n20990 = n20989 ^ n9114 ^ n5513 ;
  assign n20991 = ( n11777 & n17324 ) | ( n11777 & ~n20990 ) | ( n17324 & ~n20990 ) ;
  assign n20986 = n912 ^ n349 ^ 1'b0 ;
  assign n20987 = ~n8453 & n20986 ;
  assign n20984 = n2543 & n5147 ;
  assign n20985 = ( n6561 & n14723 ) | ( n6561 & ~n20984 ) | ( n14723 & ~n20984 ) ;
  assign n20992 = n20991 ^ n20987 ^ n20985 ;
  assign n20993 = n18246 ^ n7454 ^ n5141 ;
  assign n20994 = ( n256 & ~n6592 ) | ( n256 & n14175 ) | ( ~n6592 & n14175 ) ;
  assign n20995 = ( n2024 & ~n5313 ) | ( n2024 & n9949 ) | ( ~n5313 & n9949 ) ;
  assign n20996 = n20995 ^ n10551 ^ 1'b0 ;
  assign n20997 = n20994 & n20996 ;
  assign n20998 = ~n9626 & n10472 ;
  assign n20999 = n20998 ^ n2556 ^ 1'b0 ;
  assign n21000 = n20999 ^ n15825 ^ 1'b0 ;
  assign n21001 = x167 & n21000 ;
  assign n21002 = ( n3397 & n11932 ) | ( n3397 & n20277 ) | ( n11932 & n20277 ) ;
  assign n21003 = n470 | n21002 ;
  assign n21004 = n21003 ^ n12226 ^ 1'b0 ;
  assign n21005 = n15289 ^ n2981 ^ n674 ;
  assign n21006 = ( n3741 & n21004 ) | ( n3741 & ~n21005 ) | ( n21004 & ~n21005 ) ;
  assign n21007 = ( n9021 & n17205 ) | ( n9021 & ~n21006 ) | ( n17205 & ~n21006 ) ;
  assign n21008 = ( n3806 & n4475 ) | ( n3806 & n15663 ) | ( n4475 & n15663 ) ;
  assign n21009 = ( n1476 & n7366 ) | ( n1476 & n21008 ) | ( n7366 & n21008 ) ;
  assign n21010 = n21009 ^ n5082 ^ 1'b0 ;
  assign n21011 = n15167 | n18682 ;
  assign n21016 = n7652 ^ n7436 ^ 1'b0 ;
  assign n21017 = n3430 & ~n21016 ;
  assign n21018 = ( n1988 & n18747 ) | ( n1988 & n21017 ) | ( n18747 & n21017 ) ;
  assign n21019 = ~n6531 & n21018 ;
  assign n21020 = n21019 ^ n663 ^ 1'b0 ;
  assign n21012 = n3281 ^ n625 ^ 1'b0 ;
  assign n21013 = ~n4822 & n21012 ;
  assign n21014 = n21013 ^ n17046 ^ n2298 ;
  assign n21015 = ~n5526 & n21014 ;
  assign n21021 = n21020 ^ n21015 ^ 1'b0 ;
  assign n21022 = n6463 & n21021 ;
  assign n21023 = n3087 ^ n1266 ^ 1'b0 ;
  assign n21024 = n11238 & n18533 ;
  assign n21025 = n21023 & n21024 ;
  assign n21026 = n7553 & ~n21025 ;
  assign n21027 = n17888 & ~n21026 ;
  assign n21028 = n21027 ^ n15330 ^ 1'b0 ;
  assign n21029 = n10790 ^ n5214 ^ 1'b0 ;
  assign n21030 = ~n13212 & n21029 ;
  assign n21032 = ( n967 & n4200 ) | ( n967 & n6891 ) | ( n4200 & n6891 ) ;
  assign n21031 = n3297 & ~n4179 ;
  assign n21033 = n21032 ^ n21031 ^ 1'b0 ;
  assign n21034 = ( n3330 & ~n5622 ) | ( n3330 & n21033 ) | ( ~n5622 & n21033 ) ;
  assign n21035 = n21034 ^ n3392 ^ n1884 ;
  assign n21036 = n2637 & ~n3741 ;
  assign n21037 = n17539 | n21036 ;
  assign n21038 = n2471 & n21037 ;
  assign n21039 = n3262 & n21038 ;
  assign n21040 = n16451 | n21039 ;
  assign n21041 = n6652 & ~n21040 ;
  assign n21042 = n2270 | n21041 ;
  assign n21043 = n21042 ^ n5213 ^ 1'b0 ;
  assign n21044 = n14040 ^ x193 ^ 1'b0 ;
  assign n21046 = n15573 ^ n4476 ^ 1'b0 ;
  assign n21045 = n7388 & ~n15485 ;
  assign n21047 = n21046 ^ n21045 ^ 1'b0 ;
  assign n21051 = ~n593 & n12032 ;
  assign n21048 = n16734 ^ n4902 ^ n4241 ;
  assign n21049 = n21048 ^ n8382 ^ 1'b0 ;
  assign n21050 = ~n9150 & n21049 ;
  assign n21052 = n21051 ^ n21050 ^ 1'b0 ;
  assign n21053 = n21047 | n21052 ;
  assign n21054 = n10662 ^ n8209 ^ n2700 ;
  assign n21055 = n21054 ^ n14824 ^ 1'b0 ;
  assign n21056 = ~n12730 & n19182 ;
  assign n21057 = ( n355 & n1966 ) | ( n355 & ~n11774 ) | ( n1966 & ~n11774 ) ;
  assign n21058 = n13617 ^ n1776 ^ x145 ;
  assign n21059 = ~n11970 & n21058 ;
  assign n21060 = ( ~n11515 & n15975 ) | ( ~n11515 & n21059 ) | ( n15975 & n21059 ) ;
  assign n21064 = n11678 ^ n9720 ^ 1'b0 ;
  assign n21061 = n1067 ^ x227 ^ x159 ;
  assign n21062 = n5153 & ~n21061 ;
  assign n21063 = n21062 ^ n11944 ^ n2309 ;
  assign n21065 = n21064 ^ n21063 ^ n3061 ;
  assign n21066 = ~n2280 & n10751 ;
  assign n21067 = n20217 ^ n16349 ^ 1'b0 ;
  assign n21068 = ~n21066 & n21067 ;
  assign n21069 = n3810 | n17604 ;
  assign n21070 = n4960 ^ x173 ^ 1'b0 ;
  assign n21071 = n9204 | n21070 ;
  assign n21072 = n21071 ^ n16602 ^ n11811 ;
  assign n21073 = ~n12049 & n14712 ;
  assign n21074 = n18620 ^ n4645 ^ n1418 ;
  assign n21075 = n21074 ^ n789 ^ 1'b0 ;
  assign n21077 = ~n835 & n9225 ;
  assign n21078 = ~n3350 & n21077 ;
  assign n21079 = n5835 ^ n1173 ^ 1'b0 ;
  assign n21080 = n8173 & ~n21079 ;
  assign n21081 = n14775 & n21080 ;
  assign n21082 = ( n4249 & n21078 ) | ( n4249 & n21081 ) | ( n21078 & n21081 ) ;
  assign n21076 = n18374 ^ n12685 ^ 1'b0 ;
  assign n21083 = n21082 ^ n21076 ^ n8456 ;
  assign n21084 = n8738 & n11873 ;
  assign n21086 = n14695 ^ n13212 ^ n3538 ;
  assign n21085 = x206 & ~n7343 ;
  assign n21087 = n21086 ^ n21085 ^ 1'b0 ;
  assign n21088 = n6287 ^ n1137 ^ 1'b0 ;
  assign n21089 = n21088 ^ n19953 ^ n15579 ;
  assign n21090 = ( n14586 & n17094 ) | ( n14586 & ~n21089 ) | ( n17094 & ~n21089 ) ;
  assign n21091 = ( ~n17717 & n21087 ) | ( ~n17717 & n21090 ) | ( n21087 & n21090 ) ;
  assign n21092 = n12624 | n16519 ;
  assign n21093 = n15053 | n21092 ;
  assign n21094 = n3538 | n10373 ;
  assign n21095 = n7227 | n21094 ;
  assign n21096 = n2048 | n15822 ;
  assign n21097 = ~n6957 & n21096 ;
  assign n21098 = n21097 ^ x252 ^ 1'b0 ;
  assign n21099 = ( ~n15742 & n21095 ) | ( ~n15742 & n21098 ) | ( n21095 & n21098 ) ;
  assign n21100 = n9231 ^ n9029 ^ 1'b0 ;
  assign n21101 = n21099 | n21100 ;
  assign n21102 = n21093 | n21101 ;
  assign n21103 = n7185 | n17580 ;
  assign n21104 = n21103 ^ n270 ^ 1'b0 ;
  assign n21105 = n7461 & ~n8781 ;
  assign n21108 = n11440 ^ n840 ^ x151 ;
  assign n21106 = n9978 ^ n4577 ^ 1'b0 ;
  assign n21107 = ~n9085 & n21106 ;
  assign n21109 = n21108 ^ n21107 ^ n8665 ;
  assign n21110 = n16080 ^ n15000 ^ n4817 ;
  assign n21111 = n2829 & n21110 ;
  assign n21112 = ( n2311 & n2705 ) | ( n2311 & ~n13243 ) | ( n2705 & ~n13243 ) ;
  assign n21113 = n4139 ^ n683 ^ 1'b0 ;
  assign n21114 = ~n2198 & n21113 ;
  assign n21115 = ~n21112 & n21114 ;
  assign n21116 = ~n6990 & n21115 ;
  assign n21117 = ( ~n2141 & n6973 ) | ( ~n2141 & n21116 ) | ( n6973 & n21116 ) ;
  assign n21118 = ( n829 & ~n2302 ) | ( n829 & n21117 ) | ( ~n2302 & n21117 ) ;
  assign n21119 = n17592 ^ n15334 ^ n771 ;
  assign n21120 = ~n4728 & n21119 ;
  assign n21121 = n8417 & n21120 ;
  assign n21122 = n636 & ~n3786 ;
  assign n21123 = n8913 | n21122 ;
  assign n21124 = n21121 & ~n21123 ;
  assign n21125 = n7940 & ~n18678 ;
  assign n21126 = n13658 ^ n6207 ^ n5262 ;
  assign n21127 = n10369 & ~n21126 ;
  assign n21128 = n21127 ^ n3656 ^ 1'b0 ;
  assign n21131 = ~n2456 & n2694 ;
  assign n21132 = n6905 & n21131 ;
  assign n21133 = n19766 & ~n21132 ;
  assign n21129 = n4687 & n8072 ;
  assign n21130 = ~n8079 & n21129 ;
  assign n21134 = n21133 ^ n21130 ^ n408 ;
  assign n21135 = n12725 ^ n9108 ^ n512 ;
  assign n21136 = ( n6753 & n9548 ) | ( n6753 & ~n12634 ) | ( n9548 & ~n12634 ) ;
  assign n21137 = n15491 ^ n12778 ^ n7539 ;
  assign n21138 = ( n21135 & n21136 ) | ( n21135 & n21137 ) | ( n21136 & n21137 ) ;
  assign n21139 = n10774 ^ n1753 ^ 1'b0 ;
  assign n21143 = n10330 ^ n9940 ^ n7323 ;
  assign n21140 = ~x36 & n2006 ;
  assign n21141 = n3028 & n21140 ;
  assign n21142 = n1328 & ~n21141 ;
  assign n21144 = n21143 ^ n21142 ^ n5435 ;
  assign n21145 = n5297 | n5953 ;
  assign n21148 = n7832 & n11601 ;
  assign n21146 = n5561 ^ n4672 ^ n4222 ;
  assign n21147 = ( n13286 & n16595 ) | ( n13286 & n21146 ) | ( n16595 & n21146 ) ;
  assign n21149 = n21148 ^ n21147 ^ n9541 ;
  assign n21150 = n1172 & n1611 ;
  assign n21151 = n21150 ^ n453 ^ 1'b0 ;
  assign n21152 = n920 | n14055 ;
  assign n21153 = ( n5587 & n10343 ) | ( n5587 & n20026 ) | ( n10343 & n20026 ) ;
  assign n21154 = n14207 ^ n12927 ^ 1'b0 ;
  assign n21155 = n11206 | n21154 ;
  assign n21156 = n21153 | n21155 ;
  assign n21157 = ( n8507 & ~n21152 ) | ( n8507 & n21156 ) | ( ~n21152 & n21156 ) ;
  assign n21158 = n21151 & n21157 ;
  assign n21159 = ( n4117 & n21149 ) | ( n4117 & ~n21158 ) | ( n21149 & ~n21158 ) ;
  assign n21160 = ( n1326 & ~n1867 ) | ( n1326 & n2110 ) | ( ~n1867 & n2110 ) ;
  assign n21161 = ( n4525 & ~n14253 ) | ( n4525 & n21160 ) | ( ~n14253 & n21160 ) ;
  assign n21162 = n15514 | n21161 ;
  assign n21163 = n20948 ^ n4195 ^ n713 ;
  assign n21164 = n21163 ^ n2782 ^ 1'b0 ;
  assign n21165 = n13913 ^ n3283 ^ 1'b0 ;
  assign n21166 = n20458 & n21165 ;
  assign n21167 = n11274 | n21166 ;
  assign n21168 = n8793 & ~n21167 ;
  assign n21169 = n5428 ^ n4529 ^ x151 ;
  assign n21170 = x186 & ~n3022 ;
  assign n21171 = n21170 ^ n1063 ^ 1'b0 ;
  assign n21172 = n5005 & ~n21171 ;
  assign n21173 = ~n21169 & n21172 ;
  assign n21174 = n11653 & ~n12059 ;
  assign n21175 = n4687 & n8686 ;
  assign n21176 = n14416 & n21175 ;
  assign n21177 = ( n1254 & ~n2402 ) | ( n1254 & n21176 ) | ( ~n2402 & n21176 ) ;
  assign n21178 = ( n7867 & n21174 ) | ( n7867 & n21177 ) | ( n21174 & n21177 ) ;
  assign n21179 = n21178 ^ n17737 ^ n6379 ;
  assign n21180 = ~n10361 & n14256 ;
  assign n21181 = n21180 ^ n7369 ^ 1'b0 ;
  assign n21182 = n12559 | n21181 ;
  assign n21183 = n16077 | n21182 ;
  assign n21184 = n2033 | n5458 ;
  assign n21185 = n14976 & ~n21184 ;
  assign n21186 = n2817 | n8247 ;
  assign n21187 = n7857 | n10451 ;
  assign n21188 = n21186 & ~n21187 ;
  assign n21189 = n21188 ^ n13971 ^ n8854 ;
  assign n21190 = ( ~n569 & n4452 ) | ( ~n569 & n7899 ) | ( n4452 & n7899 ) ;
  assign n21191 = n21190 ^ n11313 ^ 1'b0 ;
  assign n21192 = n13340 | n21191 ;
  assign n21193 = ( ~n3022 & n9926 ) | ( ~n3022 & n20599 ) | ( n9926 & n20599 ) ;
  assign n21194 = ( ~n1203 & n4351 ) | ( ~n1203 & n9416 ) | ( n4351 & n9416 ) ;
  assign n21195 = n8887 ^ n7077 ^ 1'b0 ;
  assign n21196 = n9007 ^ n4904 ^ n1430 ;
  assign n21197 = n15201 & ~n21196 ;
  assign n21198 = n21197 ^ n2426 ^ 1'b0 ;
  assign n21199 = n1113 & n16903 ;
  assign n21200 = n21199 ^ n7899 ^ n3898 ;
  assign n21201 = n21200 ^ n4895 ^ 1'b0 ;
  assign n21202 = n10564 & n21201 ;
  assign n21203 = n5087 ^ n4933 ^ 1'b0 ;
  assign n21204 = ~n1972 & n21203 ;
  assign n21205 = n13884 & n21204 ;
  assign n21206 = n21205 ^ n4741 ^ 1'b0 ;
  assign n21207 = n21206 ^ n12576 ^ n3744 ;
  assign n21208 = ( n3117 & n15339 ) | ( n3117 & ~n21207 ) | ( n15339 & ~n21207 ) ;
  assign n21209 = n18298 ^ n4138 ^ n3835 ;
  assign n21210 = n21209 ^ n15129 ^ n5411 ;
  assign n21211 = n17556 ^ n10740 ^ 1'b0 ;
  assign n21212 = ( n5646 & n7343 ) | ( n5646 & n16874 ) | ( n7343 & n16874 ) ;
  assign n21213 = n4819 & ~n20366 ;
  assign n21214 = n18354 ^ n13527 ^ 1'b0 ;
  assign n21215 = n17253 & ~n21214 ;
  assign n21216 = n513 & n21215 ;
  assign n21217 = n21216 ^ n14328 ^ 1'b0 ;
  assign n21218 = n19028 ^ n11478 ^ n2142 ;
  assign n21219 = n21218 ^ n16392 ^ 1'b0 ;
  assign n21220 = n17843 | n21219 ;
  assign n21221 = ( n1465 & n8150 ) | ( n1465 & n10473 ) | ( n8150 & n10473 ) ;
  assign n21222 = ( n8782 & n11641 ) | ( n8782 & ~n17974 ) | ( n11641 & ~n17974 ) ;
  assign n21223 = n21221 | n21222 ;
  assign n21224 = ~n7992 & n11263 ;
  assign n21225 = n21223 & n21224 ;
  assign n21226 = ~n9436 & n15682 ;
  assign n21227 = n4771 ^ n4430 ^ x39 ;
  assign n21228 = n12078 ^ n11188 ^ n3603 ;
  assign n21229 = ( n8676 & n21227 ) | ( n8676 & n21228 ) | ( n21227 & n21228 ) ;
  assign n21230 = ( ~n4820 & n8138 ) | ( ~n4820 & n14848 ) | ( n8138 & n14848 ) ;
  assign n21231 = n21230 ^ n4359 ^ n1650 ;
  assign n21233 = n1282 ^ n952 ^ 1'b0 ;
  assign n21234 = n7630 | n21233 ;
  assign n21235 = ( n8205 & ~n14070 ) | ( n8205 & n21234 ) | ( ~n14070 & n21234 ) ;
  assign n21232 = n2143 | n10589 ;
  assign n21236 = n21235 ^ n21232 ^ 1'b0 ;
  assign n21237 = ~n1597 & n13210 ;
  assign n21238 = ~n1276 & n21237 ;
  assign n21239 = n14638 ^ n13427 ^ 1'b0 ;
  assign n21240 = n10638 | n21239 ;
  assign n21241 = n11180 ^ n4499 ^ x90 ;
  assign n21242 = ( n9018 & n21240 ) | ( n9018 & ~n21241 ) | ( n21240 & ~n21241 ) ;
  assign n21243 = ~n20295 & n21242 ;
  assign n21244 = n21238 & n21243 ;
  assign n21245 = ( n1235 & ~n2977 ) | ( n1235 & n4309 ) | ( ~n2977 & n4309 ) ;
  assign n21246 = n4889 ^ n1867 ^ 1'b0 ;
  assign n21247 = n18536 & ~n21246 ;
  assign n21248 = n6353 & n11534 ;
  assign n21249 = n5793 & ~n8576 ;
  assign n21250 = n16732 | n21249 ;
  assign n21251 = n2283 | n21250 ;
  assign n21252 = ( n8522 & ~n15022 ) | ( n8522 & n21251 ) | ( ~n15022 & n21251 ) ;
  assign n21257 = n7979 ^ n5638 ^ 1'b0 ;
  assign n21258 = n21257 ^ n12328 ^ n8178 ;
  assign n21253 = n3200 ^ n370 ^ 1'b0 ;
  assign n21254 = n3365 & ~n21253 ;
  assign n21255 = n4787 & n10069 ;
  assign n21256 = ~n21254 & n21255 ;
  assign n21259 = n21258 ^ n21256 ^ n14019 ;
  assign n21260 = ( ~n17644 & n19746 ) | ( ~n17644 & n21259 ) | ( n19746 & n21259 ) ;
  assign n21261 = ( n5204 & n15486 ) | ( n5204 & n20677 ) | ( n15486 & n20677 ) ;
  assign n21262 = n21261 ^ n6980 ^ n623 ;
  assign n21263 = n4075 | n12811 ;
  assign n21264 = ( n4948 & n12143 ) | ( n4948 & ~n21263 ) | ( n12143 & ~n21263 ) ;
  assign n21265 = n5629 | n21264 ;
  assign n21266 = n12098 ^ n4200 ^ n505 ;
  assign n21267 = n21266 ^ n20724 ^ n5186 ;
  assign n21268 = n1499 & ~n18664 ;
  assign n21271 = ( n1880 & n2356 ) | ( n1880 & ~n3344 ) | ( n2356 & ~n3344 ) ;
  assign n21270 = n14234 ^ n13556 ^ n1492 ;
  assign n21272 = n21271 ^ n21270 ^ n5155 ;
  assign n21269 = ( ~n8157 & n15932 ) | ( ~n8157 & n16092 ) | ( n15932 & n16092 ) ;
  assign n21273 = n21272 ^ n21269 ^ n10874 ;
  assign n21274 = n21273 ^ n5704 ^ 1'b0 ;
  assign n21275 = n4345 | n19373 ;
  assign n21276 = n19233 | n21275 ;
  assign n21277 = n21276 ^ n8847 ^ n4298 ;
  assign n21278 = ( ~n11831 & n12679 ) | ( ~n11831 & n21079 ) | ( n12679 & n21079 ) ;
  assign n21279 = ( ~n6029 & n9869 ) | ( ~n6029 & n21278 ) | ( n9869 & n21278 ) ;
  assign n21280 = n14744 ^ n7402 ^ n4793 ;
  assign n21281 = ( ~n4329 & n17341 ) | ( ~n4329 & n21280 ) | ( n17341 & n21280 ) ;
  assign n21282 = ( n17051 & ~n21279 ) | ( n17051 & n21281 ) | ( ~n21279 & n21281 ) ;
  assign n21283 = n8740 | n16964 ;
  assign n21284 = n13216 & ~n21283 ;
  assign n21285 = n14127 | n18339 ;
  assign n21286 = n21285 ^ n4322 ^ 1'b0 ;
  assign n21287 = n14041 ^ n4948 ^ 1'b0 ;
  assign n21288 = ~n3215 & n21287 ;
  assign n21289 = n9242 & n21288 ;
  assign n21290 = ~n7180 & n8344 ;
  assign n21291 = n12983 & n21290 ;
  assign n21292 = ~n18686 & n21291 ;
  assign n21293 = ~n8663 & n16791 ;
  assign n21294 = n21293 ^ n1678 ^ 1'b0 ;
  assign n21295 = ( n12654 & n21292 ) | ( n12654 & ~n21294 ) | ( n21292 & ~n21294 ) ;
  assign n21296 = ( n19971 & n21289 ) | ( n19971 & n21295 ) | ( n21289 & n21295 ) ;
  assign n21297 = ( n6285 & ~n7131 ) | ( n6285 & n12985 ) | ( ~n7131 & n12985 ) ;
  assign n21298 = ( x174 & x242 ) | ( x174 & n4559 ) | ( x242 & n4559 ) ;
  assign n21299 = ( n5980 & n20135 ) | ( n5980 & ~n21298 ) | ( n20135 & ~n21298 ) ;
  assign n21300 = n21299 ^ n17266 ^ 1'b0 ;
  assign n21301 = n5184 | n21300 ;
  assign n21303 = n1043 & n1870 ;
  assign n21302 = n15164 | n17110 ;
  assign n21304 = n21303 ^ n21302 ^ 1'b0 ;
  assign n21305 = ( ~n4434 & n14692 ) | ( ~n4434 & n21304 ) | ( n14692 & n21304 ) ;
  assign n21306 = n5206 ^ n5076 ^ 1'b0 ;
  assign n21307 = n11886 & ~n21306 ;
  assign n21308 = n5657 & n21307 ;
  assign n21309 = ( n1304 & ~n1708 ) | ( n1304 & n8457 ) | ( ~n1708 & n8457 ) ;
  assign n21310 = n21309 ^ n3188 ^ n1447 ;
  assign n21311 = n15631 | n21310 ;
  assign n21312 = n5382 | n21311 ;
  assign n21313 = n1232 | n7493 ;
  assign n21314 = n15089 & n21313 ;
  assign n21315 = n9389 ^ n418 ^ 1'b0 ;
  assign n21316 = n21315 ^ n11830 ^ n2434 ;
  assign n21317 = n21316 ^ n12351 ^ n6339 ;
  assign n21318 = n12882 ^ n3050 ^ n483 ;
  assign n21319 = n11514 ^ n2210 ^ 1'b0 ;
  assign n21320 = ~n21318 & n21319 ;
  assign n21321 = n9053 ^ n3274 ^ n1139 ;
  assign n21322 = n16625 ^ n9263 ^ 1'b0 ;
  assign n21323 = n21321 & ~n21322 ;
  assign n21324 = ( n6893 & ~n13368 ) | ( n6893 & n18179 ) | ( ~n13368 & n18179 ) ;
  assign n21325 = n20582 ^ n3121 ^ 1'b0 ;
  assign n21326 = ( n3204 & n15677 ) | ( n3204 & n17046 ) | ( n15677 & n17046 ) ;
  assign n21327 = n21326 ^ n12017 ^ n11904 ;
  assign n21328 = n21327 ^ n18612 ^ 1'b0 ;
  assign n21329 = ~n2604 & n21328 ;
  assign n21330 = n10412 ^ n1462 ^ 1'b0 ;
  assign n21331 = n21330 ^ n12500 ^ 1'b0 ;
  assign n21333 = n7973 ^ n6273 ^ 1'b0 ;
  assign n21334 = ~n14618 & n21333 ;
  assign n21335 = n21334 ^ n12323 ^ 1'b0 ;
  assign n21336 = n13144 | n21335 ;
  assign n21337 = n17258 | n21336 ;
  assign n21332 = n779 & ~n2562 ;
  assign n21338 = n21337 ^ n21332 ^ n7638 ;
  assign n21339 = n19103 ^ n13157 ^ n10774 ;
  assign n21340 = n10548 ^ n933 ^ n433 ;
  assign n21341 = n16318 ^ n13327 ^ n1279 ;
  assign n21342 = n21341 ^ n11155 ^ n1156 ;
  assign n21343 = ~n11496 & n21342 ;
  assign n21344 = ~n5475 & n21343 ;
  assign n21347 = ~n11755 & n13886 ;
  assign n21345 = n6654 & n8494 ;
  assign n21346 = n21345 ^ n11806 ^ 1'b0 ;
  assign n21348 = n21347 ^ n21346 ^ n14695 ;
  assign n21349 = ( ~n21340 & n21344 ) | ( ~n21340 & n21348 ) | ( n21344 & n21348 ) ;
  assign n21350 = n17699 ^ n8109 ^ n5738 ;
  assign n21351 = n3094 & ~n10480 ;
  assign n21352 = ~n6793 & n21351 ;
  assign n21353 = n14036 ^ n4244 ^ n3210 ;
  assign n21354 = n21352 & ~n21353 ;
  assign n21355 = ( ~n695 & n10809 ) | ( ~n695 & n15378 ) | ( n10809 & n15378 ) ;
  assign n21356 = n5952 & n21355 ;
  assign n21357 = n10172 & n21356 ;
  assign n21363 = ( n446 & n8403 ) | ( n446 & ~n17592 ) | ( n8403 & ~n17592 ) ;
  assign n21358 = n21133 ^ n19583 ^ n4721 ;
  assign n21359 = ( n1276 & ~n2183 ) | ( n1276 & n5730 ) | ( ~n2183 & n5730 ) ;
  assign n21360 = n16977 ^ n10311 ^ 1'b0 ;
  assign n21361 = n21359 & n21360 ;
  assign n21362 = ( ~n17226 & n21358 ) | ( ~n17226 & n21361 ) | ( n21358 & n21361 ) ;
  assign n21364 = n21363 ^ n21362 ^ 1'b0 ;
  assign n21365 = ~n12976 & n21364 ;
  assign n21366 = n11878 ^ n9580 ^ n4189 ;
  assign n21367 = n309 & ~n19106 ;
  assign n21368 = ( n12190 & ~n21366 ) | ( n12190 & n21367 ) | ( ~n21366 & n21367 ) ;
  assign n21369 = n21368 ^ n13347 ^ 1'b0 ;
  assign n21370 = n17912 & ~n21369 ;
  assign n21371 = n21370 ^ n13731 ^ n8895 ;
  assign n21372 = n17638 ^ n8109 ^ 1'b0 ;
  assign n21373 = n4416 & n21372 ;
  assign n21374 = n21373 ^ n18400 ^ n17783 ;
  assign n21375 = ( n2793 & n8013 ) | ( n2793 & n12243 ) | ( n8013 & n12243 ) ;
  assign n21377 = ( n6301 & n13364 ) | ( n6301 & ~n16227 ) | ( n13364 & ~n16227 ) ;
  assign n21378 = n3613 & ~n21377 ;
  assign n21376 = n16586 ^ n9498 ^ n5961 ;
  assign n21379 = n21378 ^ n21376 ^ n12147 ;
  assign n21380 = ( ~n5001 & n20313 ) | ( ~n5001 & n21379 ) | ( n20313 & n21379 ) ;
  assign n21381 = n21380 ^ n6275 ^ 1'b0 ;
  assign n21382 = ~n21375 & n21381 ;
  assign n21383 = n7203 | n17605 ;
  assign n21384 = n21383 ^ n4786 ^ 1'b0 ;
  assign n21385 = n17872 ^ n12859 ^ n9618 ;
  assign n21386 = ( n1025 & ~n1569 ) | ( n1025 & n21385 ) | ( ~n1569 & n21385 ) ;
  assign n21387 = ( ~n427 & n4760 ) | ( ~n427 & n7162 ) | ( n4760 & n7162 ) ;
  assign n21388 = ( n2014 & n7932 ) | ( n2014 & n21387 ) | ( n7932 & n21387 ) ;
  assign n21389 = n8323 & n21388 ;
  assign n21390 = n21389 ^ n9145 ^ 1'b0 ;
  assign n21391 = n21390 ^ n11868 ^ 1'b0 ;
  assign n21392 = n17905 & n21391 ;
  assign n21393 = n21392 ^ n13769 ^ n9431 ;
  assign n21394 = n21393 ^ n9667 ^ 1'b0 ;
  assign n21395 = n16790 ^ n10873 ^ n5416 ;
  assign n21396 = n6351 & ~n21395 ;
  assign n21397 = n18226 ^ n13564 ^ 1'b0 ;
  assign n21404 = ( n684 & ~n7042 ) | ( n684 & n9378 ) | ( ~n7042 & n9378 ) ;
  assign n21405 = n1505 | n21404 ;
  assign n21399 = n15505 ^ n8740 ^ 1'b0 ;
  assign n21398 = n2096 | n7139 ;
  assign n21400 = n21399 ^ n21398 ^ 1'b0 ;
  assign n21401 = n21400 ^ n7664 ^ 1'b0 ;
  assign n21402 = n9906 & n12972 ;
  assign n21403 = n21401 & n21402 ;
  assign n21406 = n21405 ^ n21403 ^ 1'b0 ;
  assign n21407 = n21406 ^ n11283 ^ n1851 ;
  assign n21408 = n18727 ^ n10850 ^ n6583 ;
  assign n21409 = ( n450 & ~n2800 ) | ( n450 & n21408 ) | ( ~n2800 & n21408 ) ;
  assign n21410 = n21409 ^ n20336 ^ n7899 ;
  assign n21411 = n9861 & n21410 ;
  assign n21412 = n9645 ^ n1052 ^ 1'b0 ;
  assign n21413 = n21412 ^ n17468 ^ 1'b0 ;
  assign n21414 = n6527 & ~n17808 ;
  assign n21415 = n21414 ^ n12272 ^ 1'b0 ;
  assign n21416 = ( n16706 & n17880 ) | ( n16706 & ~n21415 ) | ( n17880 & ~n21415 ) ;
  assign n21417 = n15465 ^ n8558 ^ 1'b0 ;
  assign n21418 = ~n21416 & n21417 ;
  assign n21419 = n2460 & n17574 ;
  assign n21421 = n10177 ^ n7354 ^ n6072 ;
  assign n21420 = n1239 & n5376 ;
  assign n21422 = n21421 ^ n21420 ^ 1'b0 ;
  assign n21423 = ( n11366 & n21419 ) | ( n11366 & ~n21422 ) | ( n21419 & ~n21422 ) ;
  assign n21424 = n494 | n3106 ;
  assign n21425 = ( ~n4245 & n9128 ) | ( ~n4245 & n20844 ) | ( n9128 & n20844 ) ;
  assign n21426 = n2475 | n16103 ;
  assign n21427 = n9336 & ~n21426 ;
  assign n21428 = n16226 ^ n2187 ^ 1'b0 ;
  assign n21430 = n17391 ^ n11642 ^ n8233 ;
  assign n21429 = n1478 & n1974 ;
  assign n21431 = n21430 ^ n21429 ^ 1'b0 ;
  assign n21432 = n21431 ^ n3801 ^ 1'b0 ;
  assign n21433 = n2604 | n21432 ;
  assign n21434 = n21428 | n21433 ;
  assign n21435 = n10858 & ~n11650 ;
  assign n21436 = ~n5781 & n21435 ;
  assign n21437 = n10274 | n21436 ;
  assign n21438 = n12346 | n21437 ;
  assign n21439 = n16296 ^ n445 ^ 1'b0 ;
  assign n21440 = n2510 | n11736 ;
  assign n21441 = n7491 | n21440 ;
  assign n21442 = ( n7899 & n17578 ) | ( n7899 & ~n21441 ) | ( n17578 & ~n21441 ) ;
  assign n21443 = ~n21439 & n21442 ;
  assign n21444 = n21443 ^ n8094 ^ 1'b0 ;
  assign n21445 = ( n5361 & n10127 ) | ( n5361 & n11982 ) | ( n10127 & n11982 ) ;
  assign n21446 = x57 | n21445 ;
  assign n21447 = n3346 | n11702 ;
  assign n21448 = n21446 | n21447 ;
  assign n21449 = n10770 ^ n10695 ^ n8397 ;
  assign n21450 = ( n20139 & n21448 ) | ( n20139 & n21449 ) | ( n21448 & n21449 ) ;
  assign n21451 = ~n3638 & n4162 ;
  assign n21452 = n19678 ^ n2864 ^ n2167 ;
  assign n21453 = n17489 & ~n21452 ;
  assign n21454 = n10786 ^ n8222 ^ 1'b0 ;
  assign n21455 = ~n21453 & n21454 ;
  assign n21456 = ( n681 & n1020 ) | ( n681 & n9230 ) | ( n1020 & n9230 ) ;
  assign n21457 = n21456 ^ n3535 ^ n257 ;
  assign n21458 = ( n1923 & ~n3440 ) | ( n1923 & n3470 ) | ( ~n3440 & n3470 ) ;
  assign n21459 = n3106 & ~n21458 ;
  assign n21460 = n11166 & n21459 ;
  assign n21461 = n21460 ^ n15552 ^ 1'b0 ;
  assign n21462 = ~n21457 & n21461 ;
  assign n21463 = n21462 ^ n10278 ^ 1'b0 ;
  assign n21464 = n21455 & ~n21463 ;
  assign n21465 = ( n6494 & n8205 ) | ( n6494 & n13080 ) | ( n8205 & n13080 ) ;
  assign n21466 = n972 & ~n1521 ;
  assign n21467 = n21466 ^ n2014 ^ 1'b0 ;
  assign n21468 = n4753 | n10897 ;
  assign n21469 = n21468 ^ n6065 ^ 1'b0 ;
  assign n21470 = ( n3402 & n6994 ) | ( n3402 & n9512 ) | ( n6994 & n9512 ) ;
  assign n21471 = n13741 ^ n11914 ^ 1'b0 ;
  assign n21472 = n5272 ^ n3483 ^ n1997 ;
  assign n21473 = ( n15213 & n21471 ) | ( n15213 & ~n21472 ) | ( n21471 & ~n21472 ) ;
  assign n21474 = ( n695 & n21470 ) | ( n695 & ~n21473 ) | ( n21470 & ~n21473 ) ;
  assign n21475 = n4365 | n15086 ;
  assign n21476 = ( n3536 & n6462 ) | ( n3536 & ~n8794 ) | ( n6462 & ~n8794 ) ;
  assign n21477 = n21476 ^ n10619 ^ 1'b0 ;
  assign n21478 = ( n15148 & ~n21475 ) | ( n15148 & n21477 ) | ( ~n21475 & n21477 ) ;
  assign n21479 = ~n533 & n3623 ;
  assign n21480 = n21479 ^ n4764 ^ 1'b0 ;
  assign n21481 = n2784 | n10500 ;
  assign n21482 = n21481 ^ n15616 ^ n7468 ;
  assign n21483 = ( n5803 & n21480 ) | ( n5803 & ~n21482 ) | ( n21480 & ~n21482 ) ;
  assign n21484 = n12513 ^ n3140 ^ n1570 ;
  assign n21485 = ( n707 & n4062 ) | ( n707 & ~n5651 ) | ( n4062 & ~n5651 ) ;
  assign n21486 = ( n14874 & n19155 ) | ( n14874 & n21485 ) | ( n19155 & n21485 ) ;
  assign n21487 = n16654 ^ n14459 ^ n485 ;
  assign n21488 = n4555 ^ n3792 ^ 1'b0 ;
  assign n21489 = ~n21487 & n21488 ;
  assign n21490 = ~n6107 & n16525 ;
  assign n21491 = n21490 ^ n3546 ^ 1'b0 ;
  assign n21492 = n21489 & n21491 ;
  assign n21493 = n454 & n21492 ;
  assign n21494 = ( n11343 & n12318 ) | ( n11343 & ~n13095 ) | ( n12318 & ~n13095 ) ;
  assign n21495 = n19812 ^ n3109 ^ 1'b0 ;
  assign n21496 = n16868 | n21495 ;
  assign n21497 = n4418 ^ n2306 ^ n1630 ;
  assign n21498 = n1638 & ~n21497 ;
  assign n21499 = n21498 ^ n11219 ^ 1'b0 ;
  assign n21500 = ( n6857 & n7527 ) | ( n6857 & ~n15719 ) | ( n7527 & ~n15719 ) ;
  assign n21501 = n5218 & ~n6033 ;
  assign n21502 = n946 ^ x159 ^ 1'b0 ;
  assign n21503 = ( n14207 & ~n14922 ) | ( n14207 & n21502 ) | ( ~n14922 & n21502 ) ;
  assign n21504 = n12890 & ~n21503 ;
  assign n21505 = ( n5702 & ~n5965 ) | ( n5702 & n10222 ) | ( ~n5965 & n10222 ) ;
  assign n21506 = ~n17032 & n21505 ;
  assign n21507 = n21506 ^ n9922 ^ 1'b0 ;
  assign n21508 = n12872 & ~n13722 ;
  assign n21509 = n21508 ^ n5146 ^ 1'b0 ;
  assign n21510 = n21509 ^ n6564 ^ n3804 ;
  assign n21511 = x150 | n21510 ;
  assign n21512 = n11478 & ~n21511 ;
  assign n21513 = n3911 | n21512 ;
  assign n21514 = n21513 ^ n7369 ^ 1'b0 ;
  assign n21515 = ~n16678 & n20563 ;
  assign n21516 = n21515 ^ n4559 ^ 1'b0 ;
  assign n21518 = ~n697 & n12055 ;
  assign n21517 = n3515 & ~n14022 ;
  assign n21519 = n21518 ^ n21517 ^ n2988 ;
  assign n21520 = ~n2520 & n14787 ;
  assign n21521 = n21520 ^ n2924 ^ 1'b0 ;
  assign n21522 = n21521 ^ n15409 ^ n10961 ;
  assign n21523 = n21522 ^ n17951 ^ 1'b0 ;
  assign n21525 = n3298 ^ n3253 ^ n1018 ;
  assign n21526 = ( ~n2407 & n10124 ) | ( ~n2407 & n21525 ) | ( n10124 & n21525 ) ;
  assign n21527 = n21526 ^ n12344 ^ n10058 ;
  assign n21524 = n9998 ^ n6523 ^ 1'b0 ;
  assign n21528 = n21527 ^ n21524 ^ n4038 ;
  assign n21529 = ( ~n1797 & n5885 ) | ( ~n1797 & n21528 ) | ( n5885 & n21528 ) ;
  assign n21530 = ( n4399 & n4771 ) | ( n4399 & n14998 ) | ( n4771 & n14998 ) ;
  assign n21531 = n11552 ^ n7221 ^ n397 ;
  assign n21532 = ( n1246 & ~n5355 ) | ( n1246 & n12466 ) | ( ~n5355 & n12466 ) ;
  assign n21533 = ( n4574 & n8719 ) | ( n4574 & ~n16882 ) | ( n8719 & ~n16882 ) ;
  assign n21534 = ( n21079 & ~n21532 ) | ( n21079 & n21533 ) | ( ~n21532 & n21533 ) ;
  assign n21535 = n387 & ~n21534 ;
  assign n21540 = ( n4061 & ~n10138 ) | ( n4061 & n18428 ) | ( ~n10138 & n18428 ) ;
  assign n21541 = ~n15998 & n20840 ;
  assign n21542 = ~n21540 & n21541 ;
  assign n21536 = n10281 ^ n7490 ^ n4458 ;
  assign n21537 = ( n14188 & n14787 ) | ( n14188 & ~n21536 ) | ( n14787 & ~n21536 ) ;
  assign n21538 = n21537 ^ n7840 ^ 1'b0 ;
  assign n21539 = n8306 & n21538 ;
  assign n21543 = n21542 ^ n21539 ^ 1'b0 ;
  assign n21544 = ( ~n3487 & n5385 ) | ( ~n3487 & n15221 ) | ( n5385 & n15221 ) ;
  assign n21545 = n7729 ^ n2337 ^ 1'b0 ;
  assign n21546 = n872 & n8266 ;
  assign n21547 = n8880 & ~n21546 ;
  assign n21548 = n21547 ^ n18420 ^ 1'b0 ;
  assign n21549 = n2355 & n11850 ;
  assign n21550 = n21549 ^ n4855 ^ 1'b0 ;
  assign n21551 = n19183 ^ n14875 ^ n14466 ;
  assign n21552 = n9176 ^ n1305 ^ 1'b0 ;
  assign n21553 = ~n2412 & n21552 ;
  assign n21554 = ~n17969 & n21553 ;
  assign n21555 = ( n5330 & n10862 ) | ( n5330 & n21554 ) | ( n10862 & n21554 ) ;
  assign n21556 = n17081 ^ n13305 ^ n9717 ;
  assign n21557 = n21556 ^ n19424 ^ n16022 ;
  assign n21558 = ( n4504 & n6748 ) | ( n4504 & n21557 ) | ( n6748 & n21557 ) ;
  assign n21559 = n9757 ^ n894 ^ 1'b0 ;
  assign n21560 = n20863 ^ n7746 ^ n2104 ;
  assign n21561 = ( ~n9189 & n12551 ) | ( ~n9189 & n21560 ) | ( n12551 & n21560 ) ;
  assign n21562 = ~n5562 & n14406 ;
  assign n21563 = n21562 ^ n2865 ^ 1'b0 ;
  assign n21564 = n21561 & ~n21563 ;
  assign n21565 = n5803 & n8695 ;
  assign n21566 = n12112 & n21565 ;
  assign n21567 = ( ~n1592 & n13979 ) | ( ~n1592 & n17414 ) | ( n13979 & n17414 ) ;
  assign n21568 = ( n2513 & n21566 ) | ( n2513 & ~n21567 ) | ( n21566 & ~n21567 ) ;
  assign n21569 = n13865 ^ n7663 ^ 1'b0 ;
  assign n21570 = ~n816 & n5245 ;
  assign n21571 = ( n4495 & n5102 ) | ( n4495 & ~n21570 ) | ( n5102 & ~n21570 ) ;
  assign n21577 = n9178 ^ n5236 ^ n386 ;
  assign n21578 = ( n1822 & ~n3097 ) | ( n1822 & n21577 ) | ( ~n3097 & n21577 ) ;
  assign n21579 = n21578 ^ n12044 ^ n9518 ;
  assign n21572 = ( n954 & ~n5468 ) | ( n954 & n9955 ) | ( ~n5468 & n9955 ) ;
  assign n21573 = n21572 ^ n7633 ^ n6637 ;
  assign n21574 = n21573 ^ n11873 ^ n4046 ;
  assign n21575 = ~n1883 & n21574 ;
  assign n21576 = n21575 ^ n16103 ^ 1'b0 ;
  assign n21580 = n21579 ^ n21576 ^ n13921 ;
  assign n21581 = n9213 ^ n7097 ^ 1'b0 ;
  assign n21582 = ~n20779 & n21581 ;
  assign n21583 = ( n12499 & n21580 ) | ( n12499 & ~n21582 ) | ( n21580 & ~n21582 ) ;
  assign n21584 = n19533 ^ n3703 ^ n1307 ;
  assign n21585 = n11616 ^ n4471 ^ n1228 ;
  assign n21586 = n17490 & n21585 ;
  assign n21587 = n21586 ^ n2139 ^ 1'b0 ;
  assign n21588 = ( n4635 & ~n8320 ) | ( n4635 & n21587 ) | ( ~n8320 & n21587 ) ;
  assign n21589 = n9005 | n21588 ;
  assign n21590 = n21589 ^ n9484 ^ 1'b0 ;
  assign n21592 = n4166 | n18466 ;
  assign n21591 = ( n2394 & n3357 ) | ( n2394 & ~n4471 ) | ( n3357 & ~n4471 ) ;
  assign n21593 = n21592 ^ n21591 ^ n12616 ;
  assign n21595 = n20926 ^ n7659 ^ 1'b0 ;
  assign n21594 = n12909 ^ n7409 ^ n2238 ;
  assign n21596 = n21595 ^ n21594 ^ n19829 ;
  assign n21597 = n18239 ^ n11637 ^ 1'b0 ;
  assign n21598 = n7193 & ~n8341 ;
  assign n21599 = n21598 ^ n13618 ^ 1'b0 ;
  assign n21600 = n1494 ^ x28 ^ 1'b0 ;
  assign n21601 = ( n4257 & n21599 ) | ( n4257 & ~n21600 ) | ( n21599 & ~n21600 ) ;
  assign n21602 = n4750 ^ n4111 ^ 1'b0 ;
  assign n21603 = n17415 ^ n3450 ^ 1'b0 ;
  assign n21604 = n16247 & n21603 ;
  assign n21605 = n5572 | n19309 ;
  assign n21606 = n4767 & ~n21605 ;
  assign n21607 = n15609 ^ n12984 ^ 1'b0 ;
  assign n21608 = ( n7329 & n21606 ) | ( n7329 & ~n21607 ) | ( n21606 & ~n21607 ) ;
  assign n21609 = ( n1002 & n17489 ) | ( n1002 & ~n21458 ) | ( n17489 & ~n21458 ) ;
  assign n21610 = n21609 ^ n10083 ^ n4927 ;
  assign n21611 = n3764 | n21610 ;
  assign n21612 = n7023 & ~n21611 ;
  assign n21613 = n19023 ^ n2812 ^ 1'b0 ;
  assign n21614 = n13863 ^ n10602 ^ 1'b0 ;
  assign n21615 = n21614 ^ n11673 ^ n4641 ;
  assign n21616 = n10318 & ~n21615 ;
  assign n21617 = ( n4298 & n12737 ) | ( n4298 & ~n21616 ) | ( n12737 & ~n21616 ) ;
  assign n21618 = n3087 | n5701 ;
  assign n21619 = n21618 ^ n12995 ^ 1'b0 ;
  assign n21620 = x213 | n7417 ;
  assign n21621 = n21620 ^ n12788 ^ n5259 ;
  assign n21622 = ~n2412 & n15933 ;
  assign n21623 = ( n12292 & n19606 ) | ( n12292 & ~n21622 ) | ( n19606 & ~n21622 ) ;
  assign n21624 = ( n2187 & ~n7198 ) | ( n2187 & n7915 ) | ( ~n7198 & n7915 ) ;
  assign n21628 = n9672 ^ n6938 ^ 1'b0 ;
  assign n21629 = n21628 ^ n18013 ^ n5791 ;
  assign n21626 = n3190 & n10481 ;
  assign n21625 = n1643 | n7888 ;
  assign n21627 = n21626 ^ n21625 ^ 1'b0 ;
  assign n21630 = n21629 ^ n21627 ^ 1'b0 ;
  assign n21631 = ~n21624 & n21630 ;
  assign n21632 = n1841 | n6230 ;
  assign n21633 = n15336 ^ n14545 ^ n5163 ;
  assign n21634 = n14386 | n18520 ;
  assign n21635 = n21634 ^ n5420 ^ 1'b0 ;
  assign n21636 = n12175 ^ n5905 ^ 1'b0 ;
  assign n21637 = n17880 | n21636 ;
  assign n21638 = n15835 ^ n5653 ^ 1'b0 ;
  assign n21639 = ( n1713 & ~n15201 ) | ( n1713 & n21638 ) | ( ~n15201 & n21638 ) ;
  assign n21640 = n21639 ^ n14980 ^ 1'b0 ;
  assign n21641 = n9500 & n21640 ;
  assign n21642 = ( n353 & n900 ) | ( n353 & n20085 ) | ( n900 & n20085 ) ;
  assign n21643 = n6374 | n12093 ;
  assign n21644 = n21643 ^ n5249 ^ 1'b0 ;
  assign n21645 = ( n14115 & ~n21642 ) | ( n14115 & n21644 ) | ( ~n21642 & n21644 ) ;
  assign n21646 = ( n10756 & n18872 ) | ( n10756 & n19519 ) | ( n18872 & n19519 ) ;
  assign n21647 = ( ~n480 & n9216 ) | ( ~n480 & n15084 ) | ( n9216 & n15084 ) ;
  assign n21648 = n21647 ^ n15393 ^ n8403 ;
  assign n21649 = n4804 ^ n2143 ^ 1'b0 ;
  assign n21650 = n21649 ^ n9467 ^ n6879 ;
  assign n21651 = n17251 ^ n6442 ^ n1783 ;
  assign n21652 = n21651 ^ n12385 ^ 1'b0 ;
  assign n21653 = ( n880 & n21650 ) | ( n880 & ~n21652 ) | ( n21650 & ~n21652 ) ;
  assign n21654 = n21653 ^ n17115 ^ 1'b0 ;
  assign n21655 = n21648 & n21654 ;
  assign n21656 = ( ~n1769 & n21646 ) | ( ~n1769 & n21655 ) | ( n21646 & n21655 ) ;
  assign n21657 = n6864 | n11025 ;
  assign n21658 = n11119 | n21657 ;
  assign n21659 = n9080 | n21658 ;
  assign n21660 = ( x78 & n3737 ) | ( x78 & n7610 ) | ( n3737 & n7610 ) ;
  assign n21661 = n21660 ^ n939 ^ 1'b0 ;
  assign n21662 = ( n347 & n10537 ) | ( n347 & ~n21661 ) | ( n10537 & ~n21661 ) ;
  assign n21663 = ~n2048 & n8794 ;
  assign n21664 = ~n21662 & n21663 ;
  assign n21665 = n4579 ^ n1703 ^ 1'b0 ;
  assign n21666 = ( n3666 & n4284 ) | ( n3666 & ~n21665 ) | ( n4284 & ~n21665 ) ;
  assign n21667 = ( ~n2782 & n6004 ) | ( ~n2782 & n11771 ) | ( n6004 & n11771 ) ;
  assign n21668 = n6863 ^ n3889 ^ 1'b0 ;
  assign n21669 = ( n12888 & ~n15182 ) | ( n12888 & n19275 ) | ( ~n15182 & n19275 ) ;
  assign n21670 = n3484 & ~n21669 ;
  assign n21671 = ~n21668 & n21670 ;
  assign n21672 = n10813 & n21671 ;
  assign n21673 = n15313 | n20031 ;
  assign n21674 = n13913 | n21673 ;
  assign n21675 = ~n12235 & n21674 ;
  assign n21676 = n1304 | n3920 ;
  assign n21677 = ~n4134 & n21676 ;
  assign n21678 = n10363 | n21677 ;
  assign n21679 = n21678 ^ n18107 ^ 1'b0 ;
  assign n21680 = n12157 ^ n311 ^ 1'b0 ;
  assign n21681 = n5270 & ~n8739 ;
  assign n21682 = ~n5906 & n21681 ;
  assign n21683 = ( n1542 & n5687 ) | ( n1542 & n21682 ) | ( n5687 & n21682 ) ;
  assign n21684 = n21683 ^ n10216 ^ 1'b0 ;
  assign n21685 = n19580 & n21684 ;
  assign n21686 = ( x94 & ~n17707 ) | ( x94 & n21685 ) | ( ~n17707 & n21685 ) ;
  assign n21687 = n5956 | n14274 ;
  assign n21688 = n21687 ^ n13902 ^ 1'b0 ;
  assign n21689 = n17964 ^ n8484 ^ 1'b0 ;
  assign n21690 = ~n3230 & n17319 ;
  assign n21691 = ~n4893 & n21690 ;
  assign n21692 = n16794 & ~n21691 ;
  assign n21694 = n8234 & ~n9677 ;
  assign n21695 = n21694 ^ n10896 ^ n631 ;
  assign n21696 = n13246 & n21695 ;
  assign n21693 = n2992 & n14197 ;
  assign n21697 = n21696 ^ n21693 ^ n4759 ;
  assign n21698 = n21697 ^ n7119 ^ n3397 ;
  assign n21699 = n21698 ^ n15243 ^ 1'b0 ;
  assign n21700 = n7987 & n21699 ;
  assign n21702 = n938 & n10350 ;
  assign n21703 = ~n1760 & n21702 ;
  assign n21701 = ~n2708 & n9039 ;
  assign n21704 = n21703 ^ n21701 ^ 1'b0 ;
  assign n21709 = ( ~n6058 & n7497 ) | ( ~n6058 & n14169 ) | ( n7497 & n14169 ) ;
  assign n21710 = n21709 ^ n2305 ^ 1'b0 ;
  assign n21705 = ~n5115 & n9606 ;
  assign n21706 = ~n858 & n21705 ;
  assign n21707 = ( n1692 & ~n5705 ) | ( n1692 & n21706 ) | ( ~n5705 & n21706 ) ;
  assign n21708 = n21707 ^ n13652 ^ n4617 ;
  assign n21711 = n21710 ^ n21708 ^ 1'b0 ;
  assign n21713 = n9010 ^ n5277 ^ 1'b0 ;
  assign n21714 = n4976 | n21713 ;
  assign n21715 = n21714 ^ n2276 ^ 1'b0 ;
  assign n21712 = n3941 ^ x87 ^ 1'b0 ;
  assign n21716 = n21715 ^ n21712 ^ 1'b0 ;
  assign n21717 = ~n21711 & n21716 ;
  assign n21718 = n21717 ^ n19141 ^ n17388 ;
  assign n21719 = n15427 ^ n2962 ^ 1'b0 ;
  assign n21720 = ~n405 & n21719 ;
  assign n21721 = n21720 ^ n15159 ^ 1'b0 ;
  assign n21722 = n5403 & n21721 ;
  assign n21723 = n21722 ^ n11959 ^ 1'b0 ;
  assign n21724 = x133 & ~n21723 ;
  assign n21725 = ( ~n1636 & n19061 ) | ( ~n1636 & n21724 ) | ( n19061 & n21724 ) ;
  assign n21726 = ( n5468 & ~n7009 ) | ( n5468 & n21256 ) | ( ~n7009 & n21256 ) ;
  assign n21727 = n13010 ^ n11419 ^ n9389 ;
  assign n21728 = n460 & ~n21346 ;
  assign n21729 = ~n8812 & n21728 ;
  assign n21730 = n12053 ^ n9557 ^ n1950 ;
  assign n21733 = x186 & ~n11122 ;
  assign n21732 = n4092 & ~n6382 ;
  assign n21734 = n21733 ^ n21732 ^ n11876 ;
  assign n21731 = ( ~n504 & n2558 ) | ( ~n504 & n10195 ) | ( n2558 & n10195 ) ;
  assign n21735 = n21734 ^ n21731 ^ 1'b0 ;
  assign n21739 = n2755 | n18194 ;
  assign n21740 = n21739 ^ n11854 ^ 1'b0 ;
  assign n21736 = ( ~n8754 & n10585 ) | ( ~n8754 & n13090 ) | ( n10585 & n13090 ) ;
  assign n21737 = ( n883 & ~n10239 ) | ( n883 & n14085 ) | ( ~n10239 & n14085 ) ;
  assign n21738 = n21736 | n21737 ;
  assign n21741 = n21740 ^ n21738 ^ 1'b0 ;
  assign n21742 = n20582 ^ n17249 ^ 1'b0 ;
  assign n21743 = ( n15276 & n19849 ) | ( n15276 & ~n21742 ) | ( n19849 & ~n21742 ) ;
  assign n21744 = ( n3759 & n21741 ) | ( n3759 & ~n21743 ) | ( n21741 & ~n21743 ) ;
  assign n21745 = n7726 ^ n733 ^ 1'b0 ;
  assign n21746 = n10210 & n21745 ;
  assign n21747 = n3264 | n13847 ;
  assign n21749 = n2250 | n4659 ;
  assign n21750 = n896 & ~n21749 ;
  assign n21748 = n10105 ^ n4266 ^ 1'b0 ;
  assign n21751 = n21750 ^ n21748 ^ n11197 ;
  assign n21752 = n21209 ^ n18728 ^ n14334 ;
  assign n21754 = n4993 ^ n3184 ^ 1'b0 ;
  assign n21753 = n11774 ^ n9942 ^ n3781 ;
  assign n21755 = n21754 ^ n21753 ^ n15414 ;
  assign n21756 = x14 & n21755 ;
  assign n21757 = n21756 ^ n8887 ^ 1'b0 ;
  assign n21758 = n13190 ^ n2195 ^ 1'b0 ;
  assign n21759 = ~n3320 & n21758 ;
  assign n21760 = ~n665 & n2374 ;
  assign n21761 = n21760 ^ n1128 ^ 1'b0 ;
  assign n21762 = n1587 ^ x236 ^ 1'b0 ;
  assign n21763 = ~n17544 & n21762 ;
  assign n21764 = n7833 & n21763 ;
  assign n21765 = n21761 & n21764 ;
  assign n21766 = n15140 ^ n13609 ^ n2594 ;
  assign n21767 = n21766 ^ n9291 ^ n7977 ;
  assign n21770 = n6284 ^ n3529 ^ 1'b0 ;
  assign n21771 = n17144 & n21770 ;
  assign n21772 = ( n3658 & n16440 ) | ( n3658 & ~n21771 ) | ( n16440 & ~n21771 ) ;
  assign n21768 = n14455 ^ n5036 ^ 1'b0 ;
  assign n21769 = ~n18827 & n21768 ;
  assign n21773 = n21772 ^ n21769 ^ 1'b0 ;
  assign n21774 = n17584 ^ n5017 ^ n494 ;
  assign n21775 = n11588 ^ n1609 ^ 1'b0 ;
  assign n21776 = n21774 & n21775 ;
  assign n21777 = n7706 ^ n5061 ^ 1'b0 ;
  assign n21778 = n5439 & n21777 ;
  assign n21779 = n21778 ^ n6121 ^ 1'b0 ;
  assign n21780 = ~n4182 & n21779 ;
  assign n21781 = ( ~n8852 & n9921 ) | ( ~n8852 & n21780 ) | ( n9921 & n21780 ) ;
  assign n21782 = ~n6519 & n21781 ;
  assign n21783 = n12938 ^ n4282 ^ n576 ;
  assign n21784 = ( n6883 & n7956 ) | ( n6883 & n21783 ) | ( n7956 & n21783 ) ;
  assign n21785 = n18624 ^ n14520 ^ n290 ;
  assign n21786 = ( ~n722 & n1137 ) | ( ~n722 & n21785 ) | ( n1137 & n21785 ) ;
  assign n21787 = ~n6164 & n14769 ;
  assign n21788 = n5783 ^ n4487 ^ 1'b0 ;
  assign n21789 = n21788 ^ n13430 ^ n4804 ;
  assign n21790 = n21789 ^ n12060 ^ n896 ;
  assign n21792 = n12712 ^ n1897 ^ 1'b0 ;
  assign n21793 = n388 & n21792 ;
  assign n21791 = n13500 ^ n12543 ^ n1856 ;
  assign n21794 = n21793 ^ n21791 ^ n10430 ;
  assign n21795 = n21794 ^ n1216 ^ 1'b0 ;
  assign n21796 = n21790 & n21795 ;
  assign n21797 = ~n710 & n21796 ;
  assign n21798 = ~n5271 & n12285 ;
  assign n21799 = n5696 ^ n1812 ^ n477 ;
  assign n21800 = ( n15406 & n17091 ) | ( n15406 & n21799 ) | ( n17091 & n21799 ) ;
  assign n21801 = n20053 ^ n18945 ^ n6925 ;
  assign n21802 = n21801 ^ n6279 ^ 1'b0 ;
  assign n21803 = n2924 & ~n6887 ;
  assign n21804 = ~n2121 & n21803 ;
  assign n21805 = n12974 & n21804 ;
  assign n21806 = ~n3677 & n4724 ;
  assign n21807 = n21806 ^ n5467 ^ 1'b0 ;
  assign n21808 = n7680 & n16408 ;
  assign n21809 = n7088 & n21808 ;
  assign n21810 = n5788 & n12740 ;
  assign n21811 = n10205 & ~n21810 ;
  assign n21812 = n21809 & n21811 ;
  assign n21813 = n4598 & ~n9577 ;
  assign n21814 = n21813 ^ n16974 ^ 1'b0 ;
  assign n21815 = ( ~n18266 & n20851 ) | ( ~n18266 & n21814 ) | ( n20851 & n21814 ) ;
  assign n21816 = n17757 ^ n10146 ^ 1'b0 ;
  assign n21817 = n16967 & n21816 ;
  assign n21818 = ~n8721 & n13961 ;
  assign n21819 = n2230 & n21818 ;
  assign n21820 = n3313 & n21819 ;
  assign n21821 = ~n2168 & n16321 ;
  assign n21822 = n21821 ^ n18485 ^ 1'b0 ;
  assign n21823 = ( n10589 & ~n21820 ) | ( n10589 & n21822 ) | ( ~n21820 & n21822 ) ;
  assign n21824 = n21817 & ~n21823 ;
  assign n21825 = ( n7360 & n12977 ) | ( n7360 & ~n16921 ) | ( n12977 & ~n16921 ) ;
  assign n21826 = n21825 ^ n20267 ^ n7099 ;
  assign n21827 = n4430 & ~n16048 ;
  assign n21828 = n893 & ~n11514 ;
  assign n21829 = n21828 ^ n7379 ^ 1'b0 ;
  assign n21830 = n8684 & n21829 ;
  assign n21832 = n4003 ^ n1424 ^ 1'b0 ;
  assign n21833 = n20343 & n21832 ;
  assign n21834 = n21833 ^ n2053 ^ n603 ;
  assign n21831 = n16314 ^ n16011 ^ 1'b0 ;
  assign n21835 = n21834 ^ n21831 ^ 1'b0 ;
  assign n21836 = n21835 ^ n15501 ^ 1'b0 ;
  assign n21837 = n9575 ^ n2953 ^ n802 ;
  assign n21838 = n2979 & n21837 ;
  assign n21841 = n6887 ^ n1401 ^ 1'b0 ;
  assign n21842 = n2126 & n21841 ;
  assign n21840 = n19776 ^ n17940 ^ 1'b0 ;
  assign n21843 = n21842 ^ n21840 ^ n2673 ;
  assign n21839 = n10829 ^ n6731 ^ 1'b0 ;
  assign n21844 = n21843 ^ n21839 ^ n16610 ;
  assign n21850 = ( x41 & n4277 ) | ( x41 & n5737 ) | ( n4277 & n5737 ) ;
  assign n21851 = n21850 ^ n2316 ^ 1'b0 ;
  assign n21852 = ~n11426 & n21851 ;
  assign n21853 = n21852 ^ n13399 ^ 1'b0 ;
  assign n21845 = n17154 ^ n2353 ^ 1'b0 ;
  assign n21846 = n7042 & n21845 ;
  assign n21847 = n21846 ^ n11758 ^ n9670 ;
  assign n21848 = n21847 ^ n14501 ^ n6201 ;
  assign n21849 = ~n3877 & n21848 ;
  assign n21854 = n21853 ^ n21849 ^ 1'b0 ;
  assign n21855 = ( ~n2022 & n8986 ) | ( ~n2022 & n15026 ) | ( n8986 & n15026 ) ;
  assign n21856 = ( ~n9042 & n13647 ) | ( ~n9042 & n21855 ) | ( n13647 & n21855 ) ;
  assign n21857 = ~n10695 & n14352 ;
  assign n21858 = n21857 ^ n19966 ^ 1'b0 ;
  assign n21859 = ~n2121 & n6274 ;
  assign n21860 = ~n15064 & n21859 ;
  assign n21861 = n21860 ^ n5714 ^ n2651 ;
  assign n21862 = ( n10071 & ~n20730 ) | ( n10071 & n21861 ) | ( ~n20730 & n21861 ) ;
  assign n21863 = n21858 & n21862 ;
  assign n21864 = n11161 ^ n3712 ^ n1495 ;
  assign n21865 = n17866 & n21864 ;
  assign n21866 = n21865 ^ n12708 ^ 1'b0 ;
  assign n21867 = ~n7080 & n21866 ;
  assign n21868 = n11243 & n21867 ;
  assign n21870 = ~n3195 & n18253 ;
  assign n21871 = n4735 | n21870 ;
  assign n21872 = n2657 & ~n21871 ;
  assign n21869 = n14854 ^ n6526 ^ n6302 ;
  assign n21873 = n21872 ^ n21869 ^ 1'b0 ;
  assign n21874 = ( n5670 & n10814 ) | ( n5670 & ~n21873 ) | ( n10814 & ~n21873 ) ;
  assign n21875 = ~n12005 & n17637 ;
  assign n21876 = ~n9185 & n12476 ;
  assign n21877 = ( n3529 & n8637 ) | ( n3529 & n21876 ) | ( n8637 & n21876 ) ;
  assign n21878 = ( ~n10508 & n15104 ) | ( ~n10508 & n15703 ) | ( n15104 & n15703 ) ;
  assign n21879 = n9374 ^ n4463 ^ 1'b0 ;
  assign n21880 = n7417 & ~n21879 ;
  assign n21881 = n16518 ^ n1826 ^ 1'b0 ;
  assign n21882 = n2740 ^ n317 ^ 1'b0 ;
  assign n21883 = n21881 | n21882 ;
  assign n21884 = n11629 | n16632 ;
  assign n21885 = n21884 ^ n13663 ^ 1'b0 ;
  assign n21886 = n21885 ^ n7704 ^ 1'b0 ;
  assign n21887 = n5810 ^ n2451 ^ 1'b0 ;
  assign n21888 = n21887 ^ n8380 ^ n6758 ;
  assign n21889 = n20611 & n21661 ;
  assign n21890 = n21888 & n21889 ;
  assign n21891 = n21890 ^ n10831 ^ n4283 ;
  assign n21892 = n21891 ^ n20918 ^ 1'b0 ;
  assign n21893 = n896 & n13097 ;
  assign n21894 = n4654 & ~n21893 ;
  assign n21895 = n17300 & n21894 ;
  assign n21896 = n1941 | n10651 ;
  assign n21897 = n17183 ^ n9231 ^ 1'b0 ;
  assign n21898 = n21896 & ~n21897 ;
  assign n21899 = ~n1076 & n2100 ;
  assign n21900 = n21899 ^ n13830 ^ 1'b0 ;
  assign n21901 = ~n4934 & n21900 ;
  assign n21902 = n21901 ^ n14913 ^ 1'b0 ;
  assign n21903 = n16046 ^ n6003 ^ 1'b0 ;
  assign n21904 = n15802 & ~n21903 ;
  assign n21905 = ( n3709 & n5244 ) | ( n3709 & ~n14069 ) | ( n5244 & ~n14069 ) ;
  assign n21906 = n7851 & n21905 ;
  assign n21907 = n21906 ^ n11201 ^ 1'b0 ;
  assign n21908 = ( ~n20389 & n21904 ) | ( ~n20389 & n21907 ) | ( n21904 & n21907 ) ;
  assign n21909 = ( n16544 & ~n21623 ) | ( n16544 & n21908 ) | ( ~n21623 & n21908 ) ;
  assign n21910 = n15040 ^ n11900 ^ n2791 ;
  assign n21911 = n21292 & n21910 ;
  assign n21912 = n21911 ^ n2799 ^ 1'b0 ;
  assign n21913 = n14980 ^ n8857 ^ 1'b0 ;
  assign n21914 = ( n2796 & n3485 ) | ( n2796 & ~n4047 ) | ( n3485 & ~n4047 ) ;
  assign n21915 = ( ~n12252 & n13729 ) | ( ~n12252 & n21914 ) | ( n13729 & n21914 ) ;
  assign n21916 = n15584 ^ n3116 ^ 1'b0 ;
  assign n21917 = ~n2807 & n21916 ;
  assign n21918 = n17740 & n21917 ;
  assign n21919 = n4584 & n21918 ;
  assign n21920 = ( ~n21913 & n21915 ) | ( ~n21913 & n21919 ) | ( n21915 & n21919 ) ;
  assign n21921 = n5065 & ~n10438 ;
  assign n21922 = ~x249 & n21921 ;
  assign n21923 = n21922 ^ n6036 ^ 1'b0 ;
  assign n21924 = n6709 | n21923 ;
  assign n21925 = n15056 | n21924 ;
  assign n21926 = n21925 ^ n3203 ^ 1'b0 ;
  assign n21927 = n2018 | n21926 ;
  assign n21928 = n21927 ^ n17713 ^ 1'b0 ;
  assign n21931 = n4774 ^ n798 ^ 1'b0 ;
  assign n21929 = n9418 | n21143 ;
  assign n21930 = n21929 ^ n3230 ^ 1'b0 ;
  assign n21932 = n21931 ^ n21930 ^ 1'b0 ;
  assign n21933 = n10052 & n21932 ;
  assign n21934 = n8126 & n19258 ;
  assign n21935 = n8819 & n21934 ;
  assign n21936 = ( n11137 & n12511 ) | ( n11137 & n21935 ) | ( n12511 & n21935 ) ;
  assign n21937 = n21936 ^ n2184 ^ x252 ;
  assign n21941 = n7262 & ~n15029 ;
  assign n21942 = ~n16464 & n21941 ;
  assign n21938 = n1394 & n17357 ;
  assign n21939 = n3601 & n21938 ;
  assign n21940 = n15687 & ~n21939 ;
  assign n21943 = n21942 ^ n21940 ^ 1'b0 ;
  assign n21944 = n20797 ^ n4612 ^ 1'b0 ;
  assign n21945 = ( n10244 & ~n17189 ) | ( n10244 & n17748 ) | ( ~n17189 & n17748 ) ;
  assign n21946 = n21945 ^ n4185 ^ 1'b0 ;
  assign n21947 = x214 | n13232 ;
  assign n21948 = ( ~n9350 & n9887 ) | ( ~n9350 & n20369 ) | ( n9887 & n20369 ) ;
  assign n21949 = ~n1289 & n7370 ;
  assign n21950 = n21949 ^ n4626 ^ n1923 ;
  assign n21951 = ~n21948 & n21950 ;
  assign n21952 = ~n1977 & n4686 ;
  assign n21953 = n4525 | n5567 ;
  assign n21954 = n5087 | n21953 ;
  assign n21955 = n8723 & n18125 ;
  assign n21956 = ~n21954 & n21955 ;
  assign n21957 = n21952 & ~n21956 ;
  assign n21958 = n17421 & ~n17769 ;
  assign n21959 = n2422 ^ n1018 ^ 1'b0 ;
  assign n21960 = n21959 ^ n3274 ^ 1'b0 ;
  assign n21961 = n7085 & ~n21960 ;
  assign n21962 = ( n1527 & ~n20504 ) | ( n1527 & n21961 ) | ( ~n20504 & n21961 ) ;
  assign n21963 = n21590 | n21668 ;
  assign n21964 = n10222 ^ n8969 ^ 1'b0 ;
  assign n21965 = n18259 | n21964 ;
  assign n21966 = n1329 | n21965 ;
  assign n21967 = n21966 ^ n17532 ^ 1'b0 ;
  assign n21968 = n12700 ^ n11991 ^ n1291 ;
  assign n21969 = n21001 ^ n7968 ^ n6877 ;
  assign n21970 = n14820 ^ n5686 ^ n4804 ;
  assign n21971 = n20202 & n21970 ;
  assign n21972 = n11319 ^ n2246 ^ 1'b0 ;
  assign n21973 = n18318 ^ n15825 ^ n12730 ;
  assign n21974 = n16348 & ~n21973 ;
  assign n21975 = n21974 ^ n10788 ^ 1'b0 ;
  assign n21976 = n19639 | n21975 ;
  assign n21977 = n21976 ^ n4914 ^ 1'b0 ;
  assign n21978 = n16247 ^ n12585 ^ n6242 ;
  assign n21979 = n4286 & n5524 ;
  assign n21980 = n7999 & n21979 ;
  assign n21981 = ( n3875 & ~n4536 ) | ( n3875 & n10138 ) | ( ~n4536 & n10138 ) ;
  assign n21982 = n21981 ^ n18033 ^ n12936 ;
  assign n21983 = n21980 | n21982 ;
  assign n21984 = n12993 | n21983 ;
  assign n21985 = n6406 | n20625 ;
  assign n21986 = n21985 ^ n12990 ^ n6393 ;
  assign n21987 = ~n1374 & n4282 ;
  assign n21988 = n8579 ^ n7013 ^ n6749 ;
  assign n21989 = n21988 ^ n7128 ^ 1'b0 ;
  assign n21990 = n4203 | n21989 ;
  assign n21991 = n10476 & n21990 ;
  assign n21992 = ~n17567 & n21991 ;
  assign n21993 = n21987 & n21992 ;
  assign n21994 = n21993 ^ n16862 ^ n10984 ;
  assign n21995 = n15710 & ~n21994 ;
  assign n21996 = n3247 & n21995 ;
  assign n21997 = ( n4828 & n6045 ) | ( n4828 & n7572 ) | ( n6045 & n7572 ) ;
  assign n21998 = n21997 ^ n2638 ^ 1'b0 ;
  assign n21999 = n4617 & n21998 ;
  assign n22000 = n17406 & n21999 ;
  assign n22001 = n2463 | n12162 ;
  assign n22002 = n7663 & ~n12337 ;
  assign n22003 = n22002 ^ n4021 ^ 1'b0 ;
  assign n22004 = ( n1717 & ~n4498 ) | ( n1717 & n22003 ) | ( ~n4498 & n22003 ) ;
  assign n22005 = ~n1294 & n22004 ;
  assign n22006 = ~n13615 & n22005 ;
  assign n22007 = n4040 | n9661 ;
  assign n22008 = n22007 ^ n7521 ^ 1'b0 ;
  assign n22009 = n22008 ^ n7725 ^ 1'b0 ;
  assign n22010 = n11655 ^ n1205 ^ x113 ;
  assign n22011 = n18243 | n22010 ;
  assign n22012 = n22011 ^ n16041 ^ n2207 ;
  assign n22013 = n22012 ^ n16280 ^ n10070 ;
  assign n22014 = n6031 & ~n18111 ;
  assign n22015 = n22014 ^ n6550 ^ 1'b0 ;
  assign n22016 = ( n2997 & n4771 ) | ( n2997 & n22015 ) | ( n4771 & n22015 ) ;
  assign n22017 = n15595 ^ n15298 ^ 1'b0 ;
  assign n22018 = n2173 & ~n22017 ;
  assign n22019 = n14380 ^ n9329 ^ n1411 ;
  assign n22020 = n22019 ^ n21088 ^ n5855 ;
  assign n22021 = n22020 ^ n14758 ^ 1'b0 ;
  assign n22022 = n5114 ^ n4426 ^ 1'b0 ;
  assign n22023 = n22022 ^ n13717 ^ n1722 ;
  assign n22024 = n2296 & n3880 ;
  assign n22025 = n22024 ^ n18527 ^ n15214 ;
  assign n22026 = n7622 & ~n9763 ;
  assign n22027 = n6752 & n22026 ;
  assign n22028 = n9601 ^ n3673 ^ 1'b0 ;
  assign n22029 = ( n8604 & n15495 ) | ( n8604 & n22028 ) | ( n15495 & n22028 ) ;
  assign n22030 = n22029 ^ n11789 ^ n3501 ;
  assign n22032 = n12214 ^ n10255 ^ n8824 ;
  assign n22031 = n20811 ^ n3408 ^ 1'b0 ;
  assign n22033 = n22032 ^ n22031 ^ n13599 ;
  assign n22034 = n12211 ^ n4811 ^ 1'b0 ;
  assign n22035 = n22034 ^ n14671 ^ 1'b0 ;
  assign n22036 = ~n10704 & n12370 ;
  assign n22037 = n22036 ^ n5963 ^ 1'b0 ;
  assign n22038 = n22037 ^ n12872 ^ 1'b0 ;
  assign n22039 = ( n2829 & ~n17372 ) | ( n2829 & n22038 ) | ( ~n17372 & n22038 ) ;
  assign n22044 = ~n12873 & n21988 ;
  assign n22043 = ~n2367 & n13263 ;
  assign n22045 = n22044 ^ n22043 ^ 1'b0 ;
  assign n22041 = n9711 ^ n4613 ^ 1'b0 ;
  assign n22042 = ( n9758 & n15159 ) | ( n9758 & ~n22041 ) | ( n15159 & ~n22041 ) ;
  assign n22046 = n22045 ^ n22042 ^ n9263 ;
  assign n22047 = n22046 ^ n8755 ^ 1'b0 ;
  assign n22040 = n11192 & n15516 ;
  assign n22048 = n22047 ^ n22040 ^ 1'b0 ;
  assign n22049 = n9341 & n12820 ;
  assign n22050 = ( n2018 & n22048 ) | ( n2018 & n22049 ) | ( n22048 & n22049 ) ;
  assign n22051 = ~n22039 & n22050 ;
  assign n22052 = ~n22035 & n22051 ;
  assign n22055 = ~n6705 & n12931 ;
  assign n22053 = n21733 ^ n20841 ^ n20126 ;
  assign n22054 = n22053 ^ n7278 ^ 1'b0 ;
  assign n22056 = n22055 ^ n22054 ^ 1'b0 ;
  assign n22057 = n6180 ^ n2178 ^ n1044 ;
  assign n22058 = n22057 ^ n3242 ^ n549 ;
  assign n22059 = ~n9429 & n22058 ;
  assign n22060 = n13368 ^ n7798 ^ 1'b0 ;
  assign n22061 = n7811 & n22060 ;
  assign n22062 = n22061 ^ n8414 ^ n5759 ;
  assign n22063 = ~n22059 & n22062 ;
  assign n22064 = n12564 ^ n6864 ^ 1'b0 ;
  assign n22065 = n2320 & ~n22064 ;
  assign n22067 = n5236 ^ n3767 ^ 1'b0 ;
  assign n22066 = n11170 ^ n7757 ^ n2145 ;
  assign n22068 = n22067 ^ n22066 ^ n1450 ;
  assign n22069 = n22068 ^ n2545 ^ 1'b0 ;
  assign n22070 = n6562 | n22069 ;
  assign n22071 = ( n13358 & n21905 ) | ( n13358 & n22070 ) | ( n21905 & n22070 ) ;
  assign n22072 = n18858 ^ n7726 ^ n868 ;
  assign n22073 = n22072 ^ n15378 ^ 1'b0 ;
  assign n22074 = n22073 ^ n15736 ^ n4662 ;
  assign n22076 = ~n5718 & n6594 ;
  assign n22077 = n5244 & n22076 ;
  assign n22075 = ( n3489 & ~n5175 ) | ( n3489 & n7402 ) | ( ~n5175 & n7402 ) ;
  assign n22078 = n22077 ^ n22075 ^ n3456 ;
  assign n22079 = n22078 ^ n2571 ^ n488 ;
  assign n22080 = n12518 | n22079 ;
  assign n22081 = n14994 | n22080 ;
  assign n22082 = ( n1368 & ~n7621 ) | ( n1368 & n22081 ) | ( ~n7621 & n22081 ) ;
  assign n22083 = n20579 ^ n13149 ^ n1895 ;
  assign n22084 = ~n758 & n18950 ;
  assign n22085 = ~n10766 & n22084 ;
  assign n22086 = ( ~n3626 & n5252 ) | ( ~n3626 & n11431 ) | ( n5252 & n11431 ) ;
  assign n22087 = ~n18564 & n22086 ;
  assign n22088 = n22087 ^ n8548 ^ 1'b0 ;
  assign n22089 = n8927 & ~n9266 ;
  assign n22090 = n22089 ^ n11039 ^ 1'b0 ;
  assign n22091 = n3215 | n22090 ;
  assign n22092 = n22091 ^ n7979 ^ n4239 ;
  assign n22093 = n16176 ^ n5387 ^ n4211 ;
  assign n22094 = n22093 ^ n21722 ^ n10585 ;
  assign n22095 = n17221 & n22094 ;
  assign n22096 = ( n9310 & n16367 ) | ( n9310 & n21870 ) | ( n16367 & n21870 ) ;
  assign n22097 = n22096 ^ n7258 ^ n1454 ;
  assign n22098 = ( ~n4523 & n10314 ) | ( ~n4523 & n16457 ) | ( n10314 & n16457 ) ;
  assign n22099 = n22098 ^ n14770 ^ n778 ;
  assign n22105 = n5962 | n10850 ;
  assign n22106 = n22105 ^ n2417 ^ 1'b0 ;
  assign n22100 = n12701 ^ n7842 ^ n4067 ;
  assign n22101 = ( x180 & ~n9516 ) | ( x180 & n22100 ) | ( ~n9516 & n22100 ) ;
  assign n22102 = ( n9485 & n18752 ) | ( n9485 & ~n22101 ) | ( n18752 & ~n22101 ) ;
  assign n22103 = n22102 ^ n16599 ^ n4138 ;
  assign n22104 = n1648 | n22103 ;
  assign n22107 = n22106 ^ n22104 ^ 1'b0 ;
  assign n22108 = ( ~n817 & n4802 ) | ( ~n817 & n11653 ) | ( n4802 & n11653 ) ;
  assign n22109 = n22108 ^ n9360 ^ 1'b0 ;
  assign n22112 = ~n8438 & n11099 ;
  assign n22113 = ~n6042 & n22112 ;
  assign n22110 = n7384 ^ n3741 ^ 1'b0 ;
  assign n22111 = n22110 ^ n6677 ^ n3071 ;
  assign n22114 = n22113 ^ n22111 ^ 1'b0 ;
  assign n22115 = n22109 & n22114 ;
  assign n22116 = n7880 & ~n8515 ;
  assign n22117 = n18411 ^ n6589 ^ n5854 ;
  assign n22118 = n8695 ^ n1243 ^ 1'b0 ;
  assign n22119 = ~n17203 & n22118 ;
  assign n22120 = n13751 & n22119 ;
  assign n22122 = n6039 & n11053 ;
  assign n22123 = ~n7494 & n22122 ;
  assign n22121 = n8306 & n8484 ;
  assign n22124 = n22123 ^ n22121 ^ n4782 ;
  assign n22125 = n14165 | n14972 ;
  assign n22126 = n13786 & ~n22125 ;
  assign n22127 = n22126 ^ n7723 ^ 1'b0 ;
  assign n22128 = x51 | n4374 ;
  assign n22130 = n5115 ^ n4510 ^ 1'b0 ;
  assign n22129 = n3803 | n11677 ;
  assign n22131 = n22130 ^ n22129 ^ 1'b0 ;
  assign n22132 = n16080 | n22131 ;
  assign n22140 = n12595 & n20295 ;
  assign n22133 = ( ~n1997 & n2261 ) | ( ~n1997 & n10530 ) | ( n2261 & n10530 ) ;
  assign n22134 = ~n2118 & n8957 ;
  assign n22135 = ( n5498 & n22133 ) | ( n5498 & ~n22134 ) | ( n22133 & ~n22134 ) ;
  assign n22136 = n22135 ^ n10010 ^ n4227 ;
  assign n22137 = ~n7395 & n9128 ;
  assign n22138 = n22137 ^ n20694 ^ 1'b0 ;
  assign n22139 = n22136 & n22138 ;
  assign n22141 = n22140 ^ n22139 ^ 1'b0 ;
  assign n22149 = n6274 ^ n4789 ^ 1'b0 ;
  assign n22150 = n2615 & ~n22149 ;
  assign n22151 = n8157 ^ n7317 ^ 1'b0 ;
  assign n22152 = n3305 | n22151 ;
  assign n22153 = n22150 & n22152 ;
  assign n22142 = n17607 ^ n13581 ^ 1'b0 ;
  assign n22143 = ~n13429 & n22142 ;
  assign n22144 = ~n1866 & n22143 ;
  assign n22145 = ~x192 & n22144 ;
  assign n22146 = n22145 ^ n22042 ^ n15622 ;
  assign n22147 = ( ~n1439 & n16272 ) | ( ~n1439 & n22146 ) | ( n16272 & n22146 ) ;
  assign n22148 = ( n2993 & n17978 ) | ( n2993 & n22147 ) | ( n17978 & n22147 ) ;
  assign n22154 = n22153 ^ n22148 ^ n20332 ;
  assign n22155 = x34 & n13918 ;
  assign n22156 = n22155 ^ n5270 ^ 1'b0 ;
  assign n22157 = n22156 ^ n20747 ^ n5451 ;
  assign n22159 = n20031 ^ n7824 ^ n1481 ;
  assign n22158 = n4846 | n9675 ;
  assign n22160 = n22159 ^ n22158 ^ 1'b0 ;
  assign n22161 = n17576 ^ n11443 ^ n4051 ;
  assign n22165 = n4057 | n5287 ;
  assign n22164 = x148 & ~n2163 ;
  assign n22166 = n22165 ^ n22164 ^ n17971 ;
  assign n22162 = x204 ^ x64 ^ 1'b0 ;
  assign n22163 = ~n13983 & n22162 ;
  assign n22167 = n22166 ^ n22163 ^ 1'b0 ;
  assign n22168 = n12608 & n17264 ;
  assign n22169 = n5460 ^ n261 ^ 1'b0 ;
  assign n22170 = n13113 & n22169 ;
  assign n22171 = ( n2257 & ~n17188 ) | ( n2257 & n17513 ) | ( ~n17188 & n17513 ) ;
  assign n22172 = n20086 ^ n9998 ^ 1'b0 ;
  assign n22173 = n22171 & ~n22172 ;
  assign n22174 = ( n12916 & ~n22170 ) | ( n12916 & n22173 ) | ( ~n22170 & n22173 ) ;
  assign n22175 = ( n8118 & ~n14017 ) | ( n8118 & n22174 ) | ( ~n14017 & n22174 ) ;
  assign n22176 = n22175 ^ x120 ^ 1'b0 ;
  assign n22177 = ( x86 & n3166 ) | ( x86 & ~n8988 ) | ( n3166 & ~n8988 ) ;
  assign n22178 = ( n2424 & n3705 ) | ( n2424 & ~n13919 ) | ( n3705 & ~n13919 ) ;
  assign n22179 = n7044 & n8163 ;
  assign n22180 = n22179 ^ n5776 ^ 1'b0 ;
  assign n22181 = n17077 & ~n22180 ;
  assign n22182 = n5451 & ~n6762 ;
  assign n22183 = n22182 ^ n11519 ^ n6934 ;
  assign n22184 = n7989 & ~n22183 ;
  assign n22185 = n22184 ^ n10230 ^ n5428 ;
  assign n22186 = n14593 ^ n13442 ^ n3950 ;
  assign n22187 = n22186 ^ n18996 ^ n10270 ;
  assign n22188 = n10345 ^ n2333 ^ n1216 ;
  assign n22189 = n9120 ^ n6532 ^ 1'b0 ;
  assign n22190 = n22188 & ~n22189 ;
  assign n22191 = n10377 ^ n6110 ^ n5808 ;
  assign n22192 = n17600 ^ n1545 ^ 1'b0 ;
  assign n22193 = n12177 & ~n22192 ;
  assign n22194 = n22191 & n22193 ;
  assign n22195 = n22194 ^ n17136 ^ n15842 ;
  assign n22196 = n16618 ^ n6359 ^ n5093 ;
  assign n22197 = n7855 & ~n11964 ;
  assign n22198 = n1489 & n22197 ;
  assign n22199 = ( n8019 & n8509 ) | ( n8019 & n22198 ) | ( n8509 & n22198 ) ;
  assign n22200 = ( n844 & n4268 ) | ( n844 & n11096 ) | ( n4268 & n11096 ) ;
  assign n22201 = n22200 ^ n8462 ^ 1'b0 ;
  assign n22202 = n10913 ^ n6302 ^ n2324 ;
  assign n22203 = n9627 ^ n4243 ^ 1'b0 ;
  assign n22204 = ( ~n21987 & n22202 ) | ( ~n21987 & n22203 ) | ( n22202 & n22203 ) ;
  assign n22205 = ( n5718 & ~n22201 ) | ( n5718 & n22204 ) | ( ~n22201 & n22204 ) ;
  assign n22206 = ~n3625 & n17791 ;
  assign n22207 = n8604 ^ n3157 ^ 1'b0 ;
  assign n22208 = ~n3285 & n22207 ;
  assign n22209 = n4779 & ~n5958 ;
  assign n22210 = ( ~n21000 & n22208 ) | ( ~n21000 & n22209 ) | ( n22208 & n22209 ) ;
  assign n22211 = n22210 ^ n6139 ^ n3092 ;
  assign n22212 = ~n1193 & n2502 ;
  assign n22213 = n8667 & n22212 ;
  assign n22214 = ~n4192 & n6030 ;
  assign n22215 = n22213 & n22214 ;
  assign n22216 = n12552 ^ n7475 ^ n2402 ;
  assign n22221 = ( n358 & n4595 ) | ( n358 & n10838 ) | ( n4595 & n10838 ) ;
  assign n22222 = ( n3344 & ~n16244 ) | ( n3344 & n22221 ) | ( ~n16244 & n22221 ) ;
  assign n22217 = n9016 | n10384 ;
  assign n22218 = n22217 ^ n9560 ^ 1'b0 ;
  assign n22219 = n15587 | n22218 ;
  assign n22220 = n273 & ~n22219 ;
  assign n22223 = n22222 ^ n22220 ^ 1'b0 ;
  assign n22224 = n12035 & n22223 ;
  assign n22225 = n7588 ^ n6497 ^ n4621 ;
  assign n22226 = n22225 ^ n4502 ^ 1'b0 ;
  assign n22227 = n5322 ^ n1317 ^ n465 ;
  assign n22228 = ~n12509 & n22227 ;
  assign n22229 = ( ~n6649 & n7398 ) | ( ~n6649 & n16604 ) | ( n7398 & n16604 ) ;
  assign n22230 = ~n22228 & n22229 ;
  assign n22231 = n22230 ^ n21858 ^ 1'b0 ;
  assign n22232 = n22231 ^ n21384 ^ 1'b0 ;
  assign n22233 = ~n16249 & n22232 ;
  assign n22234 = n14195 ^ n5378 ^ 1'b0 ;
  assign n22235 = x167 & ~n22234 ;
  assign n22236 = ~n9479 & n22235 ;
  assign n22237 = n3350 & n4584 ;
  assign n22238 = n10969 ^ n6990 ^ n1224 ;
  assign n22239 = ~n22237 & n22238 ;
  assign n22240 = n22236 & n22239 ;
  assign n22241 = n10825 ^ n10261 ^ n2360 ;
  assign n22242 = n22241 ^ n4303 ^ 1'b0 ;
  assign n22243 = n22242 ^ n17966 ^ n7220 ;
  assign n22244 = ( x84 & ~n363 ) | ( x84 & n2154 ) | ( ~n363 & n2154 ) ;
  assign n22245 = n22244 ^ n7808 ^ n2574 ;
  assign n22246 = n22015 & n22245 ;
  assign n22247 = n22246 ^ n5394 ^ 1'b0 ;
  assign n22248 = ( n16032 & ~n22243 ) | ( n16032 & n22247 ) | ( ~n22243 & n22247 ) ;
  assign n22249 = x239 & n7215 ;
  assign n22250 = n1124 & n22249 ;
  assign n22251 = n16821 & n22250 ;
  assign n22252 = n10980 ^ n6807 ^ 1'b0 ;
  assign n22253 = n8804 & n22252 ;
  assign n22254 = ( n1749 & ~n9340 ) | ( n1749 & n22253 ) | ( ~n9340 & n22253 ) ;
  assign n22255 = n22254 ^ n16766 ^ 1'b0 ;
  assign n22256 = n8917 & ~n22255 ;
  assign n22257 = n22256 ^ n18162 ^ 1'b0 ;
  assign n22258 = ~n22034 & n22257 ;
  assign n22259 = n4568 & n22258 ;
  assign n22260 = ( n1738 & n2074 ) | ( n1738 & n3556 ) | ( n2074 & n3556 ) ;
  assign n22261 = n22260 ^ n19252 ^ 1'b0 ;
  assign n22262 = ~n4942 & n22261 ;
  assign n22263 = n22262 ^ n5173 ^ 1'b0 ;
  assign n22264 = n19454 ^ n4967 ^ 1'b0 ;
  assign n22268 = n6483 & ~n10777 ;
  assign n22265 = n14188 ^ n723 ^ 1'b0 ;
  assign n22266 = n12467 & ~n22265 ;
  assign n22267 = ( n9084 & ~n16287 ) | ( n9084 & n22266 ) | ( ~n16287 & n22266 ) ;
  assign n22269 = n22268 ^ n22267 ^ n3740 ;
  assign n22270 = n22269 ^ n6423 ^ 1'b0 ;
  assign n22271 = n7352 | n22270 ;
  assign n22272 = n4611 ^ n2034 ^ 1'b0 ;
  assign n22273 = ~n18804 & n22272 ;
  assign n22276 = ( ~n12814 & n21046 ) | ( ~n12814 & n21139 ) | ( n21046 & n21139 ) ;
  assign n22274 = ~n4196 & n11578 ;
  assign n22275 = n21644 | n22274 ;
  assign n22277 = n22276 ^ n22275 ^ n16585 ;
  assign n22278 = ( n2441 & ~n2723 ) | ( n2441 & n4756 ) | ( ~n2723 & n4756 ) ;
  assign n22279 = ( n1235 & ~n12005 ) | ( n1235 & n22278 ) | ( ~n12005 & n22278 ) ;
  assign n22280 = ( ~n387 & n6226 ) | ( ~n387 & n15302 ) | ( n6226 & n15302 ) ;
  assign n22281 = n22280 ^ n4281 ^ 1'b0 ;
  assign n22282 = n2120 | n9755 ;
  assign n22283 = n22282 ^ n9331 ^ 1'b0 ;
  assign n22284 = n22283 ^ n6223 ^ 1'b0 ;
  assign n22285 = n10005 ^ n5373 ^ 1'b0 ;
  assign n22286 = n8157 & ~n22285 ;
  assign n22287 = n22286 ^ n20865 ^ n14649 ;
  assign n22288 = n22287 ^ n12035 ^ 1'b0 ;
  assign n22289 = n11945 & ~n22288 ;
  assign n22290 = n20987 ^ n10317 ^ n7097 ;
  assign n22291 = n4914 | n12641 ;
  assign n22292 = ~n1515 & n14809 ;
  assign n22295 = n1334 & ~n7263 ;
  assign n22296 = n13120 & n22295 ;
  assign n22293 = n8663 ^ n6046 ^ n2416 ;
  assign n22294 = ( n3844 & n5681 ) | ( n3844 & ~n22293 ) | ( n5681 & ~n22293 ) ;
  assign n22297 = n22296 ^ n22294 ^ n16079 ;
  assign n22298 = x82 & ~n17944 ;
  assign n22299 = n22297 & n22298 ;
  assign n22300 = ( n2271 & n3055 ) | ( n2271 & ~n22299 ) | ( n3055 & ~n22299 ) ;
  assign n22301 = n10106 & ~n15847 ;
  assign n22302 = n22301 ^ n12833 ^ 1'b0 ;
  assign n22303 = ~n6503 & n7766 ;
  assign n22304 = n10463 ^ n7061 ^ n6425 ;
  assign n22305 = n6458 & n10078 ;
  assign n22306 = n22305 ^ n13873 ^ 1'b0 ;
  assign n22307 = n22306 ^ n13499 ^ n11962 ;
  assign n22308 = n2547 & ~n5570 ;
  assign n22309 = n7726 & n22308 ;
  assign n22310 = ( n14101 & n22307 ) | ( n14101 & n22309 ) | ( n22307 & n22309 ) ;
  assign n22311 = ~n22304 & n22310 ;
  assign n22312 = n7272 ^ n6388 ^ n5279 ;
  assign n22313 = ( n2667 & n9270 ) | ( n2667 & ~n22312 ) | ( n9270 & ~n22312 ) ;
  assign n22314 = ~n609 & n22313 ;
  assign n22315 = ( ~n826 & n14757 ) | ( ~n826 & n15332 ) | ( n14757 & n15332 ) ;
  assign n22316 = n10373 | n21993 ;
  assign n22317 = n16841 & ~n22316 ;
  assign n22318 = n13713 ^ n7013 ^ 1'b0 ;
  assign n22319 = ( n5029 & n13022 ) | ( n5029 & n22318 ) | ( n13022 & n22318 ) ;
  assign n22320 = ( x23 & n12944 ) | ( x23 & n14847 ) | ( n12944 & n14847 ) ;
  assign n22321 = n615 & ~n14103 ;
  assign n22322 = n1422 & ~n3472 ;
  assign n22323 = ( n1209 & n18087 ) | ( n1209 & n22322 ) | ( n18087 & n22322 ) ;
  assign n22324 = n22321 | n22323 ;
  assign n22325 = ( n1355 & n5092 ) | ( n1355 & n7822 ) | ( n5092 & n7822 ) ;
  assign n22326 = n11705 & ~n22325 ;
  assign n22327 = n22326 ^ n8372 ^ 1'b0 ;
  assign n22328 = n22324 & ~n22327 ;
  assign n22333 = n5782 | n14303 ;
  assign n22329 = n5385 | n10025 ;
  assign n22330 = n2619 | n22329 ;
  assign n22331 = ( ~n4301 & n12266 ) | ( ~n4301 & n22330 ) | ( n12266 & n22330 ) ;
  assign n22332 = ( x143 & n13059 ) | ( x143 & ~n22331 ) | ( n13059 & ~n22331 ) ;
  assign n22334 = n22333 ^ n22332 ^ n5093 ;
  assign n22335 = ( ~n3804 & n12813 ) | ( ~n3804 & n13984 ) | ( n12813 & n13984 ) ;
  assign n22336 = n1570 ^ n1546 ^ 1'b0 ;
  assign n22337 = x34 & n22336 ;
  assign n22340 = n585 & ~n973 ;
  assign n22341 = n973 & n22340 ;
  assign n22342 = n19104 | n22341 ;
  assign n22338 = n10187 ^ n4325 ^ 1'b0 ;
  assign n22339 = n13067 | n22338 ;
  assign n22343 = n22342 ^ n22339 ^ 1'b0 ;
  assign n22344 = n22337 & n22343 ;
  assign n22345 = n13867 ^ n1427 ^ 1'b0 ;
  assign n22347 = n7171 ^ n5738 ^ 1'b0 ;
  assign n22346 = n4226 & ~n9919 ;
  assign n22348 = n22347 ^ n22346 ^ n6167 ;
  assign n22352 = ~n625 & n3883 ;
  assign n22353 = n15895 & n22352 ;
  assign n22354 = n22353 ^ n1250 ^ 1'b0 ;
  assign n22349 = n10396 ^ n3577 ^ 1'b0 ;
  assign n22350 = n4936 & ~n22349 ;
  assign n22351 = ~n4011 & n22350 ;
  assign n22355 = n22354 ^ n22351 ^ 1'b0 ;
  assign n22356 = n11381 | n22355 ;
  assign n22357 = n22356 ^ n20483 ^ 1'b0 ;
  assign n22360 = ( n1796 & n5231 ) | ( n1796 & n5418 ) | ( n5231 & n5418 ) ;
  assign n22359 = n11533 ^ n6628 ^ n6298 ;
  assign n22361 = n22360 ^ n22359 ^ n6443 ;
  assign n22362 = ( ~n1791 & n3449 ) | ( ~n1791 & n22361 ) | ( n3449 & n22361 ) ;
  assign n22363 = n13729 & ~n22362 ;
  assign n22358 = n4009 & n18539 ;
  assign n22364 = n22363 ^ n22358 ^ 1'b0 ;
  assign n22365 = n5546 ^ n5273 ^ 1'b0 ;
  assign n22366 = ~n2930 & n22365 ;
  assign n22367 = n22366 ^ n12479 ^ 1'b0 ;
  assign n22368 = ~n5734 & n19279 ;
  assign n22369 = n22368 ^ n3709 ^ 1'b0 ;
  assign n22370 = n11341 & ~n22369 ;
  assign n22371 = n22370 ^ n11564 ^ n4761 ;
  assign n22372 = n312 & n736 ;
  assign n22373 = n13318 & n22372 ;
  assign n22375 = ( n3319 & ~n18505 ) | ( n3319 & n19920 ) | ( ~n18505 & n19920 ) ;
  assign n22374 = ~n2503 & n9385 ;
  assign n22376 = n22375 ^ n22374 ^ 1'b0 ;
  assign n22377 = ( x95 & ~n936 ) | ( x95 & n6822 ) | ( ~n936 & n6822 ) ;
  assign n22378 = x222 & n3904 ;
  assign n22379 = n4536 & n22378 ;
  assign n22380 = n22377 | n22379 ;
  assign n22381 = n6068 ^ n1315 ^ x234 ;
  assign n22382 = ( n2388 & n11749 ) | ( n2388 & ~n22381 ) | ( n11749 & ~n22381 ) ;
  assign n22383 = n22382 ^ n21234 ^ n13816 ;
  assign n22384 = ( ~n8602 & n11570 ) | ( ~n8602 & n21576 ) | ( n11570 & n21576 ) ;
  assign n22385 = ( n2065 & n14931 ) | ( n2065 & n22384 ) | ( n14931 & n22384 ) ;
  assign n22386 = n5170 & ~n20130 ;
  assign n22387 = n9402 & n22386 ;
  assign n22388 = ( n1738 & ~n7794 ) | ( n1738 & n13346 ) | ( ~n7794 & n13346 ) ;
  assign n22391 = n2387 ^ n887 ^ 1'b0 ;
  assign n22392 = ~n9342 & n22391 ;
  assign n22393 = n22392 ^ n304 ^ 1'b0 ;
  assign n22389 = x22 & ~n20382 ;
  assign n22390 = n22389 ^ n10424 ^ 1'b0 ;
  assign n22394 = n22393 ^ n22390 ^ n7244 ;
  assign n22396 = n4897 ^ n4368 ^ n1511 ;
  assign n22395 = ~n1981 & n5604 ;
  assign n22397 = n22396 ^ n22395 ^ 1'b0 ;
  assign n22398 = n6666 | n22397 ;
  assign n22399 = n10743 ^ n6541 ^ n2717 ;
  assign n22400 = n4020 & n22399 ;
  assign n22401 = n22400 ^ n734 ^ 1'b0 ;
  assign n22402 = n3968 & ~n22401 ;
  assign n22403 = n22402 ^ n14074 ^ 1'b0 ;
  assign n22404 = n664 | n16737 ;
  assign n22405 = ~n9172 & n22404 ;
  assign n22406 = n8983 ^ n8546 ^ n5086 ;
  assign n22407 = n22405 | n22406 ;
  assign n22408 = ( n2002 & n3189 ) | ( n2002 & ~n5670 ) | ( n3189 & ~n5670 ) ;
  assign n22409 = ( n9320 & ~n9754 ) | ( n9320 & n9955 ) | ( ~n9754 & n9955 ) ;
  assign n22410 = ( n10740 & n22408 ) | ( n10740 & n22409 ) | ( n22408 & n22409 ) ;
  assign n22411 = ( ~n6762 & n16528 ) | ( ~n6762 & n22410 ) | ( n16528 & n22410 ) ;
  assign n22412 = n20942 ^ n7036 ^ 1'b0 ;
  assign n22418 = n3939 & ~n15250 ;
  assign n22417 = n9146 ^ n7971 ^ n1310 ;
  assign n22419 = n22418 ^ n22417 ^ n14116 ;
  assign n22414 = n15965 ^ n11446 ^ n9567 ;
  assign n22413 = ~n12707 & n21991 ;
  assign n22415 = n22414 ^ n22413 ^ 1'b0 ;
  assign n22416 = n10070 & n22415 ;
  assign n22420 = n22419 ^ n22416 ^ n2492 ;
  assign n22421 = n4635 ^ n3303 ^ n2909 ;
  assign n22422 = n22421 ^ n16311 ^ 1'b0 ;
  assign n22423 = n9503 & ~n22422 ;
  assign n22424 = n12919 ^ x193 ^ x104 ;
  assign n22425 = n9220 | n22424 ;
  assign n22426 = n22423 | n22425 ;
  assign n22427 = ( n849 & n7442 ) | ( n849 & ~n8822 ) | ( n7442 & ~n8822 ) ;
  assign n22428 = n22427 ^ n5146 ^ 1'b0 ;
  assign n22429 = n6197 ^ n2746 ^ 1'b0 ;
  assign n22430 = ( n15157 & ~n17391 ) | ( n15157 & n22429 ) | ( ~n17391 & n22429 ) ;
  assign n22433 = n1538 | n1563 ;
  assign n22434 = n926 & ~n22433 ;
  assign n22435 = n2185 | n12373 ;
  assign n22436 = n22434 & ~n22435 ;
  assign n22431 = n18620 ^ n3761 ^ 1'b0 ;
  assign n22432 = ~n1550 & n22431 ;
  assign n22437 = n22436 ^ n22432 ^ n15298 ;
  assign n22438 = ~n21280 & n22437 ;
  assign n22439 = ( n5198 & n6277 ) | ( n5198 & ~n11189 ) | ( n6277 & ~n11189 ) ;
  assign n22440 = ( n326 & ~n2619 ) | ( n326 & n22439 ) | ( ~n2619 & n22439 ) ;
  assign n22441 = ( n18487 & n21840 ) | ( n18487 & n22324 ) | ( n21840 & n22324 ) ;
  assign n22442 = n11438 ^ n6673 ^ n6485 ;
  assign n22443 = n1987 | n16773 ;
  assign n22444 = ( n18728 & n22442 ) | ( n18728 & ~n22443 ) | ( n22442 & ~n22443 ) ;
  assign n22445 = n10788 & n13296 ;
  assign n22446 = n22445 ^ n701 ^ 1'b0 ;
  assign n22449 = n1166 | n2959 ;
  assign n22447 = n12753 ^ n9451 ^ 1'b0 ;
  assign n22448 = n2415 & n22447 ;
  assign n22450 = n22449 ^ n22448 ^ 1'b0 ;
  assign n22451 = n15475 ^ n14175 ^ 1'b0 ;
  assign n22452 = n15072 & n22451 ;
  assign n22453 = ( n3409 & n13200 ) | ( n3409 & n20424 ) | ( n13200 & n20424 ) ;
  assign n22454 = n21606 ^ n12626 ^ n9467 ;
  assign n22455 = n22454 ^ n7758 ^ 1'b0 ;
  assign n22456 = ~n1862 & n9692 ;
  assign n22457 = n22455 & n22456 ;
  assign n22458 = ( n2708 & ~n3133 ) | ( n2708 & n6517 ) | ( ~n3133 & n6517 ) ;
  assign n22459 = ~n3203 & n22458 ;
  assign n22460 = ~n556 & n4519 ;
  assign n22461 = n22460 ^ n11829 ^ 1'b0 ;
  assign n22462 = n17570 ^ n17462 ^ n8224 ;
  assign n22463 = ( n8002 & ~n22461 ) | ( n8002 & n22462 ) | ( ~n22461 & n22462 ) ;
  assign n22464 = n2208 | n4958 ;
  assign n22465 = n4961 & ~n22464 ;
  assign n22466 = n17623 & ~n22465 ;
  assign n22467 = n22466 ^ n5697 ^ 1'b0 ;
  assign n22468 = ( n6857 & ~n10943 ) | ( n6857 & n16108 ) | ( ~n10943 & n16108 ) ;
  assign n22469 = n9583 ^ n4640 ^ 1'b0 ;
  assign n22470 = n7342 | n22469 ;
  assign n22471 = ( n4043 & n9511 ) | ( n4043 & n22470 ) | ( n9511 & n22470 ) ;
  assign n22474 = n3853 & ~n11292 ;
  assign n22475 = n3430 ^ n2720 ^ 1'b0 ;
  assign n22476 = n7642 | n22475 ;
  assign n22477 = ( n8454 & n19247 ) | ( n8454 & n22476 ) | ( n19247 & n22476 ) ;
  assign n22478 = n22474 & n22477 ;
  assign n22479 = n22478 ^ n19891 ^ n2386 ;
  assign n22472 = n5989 ^ n5245 ^ 1'b0 ;
  assign n22473 = ( n7129 & n15277 ) | ( n7129 & ~n22472 ) | ( n15277 & ~n22472 ) ;
  assign n22480 = n22479 ^ n22473 ^ 1'b0 ;
  assign n22481 = ( n21817 & ~n22471 ) | ( n21817 & n22480 ) | ( ~n22471 & n22480 ) ;
  assign n22482 = n4484 | n18513 ;
  assign n22483 = n22482 ^ n1188 ^ 1'b0 ;
  assign n22484 = n22483 ^ n12483 ^ 1'b0 ;
  assign n22485 = n5158 | n10256 ;
  assign n22486 = n293 & ~n15913 ;
  assign n22487 = n22486 ^ n11407 ^ 1'b0 ;
  assign n22488 = ~n22485 & n22487 ;
  assign n22489 = ( ~n2337 & n22484 ) | ( ~n2337 & n22488 ) | ( n22484 & n22488 ) ;
  assign n22491 = n1452 & n5455 ;
  assign n22490 = n1952 & ~n2009 ;
  assign n22492 = n22491 ^ n22490 ^ 1'b0 ;
  assign n22497 = x235 & n1881 ;
  assign n22498 = n12605 & n22497 ;
  assign n22499 = ( n6106 & n8895 ) | ( n6106 & n22498 ) | ( n8895 & n22498 ) ;
  assign n22493 = ~n8773 & n20056 ;
  assign n22494 = ~n17594 & n22493 ;
  assign n22495 = n22494 ^ n10153 ^ 1'b0 ;
  assign n22496 = n18512 & n22495 ;
  assign n22500 = n22499 ^ n22496 ^ 1'b0 ;
  assign n22501 = n5569 & n15634 ;
  assign n22502 = n22501 ^ n4760 ^ 1'b0 ;
  assign n22503 = n11084 & ~n22502 ;
  assign n22504 = n22503 ^ n19049 ^ 1'b0 ;
  assign n22505 = n2040 | n7089 ;
  assign n22506 = n22505 ^ n3527 ^ 1'b0 ;
  assign n22507 = n22506 ^ n1980 ^ 1'b0 ;
  assign n22508 = n1631 & ~n11819 ;
  assign n22509 = n10048 & n22508 ;
  assign n22510 = n22091 | n22509 ;
  assign n22511 = n22510 ^ n19393 ^ 1'b0 ;
  assign n22512 = n22511 ^ n13129 ^ 1'b0 ;
  assign n22513 = ( n10277 & n22322 ) | ( n10277 & ~n22512 ) | ( n22322 & ~n22512 ) ;
  assign n22514 = n22028 ^ n15023 ^ n8032 ;
  assign n22515 = ( n4930 & n12680 ) | ( n4930 & ~n22514 ) | ( n12680 & ~n22514 ) ;
  assign n22516 = n11329 ^ n1211 ^ 1'b0 ;
  assign n22517 = n8276 & ~n22516 ;
  assign n22518 = n22517 ^ n9308 ^ 1'b0 ;
  assign n22519 = n7924 & n21194 ;
  assign n22521 = n11725 & n18604 ;
  assign n22522 = ( n461 & n7347 ) | ( n461 & ~n22521 ) | ( n7347 & ~n22521 ) ;
  assign n22520 = n1235 & ~n3741 ;
  assign n22523 = n22522 ^ n22520 ^ n4263 ;
  assign n22524 = ~n4141 & n13396 ;
  assign n22525 = n22524 ^ n2445 ^ 1'b0 ;
  assign n22526 = ( n8397 & n14494 ) | ( n8397 & n18727 ) | ( n14494 & n18727 ) ;
  assign n22527 = n17151 ^ n6036 ^ 1'b0 ;
  assign n22528 = n5542 & ~n22527 ;
  assign n22529 = n14296 ^ n11677 ^ 1'b0 ;
  assign n22530 = n19002 ^ n7309 ^ 1'b0 ;
  assign n22531 = n5832 & ~n22530 ;
  assign n22532 = ( n16971 & n18004 ) | ( n16971 & n22323 ) | ( n18004 & n22323 ) ;
  assign n22533 = n22532 ^ n8189 ^ 1'b0 ;
  assign n22534 = ~n21241 & n22533 ;
  assign n22535 = n19229 ^ n6432 ^ n1519 ;
  assign n22536 = ( n6977 & n11108 ) | ( n6977 & ~n12064 ) | ( n11108 & ~n12064 ) ;
  assign n22537 = n16793 ^ n10196 ^ 1'b0 ;
  assign n22538 = ~n17213 & n22537 ;
  assign n22539 = n21917 & ~n22538 ;
  assign n22540 = ( n22535 & n22536 ) | ( n22535 & ~n22539 ) | ( n22536 & ~n22539 ) ;
  assign n22541 = n9996 ^ n2538 ^ 1'b0 ;
  assign n22542 = n16451 | n22541 ;
  assign n22543 = n21485 ^ n8166 ^ n5293 ;
  assign n22544 = n16570 | n22543 ;
  assign n22545 = n4058 ^ n723 ^ 1'b0 ;
  assign n22546 = ( n4151 & ~n11470 ) | ( n4151 & n22545 ) | ( ~n11470 & n22545 ) ;
  assign n22547 = n22546 ^ n5314 ^ n461 ;
  assign n22548 = n9686 | n22547 ;
  assign n22549 = n22548 ^ n8864 ^ 1'b0 ;
  assign n22550 = n13580 ^ n12574 ^ n5646 ;
  assign n22551 = n22550 ^ n14428 ^ n11616 ;
  assign n22552 = n22551 ^ n11497 ^ n9192 ;
  assign n22553 = n5524 ^ n554 ^ 1'b0 ;
  assign n22554 = n5619 ^ n3748 ^ n1518 ;
  assign n22555 = n22554 ^ n1294 ^ 1'b0 ;
  assign n22556 = n7349 & n22555 ;
  assign n22557 = ( n1440 & ~n2702 ) | ( n1440 & n2799 ) | ( ~n2702 & n2799 ) ;
  assign n22558 = n22557 ^ n19927 ^ 1'b0 ;
  assign n22559 = n8109 & n22558 ;
  assign n22561 = ( ~n9769 & n10030 ) | ( ~n9769 & n13622 ) | ( n10030 & n13622 ) ;
  assign n22560 = n350 & n7310 ;
  assign n22562 = n22561 ^ n22560 ^ 1'b0 ;
  assign n22563 = n16313 ^ n9027 ^ n8828 ;
  assign n22564 = ( n2194 & ~n4349 ) | ( n2194 & n11968 ) | ( ~n4349 & n11968 ) ;
  assign n22565 = n10284 ^ n4078 ^ 1'b0 ;
  assign n22566 = ~n9012 & n22565 ;
  assign n22567 = n17232 ^ n8772 ^ 1'b0 ;
  assign n22568 = n22566 & n22567 ;
  assign n22569 = n15825 ^ n11529 ^ n4962 ;
  assign n22571 = ( ~n818 & n2256 ) | ( ~n818 & n7761 ) | ( n2256 & n7761 ) ;
  assign n22570 = ( n3073 & n6227 ) | ( n3073 & ~n11147 ) | ( n6227 & ~n11147 ) ;
  assign n22572 = n22571 ^ n22570 ^ n7065 ;
  assign n22573 = n20450 ^ n17313 ^ 1'b0 ;
  assign n22574 = ~n22572 & n22573 ;
  assign n22575 = n22574 ^ n21521 ^ 1'b0 ;
  assign n22576 = n638 | n3885 ;
  assign n22577 = n22576 ^ n1796 ^ 1'b0 ;
  assign n22578 = n4130 & n20405 ;
  assign n22579 = ( ~n6261 & n22577 ) | ( ~n6261 & n22578 ) | ( n22577 & n22578 ) ;
  assign n22580 = n12753 ^ n6238 ^ n5221 ;
  assign n22583 = ( n1666 & n4161 ) | ( n1666 & ~n4629 ) | ( n4161 & ~n4629 ) ;
  assign n22584 = n22583 ^ n6532 ^ n1125 ;
  assign n22581 = ( n9655 & n10465 ) | ( n9655 & n21064 ) | ( n10465 & n21064 ) ;
  assign n22582 = n14807 | n22581 ;
  assign n22585 = n22584 ^ n22582 ^ 1'b0 ;
  assign n22587 = n2631 & n5192 ;
  assign n22588 = n5773 & n22587 ;
  assign n22586 = n622 & n1304 ;
  assign n22589 = n22588 ^ n22586 ^ 1'b0 ;
  assign n22590 = n11883 ^ n10139 ^ 1'b0 ;
  assign n22596 = ~n9654 & n19777 ;
  assign n22597 = ~n10460 & n22596 ;
  assign n22591 = ~n4139 & n4142 ;
  assign n22592 = n815 | n22591 ;
  assign n22593 = n22592 ^ n4152 ^ 1'b0 ;
  assign n22594 = n22593 ^ n6104 ^ 1'b0 ;
  assign n22595 = ~n11371 & n22594 ;
  assign n22598 = n22597 ^ n22595 ^ n21148 ;
  assign n22599 = n20040 ^ n18375 ^ 1'b0 ;
  assign n22600 = n8957 ^ n5394 ^ 1'b0 ;
  assign n22601 = n20999 | n22600 ;
  assign n22602 = n22601 ^ n7776 ^ n5749 ;
  assign n22603 = n11466 ^ n9744 ^ 1'b0 ;
  assign n22604 = n2676 ^ x136 ^ 1'b0 ;
  assign n22605 = ( n9178 & n9376 ) | ( n9178 & n22604 ) | ( n9376 & n22604 ) ;
  assign n22606 = n5417 | n10100 ;
  assign n22607 = ~n3050 & n4563 ;
  assign n22608 = ~n1315 & n22607 ;
  assign n22609 = ( n5664 & ~n7763 ) | ( n5664 & n17946 ) | ( ~n7763 & n17946 ) ;
  assign n22610 = n2087 | n2947 ;
  assign n22611 = n576 | n3762 ;
  assign n22612 = n3181 | n22611 ;
  assign n22613 = n22612 ^ n20225 ^ n14087 ;
  assign n22614 = ~n22610 & n22613 ;
  assign n22615 = n22609 & n22614 ;
  assign n22616 = ( n9189 & ~n22608 ) | ( n9189 & n22615 ) | ( ~n22608 & n22615 ) ;
  assign n22621 = ( x169 & n1241 ) | ( x169 & n3348 ) | ( n1241 & n3348 ) ;
  assign n22622 = n22621 ^ n6196 ^ n2475 ;
  assign n22617 = n2639 ^ n1165 ^ 1'b0 ;
  assign n22618 = n4864 | n22617 ;
  assign n22619 = n22618 ^ n15994 ^ n7464 ;
  assign n22620 = n22619 ^ n9118 ^ n3226 ;
  assign n22623 = n22622 ^ n22620 ^ 1'b0 ;
  assign n22624 = ~n22616 & n22623 ;
  assign n22625 = n4782 & n10223 ;
  assign n22626 = n19105 ^ n4936 ^ 1'b0 ;
  assign n22627 = n2178 & ~n6421 ;
  assign n22628 = n22627 ^ n22032 ^ n7798 ;
  assign n22629 = ( x39 & n8460 ) | ( x39 & n15078 ) | ( n8460 & n15078 ) ;
  assign n22630 = n4060 | n5642 ;
  assign n22631 = n22630 ^ n12475 ^ 1'b0 ;
  assign n22632 = n22631 ^ n2896 ^ x144 ;
  assign n22633 = ( n3874 & ~n8301 ) | ( n3874 & n22632 ) | ( ~n8301 & n22632 ) ;
  assign n22634 = n19472 ^ n1302 ^ 1'b0 ;
  assign n22635 = ~n22633 & n22634 ;
  assign n22636 = ~n22629 & n22635 ;
  assign n22637 = n2324 & n22636 ;
  assign n22638 = ( n9562 & n11123 ) | ( n9562 & ~n20755 ) | ( n11123 & ~n20755 ) ;
  assign n22639 = n22638 ^ n15244 ^ 1'b0 ;
  assign n22643 = n3242 ^ n1957 ^ 1'b0 ;
  assign n22644 = n2592 & n22643 ;
  assign n22640 = n13353 ^ n4978 ^ 1'b0 ;
  assign n22641 = ~n6227 & n22640 ;
  assign n22642 = ~n7480 & n22641 ;
  assign n22645 = n22644 ^ n22642 ^ 1'b0 ;
  assign n22646 = n1472 ^ n871 ^ 1'b0 ;
  assign n22647 = ( n5188 & n11192 ) | ( n5188 & n22646 ) | ( n11192 & n22646 ) ;
  assign n22648 = n15362 & n22647 ;
  assign n22649 = n22648 ^ n3592 ^ 1'b0 ;
  assign n22650 = n9319 ^ n9277 ^ n4121 ;
  assign n22651 = n15449 ^ n9658 ^ 1'b0 ;
  assign n22652 = n22651 ^ n20414 ^ n5863 ;
  assign n22653 = n5002 | n22652 ;
  assign n22654 = n22653 ^ n5108 ^ 1'b0 ;
  assign n22655 = n12186 | n20240 ;
  assign n22656 = n9248 ^ n3080 ^ n3010 ;
  assign n22657 = n2243 & ~n22656 ;
  assign n22658 = n22657 ^ n4145 ^ 1'b0 ;
  assign n22659 = n22658 ^ n2067 ^ 1'b0 ;
  assign n22660 = ~n7810 & n22659 ;
  assign n22661 = ( n3114 & ~n22081 ) | ( n3114 & n22660 ) | ( ~n22081 & n22660 ) ;
  assign n22662 = n2424 ^ n2109 ^ 1'b0 ;
  assign n22663 = ~n7669 & n22662 ;
  assign n22664 = n22663 ^ n5340 ^ 1'b0 ;
  assign n22665 = n22664 ^ n13829 ^ 1'b0 ;
  assign n22666 = n22256 ^ n18401 ^ n11866 ;
  assign n22667 = n17221 ^ n14683 ^ 1'b0 ;
  assign n22668 = ( n20406 & ~n22666 ) | ( n20406 & n22667 ) | ( ~n22666 & n22667 ) ;
  assign n22669 = n14690 ^ n4642 ^ 1'b0 ;
  assign n22670 = n9570 & n22669 ;
  assign n22671 = n22670 ^ n679 ^ 1'b0 ;
  assign n22672 = ( ~n2163 & n9520 ) | ( ~n2163 & n18679 ) | ( n9520 & n18679 ) ;
  assign n22674 = n5419 ^ n4776 ^ n4326 ;
  assign n22673 = n18471 ^ n8262 ^ n5279 ;
  assign n22675 = n22674 ^ n22673 ^ 1'b0 ;
  assign n22676 = ~n6739 & n13196 ;
  assign n22677 = n8671 & ~n9597 ;
  assign n22678 = n22677 ^ n8915 ^ 1'b0 ;
  assign n22679 = ( n7588 & ~n22676 ) | ( n7588 & n22678 ) | ( ~n22676 & n22678 ) ;
  assign n22680 = n12214 ^ n12168 ^ n3845 ;
  assign n22681 = n22680 ^ n4042 ^ 1'b0 ;
  assign n22682 = n9976 ^ n5038 ^ x183 ;
  assign n22683 = n22682 ^ n7936 ^ 1'b0 ;
  assign n22684 = n13217 | n22683 ;
  assign n22685 = n3535 ^ n2147 ^ n1727 ;
  assign n22686 = n5966 & n22685 ;
  assign n22687 = ~n352 & n22686 ;
  assign n22688 = n22687 ^ n11962 ^ n1524 ;
  assign n22689 = n11868 ^ n1950 ^ 1'b0 ;
  assign n22690 = ~n16317 & n22689 ;
  assign n22691 = ~n13279 & n14087 ;
  assign n22692 = n17693 & n22691 ;
  assign n22693 = ( n7929 & n18071 ) | ( n7929 & n22692 ) | ( n18071 & n22692 ) ;
  assign n22694 = ( n4399 & n22690 ) | ( n4399 & ~n22693 ) | ( n22690 & ~n22693 ) ;
  assign n22697 = n7595 ^ n3241 ^ n1358 ;
  assign n22698 = n22697 ^ n15498 ^ 1'b0 ;
  assign n22695 = ~n296 & n11226 ;
  assign n22696 = n22695 ^ n9122 ^ 1'b0 ;
  assign n22699 = n22698 ^ n22696 ^ n346 ;
  assign n22700 = ( n1593 & ~n16160 ) | ( n1593 & n19897 ) | ( ~n16160 & n19897 ) ;
  assign n22701 = ( n711 & n3441 ) | ( n711 & ~n7958 ) | ( n3441 & ~n7958 ) ;
  assign n22704 = n15045 ^ n4693 ^ n1723 ;
  assign n22702 = n21525 ^ n17639 ^ 1'b0 ;
  assign n22703 = n22702 ^ n11139 ^ 1'b0 ;
  assign n22705 = n22704 ^ n22703 ^ n12263 ;
  assign n22706 = ( n1893 & n8514 ) | ( n1893 & ~n20464 ) | ( n8514 & ~n20464 ) ;
  assign n22707 = n21294 ^ n17203 ^ n11929 ;
  assign n22708 = ( ~x229 & n2797 ) | ( ~x229 & n6565 ) | ( n2797 & n6565 ) ;
  assign n22709 = n14146 | n22708 ;
  assign n22710 = n22709 ^ n1725 ^ 1'b0 ;
  assign n22711 = ( ~n1351 & n1390 ) | ( ~n1351 & n3554 ) | ( n1390 & n3554 ) ;
  assign n22712 = n22711 ^ n20310 ^ 1'b0 ;
  assign n22713 = n22712 ^ n18415 ^ 1'b0 ;
  assign n22714 = n22710 & ~n22713 ;
  assign n22715 = n19527 & n22347 ;
  assign n22716 = ~n17700 & n22715 ;
  assign n22717 = n16742 ^ n14360 ^ n6266 ;
  assign n22718 = n14148 ^ n7108 ^ 1'b0 ;
  assign n22719 = ~n22717 & n22718 ;
  assign n22720 = n16332 ^ n7581 ^ n5642 ;
  assign n22721 = ( n858 & n6678 ) | ( n858 & n22720 ) | ( n6678 & n22720 ) ;
  assign n22722 = n6639 & n9788 ;
  assign n22723 = n22722 ^ n3070 ^ n1442 ;
  assign n22724 = n11380 ^ n7222 ^ 1'b0 ;
  assign n22725 = ( ~n2627 & n13130 ) | ( ~n2627 & n19561 ) | ( n13130 & n19561 ) ;
  assign n22726 = n16487 & ~n17822 ;
  assign n22727 = n12429 ^ n4654 ^ 1'b0 ;
  assign n22728 = n10418 ^ n6320 ^ 1'b0 ;
  assign n22729 = n5057 ^ n3784 ^ 1'b0 ;
  assign n22730 = n11617 & ~n22729 ;
  assign n22731 = ~n4980 & n22730 ;
  assign n22732 = ( n910 & n7211 ) | ( n910 & ~n22731 ) | ( n7211 & ~n22731 ) ;
  assign n22733 = ( n10616 & n12331 ) | ( n10616 & n22732 ) | ( n12331 & n22732 ) ;
  assign n22736 = ( ~n6468 & n9205 ) | ( ~n6468 & n12461 ) | ( n9205 & n12461 ) ;
  assign n22735 = n5949 ^ n4462 ^ n3420 ;
  assign n22734 = n8017 ^ n6006 ^ n883 ;
  assign n22737 = n22736 ^ n22735 ^ n22734 ;
  assign n22738 = n22737 ^ n16670 ^ n8429 ;
  assign n22739 = n6214 | n8883 ;
  assign n22740 = ( ~n5435 & n16929 ) | ( ~n5435 & n22739 ) | ( n16929 & n22739 ) ;
  assign n22741 = n10560 & ~n14147 ;
  assign n22742 = ~n11881 & n22741 ;
  assign n22743 = n19340 ^ n7801 ^ 1'b0 ;
  assign n22744 = x235 & ~n22743 ;
  assign n22747 = n12585 ^ n7689 ^ n3931 ;
  assign n22748 = n22747 ^ n19535 ^ n2154 ;
  assign n22745 = n2960 & n19142 ;
  assign n22746 = n22745 ^ n7171 ^ 1'b0 ;
  assign n22749 = n22748 ^ n22746 ^ n3626 ;
  assign n22750 = ( ~n722 & n22744 ) | ( ~n722 & n22749 ) | ( n22744 & n22749 ) ;
  assign n22751 = n22750 ^ n14730 ^ 1'b0 ;
  assign n22752 = n10550 ^ n4636 ^ 1'b0 ;
  assign n22753 = n17954 & n22752 ;
  assign n22754 = n22753 ^ n6633 ^ 1'b0 ;
  assign n22758 = ( ~n4052 & n11975 ) | ( ~n4052 & n16825 ) | ( n11975 & n16825 ) ;
  assign n22755 = n5380 ^ n2562 ^ 1'b0 ;
  assign n22756 = n5643 & n22755 ;
  assign n22757 = n22756 ^ n19280 ^ 1'b0 ;
  assign n22759 = n22758 ^ n22757 ^ n11473 ;
  assign n22760 = n13118 ^ n5580 ^ n1710 ;
  assign n22761 = ~n6550 & n22760 ;
  assign n22762 = n22761 ^ n1675 ^ 1'b0 ;
  assign n22763 = n18545 ^ n13932 ^ n610 ;
  assign n22764 = ~n8074 & n12076 ;
  assign n22765 = n22764 ^ n3942 ^ 1'b0 ;
  assign n22766 = n13603 ^ n9203 ^ 1'b0 ;
  assign n22767 = ( n3416 & n22765 ) | ( n3416 & ~n22766 ) | ( n22765 & ~n22766 ) ;
  assign n22768 = n1620 | n5126 ;
  assign n22769 = ( n11895 & ~n13590 ) | ( n11895 & n22768 ) | ( ~n13590 & n22768 ) ;
  assign n22770 = n9983 | n22769 ;
  assign n22771 = n13069 ^ n7828 ^ 1'b0 ;
  assign n22772 = n22770 & n22771 ;
  assign n22773 = n17799 ^ n871 ^ 1'b0 ;
  assign n22774 = n12356 & ~n22773 ;
  assign n22775 = n14507 & n22774 ;
  assign n22776 = n15258 ^ n9848 ^ n8927 ;
  assign n22777 = n19991 | n22776 ;
  assign n22778 = n12600 & ~n22777 ;
  assign n22779 = n22778 ^ n8526 ^ 1'b0 ;
  assign n22780 = n22779 ^ n1086 ^ 1'b0 ;
  assign n22781 = n19584 & ~n22780 ;
  assign n22782 = ( n17957 & n21004 ) | ( n17957 & ~n22781 ) | ( n21004 & ~n22781 ) ;
  assign n22783 = n4139 ^ n1254 ^ 1'b0 ;
  assign n22784 = n9052 & n13435 ;
  assign n22785 = n22784 ^ n8802 ^ 1'b0 ;
  assign n22786 = n6917 ^ n2510 ^ 1'b0 ;
  assign n22787 = n12082 | n22786 ;
  assign n22788 = n10460 | n22787 ;
  assign n22789 = n22788 ^ n4646 ^ 1'b0 ;
  assign n22790 = n6920 & ~n10587 ;
  assign n22791 = ~x139 & n22790 ;
  assign n22792 = ( n1086 & ~n5918 ) | ( n1086 & n22791 ) | ( ~n5918 & n22791 ) ;
  assign n22793 = n22792 ^ n13820 ^ n695 ;
  assign n22794 = n20203 ^ n17765 ^ n12338 ;
  assign n22795 = n19324 ^ n12240 ^ n12106 ;
  assign n22796 = n15184 ^ n1262 ^ 1'b0 ;
  assign n22797 = ~n22795 & n22796 ;
  assign n22798 = n9983 ^ n6787 ^ 1'b0 ;
  assign n22799 = n9176 & n22798 ;
  assign n22801 = ~n6031 & n14790 ;
  assign n22800 = n9399 ^ n8282 ^ n3880 ;
  assign n22802 = n22801 ^ n22800 ^ n6330 ;
  assign n22803 = n15508 & ~n22802 ;
  assign n22804 = ~n22799 & n22803 ;
  assign n22805 = n15368 ^ n8212 ^ 1'b0 ;
  assign n22806 = n11455 & n22805 ;
  assign n22807 = n5200 ^ n3643 ^ 1'b0 ;
  assign n22808 = n9620 ^ n370 ^ 1'b0 ;
  assign n22809 = ~n7021 & n22808 ;
  assign n22810 = n6337 & n22809 ;
  assign n22811 = n20925 & n22810 ;
  assign n22812 = n22807 | n22811 ;
  assign n22813 = n22812 ^ x147 ^ 1'b0 ;
  assign n22814 = n16509 & n17513 ;
  assign n22815 = ( n6743 & ~n8451 ) | ( n6743 & n14679 ) | ( ~n8451 & n14679 ) ;
  assign n22816 = n22815 ^ n9365 ^ n474 ;
  assign n22817 = n1264 & ~n9104 ;
  assign n22818 = ( ~n2538 & n11868 ) | ( ~n2538 & n17979 ) | ( n11868 & n17979 ) ;
  assign n22820 = n3010 | n11105 ;
  assign n22821 = n22820 ^ n14423 ^ n341 ;
  assign n22819 = ~n5006 & n7365 ;
  assign n22822 = n22821 ^ n22819 ^ 1'b0 ;
  assign n22823 = ( ~n520 & n11607 ) | ( ~n520 & n22822 ) | ( n11607 & n22822 ) ;
  assign n22824 = ~n3621 & n13502 ;
  assign n22825 = ( n1617 & n9945 ) | ( n1617 & ~n22824 ) | ( n9945 & ~n22824 ) ;
  assign n22826 = ~n11012 & n22825 ;
  assign n22827 = ~n12890 & n22826 ;
  assign n22828 = ( n21788 & ~n21790 ) | ( n21788 & n22827 ) | ( ~n21790 & n22827 ) ;
  assign n22829 = ( n617 & ~n2306 ) | ( n617 & n6220 ) | ( ~n2306 & n6220 ) ;
  assign n22830 = n22829 ^ n15518 ^ 1'b0 ;
  assign n22831 = ( ~n2634 & n10587 ) | ( ~n2634 & n22830 ) | ( n10587 & n22830 ) ;
  assign n22832 = n17653 ^ n10500 ^ 1'b0 ;
  assign n22833 = ~n327 & n22832 ;
  assign n22836 = ~n6307 & n10617 ;
  assign n22834 = n11721 ^ n10773 ^ n8384 ;
  assign n22835 = n13580 & n22834 ;
  assign n22837 = n22836 ^ n22835 ^ 1'b0 ;
  assign n22838 = n6769 & ~n15513 ;
  assign n22846 = ( n2310 & ~n4612 ) | ( n2310 & n9713 ) | ( ~n4612 & n9713 ) ;
  assign n22839 = ( n1415 & n3987 ) | ( n1415 & n5316 ) | ( n3987 & n5316 ) ;
  assign n22840 = n22839 ^ n4153 ^ 1'b0 ;
  assign n22841 = n2492 | n22840 ;
  assign n22842 = n22841 ^ n14903 ^ 1'b0 ;
  assign n22843 = n22842 ^ n21439 ^ n12947 ;
  assign n22844 = n16330 | n22843 ;
  assign n22845 = n4981 & ~n22844 ;
  assign n22847 = n22846 ^ n22845 ^ 1'b0 ;
  assign n22848 = ~n22838 & n22847 ;
  assign n22852 = n3729 & n15651 ;
  assign n22853 = n22852 ^ n8693 ^ 1'b0 ;
  assign n22854 = n22853 ^ n13209 ^ n5367 ;
  assign n22849 = n8369 ^ n6674 ^ n5842 ;
  assign n22850 = ( n11239 & n15300 ) | ( n11239 & ~n22849 ) | ( n15300 & ~n22849 ) ;
  assign n22851 = ~n14980 & n22850 ;
  assign n22855 = n22854 ^ n22851 ^ 1'b0 ;
  assign n22856 = ( n1589 & n5217 ) | ( n1589 & n20066 ) | ( n5217 & n20066 ) ;
  assign n22857 = n22856 ^ n20937 ^ n10230 ;
  assign n22858 = ( ~x127 & n6232 ) | ( ~x127 & n18779 ) | ( n6232 & n18779 ) ;
  assign n22864 = n9206 ^ n4876 ^ 1'b0 ;
  assign n22859 = n5400 | n5990 ;
  assign n22860 = n735 & n7008 ;
  assign n22861 = ~n11848 & n22860 ;
  assign n22862 = ( n2728 & n22859 ) | ( n2728 & ~n22861 ) | ( n22859 & ~n22861 ) ;
  assign n22863 = n13367 & n22862 ;
  assign n22865 = n22864 ^ n22863 ^ n1548 ;
  assign n22871 = n801 & n21693 ;
  assign n22872 = n22871 ^ n6298 ^ 1'b0 ;
  assign n22866 = ( n3430 & n3908 ) | ( n3430 & n15078 ) | ( n3908 & n15078 ) ;
  assign n22867 = n10153 | n22866 ;
  assign n22868 = n10408 | n22867 ;
  assign n22869 = n22868 ^ n5305 ^ n1040 ;
  assign n22870 = n4638 | n22869 ;
  assign n22873 = n22872 ^ n22870 ^ 1'b0 ;
  assign n22874 = n20432 ^ n5725 ^ 1'b0 ;
  assign n22875 = n4303 & n22874 ;
  assign n22876 = n22875 ^ n8684 ^ n5543 ;
  assign n22877 = ( x39 & n18630 ) | ( x39 & ~n22876 ) | ( n18630 & ~n22876 ) ;
  assign n22878 = ( n866 & n5539 ) | ( n866 & n22877 ) | ( n5539 & n22877 ) ;
  assign n22879 = n549 | n1337 ;
  assign n22880 = n16063 | n22879 ;
  assign n22881 = ( n2458 & n9286 ) | ( n2458 & n22880 ) | ( n9286 & n22880 ) ;
  assign n22882 = ( n1890 & n8996 ) | ( n1890 & n9895 ) | ( n8996 & n9895 ) ;
  assign n22883 = n22882 ^ n8074 ^ 1'b0 ;
  assign n22884 = n12974 & ~n22883 ;
  assign n22885 = n22884 ^ n10182 ^ n514 ;
  assign n22886 = ( ~n9160 & n10068 ) | ( ~n9160 & n16230 ) | ( n10068 & n16230 ) ;
  assign n22887 = ( n3718 & ~n4454 ) | ( n3718 & n22886 ) | ( ~n4454 & n22886 ) ;
  assign n22888 = n19730 ^ n13939 ^ 1'b0 ;
  assign n22889 = n14178 | n22888 ;
  assign n22890 = ( n13796 & n15601 ) | ( n13796 & n22889 ) | ( n15601 & n22889 ) ;
  assign n22891 = n8247 ^ n4076 ^ n3821 ;
  assign n22892 = n1697 | n22891 ;
  assign n22893 = n13164 | n22892 ;
  assign n22894 = n22890 | n22893 ;
  assign n22895 = n15045 ^ n1336 ^ 1'b0 ;
  assign n22896 = n1968 & ~n22895 ;
  assign n22897 = n22896 ^ x14 ^ 1'b0 ;
  assign n22898 = n13678 & n22897 ;
  assign n22899 = n555 & ~n3772 ;
  assign n22900 = n22899 ^ n16473 ^ 1'b0 ;
  assign n22902 = ~n1524 & n3675 ;
  assign n22903 = n9012 ^ n6647 ^ n2513 ;
  assign n22904 = ( n11704 & n22902 ) | ( n11704 & ~n22903 ) | ( n22902 & ~n22903 ) ;
  assign n22901 = n5876 | n11965 ;
  assign n22905 = n22904 ^ n22901 ^ n11106 ;
  assign n22906 = n282 & ~n9267 ;
  assign n22907 = n19341 ^ n4319 ^ 1'b0 ;
  assign n22908 = ( n3370 & ~n22638 ) | ( n3370 & n22907 ) | ( ~n22638 & n22907 ) ;
  assign n22909 = n6628 | n10570 ;
  assign n22910 = n22909 ^ n2582 ^ 1'b0 ;
  assign n22911 = n9938 ^ n665 ^ n654 ;
  assign n22912 = n22910 | n22911 ;
  assign n22913 = ~n3623 & n4612 ;
  assign n22914 = n20441 ^ n5408 ^ 1'b0 ;
  assign n22915 = n22914 ^ n6495 ^ n1228 ;
  assign n22916 = n14347 ^ n800 ^ 1'b0 ;
  assign n22917 = n13694 ^ n7990 ^ 1'b0 ;
  assign n22918 = n22917 ^ n3807 ^ 1'b0 ;
  assign n22919 = ( n10177 & n20691 ) | ( n10177 & ~n22223 ) | ( n20691 & ~n22223 ) ;
  assign n22920 = ( n2778 & n3482 ) | ( n2778 & n9601 ) | ( n3482 & n9601 ) ;
  assign n22921 = ( n1693 & n6864 ) | ( n1693 & ~n10976 ) | ( n6864 & ~n10976 ) ;
  assign n22922 = n6783 ^ n5643 ^ n2753 ;
  assign n22923 = n7547 ^ n6440 ^ n3847 ;
  assign n22924 = ~n22922 & n22923 ;
  assign n22925 = n22921 & n22924 ;
  assign n22926 = ( n19777 & n22920 ) | ( n19777 & n22925 ) | ( n22920 & n22925 ) ;
  assign n22927 = n3283 ^ n577 ^ n463 ;
  assign n22928 = ( n4336 & ~n21793 ) | ( n4336 & n22927 ) | ( ~n21793 & n22927 ) ;
  assign n22929 = n9658 | n22928 ;
  assign n22930 = ( n772 & n8491 ) | ( n772 & n12032 ) | ( n8491 & n12032 ) ;
  assign n22931 = n723 & n3643 ;
  assign n22932 = ( n20483 & n22930 ) | ( n20483 & ~n22931 ) | ( n22930 & ~n22931 ) ;
  assign n22933 = n18893 ^ n2407 ^ 1'b0 ;
  assign n22934 = ( ~n4032 & n5676 ) | ( ~n4032 & n22933 ) | ( n5676 & n22933 ) ;
  assign n22937 = n595 & n662 ;
  assign n22938 = n22937 ^ n1597 ^ 1'b0 ;
  assign n22939 = n22938 ^ n4606 ^ n1781 ;
  assign n22935 = n12334 ^ n6797 ^ 1'b0 ;
  assign n22936 = n18197 & ~n22935 ;
  assign n22940 = n22939 ^ n22936 ^ n15538 ;
  assign n22941 = ~n2515 & n4298 ;
  assign n22942 = n22941 ^ n19948 ^ 1'b0 ;
  assign n22943 = n14619 ^ n508 ^ 1'b0 ;
  assign n22944 = n22943 ^ n19801 ^ 1'b0 ;
  assign n22945 = n5475 & n22944 ;
  assign n22946 = n22945 ^ n7682 ^ 1'b0 ;
  assign n22947 = n22942 | n22946 ;
  assign n22948 = ~n2480 & n17035 ;
  assign n22949 = n21706 ^ n6353 ^ 1'b0 ;
  assign n22950 = ~n13354 & n22949 ;
  assign n22951 = ( n1978 & n2270 ) | ( n1978 & n10222 ) | ( n2270 & n10222 ) ;
  assign n22960 = n701 & ~n18590 ;
  assign n22961 = n684 & n7219 ;
  assign n22962 = n22961 ^ n1534 ^ 1'b0 ;
  assign n22963 = ~n22960 & n22962 ;
  assign n22956 = ~n9686 & n10881 ;
  assign n22957 = ~n4317 & n22956 ;
  assign n22958 = n21119 & ~n22957 ;
  assign n22959 = n9204 & n22958 ;
  assign n22952 = n14462 | n22921 ;
  assign n22953 = n22952 ^ n10118 ^ 1'b0 ;
  assign n22954 = n562 | n22953 ;
  assign n22955 = n4391 | n22954 ;
  assign n22964 = n22963 ^ n22959 ^ n22955 ;
  assign n22965 = n22964 ^ n20522 ^ n19123 ;
  assign n22966 = ( ~n19621 & n22951 ) | ( ~n19621 & n22965 ) | ( n22951 & n22965 ) ;
  assign n22967 = n16095 & ~n21406 ;
  assign n22968 = ( ~n5459 & n8955 ) | ( ~n5459 & n18402 ) | ( n8955 & n18402 ) ;
  assign n22969 = n8320 ^ n811 ^ 1'b0 ;
  assign n22970 = n7541 & ~n22969 ;
  assign n22971 = n10814 & ~n22970 ;
  assign n22972 = ~n2020 & n15398 ;
  assign n22973 = ( n5152 & n19045 ) | ( n5152 & n22972 ) | ( n19045 & n22972 ) ;
  assign n22974 = ( n1211 & n2030 ) | ( n1211 & n16079 ) | ( n2030 & n16079 ) ;
  assign n22975 = n5890 ^ n900 ^ n793 ;
  assign n22976 = ~n3346 & n22975 ;
  assign n22977 = n3353 & n22976 ;
  assign n22978 = n22974 | n22977 ;
  assign n22979 = n1558 & n11917 ;
  assign n22980 = n22979 ^ n8203 ^ 1'b0 ;
  assign n22981 = n22980 ^ n5833 ^ 1'b0 ;
  assign n22982 = n8487 & n22981 ;
  assign n22983 = ( ~n378 & n7230 ) | ( ~n378 & n19566 ) | ( n7230 & n19566 ) ;
  assign n22984 = n4826 | n22983 ;
  assign n22985 = n6356 | n22984 ;
  assign n22986 = ~n7665 & n22985 ;
  assign n22987 = n12532 ^ n12219 ^ 1'b0 ;
  assign n22988 = ~n19564 & n22987 ;
  assign n22989 = n2443 & ~n22988 ;
  assign n22990 = n20466 & n20956 ;
  assign n22991 = n4908 & n22990 ;
  assign n22992 = ( n5430 & ~n19882 ) | ( n5430 & n22991 ) | ( ~n19882 & n22991 ) ;
  assign n22993 = n14090 ^ n8602 ^ 1'b0 ;
  assign n22994 = ( ~n8524 & n14682 ) | ( ~n8524 & n20160 ) | ( n14682 & n20160 ) ;
  assign n22995 = n22957 ^ n18861 ^ n18471 ;
  assign n22996 = ( ~n5277 & n5328 ) | ( ~n5277 & n22182 ) | ( n5328 & n22182 ) ;
  assign n22997 = n22996 ^ n14319 ^ n2743 ;
  assign n22998 = n22997 ^ n15620 ^ 1'b0 ;
  assign n22999 = n6828 & ~n22998 ;
  assign n23002 = n2048 | n8239 ;
  assign n23000 = n12151 | n13163 ;
  assign n23001 = ( n4024 & n15328 ) | ( n4024 & n23000 ) | ( n15328 & n23000 ) ;
  assign n23003 = n23002 ^ n23001 ^ n18934 ;
  assign n23004 = n21986 ^ n2874 ^ 1'b0 ;
  assign n23005 = n23003 & ~n23004 ;
  assign n23006 = n14374 ^ n6884 ^ 1'b0 ;
  assign n23007 = n8888 ^ n2756 ^ 1'b0 ;
  assign n23008 = n23007 ^ n21456 ^ 1'b0 ;
  assign n23009 = n740 | n23008 ;
  assign n23010 = n23009 ^ n22970 ^ n3160 ;
  assign n23011 = n4040 ^ n2259 ^ 1'b0 ;
  assign n23012 = n2609 & n23011 ;
  assign n23013 = ( n11160 & n12125 ) | ( n11160 & n23012 ) | ( n12125 & n23012 ) ;
  assign n23014 = n23013 ^ n2444 ^ n1839 ;
  assign n23015 = ( n395 & ~n11390 ) | ( n395 & n12123 ) | ( ~n11390 & n12123 ) ;
  assign n23016 = ( n8728 & n23014 ) | ( n8728 & n23015 ) | ( n23014 & n23015 ) ;
  assign n23017 = n11578 ^ n5383 ^ 1'b0 ;
  assign n23018 = n13335 ^ n2944 ^ 1'b0 ;
  assign n23019 = n1590 & n22330 ;
  assign n23020 = n23019 ^ n4014 ^ 1'b0 ;
  assign n23021 = n23020 ^ n2930 ^ 1'b0 ;
  assign n23022 = ~n920 & n5504 ;
  assign n23023 = n18937 ^ n3274 ^ 1'b0 ;
  assign n23024 = n11035 ^ n10596 ^ 1'b0 ;
  assign n23025 = ~n14150 & n23024 ;
  assign n23026 = ( n12338 & n23023 ) | ( n12338 & n23025 ) | ( n23023 & n23025 ) ;
  assign n23027 = n23026 ^ n12578 ^ n6863 ;
  assign n23028 = ( ~n14384 & n23022 ) | ( ~n14384 & n23027 ) | ( n23022 & n23027 ) ;
  assign n23029 = n19831 ^ n12070 ^ n437 ;
  assign n23030 = n23029 ^ n16328 ^ n9496 ;
  assign n23033 = n10626 | n22680 ;
  assign n23034 = n15008 & ~n23033 ;
  assign n23031 = n12070 ^ n4709 ^ 1'b0 ;
  assign n23032 = ~n6990 & n23031 ;
  assign n23035 = n23034 ^ n23032 ^ n14697 ;
  assign n23037 = ( n2556 & n4194 ) | ( n2556 & n14451 ) | ( n4194 & n14451 ) ;
  assign n23038 = ( n6917 & n9675 ) | ( n6917 & ~n23037 ) | ( n9675 & ~n23037 ) ;
  assign n23036 = n7899 & n13856 ;
  assign n23039 = n23038 ^ n23036 ^ 1'b0 ;
  assign n23040 = n23039 ^ n3076 ^ 1'b0 ;
  assign n23041 = n7207 ^ n3109 ^ 1'b0 ;
  assign n23042 = ~n5282 & n13100 ;
  assign n23043 = n6160 & n23042 ;
  assign n23044 = n23043 ^ n16431 ^ n8214 ;
  assign n23045 = n16408 ^ n14537 ^ n11633 ;
  assign n23046 = ( n1025 & ~n3154 ) | ( n1025 & n11740 ) | ( ~n3154 & n11740 ) ;
  assign n23047 = n23046 ^ n18266 ^ 1'b0 ;
  assign n23048 = n23047 ^ n16625 ^ 1'b0 ;
  assign n23049 = n19849 ^ n16174 ^ 1'b0 ;
  assign n23050 = n9996 & n23049 ;
  assign n23051 = ~n1961 & n23050 ;
  assign n23052 = ~n11192 & n23051 ;
  assign n23053 = n8494 & ~n23052 ;
  assign n23054 = ( ~n2973 & n6784 ) | ( ~n2973 & n12647 ) | ( n6784 & n12647 ) ;
  assign n23055 = ~n22842 & n23054 ;
  assign n23056 = n12708 | n23055 ;
  assign n23057 = n6328 & ~n23056 ;
  assign n23058 = n3106 & ~n3650 ;
  assign n23059 = n23058 ^ n930 ^ 1'b0 ;
  assign n23060 = n23059 ^ n13345 ^ 1'b0 ;
  assign n23061 = ~n13737 & n23060 ;
  assign n23062 = n14211 ^ n11974 ^ 1'b0 ;
  assign n23063 = n19161 & n23062 ;
  assign n23064 = n9320 ^ n2592 ^ 1'b0 ;
  assign n23065 = n17643 ^ n16428 ^ 1'b0 ;
  assign n23066 = n10058 | n17336 ;
  assign n23067 = ( n9713 & n11620 ) | ( n9713 & ~n23066 ) | ( n11620 & ~n23066 ) ;
  assign n23068 = n16013 | n23067 ;
  assign n23069 = n23068 ^ n10935 ^ 1'b0 ;
  assign n23070 = ( ~n1198 & n4568 ) | ( ~n1198 & n6064 ) | ( n4568 & n6064 ) ;
  assign n23071 = n7356 | n23070 ;
  assign n23072 = n8270 & ~n23071 ;
  assign n23073 = n23072 ^ n15207 ^ 1'b0 ;
  assign n23074 = n10228 ^ n8753 ^ n3005 ;
  assign n23075 = n23074 ^ n11579 ^ n2927 ;
  assign n23076 = n13030 ^ n2592 ^ 1'b0 ;
  assign n23077 = n10086 | n23076 ;
  assign n23078 = n23077 ^ n16268 ^ n7535 ;
  assign n23079 = n13259 ^ n5162 ^ 1'b0 ;
  assign n23080 = n21442 & n23079 ;
  assign n23081 = n10681 & n23080 ;
  assign n23082 = n11995 ^ n3068 ^ 1'b0 ;
  assign n23083 = ~n23081 & n23082 ;
  assign n23084 = n1065 & n11542 ;
  assign n23085 = n23084 ^ n18269 ^ 1'b0 ;
  assign n23088 = ( ~n636 & n14035 ) | ( ~n636 & n16177 ) | ( n14035 & n16177 ) ;
  assign n23086 = n15382 ^ n9555 ^ 1'b0 ;
  assign n23087 = ~n12352 & n23086 ;
  assign n23089 = n23088 ^ n23087 ^ n13929 ;
  assign n23090 = ( n5396 & n16691 ) | ( n5396 & ~n22561 ) | ( n16691 & ~n22561 ) ;
  assign n23091 = n15739 ^ n5377 ^ 1'b0 ;
  assign n23092 = n15986 ^ n14799 ^ n6934 ;
  assign n23093 = ( n11438 & n12872 ) | ( n11438 & n23092 ) | ( n12872 & n23092 ) ;
  assign n23094 = n23091 & n23093 ;
  assign n23095 = n23029 & n23094 ;
  assign n23096 = ( n6249 & n23090 ) | ( n6249 & ~n23095 ) | ( n23090 & ~n23095 ) ;
  assign n23097 = n21385 ^ x152 ^ 1'b0 ;
  assign n23098 = ~n7542 & n23097 ;
  assign n23099 = ( ~n3831 & n4197 ) | ( ~n3831 & n4506 ) | ( n4197 & n4506 ) ;
  assign n23100 = n17381 ^ n6430 ^ 1'b0 ;
  assign n23101 = ( ~n437 & n5831 ) | ( ~n437 & n23100 ) | ( n5831 & n23100 ) ;
  assign n23102 = n17937 ^ n7047 ^ 1'b0 ;
  assign n23103 = n23102 ^ n974 ^ 1'b0 ;
  assign n23104 = ~n19178 & n23103 ;
  assign n23105 = x9 & n23104 ;
  assign n23106 = n11727 & n23105 ;
  assign n23107 = ( ~n23099 & n23101 ) | ( ~n23099 & n23106 ) | ( n23101 & n23106 ) ;
  assign n23113 = ( n3294 & n3320 ) | ( n3294 & n10974 ) | ( n3320 & n10974 ) ;
  assign n23108 = ~n7966 & n15889 ;
  assign n23109 = ~n10170 & n23108 ;
  assign n23110 = n5032 & ~n23109 ;
  assign n23111 = ( ~n392 & n14325 ) | ( ~n392 & n23110 ) | ( n14325 & n23110 ) ;
  assign n23112 = ( n12887 & n19931 ) | ( n12887 & n23111 ) | ( n19931 & n23111 ) ;
  assign n23114 = n23113 ^ n23112 ^ n1278 ;
  assign n23115 = ( n9404 & n20377 ) | ( n9404 & n20639 ) | ( n20377 & n20639 ) ;
  assign n23116 = ~n799 & n5391 ;
  assign n23117 = n23116 ^ n6330 ^ 1'b0 ;
  assign n23118 = n12239 ^ n10195 ^ n625 ;
  assign n23123 = n16891 ^ n9277 ^ 1'b0 ;
  assign n23119 = n3630 ^ n1109 ^ 1'b0 ;
  assign n23120 = ~n2000 & n23119 ;
  assign n23121 = ( ~n2779 & n5865 ) | ( ~n2779 & n23120 ) | ( n5865 & n23120 ) ;
  assign n23122 = n6055 & n23121 ;
  assign n23124 = n23123 ^ n23122 ^ 1'b0 ;
  assign n23125 = n18040 ^ n11149 ^ 1'b0 ;
  assign n23126 = ( n8321 & n17107 ) | ( n8321 & n23125 ) | ( n17107 & n23125 ) ;
  assign n23127 = n15036 ^ n14239 ^ n7493 ;
  assign n23128 = n3563 | n8319 ;
  assign n23129 = n5723 & ~n23128 ;
  assign n23130 = ( x92 & n12244 ) | ( x92 & ~n23129 ) | ( n12244 & ~n23129 ) ;
  assign n23131 = ( ~n10828 & n17156 ) | ( ~n10828 & n23130 ) | ( n17156 & n23130 ) ;
  assign n23132 = n6509 | n13756 ;
  assign n23133 = n21861 ^ n19564 ^ n15034 ;
  assign n23134 = ( ~n12303 & n23132 ) | ( ~n12303 & n23133 ) | ( n23132 & n23133 ) ;
  assign n23137 = n988 ^ n824 ^ x25 ;
  assign n23138 = n23137 ^ n17012 ^ n12415 ;
  assign n23135 = n22545 ^ n6255 ^ 1'b0 ;
  assign n23136 = n23135 ^ n22923 ^ n5620 ;
  assign n23139 = n23138 ^ n23136 ^ 1'b0 ;
  assign n23140 = n8466 ^ n5753 ^ 1'b0 ;
  assign n23141 = n7736 & n23140 ;
  assign n23142 = n4618 | n23141 ;
  assign n23143 = n2889 & ~n23142 ;
  assign n23144 = ( n1372 & ~n2461 ) | ( n1372 & n4231 ) | ( ~n2461 & n4231 ) ;
  assign n23145 = ( n3264 & ~n18835 ) | ( n3264 & n23144 ) | ( ~n18835 & n23144 ) ;
  assign n23146 = n502 | n13158 ;
  assign n23147 = n23146 ^ n4402 ^ 1'b0 ;
  assign n23148 = ( n11645 & n23145 ) | ( n11645 & ~n23147 ) | ( n23145 & ~n23147 ) ;
  assign n23149 = n5908 & ~n6151 ;
  assign n23150 = n23149 ^ n6575 ^ 1'b0 ;
  assign n23151 = n23150 ^ n5382 ^ n857 ;
  assign n23152 = n23151 ^ n17013 ^ n14071 ;
  assign n23153 = n23152 ^ n3667 ^ 1'b0 ;
  assign n23154 = n11113 | n17455 ;
  assign n23155 = n23154 ^ n12231 ^ 1'b0 ;
  assign n23156 = n9580 ^ n3582 ^ n3160 ;
  assign n23157 = n23156 ^ n12392 ^ n4161 ;
  assign n23158 = n19502 ^ n15738 ^ 1'b0 ;
  assign n23159 = n23157 & n23158 ;
  assign n23160 = n17376 ^ n4988 ^ 1'b0 ;
  assign n23161 = n16053 & n23160 ;
  assign n23162 = n20709 ^ n18342 ^ n1515 ;
  assign n23163 = n18936 ^ n12967 ^ n2495 ;
  assign n23164 = n15235 ^ n6625 ^ n5700 ;
  assign n23165 = n7543 & n23164 ;
  assign n23166 = n1896 ^ n1313 ^ 1'b0 ;
  assign n23167 = n14360 & n23166 ;
  assign n23168 = n23167 ^ n16741 ^ 1'b0 ;
  assign n23169 = ( n779 & n7448 ) | ( n779 & n23168 ) | ( n7448 & n23168 ) ;
  assign n23170 = n9673 & ~n23169 ;
  assign n23177 = n12435 ^ n2791 ^ 1'b0 ;
  assign n23178 = n5512 | n23177 ;
  assign n23179 = n23178 ^ n1848 ^ 1'b0 ;
  assign n23171 = ~n4850 & n6030 ;
  assign n23172 = ~n1822 & n23171 ;
  assign n23173 = n23172 ^ n2418 ^ 1'b0 ;
  assign n23174 = ~n3732 & n23173 ;
  assign n23175 = ~n21098 & n23174 ;
  assign n23176 = n4546 & n23175 ;
  assign n23180 = n23179 ^ n23176 ^ 1'b0 ;
  assign n23181 = ~n23170 & n23180 ;
  assign n23182 = n4247 & n9916 ;
  assign n23183 = n23182 ^ n7479 ^ 1'b0 ;
  assign n23184 = ~n9599 & n23183 ;
  assign n23185 = ( ~n959 & n3762 ) | ( ~n959 & n10411 ) | ( n3762 & n10411 ) ;
  assign n23186 = n12141 | n23185 ;
  assign n23187 = n20564 ^ n17592 ^ 1'b0 ;
  assign n23188 = n11757 | n23187 ;
  assign n23189 = ~n2424 & n6706 ;
  assign n23190 = n23189 ^ n21299 ^ 1'b0 ;
  assign n23191 = ~n14906 & n23190 ;
  assign n23192 = ( n5718 & n7783 ) | ( n5718 & n12147 ) | ( n7783 & n12147 ) ;
  assign n23193 = ( ~n9290 & n10602 ) | ( ~n9290 & n23192 ) | ( n10602 & n23192 ) ;
  assign n23194 = n23193 ^ n10903 ^ 1'b0 ;
  assign n23195 = n3844 & n23194 ;
  assign n23196 = x15 & ~n23195 ;
  assign n23197 = ~n6022 & n7469 ;
  assign n23198 = n1919 & ~n23197 ;
  assign n23199 = n8958 & n23198 ;
  assign n23200 = ~n23196 & n23199 ;
  assign n23201 = n6149 & ~n23022 ;
  assign n23202 = n23201 ^ n2160 ^ 1'b0 ;
  assign n23203 = n5913 & n23202 ;
  assign n23204 = n23203 ^ n10811 ^ 1'b0 ;
  assign n23205 = n23204 ^ n21510 ^ n1044 ;
  assign n23206 = ~n3420 & n21321 ;
  assign n23207 = n23206 ^ n4692 ^ 1'b0 ;
  assign n23208 = n23207 ^ n18464 ^ n17333 ;
  assign n23209 = n6167 ^ n2271 ^ 1'b0 ;
  assign n23210 = n4111 ^ n587 ^ 1'b0 ;
  assign n23211 = n5063 | n23210 ;
  assign n23212 = n23209 & ~n23211 ;
  assign n23213 = ( n15707 & n16074 ) | ( n15707 & ~n23212 ) | ( n16074 & ~n23212 ) ;
  assign n23215 = n20925 ^ n2835 ^ 1'b0 ;
  assign n23216 = n6449 | n23215 ;
  assign n23214 = n1086 & ~n21742 ;
  assign n23217 = n23216 ^ n23214 ^ n21455 ;
  assign n23218 = n19661 ^ n14741 ^ 1'b0 ;
  assign n23219 = n23218 ^ n9989 ^ 1'b0 ;
  assign n23220 = ( n13557 & ~n16410 ) | ( n13557 & n16547 ) | ( ~n16410 & n16547 ) ;
  assign n23221 = n5084 & ~n23220 ;
  assign n23222 = n18867 ^ n8524 ^ 1'b0 ;
  assign n23223 = ( x31 & n4653 ) | ( x31 & ~n11022 ) | ( n4653 & ~n11022 ) ;
  assign n23224 = n23223 ^ n732 ^ 1'b0 ;
  assign n23225 = n10989 | n23224 ;
  assign n23227 = n1388 | n11040 ;
  assign n23228 = n4010 & ~n23227 ;
  assign n23226 = n18542 ^ n16287 ^ n2131 ;
  assign n23229 = n23228 ^ n23226 ^ n15301 ;
  assign n23230 = ~n14842 & n15835 ;
  assign n23231 = n1401 & ~n10021 ;
  assign n23232 = n23231 ^ n2260 ^ n675 ;
  assign n23233 = ( ~n636 & n4877 ) | ( ~n636 & n10830 ) | ( n4877 & n10830 ) ;
  assign n23234 = n23233 ^ n325 ^ 1'b0 ;
  assign n23235 = n23232 & ~n23234 ;
  assign n23236 = n19983 ^ n4702 ^ 1'b0 ;
  assign n23237 = n12962 & ~n17288 ;
  assign n23238 = n9187 ^ n3507 ^ 1'b0 ;
  assign n23239 = ( n1304 & ~n5619 ) | ( n1304 & n23238 ) | ( ~n5619 & n23238 ) ;
  assign n23240 = ( n342 & ~n18401 ) | ( n342 & n23239 ) | ( ~n18401 & n23239 ) ;
  assign n23241 = n15571 ^ n4965 ^ 1'b0 ;
  assign n23242 = n12426 & n23241 ;
  assign n23243 = n23242 ^ n18443 ^ 1'b0 ;
  assign n23244 = ( n12186 & ~n23240 ) | ( n12186 & n23243 ) | ( ~n23240 & n23243 ) ;
  assign n23245 = n10611 & n17759 ;
  assign n23246 = n23245 ^ n936 ^ 1'b0 ;
  assign n23247 = ( n5082 & ~n11507 ) | ( n5082 & n23246 ) | ( ~n11507 & n23246 ) ;
  assign n23248 = n4990 ^ n663 ^ 1'b0 ;
  assign n23249 = n14063 | n23248 ;
  assign n23251 = n13195 ^ n11490 ^ 1'b0 ;
  assign n23252 = n23251 ^ n16841 ^ 1'b0 ;
  assign n23253 = ~n22891 & n23252 ;
  assign n23250 = ~n514 & n6136 ;
  assign n23254 = n23253 ^ n23250 ^ 1'b0 ;
  assign n23255 = n23254 ^ n18450 ^ n7352 ;
  assign n23259 = n5606 | n10786 ;
  assign n23260 = n9770 | n23259 ;
  assign n23256 = n3498 ^ n2580 ^ 1'b0 ;
  assign n23257 = ( n5809 & n20382 ) | ( n5809 & ~n23256 ) | ( n20382 & ~n23256 ) ;
  assign n23258 = ( ~n2402 & n6960 ) | ( ~n2402 & n23257 ) | ( n6960 & n23257 ) ;
  assign n23261 = n23260 ^ n23258 ^ n6542 ;
  assign n23262 = n20601 & ~n23261 ;
  assign n23263 = n23262 ^ n508 ^ 1'b0 ;
  assign n23264 = n6234 ^ n1665 ^ 1'b0 ;
  assign n23265 = n10825 & ~n23264 ;
  assign n23266 = ~n17880 & n23265 ;
  assign n23267 = ~n385 & n23266 ;
  assign n23268 = n17404 | n20984 ;
  assign n23269 = n23268 ^ n12208 ^ 1'b0 ;
  assign n23270 = ( n1545 & ~n5305 ) | ( n1545 & n7452 ) | ( ~n5305 & n7452 ) ;
  assign n23271 = n11273 & n23270 ;
  assign n23272 = n23269 & n23271 ;
  assign n23273 = ( n871 & ~n21922 ) | ( n871 & n23272 ) | ( ~n21922 & n23272 ) ;
  assign n23274 = ( n3844 & n7306 ) | ( n3844 & n11105 ) | ( n7306 & n11105 ) ;
  assign n23275 = n22484 & n23274 ;
  assign n23276 = n22208 ^ n2927 ^ n2162 ;
  assign n23277 = n6607 & n23276 ;
  assign n23278 = n18710 ^ n9983 ^ 1'b0 ;
  assign n23279 = ~n10281 & n23278 ;
  assign n23280 = n16918 | n23279 ;
  assign n23281 = n8501 ^ n4815 ^ 1'b0 ;
  assign n23282 = n23280 & n23281 ;
  assign n23283 = n3618 | n5004 ;
  assign n23284 = n2469 ^ n2126 ^ n626 ;
  assign n23285 = ~n9780 & n23284 ;
  assign n23286 = n687 & n23285 ;
  assign n23287 = n14061 | n17159 ;
  assign n23288 = n23286 | n23287 ;
  assign n23289 = n1893 & ~n23288 ;
  assign n23290 = ( n15106 & n19412 ) | ( n15106 & ~n23289 ) | ( n19412 & ~n23289 ) ;
  assign n23291 = n8699 ^ n4932 ^ n2089 ;
  assign n23292 = n17905 ^ n10859 ^ n10432 ;
  assign n23293 = n23292 ^ n14420 ^ n5714 ;
  assign n23294 = ~n18885 & n23293 ;
  assign n23295 = ( ~n8356 & n23291 ) | ( ~n8356 & n23294 ) | ( n23291 & n23294 ) ;
  assign n23296 = n632 & ~n6856 ;
  assign n23297 = n23296 ^ n3471 ^ 1'b0 ;
  assign n23298 = ( n5352 & ~n11193 ) | ( n5352 & n23297 ) | ( ~n11193 & n23297 ) ;
  assign n23303 = ( n3247 & n11529 ) | ( n3247 & ~n13849 ) | ( n11529 & ~n13849 ) ;
  assign n23304 = n23303 ^ n7510 ^ 1'b0 ;
  assign n23302 = n3793 & ~n21146 ;
  assign n23305 = n23304 ^ n23302 ^ n16813 ;
  assign n23299 = n2943 & ~n9776 ;
  assign n23300 = n23299 ^ n6114 ^ 1'b0 ;
  assign n23301 = n23300 ^ n17678 ^ n12604 ;
  assign n23306 = n23305 ^ n23301 ^ 1'b0 ;
  assign n23307 = ( ~x186 & n3204 ) | ( ~x186 & n5944 ) | ( n3204 & n5944 ) ;
  assign n23308 = ( n8092 & ~n18132 ) | ( n8092 & n23307 ) | ( ~n18132 & n23307 ) ;
  assign n23309 = n3658 | n14029 ;
  assign n23310 = n23308 & ~n23309 ;
  assign n23311 = n5232 & ~n23310 ;
  assign n23312 = n23311 ^ n10373 ^ 1'b0 ;
  assign n23313 = ~n341 & n6319 ;
  assign n23314 = n7411 | n15328 ;
  assign n23315 = ( n21033 & n23313 ) | ( n21033 & ~n23314 ) | ( n23313 & ~n23314 ) ;
  assign n23316 = ~n2766 & n9350 ;
  assign n23317 = ( ~n5981 & n15571 ) | ( ~n5981 & n22408 ) | ( n15571 & n22408 ) ;
  assign n23318 = ~n19794 & n23317 ;
  assign n23319 = n10966 & n23318 ;
  assign n23320 = n23319 ^ n6984 ^ 1'b0 ;
  assign n23321 = ~n21008 & n23320 ;
  assign n23322 = n23321 ^ n2837 ^ 1'b0 ;
  assign n23323 = ( n23315 & n23316 ) | ( n23315 & ~n23322 ) | ( n23316 & ~n23322 ) ;
  assign n23324 = n13902 | n22010 ;
  assign n23325 = n23324 ^ n17249 ^ n5660 ;
  assign n23326 = n23325 ^ n15001 ^ 1'b0 ;
  assign n23327 = n14024 & n23326 ;
  assign n23328 = n23327 ^ n6080 ^ 1'b0 ;
  assign n23329 = n2887 | n23328 ;
  assign n23330 = n1749 | n5340 ;
  assign n23331 = n4408 & ~n23330 ;
  assign n23332 = n15120 ^ n6575 ^ n2858 ;
  assign n23333 = n23332 ^ n23239 ^ n7792 ;
  assign n23334 = n23331 | n23333 ;
  assign n23335 = n23334 ^ n19027 ^ 1'b0 ;
  assign n23336 = n8827 ^ n5495 ^ n502 ;
  assign n23337 = ( n15217 & ~n15454 ) | ( n15217 & n23336 ) | ( ~n15454 & n23336 ) ;
  assign n23339 = n4525 ^ n2261 ^ 1'b0 ;
  assign n23338 = ~n10104 & n11456 ;
  assign n23340 = n23339 ^ n23338 ^ 1'b0 ;
  assign n23341 = ( n3917 & ~n4137 ) | ( n3917 & n23340 ) | ( ~n4137 & n23340 ) ;
  assign n23342 = ( n10019 & ~n10364 ) | ( n10019 & n17313 ) | ( ~n10364 & n17313 ) ;
  assign n23343 = n4533 ^ n2352 ^ 1'b0 ;
  assign n23344 = ~n12991 & n23343 ;
  assign n23345 = ~n18998 & n23344 ;
  assign n23346 = n23345 ^ n5619 ^ 1'b0 ;
  assign n23347 = n23346 ^ n7934 ^ 1'b0 ;
  assign n23348 = n23347 ^ n6551 ^ 1'b0 ;
  assign n23349 = x26 & ~n23348 ;
  assign n23350 = n23342 & n23349 ;
  assign n23351 = n22788 ^ n20085 ^ 1'b0 ;
  assign n23352 = n16873 ^ n13886 ^ 1'b0 ;
  assign n23353 = n17594 ^ n7574 ^ n2127 ;
  assign n23354 = ( n14401 & n20067 ) | ( n14401 & n23353 ) | ( n20067 & n23353 ) ;
  assign n23355 = ( ~n8600 & n9943 ) | ( ~n8600 & n13978 ) | ( n9943 & n13978 ) ;
  assign n23356 = n1968 & n9511 ;
  assign n23357 = ( n3436 & n18576 ) | ( n3436 & n23356 ) | ( n18576 & n23356 ) ;
  assign n23358 = n23357 ^ n16664 ^ n7782 ;
  assign n23359 = ~n18268 & n23358 ;
  assign n23360 = n23355 & n23359 ;
  assign n23361 = ~n16895 & n22904 ;
  assign n23362 = n16177 ^ n10647 ^ 1'b0 ;
  assign n23363 = n23362 ^ n12106 ^ 1'b0 ;
  assign n23364 = n3504 & ~n23363 ;
  assign n23365 = ( n6284 & n13984 ) | ( n6284 & n23364 ) | ( n13984 & n23364 ) ;
  assign n23366 = ( n6006 & ~n7671 ) | ( n6006 & n16490 ) | ( ~n7671 & n16490 ) ;
  assign n23367 = ~n4658 & n14100 ;
  assign n23368 = n1930 & n23367 ;
  assign n23369 = ( n847 & n3457 ) | ( n847 & n12581 ) | ( n3457 & n12581 ) ;
  assign n23370 = n15618 ^ n7806 ^ n4917 ;
  assign n23371 = n613 | n5241 ;
  assign n23372 = n23371 ^ n10373 ^ 1'b0 ;
  assign n23373 = ( ~n2895 & n15301 ) | ( ~n2895 & n19626 ) | ( n15301 & n19626 ) ;
  assign n23374 = n2131 | n23373 ;
  assign n23375 = n23372 & ~n23374 ;
  assign n23376 = n18123 ^ n893 ^ 1'b0 ;
  assign n23377 = ( ~n9770 & n11812 ) | ( ~n9770 & n23376 ) | ( n11812 & n23376 ) ;
  assign n23378 = ( n11251 & ~n12552 ) | ( n11251 & n12772 ) | ( ~n12552 & n12772 ) ;
  assign n23379 = ( n1294 & ~n10531 ) | ( n1294 & n18991 ) | ( ~n10531 & n18991 ) ;
  assign n23380 = n3821 | n21682 ;
  assign n23381 = n9658 & n17311 ;
  assign n23382 = ( n3132 & n9206 ) | ( n3132 & n17839 ) | ( n9206 & n17839 ) ;
  assign n23383 = n23382 ^ n2532 ^ 1'b0 ;
  assign n23389 = n4358 | n14279 ;
  assign n23384 = n1822 & ~n4908 ;
  assign n23385 = n23384 ^ n8053 ^ 1'b0 ;
  assign n23386 = n23385 ^ n8360 ^ n5828 ;
  assign n23387 = n17469 ^ n8455 ^ 1'b0 ;
  assign n23388 = n23386 | n23387 ;
  assign n23390 = n23389 ^ n23388 ^ n2362 ;
  assign n23391 = n16371 ^ n8579 ^ 1'b0 ;
  assign n23392 = n23390 | n23391 ;
  assign n23393 = ( n592 & ~n11572 ) | ( n592 & n23392 ) | ( ~n11572 & n23392 ) ;
  assign n23394 = ~n639 & n8684 ;
  assign n23395 = n1856 | n13742 ;
  assign n23396 = n16543 & ~n23395 ;
  assign n23397 = n3699 & ~n14249 ;
  assign n23398 = n23397 ^ n10837 ^ n4141 ;
  assign n23399 = ( ~n16696 & n22084 ) | ( ~n16696 & n23398 ) | ( n22084 & n23398 ) ;
  assign n23400 = n11001 ^ n9431 ^ 1'b0 ;
  assign n23403 = n4185 | n15511 ;
  assign n23401 = ( n1804 & n9883 ) | ( n1804 & n12840 ) | ( n9883 & n12840 ) ;
  assign n23402 = n23401 ^ n22414 ^ 1'b0 ;
  assign n23404 = n23403 ^ n23402 ^ n11118 ;
  assign n23405 = ( n6718 & ~n9691 ) | ( n6718 & n10969 ) | ( ~n9691 & n10969 ) ;
  assign n23406 = ( n6883 & n17770 ) | ( n6883 & ~n23405 ) | ( n17770 & ~n23405 ) ;
  assign n23407 = ~n2785 & n23406 ;
  assign n23408 = n11478 ^ n11186 ^ n4010 ;
  assign n23409 = n23113 ^ x86 ^ 1'b0 ;
  assign n23410 = n13796 & n23409 ;
  assign n23411 = ( n8101 & n9160 ) | ( n8101 & ~n23410 ) | ( n9160 & ~n23410 ) ;
  assign n23412 = n23411 ^ n8673 ^ n8480 ;
  assign n23413 = ( ~n566 & n11965 ) | ( ~n566 & n23412 ) | ( n11965 & n23412 ) ;
  assign n23414 = ( n17539 & n23408 ) | ( n17539 & n23413 ) | ( n23408 & n23413 ) ;
  assign n23415 = n314 | n23414 ;
  assign n23416 = n17251 ^ n10602 ^ n7146 ;
  assign n23417 = n9605 | n23416 ;
  assign n23418 = n8160 & ~n23417 ;
  assign n23419 = n16400 ^ n10388 ^ n4596 ;
  assign n23420 = ~n1632 & n7625 ;
  assign n23421 = n5446 & ~n23420 ;
  assign n23422 = n20344 & n23421 ;
  assign n23423 = n19891 ^ n7690 ^ n6735 ;
  assign n23424 = n23423 ^ n13269 ^ n12313 ;
  assign n23425 = n3704 ^ n1979 ^ 1'b0 ;
  assign n23426 = ~n23424 & n23425 ;
  assign n23427 = n4133 | n12315 ;
  assign n23428 = n8832 ^ n7439 ^ n3934 ;
  assign n23429 = n23428 ^ n18922 ^ x94 ;
  assign n23430 = ( n9370 & n11997 ) | ( n9370 & ~n23429 ) | ( n11997 & ~n23429 ) ;
  assign n23433 = n14437 ^ n7181 ^ 1'b0 ;
  assign n23434 = n7456 | n23433 ;
  assign n23431 = n20711 ^ n14641 ^ n5338 ;
  assign n23432 = ( n3726 & n13481 ) | ( n3726 & n23431 ) | ( n13481 & n23431 ) ;
  assign n23435 = n23434 ^ n23432 ^ n15312 ;
  assign n23439 = n6181 ^ n1526 ^ n1491 ;
  assign n23440 = n23439 ^ n4478 ^ n601 ;
  assign n23441 = ( n725 & n11454 ) | ( n725 & ~n23440 ) | ( n11454 & ~n23440 ) ;
  assign n23442 = n23441 ^ n8514 ^ n6678 ;
  assign n23443 = n13496 | n23442 ;
  assign n23444 = n23443 ^ n7948 ^ 1'b0 ;
  assign n23436 = n6671 & ~n15813 ;
  assign n23437 = n23436 ^ n8949 ^ 1'b0 ;
  assign n23438 = n1407 & ~n23437 ;
  assign n23445 = n23444 ^ n23438 ^ 1'b0 ;
  assign n23446 = n14497 ^ n10091 ^ n1874 ;
  assign n23447 = n23446 ^ n21525 ^ 1'b0 ;
  assign n23448 = n1543 & n19643 ;
  assign n23449 = n23447 & n23448 ;
  assign n23450 = n4591 & ~n7750 ;
  assign n23451 = ( ~n3908 & n4638 ) | ( ~n3908 & n11158 ) | ( n4638 & n11158 ) ;
  assign n23452 = n23451 ^ n12260 ^ 1'b0 ;
  assign n23453 = ( n13905 & n23450 ) | ( n13905 & n23452 ) | ( n23450 & n23452 ) ;
  assign n23454 = n18858 ^ n7283 ^ 1'b0 ;
  assign n23455 = n3325 | n23454 ;
  assign n23456 = n23455 ^ n12420 ^ n4084 ;
  assign n23462 = n3917 ^ n3837 ^ 1'b0 ;
  assign n23463 = ~n2212 & n23462 ;
  assign n23464 = n23463 ^ n4566 ^ 1'b0 ;
  assign n23465 = n1042 & ~n23464 ;
  assign n23461 = n15426 & ~n19017 ;
  assign n23466 = n23465 ^ n23461 ^ 1'b0 ;
  assign n23460 = ( n347 & n5024 ) | ( n347 & n5417 ) | ( n5024 & n5417 ) ;
  assign n23457 = n13718 ^ n297 ^ 1'b0 ;
  assign n23458 = n12661 & n23457 ;
  assign n23459 = n5728 & n23458 ;
  assign n23467 = n23466 ^ n23460 ^ n23459 ;
  assign n23468 = n23456 & n23467 ;
  assign n23469 = ( ~n10435 & n21557 ) | ( ~n10435 & n22228 ) | ( n21557 & n22228 ) ;
  assign n23470 = n12897 ^ n492 ^ 1'b0 ;
  assign n23471 = ( ~n17987 & n23469 ) | ( ~n17987 & n23470 ) | ( n23469 & n23470 ) ;
  assign n23472 = n13728 ^ n8103 ^ 1'b0 ;
  assign n23473 = n5549 & ~n5681 ;
  assign n23474 = ~n23472 & n23473 ;
  assign n23475 = n23474 ^ n3994 ^ 1'b0 ;
  assign n23476 = n21296 ^ n8138 ^ n1714 ;
  assign n23477 = n10256 ^ n1298 ^ 1'b0 ;
  assign n23478 = ( ~n1982 & n17219 ) | ( ~n1982 & n23477 ) | ( n17219 & n23477 ) ;
  assign n23479 = n19151 | n23478 ;
  assign n23481 = n990 & ~n4277 ;
  assign n23482 = n23481 ^ n6399 ^ 1'b0 ;
  assign n23483 = n11440 ^ n8408 ^ 1'b0 ;
  assign n23484 = n23482 | n23483 ;
  assign n23480 = ~n5490 & n7566 ;
  assign n23485 = n23484 ^ n23480 ^ 1'b0 ;
  assign n23486 = ( n5720 & n14227 ) | ( n5720 & ~n15535 ) | ( n14227 & ~n15535 ) ;
  assign n23487 = n2996 ^ n2272 ^ 1'b0 ;
  assign n23488 = n3368 | n23487 ;
  assign n23489 = n6330 & ~n23488 ;
  assign n23490 = n23489 ^ n20344 ^ 1'b0 ;
  assign n23491 = ( ~n9801 & n23486 ) | ( ~n9801 & n23490 ) | ( n23486 & n23490 ) ;
  assign n23492 = ( n1831 & n10701 ) | ( n1831 & ~n11378 ) | ( n10701 & ~n11378 ) ;
  assign n23493 = n23492 ^ n6973 ^ 1'b0 ;
  assign n23494 = n8538 | n23493 ;
  assign n23497 = n3781 & n18473 ;
  assign n23498 = n23497 ^ n7350 ^ 1'b0 ;
  assign n23495 = n1062 ^ n1030 ^ 1'b0 ;
  assign n23496 = n16374 | n23495 ;
  assign n23499 = n23498 ^ n23496 ^ 1'b0 ;
  assign n23500 = n1865 & n6698 ;
  assign n23501 = n23500 ^ n4479 ^ 1'b0 ;
  assign n23502 = n16776 ^ n1414 ^ 1'b0 ;
  assign n23503 = n23501 & ~n23502 ;
  assign n23504 = n23503 ^ n3764 ^ 1'b0 ;
  assign n23505 = n2851 & ~n23504 ;
  assign n23506 = n23505 ^ n11066 ^ 1'b0 ;
  assign n23507 = n4204 ^ n2715 ^ 1'b0 ;
  assign n23508 = n14227 & ~n23507 ;
  assign n23509 = n2943 ^ n776 ^ 1'b0 ;
  assign n23510 = ~n20741 & n23509 ;
  assign n23511 = n23510 ^ n1702 ^ 1'b0 ;
  assign n23512 = n23508 & n23511 ;
  assign n23513 = ~n16567 & n23512 ;
  assign n23514 = ( n2311 & ~n6449 ) | ( n2311 & n14153 ) | ( ~n6449 & n14153 ) ;
  assign n23515 = n12341 & n23514 ;
  assign n23520 = n11579 ^ n3941 ^ n1249 ;
  assign n23516 = n2117 & n20106 ;
  assign n23517 = ( ~n4100 & n13406 ) | ( ~n4100 & n13499 ) | ( n13406 & n13499 ) ;
  assign n23518 = n23517 ^ n19777 ^ n17427 ;
  assign n23519 = n23516 | n23518 ;
  assign n23521 = n23520 ^ n23519 ^ 1'b0 ;
  assign n23522 = n23521 ^ n1526 ^ n458 ;
  assign n23523 = n14619 & n21917 ;
  assign n23524 = ~n7677 & n23523 ;
  assign n23525 = n19832 | n23524 ;
  assign n23526 = n13981 & ~n23525 ;
  assign n23527 = n23526 ^ n2426 ^ n1161 ;
  assign n23528 = ( n7167 & n8957 ) | ( n7167 & n14387 ) | ( n8957 & n14387 ) ;
  assign n23529 = ~n14086 & n23528 ;
  assign n23530 = ~n16927 & n23529 ;
  assign n23531 = n23530 ^ n22513 ^ n14874 ;
  assign n23532 = n20136 ^ n18537 ^ 1'b0 ;
  assign n23535 = ( ~n7579 & n8988 ) | ( ~n7579 & n12230 ) | ( n8988 & n12230 ) ;
  assign n23536 = n23535 ^ n2724 ^ 1'b0 ;
  assign n23533 = ~n18560 & n20818 ;
  assign n23534 = n23533 ^ n14874 ^ 1'b0 ;
  assign n23537 = n23536 ^ n23534 ^ 1'b0 ;
  assign n23538 = ( ~n2558 & n7263 ) | ( ~n2558 & n16472 ) | ( n7263 & n16472 ) ;
  assign n23539 = n23538 ^ n22451 ^ n9066 ;
  assign n23540 = n9757 ^ n1326 ^ 1'b0 ;
  assign n23541 = n23540 ^ n17602 ^ 1'b0 ;
  assign n23542 = n18374 & n23541 ;
  assign n23544 = n14468 ^ n10865 ^ 1'b0 ;
  assign n23545 = n23544 ^ n23373 ^ n14396 ;
  assign n23543 = n14849 | n15526 ;
  assign n23546 = n23545 ^ n23543 ^ 1'b0 ;
  assign n23547 = n12874 ^ n1144 ^ 1'b0 ;
  assign n23548 = n13810 ^ n393 ^ 1'b0 ;
  assign n23549 = n679 | n23548 ;
  assign n23550 = n6468 & ~n23549 ;
  assign n23551 = ~n11617 & n23550 ;
  assign n23552 = n18640 & ~n23551 ;
  assign n23553 = ~n655 & n23552 ;
  assign n23554 = n19378 & n23553 ;
  assign n23555 = n16095 ^ n4358 ^ 1'b0 ;
  assign n23556 = n3313 ^ n674 ^ 1'b0 ;
  assign n23557 = n7479 & ~n23556 ;
  assign n23558 = n23557 ^ n14656 ^ 1'b0 ;
  assign n23559 = n1431 & ~n23558 ;
  assign n23560 = n2657 & n22886 ;
  assign n23561 = n19128 ^ n8318 ^ 1'b0 ;
  assign n23562 = n315 | n23561 ;
  assign n23563 = n1326 & n6567 ;
  assign n23564 = n23563 ^ n11527 ^ 1'b0 ;
  assign n23565 = n23564 ^ n3625 ^ n3446 ;
  assign n23566 = n3977 & n7419 ;
  assign n23567 = n17368 ^ n2416 ^ 1'b0 ;
  assign n23568 = ( n16391 & ~n16441 ) | ( n16391 & n23567 ) | ( ~n16441 & n23567 ) ;
  assign n23569 = n6307 & n10830 ;
  assign n23570 = n23569 ^ n12442 ^ 1'b0 ;
  assign n23571 = n23570 ^ n10128 ^ 1'b0 ;
  assign n23572 = n573 & ~n17087 ;
  assign n23573 = n1091 & n3689 ;
  assign n23574 = ( x156 & n11001 ) | ( x156 & ~n18686 ) | ( n11001 & ~n18686 ) ;
  assign n23575 = ( n1572 & n13195 ) | ( n1572 & n23574 ) | ( n13195 & n23574 ) ;
  assign n23576 = ( n12412 & n14620 ) | ( n12412 & n23575 ) | ( n14620 & n23575 ) ;
  assign n23577 = ( ~n4340 & n6989 ) | ( ~n4340 & n15560 ) | ( n6989 & n15560 ) ;
  assign n23578 = n2086 & ~n23577 ;
  assign n23579 = ( n2460 & n20364 ) | ( n2460 & ~n23578 ) | ( n20364 & ~n23578 ) ;
  assign n23580 = n23579 ^ n5885 ^ 1'b0 ;
  assign n23581 = n23576 | n23580 ;
  assign n23582 = n7487 ^ n4477 ^ 1'b0 ;
  assign n23583 = ~n3557 & n23582 ;
  assign n23584 = n23583 ^ n21200 ^ n10492 ;
  assign n23587 = ( n5431 & n9932 ) | ( n5431 & ~n11901 ) | ( n9932 & ~n11901 ) ;
  assign n23585 = n4178 & ~n6512 ;
  assign n23586 = n10849 & n23585 ;
  assign n23588 = n23587 ^ n23586 ^ n20911 ;
  assign n23589 = ( n6168 & ~n6332 ) | ( n6168 & n23588 ) | ( ~n6332 & n23588 ) ;
  assign n23590 = n920 | n4451 ;
  assign n23591 = n23589 & ~n23590 ;
  assign n23592 = n23591 ^ n16684 ^ n4846 ;
  assign n23593 = ( n730 & n6198 ) | ( n730 & n14040 ) | ( n6198 & n14040 ) ;
  assign n23594 = n23593 ^ n17285 ^ n5164 ;
  assign n23595 = ~n8170 & n21096 ;
  assign n23596 = n23594 & n23595 ;
  assign n23597 = n8991 ^ n6661 ^ 1'b0 ;
  assign n23598 = n11376 ^ n10826 ^ n4017 ;
  assign n23599 = ( n4469 & n8278 ) | ( n4469 & ~n13141 ) | ( n8278 & ~n13141 ) ;
  assign n23600 = n23599 ^ n15276 ^ n1291 ;
  assign n23601 = n23598 & ~n23600 ;
  assign n23602 = ~n10886 & n23601 ;
  assign n23603 = n9769 & n14385 ;
  assign n23604 = ~n6911 & n23603 ;
  assign n23605 = n9728 ^ n712 ^ 1'b0 ;
  assign n23606 = ( ~n8911 & n23604 ) | ( ~n8911 & n23605 ) | ( n23604 & n23605 ) ;
  assign n23607 = n6598 | n16632 ;
  assign n23608 = n17526 | n23607 ;
  assign n23609 = n14221 ^ n9197 ^ n6347 ;
  assign n23610 = n2070 & n2623 ;
  assign n23611 = n23610 ^ n2083 ^ 1'b0 ;
  assign n23612 = ( n8509 & ~n13241 ) | ( n8509 & n23611 ) | ( ~n13241 & n23611 ) ;
  assign n23613 = ( n23608 & ~n23609 ) | ( n23608 & n23612 ) | ( ~n23609 & n23612 ) ;
  assign n23616 = n1714 ^ x22 ^ 1'b0 ;
  assign n23617 = n16662 | n23616 ;
  assign n23614 = n6174 ^ n3833 ^ n2641 ;
  assign n23615 = ( n1355 & n4407 ) | ( n1355 & ~n23614 ) | ( n4407 & ~n23614 ) ;
  assign n23618 = n23617 ^ n23615 ^ n18080 ;
  assign n23619 = ( ~n3942 & n18744 ) | ( ~n3942 & n23355 ) | ( n18744 & n23355 ) ;
  assign n23620 = n4651 & ~n6282 ;
  assign n23621 = ( n1155 & n8236 ) | ( n1155 & ~n23620 ) | ( n8236 & ~n23620 ) ;
  assign n23622 = n13123 ^ n10404 ^ 1'b0 ;
  assign n23623 = n23622 ^ n4199 ^ n4007 ;
  assign n23624 = n7631 ^ n6059 ^ 1'b0 ;
  assign n23625 = ~n4346 & n23624 ;
  assign n23627 = n4599 ^ n4113 ^ n2110 ;
  assign n23628 = n23627 ^ n6367 ^ n2501 ;
  assign n23626 = n1111 | n3763 ;
  assign n23629 = n23628 ^ n23626 ^ 1'b0 ;
  assign n23630 = n15121 ^ n14085 ^ n2992 ;
  assign n23631 = n9023 & n23630 ;
  assign n23632 = n2024 & n23631 ;
  assign n23633 = ( n3210 & n21327 ) | ( n3210 & n23632 ) | ( n21327 & n23632 ) ;
  assign n23634 = n23633 ^ n2627 ^ 1'b0 ;
  assign n23635 = n3914 | n13087 ;
  assign n23636 = n2696 | n5697 ;
  assign n23637 = n23636 ^ n9063 ^ n4138 ;
  assign n23638 = ( n6848 & n11560 ) | ( n6848 & ~n23637 ) | ( n11560 & ~n23637 ) ;
  assign n23639 = n23638 ^ n19530 ^ n19346 ;
  assign n23640 = n14291 & n16307 ;
  assign n23641 = n12007 ^ n4873 ^ 1'b0 ;
  assign n23642 = n445 & ~n23641 ;
  assign n23643 = n18078 & ~n23642 ;
  assign n23644 = n11579 ^ n9669 ^ 1'b0 ;
  assign n23645 = ( n7504 & n8593 ) | ( n7504 & n23644 ) | ( n8593 & n23644 ) ;
  assign n23646 = n8354 ^ n2407 ^ n2327 ;
  assign n23647 = n9502 | n14523 ;
  assign n23648 = ( n9900 & ~n15465 ) | ( n9900 & n23647 ) | ( ~n15465 & n23647 ) ;
  assign n23650 = n4431 ^ n4373 ^ 1'b0 ;
  assign n23649 = ( ~n2606 & n5606 ) | ( ~n2606 & n9544 ) | ( n5606 & n9544 ) ;
  assign n23651 = n23650 ^ n23649 ^ n7924 ;
  assign n23652 = n19209 & n23651 ;
  assign n23653 = n12261 ^ n2442 ^ 1'b0 ;
  assign n23654 = n23653 ^ n8363 ^ 1'b0 ;
  assign n23655 = ~n23277 & n23654 ;
  assign n23656 = n8987 & n12888 ;
  assign n23657 = n23656 ^ n3375 ^ 1'b0 ;
  assign n23658 = n5350 & n23657 ;
  assign n23659 = n19577 ^ n13321 ^ n10155 ;
  assign n23660 = ( n4087 & ~n6887 ) | ( n4087 & n8878 ) | ( ~n6887 & n8878 ) ;
  assign n23661 = ( n11627 & n16458 ) | ( n11627 & n23660 ) | ( n16458 & n23660 ) ;
  assign n23662 = n22084 ^ n11855 ^ n9972 ;
  assign n23663 = n1760 & n14572 ;
  assign n23664 = n23663 ^ n2238 ^ 1'b0 ;
  assign n23665 = n14418 ^ n9489 ^ 1'b0 ;
  assign n23666 = n1390 & n23665 ;
  assign n23667 = ( n687 & ~n12714 ) | ( n687 & n23666 ) | ( ~n12714 & n23666 ) ;
  assign n23668 = n5281 ^ n5224 ^ n3516 ;
  assign n23669 = n23668 ^ n23020 ^ 1'b0 ;
  assign n23670 = n23669 ^ n10641 ^ n813 ;
  assign n23671 = n5739 ^ n5708 ^ n933 ;
  assign n23672 = ( n2273 & n7590 ) | ( n2273 & ~n23671 ) | ( n7590 & ~n23671 ) ;
  assign n23673 = n2943 & ~n14455 ;
  assign n23674 = n23673 ^ n12605 ^ 1'b0 ;
  assign n23681 = ( ~n2722 & n6575 ) | ( ~n2722 & n12621 ) | ( n6575 & n12621 ) ;
  assign n23675 = n8002 ^ n7884 ^ n3448 ;
  assign n23677 = n5008 ^ n4746 ^ n2999 ;
  assign n23676 = n2006 & n2749 ;
  assign n23678 = n23677 ^ n23676 ^ 1'b0 ;
  assign n23679 = n11774 & n23678 ;
  assign n23680 = ~n23675 & n23679 ;
  assign n23682 = n23681 ^ n23680 ^ 1'b0 ;
  assign n23683 = n8594 | n23682 ;
  assign n23684 = ( ~n8117 & n19901 ) | ( ~n8117 & n23683 ) | ( n19901 & n23683 ) ;
  assign n23689 = n8196 ^ n3983 ^ 1'b0 ;
  assign n23690 = n18297 & n23689 ;
  assign n23691 = ~n16151 & n23690 ;
  assign n23692 = n3357 & n23691 ;
  assign n23693 = ~n6815 & n16898 ;
  assign n23694 = n23692 & n23693 ;
  assign n23685 = n11092 ^ n1396 ^ 1'b0 ;
  assign n23686 = n16936 | n23685 ;
  assign n23687 = n6678 & ~n23686 ;
  assign n23688 = n23687 ^ n17606 ^ 1'b0 ;
  assign n23695 = n23694 ^ n23688 ^ 1'b0 ;
  assign n23696 = x91 & ~n11698 ;
  assign n23697 = n23696 ^ n1797 ^ 1'b0 ;
  assign n23698 = n23697 ^ n16276 ^ n15139 ;
  assign n23699 = n14739 ^ n8112 ^ 1'b0 ;
  assign n23701 = n22152 ^ n6893 ^ 1'b0 ;
  assign n23702 = n1659 & ~n23701 ;
  assign n23700 = n946 & ~n18753 ;
  assign n23703 = n23702 ^ n23700 ^ 1'b0 ;
  assign n23704 = ~n10473 & n19348 ;
  assign n23705 = n18934 & n23704 ;
  assign n23706 = n23705 ^ n12162 ^ 1'b0 ;
  assign n23707 = n14917 & ~n23706 ;
  assign n23708 = n1446 | n15498 ;
  assign n23709 = n4307 | n23708 ;
  assign n23710 = n23709 ^ n11492 ^ n6879 ;
  assign n23711 = ( n7705 & n15109 ) | ( n7705 & n15945 ) | ( n15109 & n15945 ) ;
  assign n23712 = n18074 ^ n1955 ^ 1'b0 ;
  assign n23713 = n23711 & ~n23712 ;
  assign n23716 = n3516 ^ n2867 ^ 1'b0 ;
  assign n23714 = n8333 ^ n2864 ^ n264 ;
  assign n23715 = ~n19746 & n23714 ;
  assign n23717 = n23716 ^ n23715 ^ n4612 ;
  assign n23718 = ~n4288 & n7940 ;
  assign n23724 = n22272 ^ n6275 ^ 1'b0 ;
  assign n23725 = ~n2944 & n23724 ;
  assign n23726 = n23725 ^ n16789 ^ 1'b0 ;
  assign n23719 = ~n4398 & n8222 ;
  assign n23720 = n19434 ^ n4732 ^ n3287 ;
  assign n23721 = n23719 | n23720 ;
  assign n23722 = n23721 ^ n20058 ^ 1'b0 ;
  assign n23723 = n6368 | n23722 ;
  assign n23727 = n23726 ^ n23723 ^ 1'b0 ;
  assign n23728 = ( x79 & n1440 ) | ( x79 & n12388 ) | ( n1440 & n12388 ) ;
  assign n23729 = n23728 ^ n14489 ^ n2337 ;
  assign n23730 = n7553 ^ n7213 ^ 1'b0 ;
  assign n23731 = ( n15738 & n23729 ) | ( n15738 & n23730 ) | ( n23729 & n23730 ) ;
  assign n23732 = n13385 ^ n4779 ^ n2705 ;
  assign n23733 = ( ~n4807 & n15552 ) | ( ~n4807 & n23732 ) | ( n15552 & n23732 ) ;
  assign n23734 = ( ~n2722 & n9469 ) | ( ~n2722 & n23733 ) | ( n9469 & n23733 ) ;
  assign n23735 = n3335 | n11077 ;
  assign n23736 = n8243 ^ n8059 ^ n2563 ;
  assign n23737 = n23736 ^ n13496 ^ 1'b0 ;
  assign n23738 = n12321 & n23737 ;
  assign n23739 = ~n23735 & n23738 ;
  assign n23740 = n23156 ^ n3201 ^ 1'b0 ;
  assign n23741 = n1430 ^ n324 ^ 1'b0 ;
  assign n23742 = n8393 | n23741 ;
  assign n23743 = n19838 & ~n23742 ;
  assign n23744 = ~n1093 & n23743 ;
  assign n23745 = n23744 ^ n11994 ^ n1201 ;
  assign n23746 = x86 & ~n18334 ;
  assign n23747 = n23746 ^ n20673 ^ 1'b0 ;
  assign n23748 = n12032 & n23747 ;
  assign n23749 = ( n10677 & n12520 ) | ( n10677 & ~n23748 ) | ( n12520 & ~n23748 ) ;
  assign n23750 = n10216 & n21980 ;
  assign n23751 = n23750 ^ n1975 ^ 1'b0 ;
  assign n23752 = n23640 | n23751 ;
  assign n23753 = n9204 & ~n23026 ;
  assign n23754 = n8045 & n11473 ;
  assign n23755 = ~n7390 & n23754 ;
  assign n23756 = n23755 ^ n4705 ^ 1'b0 ;
  assign n23757 = n13972 ^ n6731 ^ 1'b0 ;
  assign n23758 = n6017 & ~n23757 ;
  assign n23759 = n23758 ^ n10222 ^ 1'b0 ;
  assign n23760 = n5321 & n23759 ;
  assign n23761 = n23115 ^ n6765 ^ 1'b0 ;
  assign n23762 = n23760 & ~n23761 ;
  assign n23763 = n2904 & n3223 ;
  assign n23764 = ( ~n1700 & n10930 ) | ( ~n1700 & n23763 ) | ( n10930 & n23763 ) ;
  assign n23765 = n17264 ^ n9310 ^ 1'b0 ;
  assign n23766 = n18504 & ~n23765 ;
  assign n23767 = n23766 ^ n15827 ^ n13648 ;
  assign n23768 = ~n11905 & n23767 ;
  assign n23769 = n6050 & n23768 ;
  assign n23770 = n15586 ^ n13387 ^ n8848 ;
  assign n23771 = n18933 | n23770 ;
  assign n23772 = n18442 ^ n6468 ^ 1'b0 ;
  assign n23773 = n1015 | n12145 ;
  assign n23774 = ( ~n2954 & n23463 ) | ( ~n2954 & n23773 ) | ( n23463 & n23773 ) ;
  assign n23775 = ~n23772 & n23774 ;
  assign n23776 = ~n11055 & n23775 ;
  assign n23777 = n13544 ^ n6266 ^ 1'b0 ;
  assign n23778 = x213 & ~n23777 ;
  assign n23779 = n13120 | n23192 ;
  assign n23780 = n23779 ^ n6007 ^ 1'b0 ;
  assign n23781 = n13027 ^ n11727 ^ 1'b0 ;
  assign n23782 = ( n11506 & ~n14577 ) | ( n11506 & n23781 ) | ( ~n14577 & n23781 ) ;
  assign n23783 = n9662 ^ n3838 ^ 1'b0 ;
  assign n23784 = ( ~n12912 & n22034 ) | ( ~n12912 & n23783 ) | ( n22034 & n23783 ) ;
  assign n23785 = n23784 ^ n21954 ^ n4804 ;
  assign n23786 = n21616 ^ n1485 ^ 1'b0 ;
  assign n23787 = n19542 ^ n1346 ^ 1'b0 ;
  assign n23788 = n6720 & ~n11666 ;
  assign n23789 = n22693 ^ n21078 ^ n15339 ;
  assign n23790 = n1686 & ~n15301 ;
  assign n23791 = n23790 ^ n18627 ^ 1'b0 ;
  assign n23792 = n23791 ^ n7860 ^ n2634 ;
  assign n23793 = n23792 ^ n12162 ^ n9919 ;
  assign n23794 = n23793 ^ n9625 ^ n1203 ;
  assign n23795 = ( n1901 & n12233 ) | ( n1901 & ~n18588 ) | ( n12233 & ~n18588 ) ;
  assign n23797 = n8984 ^ n2899 ^ 1'b0 ;
  assign n23798 = n23797 ^ n1530 ^ n1474 ;
  assign n23796 = n13492 ^ n7616 ^ n7217 ;
  assign n23799 = n23798 ^ n23796 ^ n8568 ;
  assign n23800 = n23799 ^ n9269 ^ 1'b0 ;
  assign n23801 = n12145 & n14067 ;
  assign n23802 = n16245 ^ n13360 ^ 1'b0 ;
  assign n23803 = ( n4080 & n14861 ) | ( n4080 & n23802 ) | ( n14861 & n23802 ) ;
  assign n23804 = n22620 ^ n13587 ^ 1'b0 ;
  assign n23805 = n23804 ^ n15655 ^ n8617 ;
  assign n23806 = ( ~n22377 & n23590 ) | ( ~n22377 & n23805 ) | ( n23590 & n23805 ) ;
  assign n23807 = n8792 ^ n3941 ^ 1'b0 ;
  assign n23808 = n3692 & ~n23807 ;
  assign n23809 = n1897 | n21151 ;
  assign n23810 = ~n962 & n7410 ;
  assign n23811 = n23810 ^ n19347 ^ 1'b0 ;
  assign n23812 = n17224 & ~n23811 ;
  assign n23813 = ~n21538 & n23812 ;
  assign n23814 = ( n23808 & ~n23809 ) | ( n23808 & n23813 ) | ( ~n23809 & n23813 ) ;
  assign n23815 = n11366 ^ n5387 ^ n5015 ;
  assign n23816 = n5711 & ~n23815 ;
  assign n23817 = n23816 ^ n7223 ^ 1'b0 ;
  assign n23818 = n4794 & ~n6033 ;
  assign n23819 = n23818 ^ n16410 ^ 1'b0 ;
  assign n23820 = n10065 & n23819 ;
  assign n23822 = n1416 & ~n4339 ;
  assign n23823 = n6056 & n23822 ;
  assign n23824 = ~n11994 & n15950 ;
  assign n23825 = ( ~n12359 & n23823 ) | ( ~n12359 & n23824 ) | ( n23823 & n23824 ) ;
  assign n23827 = ( ~n436 & n3452 ) | ( ~n436 & n4764 ) | ( n3452 & n4764 ) ;
  assign n23826 = n23501 ^ n8774 ^ n6285 ;
  assign n23828 = n23827 ^ n23826 ^ n16985 ;
  assign n23829 = ( n10834 & n23825 ) | ( n10834 & ~n23828 ) | ( n23825 & ~n23828 ) ;
  assign n23821 = n7672 | n17928 ;
  assign n23830 = n23829 ^ n23821 ^ 1'b0 ;
  assign n23831 = ( ~n12813 & n13229 ) | ( ~n12813 & n21093 ) | ( n13229 & n21093 ) ;
  assign n23832 = n18655 ^ n16770 ^ n2187 ;
  assign n23833 = n19892 ^ n16762 ^ 1'b0 ;
  assign n23834 = n11198 & ~n23833 ;
  assign n23835 = n23834 ^ n6267 ^ 1'b0 ;
  assign n23836 = ( ~n1177 & n6847 ) | ( ~n1177 & n21254 ) | ( n6847 & n21254 ) ;
  assign n23837 = n23836 ^ n6797 ^ 1'b0 ;
  assign n23838 = n4229 & n7992 ;
  assign n23839 = n8607 ^ n7389 ^ n1833 ;
  assign n23840 = n23839 ^ n13742 ^ 1'b0 ;
  assign n23841 = n15531 ^ n1472 ^ n654 ;
  assign n23842 = ( n1184 & n2464 ) | ( n1184 & n23841 ) | ( n2464 & n23841 ) ;
  assign n23843 = ( n8942 & ~n13581 ) | ( n8942 & n23842 ) | ( ~n13581 & n23842 ) ;
  assign n23844 = n11429 ^ n5183 ^ 1'b0 ;
  assign n23845 = ( n6091 & n23843 ) | ( n6091 & ~n23844 ) | ( n23843 & ~n23844 ) ;
  assign n23846 = n7233 | n20531 ;
  assign n23847 = n17266 ^ n2947 ^ 1'b0 ;
  assign n23848 = ~n6523 & n23847 ;
  assign n23849 = n23848 ^ n22988 ^ n7404 ;
  assign n23850 = n425 & ~n23849 ;
  assign n23851 = n12589 & n23850 ;
  assign n23853 = ~n6881 & n8109 ;
  assign n23854 = n23853 ^ x97 ^ 1'b0 ;
  assign n23852 = ( n982 & n5835 ) | ( n982 & n9096 ) | ( n5835 & n9096 ) ;
  assign n23855 = n23854 ^ n23852 ^ 1'b0 ;
  assign n23856 = n4971 ^ n3592 ^ n3452 ;
  assign n23857 = n8545 | n18243 ;
  assign n23858 = n23856 & ~n23857 ;
  assign n23859 = n23855 & ~n23858 ;
  assign n23860 = n13634 ^ n11038 ^ n7605 ;
  assign n23861 = ~n10922 & n17546 ;
  assign n23862 = n5542 & n12046 ;
  assign n23863 = ~n23861 & n23862 ;
  assign n23864 = n23863 ^ n8826 ^ n1797 ;
  assign n23865 = n18653 ^ n14485 ^ n8771 ;
  assign n23873 = ( x68 & ~n2976 ) | ( x68 & n9627 ) | ( ~n2976 & n9627 ) ;
  assign n23866 = n12595 ^ n7746 ^ 1'b0 ;
  assign n23867 = n11772 | n23866 ;
  assign n23868 = ( n831 & n14300 ) | ( n831 & ~n17826 ) | ( n14300 & ~n17826 ) ;
  assign n23869 = n6682 ^ n5517 ^ 1'b0 ;
  assign n23870 = n23869 ^ n7850 ^ 1'b0 ;
  assign n23871 = n23868 & ~n23870 ;
  assign n23872 = ( ~n17900 & n23867 ) | ( ~n17900 & n23871 ) | ( n23867 & n23871 ) ;
  assign n23874 = n23873 ^ n23872 ^ n9096 ;
  assign n23875 = n21737 ^ n6913 ^ n6023 ;
  assign n23876 = n23875 ^ n14497 ^ 1'b0 ;
  assign n23877 = ~n23874 & n23876 ;
  assign n23878 = n9515 | n16552 ;
  assign n23879 = n15170 | n23878 ;
  assign n23880 = n5177 | n13345 ;
  assign n23881 = ~n4399 & n11536 ;
  assign n23882 = n23881 ^ n3039 ^ 1'b0 ;
  assign n23883 = ( n6189 & n21387 ) | ( n6189 & n23564 ) | ( n21387 & n23564 ) ;
  assign n23884 = n949 | n23883 ;
  assign n23885 = n23884 ^ n2503 ^ 1'b0 ;
  assign n23886 = ( n21442 & n23882 ) | ( n21442 & n23885 ) | ( n23882 & n23885 ) ;
  assign n23887 = n23886 ^ n14007 ^ n11105 ;
  assign n23892 = n15494 ^ n3130 ^ n508 ;
  assign n23891 = n7363 & n10229 ;
  assign n23893 = n23892 ^ n23891 ^ 1'b0 ;
  assign n23894 = ~n16587 & n23893 ;
  assign n23888 = x56 & ~n16237 ;
  assign n23889 = ~n21439 & n23510 ;
  assign n23890 = n23888 & n23889 ;
  assign n23895 = n23894 ^ n23890 ^ 1'b0 ;
  assign n23896 = n4332 & n4580 ;
  assign n23897 = n23896 ^ n23401 ^ n14337 ;
  assign n23898 = n23897 ^ n11074 ^ 1'b0 ;
  assign n23899 = ( x75 & n4015 ) | ( x75 & n21342 ) | ( n4015 & n21342 ) ;
  assign n23900 = n23899 ^ n20748 ^ 1'b0 ;
  assign n23901 = n22687 ^ n10439 ^ n2739 ;
  assign n23902 = n23446 ^ n5426 ^ 1'b0 ;
  assign n23903 = ~n4460 & n7759 ;
  assign n23904 = n23903 ^ n8978 ^ 1'b0 ;
  assign n23905 = n23904 ^ n18883 ^ n642 ;
  assign n23906 = n11402 ^ n6275 ^ 1'b0 ;
  assign n23907 = n3294 & ~n6200 ;
  assign n23908 = n23907 ^ n21872 ^ 1'b0 ;
  assign n23909 = n6657 | n23908 ;
  assign n23910 = ( n1314 & n18374 ) | ( n1314 & n23909 ) | ( n18374 & n23909 ) ;
  assign n23911 = n23906 & n23910 ;
  assign n23912 = n23911 ^ n14156 ^ 1'b0 ;
  assign n23913 = n23912 ^ n22108 ^ n11091 ;
  assign n23914 = n6561 ^ n1160 ^ 1'b0 ;
  assign n23915 = n23405 | n23914 ;
  assign n23920 = n894 & ~n4732 ;
  assign n23921 = n8231 & n23920 ;
  assign n23922 = ( n3763 & n11000 ) | ( n3763 & ~n11992 ) | ( n11000 & ~n11992 ) ;
  assign n23923 = ( n20246 & n23921 ) | ( n20246 & n23922 ) | ( n23921 & n23922 ) ;
  assign n23917 = n3409 & ~n19502 ;
  assign n23918 = n23917 ^ n10349 ^ 1'b0 ;
  assign n23916 = ( ~n483 & n796 ) | ( ~n483 & n1304 ) | ( n796 & n1304 ) ;
  assign n23919 = n23918 ^ n23916 ^ n4725 ;
  assign n23924 = n23923 ^ n23919 ^ n1544 ;
  assign n23926 = ( n7195 & n7453 ) | ( n7195 & n11316 ) | ( n7453 & n11316 ) ;
  assign n23925 = ( x105 & n576 ) | ( x105 & n7411 ) | ( n576 & n7411 ) ;
  assign n23927 = n23926 ^ n23925 ^ n10258 ;
  assign n23928 = n9312 ^ n1281 ^ 1'b0 ;
  assign n23929 = ( n7128 & n23818 ) | ( n7128 & n23928 ) | ( n23818 & n23928 ) ;
  assign n23930 = n19178 ^ n12633 ^ 1'b0 ;
  assign n23931 = ( ~n2247 & n23929 ) | ( ~n2247 & n23930 ) | ( n23929 & n23930 ) ;
  assign n23932 = n7407 | n11841 ;
  assign n23933 = n13926 | n23932 ;
  assign n23934 = n23933 ^ n4818 ^ 1'b0 ;
  assign n23935 = n5373 & n16581 ;
  assign n23936 = n23935 ^ n14452 ^ 1'b0 ;
  assign n23937 = n18090 & ~n23466 ;
  assign n23938 = ( n6488 & ~n9785 ) | ( n6488 & n12808 ) | ( ~n9785 & n12808 ) ;
  assign n23939 = n23938 ^ n9530 ^ 1'b0 ;
  assign n23940 = n20688 ^ n20434 ^ n5609 ;
  assign n23941 = ~n8150 & n23117 ;
  assign n23942 = ~n13709 & n23941 ;
  assign n23943 = n20423 ^ n11759 ^ 1'b0 ;
  assign n23944 = n12411 | n23943 ;
  assign n23951 = ( ~x46 & n6634 ) | ( ~x46 & n9187 ) | ( n6634 & n9187 ) ;
  assign n23948 = n8843 & n21840 ;
  assign n23949 = n21907 ^ n5129 ^ 1'b0 ;
  assign n23950 = n23948 | n23949 ;
  assign n23945 = ( ~n3348 & n8438 ) | ( ~n3348 & n9509 ) | ( n8438 & n9509 ) ;
  assign n23946 = n12328 & n23945 ;
  assign n23947 = ( n3633 & ~n23594 ) | ( n3633 & n23946 ) | ( ~n23594 & n23946 ) ;
  assign n23952 = n23951 ^ n23950 ^ n23947 ;
  assign n23953 = n6676 & ~n8260 ;
  assign n23954 = ( n6832 & n11467 ) | ( n6832 & ~n23953 ) | ( n11467 & ~n23953 ) ;
  assign n23962 = n326 & ~n13915 ;
  assign n23961 = n19341 ^ n17122 ^ 1'b0 ;
  assign n23958 = n894 & n18690 ;
  assign n23959 = ~n11730 & n23958 ;
  assign n23960 = ~n22944 & n23959 ;
  assign n23963 = n23962 ^ n23961 ^ n23960 ;
  assign n23955 = n15829 ^ n11406 ^ n1994 ;
  assign n23956 = n15349 & n23955 ;
  assign n23957 = n9437 & ~n23956 ;
  assign n23964 = n23963 ^ n23957 ^ 1'b0 ;
  assign n23965 = ( n936 & n2875 ) | ( n936 & n6608 ) | ( n2875 & n6608 ) ;
  assign n23966 = n17891 ^ n16532 ^ n6604 ;
  assign n23967 = n23966 ^ n10911 ^ n8723 ;
  assign n23968 = n23967 ^ n15323 ^ n640 ;
  assign n23969 = n5523 & n9685 ;
  assign n23970 = n1639 & n23969 ;
  assign n23971 = n11677 ^ n7127 ^ 1'b0 ;
  assign n23972 = ~n2017 & n23971 ;
  assign n23973 = ~n3703 & n23972 ;
  assign n23974 = n23973 ^ n7814 ^ 1'b0 ;
  assign n23975 = n12938 & ~n15234 ;
  assign n23976 = n23975 ^ n4789 ^ 1'b0 ;
  assign n23977 = ( n16024 & n22297 ) | ( n16024 & n23976 ) | ( n22297 & n23976 ) ;
  assign n23978 = ( n1054 & n7758 ) | ( n1054 & ~n15162 ) | ( n7758 & ~n15162 ) ;
  assign n23979 = ( n13019 & ~n15868 ) | ( n13019 & n23978 ) | ( ~n15868 & n23978 ) ;
  assign n23980 = ~n10593 & n11452 ;
  assign n23981 = ~n23979 & n23980 ;
  assign n23982 = ~n4618 & n6044 ;
  assign n23983 = n23981 & n23982 ;
  assign n23984 = ~n6551 & n15696 ;
  assign n23985 = n23984 ^ n1270 ^ 1'b0 ;
  assign n23986 = n17528 ^ n910 ^ 1'b0 ;
  assign n23987 = ~n384 & n23986 ;
  assign n23988 = n23987 ^ n20243 ^ n733 ;
  assign n23989 = n12288 ^ n5352 ^ 1'b0 ;
  assign n23990 = x54 & n23989 ;
  assign n23991 = x91 & ~n23990 ;
  assign n23992 = ~n8493 & n13288 ;
  assign n23993 = n23992 ^ n18013 ^ 1'b0 ;
  assign n23994 = n17732 ^ n8937 ^ n5773 ;
  assign n23995 = n9010 & n23994 ;
  assign n23996 = n23993 & ~n23995 ;
  assign n23997 = n13986 ^ n6880 ^ n1200 ;
  assign n23998 = n23997 ^ n20557 ^ n18987 ;
  assign n24005 = n7228 ^ n2353 ^ 1'b0 ;
  assign n24003 = ( x134 & ~n6120 ) | ( x134 & n6286 ) | ( ~n6120 & n6286 ) ;
  assign n24004 = ( ~n11083 & n20449 ) | ( ~n11083 & n24003 ) | ( n20449 & n24003 ) ;
  assign n24000 = n14595 ^ n13692 ^ 1'b0 ;
  assign n24001 = n3246 | n24000 ;
  assign n23999 = n1022 | n23185 ;
  assign n24002 = n24001 ^ n23999 ^ 1'b0 ;
  assign n24006 = n24005 ^ n24004 ^ n24002 ;
  assign n24007 = n24006 ^ n23303 ^ n8589 ;
  assign n24008 = ( n4574 & ~n8374 ) | ( n4574 & n8857 ) | ( ~n8374 & n8857 ) ;
  assign n24009 = x156 & n24008 ;
  assign n24010 = n24009 ^ n9204 ^ 1'b0 ;
  assign n24011 = n3518 | n4728 ;
  assign n24012 = n12193 & ~n24011 ;
  assign n24013 = ( n10709 & n17460 ) | ( n10709 & ~n24012 ) | ( n17460 & ~n24012 ) ;
  assign n24014 = n22965 & n24013 ;
  assign n24015 = ( ~n3661 & n24010 ) | ( ~n3661 & n24014 ) | ( n24010 & n24014 ) ;
  assign n24016 = n6131 ^ n1621 ^ 1'b0 ;
  assign n24017 = n10773 & ~n24016 ;
  assign n24018 = n24017 ^ n541 ^ 1'b0 ;
  assign n24019 = n24018 ^ n12337 ^ n9799 ;
  assign n24020 = n15246 & ~n18404 ;
  assign n24021 = n4908 ^ n1023 ^ 1'b0 ;
  assign n24022 = n19293 | n24021 ;
  assign n24023 = n22134 | n24022 ;
  assign n24024 = n15053 ^ n9096 ^ n4967 ;
  assign n24025 = ~n2791 & n6314 ;
  assign n24026 = ~n3575 & n24025 ;
  assign n24027 = n15129 & ~n24026 ;
  assign n24028 = ~n16753 & n24027 ;
  assign n24029 = n10620 ^ n10169 ^ 1'b0 ;
  assign n24030 = n22391 & ~n24029 ;
  assign n24032 = n2071 & ~n18651 ;
  assign n24031 = ~n2140 & n10544 ;
  assign n24033 = n24032 ^ n24031 ^ 1'b0 ;
  assign n24034 = n24033 ^ n2000 ^ 1'b0 ;
  assign n24035 = n1156 & ~n24034 ;
  assign n24036 = n19391 ^ n14700 ^ 1'b0 ;
  assign n24037 = n12385 ^ n10723 ^ 1'b0 ;
  assign n24038 = n24037 ^ n13455 ^ 1'b0 ;
  assign n24039 = n24036 & n24038 ;
  assign n24040 = n10748 ^ n9586 ^ 1'b0 ;
  assign n24041 = n15929 ^ n2594 ^ x206 ;
  assign n24042 = n24040 & n24041 ;
  assign n24044 = ( ~n4094 & n14966 ) | ( ~n4094 & n14998 ) | ( n14966 & n14998 ) ;
  assign n24043 = n6756 & ~n13447 ;
  assign n24045 = n24044 ^ n24043 ^ n17234 ;
  assign n24047 = n18870 ^ n6001 ^ 1'b0 ;
  assign n24046 = n11234 & ~n14697 ;
  assign n24048 = n24047 ^ n24046 ^ n8487 ;
  assign n24049 = ( n5386 & ~n10908 ) | ( n5386 & n14223 ) | ( ~n10908 & n14223 ) ;
  assign n24050 = n19086 ^ n11137 ^ n3535 ;
  assign n24051 = n5036 & n24050 ;
  assign n24052 = ( n20588 & n24049 ) | ( n20588 & ~n24051 ) | ( n24049 & ~n24051 ) ;
  assign n24053 = n24052 ^ n5963 ^ 1'b0 ;
  assign n24054 = ~n2441 & n5313 ;
  assign n24055 = n2113 & n24054 ;
  assign n24056 = n7563 | n23892 ;
  assign n24057 = n13072 | n24056 ;
  assign n24058 = ( ~x161 & n1139 ) | ( ~x161 & n24057 ) | ( n1139 & n24057 ) ;
  assign n24059 = n13841 ^ n6899 ^ n6260 ;
  assign n24060 = n24059 ^ n17424 ^ 1'b0 ;
  assign n24061 = n24060 ^ n21660 ^ n12413 ;
  assign n24062 = n18801 ^ n11123 ^ n8330 ;
  assign n24063 = n18004 ^ n11606 ^ 1'b0 ;
  assign n24064 = n5700 & n24063 ;
  assign n24065 = n24064 ^ n10765 ^ n342 ;
  assign n24066 = n3760 ^ n1841 ^ 1'b0 ;
  assign n24067 = n8000 & ~n24066 ;
  assign n24068 = ( ~n11630 & n24065 ) | ( ~n11630 & n24067 ) | ( n24065 & n24067 ) ;
  assign n24069 = n19218 ^ n8326 ^ 1'b0 ;
  assign n24070 = n5237 & ~n15226 ;
  assign n24071 = n24070 ^ n20058 ^ 1'b0 ;
  assign n24072 = ~n23581 & n24071 ;
  assign n24073 = ~n12998 & n24072 ;
  assign n24074 = ( n2337 & ~n9073 ) | ( n2337 & n21708 ) | ( ~n9073 & n21708 ) ;
  assign n24075 = n12274 & ~n15228 ;
  assign n24076 = n24075 ^ n8324 ^ 1'b0 ;
  assign n24077 = n9156 | n24076 ;
  assign n24078 = n8118 ^ n1772 ^ 1'b0 ;
  assign n24079 = n15063 & ~n24078 ;
  assign n24080 = n21790 ^ n6737 ^ 1'b0 ;
  assign n24081 = n15766 & ~n24080 ;
  assign n24082 = n11800 & n18898 ;
  assign n24083 = n24081 & n24082 ;
  assign n24084 = n12940 ^ x137 ^ 1'b0 ;
  assign n24085 = ( n1630 & n5646 ) | ( n1630 & n24084 ) | ( n5646 & n24084 ) ;
  assign n24086 = n465 & ~n24085 ;
  assign n24087 = ~n11297 & n24086 ;
  assign n24088 = n9719 & n23120 ;
  assign n24089 = n2545 & n24088 ;
  assign n24090 = n16597 | n24089 ;
  assign n24091 = n24087 & ~n24090 ;
  assign n24092 = n776 | n12768 ;
  assign n24093 = n2025 | n7453 ;
  assign n24094 = n870 | n10160 ;
  assign n24095 = n24093 | n24094 ;
  assign n24096 = n3906 & n24095 ;
  assign n24097 = ~n24092 & n24096 ;
  assign n24098 = n24097 ^ n20393 ^ 1'b0 ;
  assign n24099 = n3561 & n15847 ;
  assign n24100 = n10961 & n17515 ;
  assign n24101 = n7168 & ~n8735 ;
  assign n24102 = n24101 ^ n1666 ^ 1'b0 ;
  assign n24105 = ( x81 & n585 ) | ( x81 & n4491 ) | ( n585 & n4491 ) ;
  assign n24104 = n10571 | n19798 ;
  assign n24106 = n24105 ^ n24104 ^ 1'b0 ;
  assign n24107 = n24106 ^ n4087 ^ 1'b0 ;
  assign n24108 = ( n3271 & n5114 ) | ( n3271 & n24107 ) | ( n5114 & n24107 ) ;
  assign n24103 = n6367 | n10949 ;
  assign n24109 = n24108 ^ n24103 ^ n1864 ;
  assign n24110 = n24109 ^ n3864 ^ 1'b0 ;
  assign n24111 = ( ~n4445 & n19518 ) | ( ~n4445 & n20079 ) | ( n19518 & n20079 ) ;
  assign n24112 = n24111 ^ n15022 ^ 1'b0 ;
  assign n24113 = n24112 ^ n9865 ^ 1'b0 ;
  assign n24114 = ( n2443 & ~n16095 ) | ( n2443 & n20077 ) | ( ~n16095 & n20077 ) ;
  assign n24115 = n15632 ^ n3919 ^ 1'b0 ;
  assign n24116 = ~n23179 & n24115 ;
  assign n24117 = n14822 & n24116 ;
  assign n24118 = n23649 ^ n11242 ^ n5309 ;
  assign n24120 = n18174 ^ n2018 ^ 1'b0 ;
  assign n24119 = n8109 & ~n16642 ;
  assign n24121 = n24120 ^ n24119 ^ 1'b0 ;
  assign n24123 = n11458 ^ n2681 ^ 1'b0 ;
  assign n24124 = n24123 ^ n9787 ^ n6811 ;
  assign n24122 = n1513 & n16960 ;
  assign n24125 = n24124 ^ n24122 ^ 1'b0 ;
  assign n24130 = n10097 ^ n6859 ^ 1'b0 ;
  assign n24126 = n8945 ^ n8281 ^ 1'b0 ;
  assign n24127 = n7790 | n24126 ;
  assign n24128 = n12320 | n24127 ;
  assign n24129 = n24128 ^ n1125 ^ 1'b0 ;
  assign n24131 = n24130 ^ n24129 ^ 1'b0 ;
  assign n24132 = ~n1958 & n14590 ;
  assign n24133 = n18386 & n24132 ;
  assign n24134 = n24133 ^ n9019 ^ 1'b0 ;
  assign n24140 = n19828 ^ n2335 ^ n1705 ;
  assign n24136 = ( ~n1646 & n2492 ) | ( ~n1646 & n9490 ) | ( n2492 & n9490 ) ;
  assign n24135 = ~n2357 & n12897 ;
  assign n24137 = n24136 ^ n24135 ^ 1'b0 ;
  assign n24138 = n9312 & ~n11766 ;
  assign n24139 = ~n24137 & n24138 ;
  assign n24141 = n24140 ^ n24139 ^ n14873 ;
  assign n24142 = n3668 & ~n9787 ;
  assign n24143 = n24142 ^ n5634 ^ 1'b0 ;
  assign n24144 = n5125 ^ n1140 ^ n425 ;
  assign n24145 = n18772 ^ n5734 ^ 1'b0 ;
  assign n24146 = n24144 & ~n24145 ;
  assign n24147 = ( ~n6224 & n8654 ) | ( ~n6224 & n10152 ) | ( n8654 & n10152 ) ;
  assign n24148 = n24147 ^ n12055 ^ n6885 ;
  assign n24150 = n5776 ^ n4640 ^ 1'b0 ;
  assign n24151 = ~n2874 & n24150 ;
  assign n24149 = n23340 ^ n21280 ^ n6968 ;
  assign n24152 = n24151 ^ n24149 ^ n4467 ;
  assign n24153 = ~n3129 & n4499 ;
  assign n24154 = n24153 ^ n3770 ^ 1'b0 ;
  assign n24155 = n24154 ^ n8403 ^ 1'b0 ;
  assign n24156 = ~n8077 & n24155 ;
  assign n24157 = n24156 ^ n2731 ^ n2551 ;
  assign n24158 = n24157 ^ n8985 ^ 1'b0 ;
  assign n24159 = n1113 & n24158 ;
  assign n24162 = n1111 & ~n19360 ;
  assign n24163 = n7920 & ~n10086 ;
  assign n24164 = n24162 & n24163 ;
  assign n24160 = n2744 & n23951 ;
  assign n24161 = n24160 ^ n16192 ^ 1'b0 ;
  assign n24165 = n24164 ^ n24161 ^ n1068 ;
  assign n24168 = n6992 | n23728 ;
  assign n24166 = n13025 ^ n7699 ^ 1'b0 ;
  assign n24167 = n24166 ^ n17433 ^ n5257 ;
  assign n24169 = n24168 ^ n24167 ^ n11634 ;
  assign n24170 = ( n2521 & n3808 ) | ( n2521 & ~n24169 ) | ( n3808 & ~n24169 ) ;
  assign n24171 = n20875 ^ n17161 ^ n11278 ;
  assign n24172 = n23825 ^ n16873 ^ n3308 ;
  assign n24173 = ( n17123 & n18929 ) | ( n17123 & n21696 ) | ( n18929 & n21696 ) ;
  assign n24174 = ( n2012 & n4841 ) | ( n2012 & n6304 ) | ( n4841 & n6304 ) ;
  assign n24175 = n24174 ^ n7309 ^ 1'b0 ;
  assign n24176 = ( n5215 & n8832 ) | ( n5215 & n10151 ) | ( n8832 & n10151 ) ;
  assign n24177 = n24176 ^ n12198 ^ 1'b0 ;
  assign n24178 = ~n2118 & n24177 ;
  assign n24180 = ~n2769 & n16587 ;
  assign n24181 = n24180 ^ n12868 ^ 1'b0 ;
  assign n24179 = n6785 & ~n6787 ;
  assign n24182 = n24181 ^ n24179 ^ 1'b0 ;
  assign n24183 = ( n261 & ~n16160 ) | ( n261 & n24182 ) | ( ~n16160 & n24182 ) ;
  assign n24184 = n14568 ^ n3413 ^ 1'b0 ;
  assign n24185 = ~n17288 & n23620 ;
  assign n24186 = n24185 ^ n20081 ^ n1457 ;
  assign n24187 = ( n2482 & ~n17033 ) | ( n2482 & n24186 ) | ( ~n17033 & n24186 ) ;
  assign n24188 = n10654 ^ n4649 ^ 1'b0 ;
  assign n24189 = n6928 & ~n24188 ;
  assign n24190 = n24189 ^ n4716 ^ 1'b0 ;
  assign n24191 = n662 & n6401 ;
  assign n24192 = ~n22734 & n24191 ;
  assign n24193 = n8169 & n24192 ;
  assign n24194 = n11530 ^ n7199 ^ n834 ;
  assign n24195 = n24194 ^ n12929 ^ 1'b0 ;
  assign n24196 = n24193 & ~n24195 ;
  assign n24197 = n14537 ^ n10255 ^ 1'b0 ;
  assign n24198 = n24196 & n24197 ;
  assign n24201 = n11937 | n14188 ;
  assign n24199 = ~n11905 & n17144 ;
  assign n24200 = ~n10193 & n24199 ;
  assign n24202 = n24201 ^ n24200 ^ 1'b0 ;
  assign n24203 = n16490 ^ n13247 ^ n3948 ;
  assign n24204 = n16407 ^ n11035 ^ 1'b0 ;
  assign n24205 = n9166 & n13547 ;
  assign n24206 = n5761 & n24205 ;
  assign n24207 = n18209 ^ n10815 ^ n7098 ;
  assign n24208 = n16513 | n24207 ;
  assign n24209 = n24206 & ~n24208 ;
  assign n24210 = ~n14070 & n14669 ;
  assign n24211 = n24210 ^ n19898 ^ 1'b0 ;
  assign n24212 = n7672 | n23974 ;
  assign n24213 = n11166 ^ n1367 ^ 1'b0 ;
  assign n24214 = n24213 ^ n12401 ^ n12030 ;
  assign n24215 = n7908 & ~n10701 ;
  assign n24216 = ( n5004 & ~n21133 ) | ( n5004 & n24215 ) | ( ~n21133 & n24215 ) ;
  assign n24217 = n14683 & n22233 ;
  assign n24218 = n24217 ^ n6263 ^ 1'b0 ;
  assign n24219 = n9574 | n15650 ;
  assign n24220 = n15929 & ~n24219 ;
  assign n24221 = n1370 & ~n24220 ;
  assign n24222 = n24221 ^ n1237 ^ 1'b0 ;
  assign n24223 = n3059 | n24215 ;
  assign n24224 = n11966 ^ n4012 ^ x118 ;
  assign n24225 = n16732 ^ n9842 ^ n2714 ;
  assign n24226 = ~n979 & n7858 ;
  assign n24227 = ~n8633 & n24226 ;
  assign n24228 = ( n1466 & ~n24225 ) | ( n1466 & n24227 ) | ( ~n24225 & n24227 ) ;
  assign n24229 = ( n2421 & n11906 ) | ( n2421 & ~n12643 ) | ( n11906 & ~n12643 ) ;
  assign n24230 = ~n14970 & n24229 ;
  assign n24234 = n9277 ^ n5433 ^ 1'b0 ;
  assign n24235 = ~n16583 & n24234 ;
  assign n24231 = n12278 ^ n4654 ^ 1'b0 ;
  assign n24232 = ( n8489 & n13654 ) | ( n8489 & ~n24231 ) | ( n13654 & ~n24231 ) ;
  assign n24233 = n24232 ^ n24104 ^ n3408 ;
  assign n24236 = n24235 ^ n24233 ^ n20257 ;
  assign n24237 = ( n3601 & ~n4625 ) | ( n3601 & n12052 ) | ( ~n4625 & n12052 ) ;
  assign n24238 = n4277 | n6392 ;
  assign n24239 = n24237 | n24238 ;
  assign n24240 = n4822 ^ n1978 ^ n1258 ;
  assign n24241 = n24240 ^ n5832 ^ n3993 ;
  assign n24242 = n24241 ^ n21548 ^ 1'b0 ;
  assign n24243 = n19201 & n24242 ;
  assign n24244 = ( n6666 & ~n24239 ) | ( n6666 & n24243 ) | ( ~n24239 & n24243 ) ;
  assign n24245 = n11852 | n13272 ;
  assign n24246 = n12446 | n24245 ;
  assign n24247 = ( n5664 & n18195 ) | ( n5664 & n24246 ) | ( n18195 & n24246 ) ;
  assign n24248 = n14848 & ~n21532 ;
  assign n24249 = n21358 ^ n6413 ^ 1'b0 ;
  assign n24250 = n3103 & ~n24249 ;
  assign n24251 = n7397 ^ n2147 ^ n1692 ;
  assign n24252 = n11729 ^ n8982 ^ 1'b0 ;
  assign n24253 = ~n21142 & n24252 ;
  assign n24254 = ~n7994 & n24253 ;
  assign n24255 = n24251 & ~n24254 ;
  assign n24256 = n13863 ^ n4285 ^ 1'b0 ;
  assign n24257 = n22883 ^ n11355 ^ 1'b0 ;
  assign n24258 = n24257 ^ n10337 ^ 1'b0 ;
  assign n24259 = ~n24256 & n24258 ;
  assign n24260 = n14142 & n24259 ;
  assign n24261 = n24260 ^ n11931 ^ 1'b0 ;
  assign n24262 = n20500 ^ n16796 ^ 1'b0 ;
  assign n24263 = ~n12450 & n24262 ;
  assign n24264 = n14702 ^ n11123 ^ n8082 ;
  assign n24265 = n24264 ^ n21970 ^ n2828 ;
  assign n24266 = n13055 ^ n10974 ^ n2183 ;
  assign n24267 = ~n5353 & n24266 ;
  assign n24268 = ( n8608 & ~n12332 ) | ( n8608 & n18206 ) | ( ~n12332 & n18206 ) ;
  assign n24269 = n6017 & ~n10215 ;
  assign n24270 = n24268 & n24269 ;
  assign n24271 = n13544 & n24270 ;
  assign n24272 = n1700 & n8139 ;
  assign n24273 = n2901 | n24272 ;
  assign n24274 = n4878 & ~n10480 ;
  assign n24275 = ( n3861 & n9969 ) | ( n3861 & ~n11544 ) | ( n9969 & ~n11544 ) ;
  assign n24276 = n24275 ^ n20421 ^ n2551 ;
  assign n24277 = ( n1803 & ~n8453 ) | ( n1803 & n12841 ) | ( ~n8453 & n12841 ) ;
  assign n24278 = n18980 ^ n1157 ^ 1'b0 ;
  assign n24279 = n24277 & ~n24278 ;
  assign n24280 = n9191 ^ n6520 ^ n3647 ;
  assign n24281 = n13848 & n24280 ;
  assign n24282 = n24281 ^ n15062 ^ 1'b0 ;
  assign n24283 = n6010 & ~n24282 ;
  assign n24284 = ~n18264 & n24283 ;
  assign n24288 = n12337 ^ n6599 ^ n2240 ;
  assign n24285 = n2910 & n12205 ;
  assign n24286 = n12219 & n24285 ;
  assign n24287 = ~n15674 & n24286 ;
  assign n24289 = n24288 ^ n24287 ^ n14136 ;
  assign n24290 = n5145 ^ n3403 ^ x160 ;
  assign n24291 = n4468 & ~n24290 ;
  assign n24292 = ~n14851 & n16372 ;
  assign n24293 = n24291 & n24292 ;
  assign n24294 = ( n7097 & ~n24289 ) | ( n7097 & n24293 ) | ( ~n24289 & n24293 ) ;
  assign n24295 = n23221 ^ n15510 ^ 1'b0 ;
  assign n24296 = n4240 & ~n24295 ;
  assign n24297 = ( n1567 & ~n5480 ) | ( n1567 & n20643 ) | ( ~n5480 & n20643 ) ;
  assign n24298 = ( n9767 & n23897 ) | ( n9767 & ~n24297 ) | ( n23897 & ~n24297 ) ;
  assign n24299 = ( ~n7650 & n10364 ) | ( ~n7650 & n12046 ) | ( n10364 & n12046 ) ;
  assign n24300 = ( n3924 & n23170 ) | ( n3924 & ~n24299 ) | ( n23170 & ~n24299 ) ;
  assign n24301 = n4875 | n24300 ;
  assign n24302 = n13894 & n22825 ;
  assign n24303 = n22767 ^ n20396 ^ n9401 ;
  assign n24304 = n16770 ^ n5850 ^ 1'b0 ;
  assign n24305 = n24304 ^ n21037 ^ n10375 ;
  assign n24306 = n6329 & n22278 ;
  assign n24307 = n24306 ^ n10748 ^ 1'b0 ;
  assign n24308 = n16621 ^ n8677 ^ n6957 ;
  assign n24309 = ~n1580 & n6149 ;
  assign n24310 = n3916 & n24309 ;
  assign n24311 = n24310 ^ n8480 ^ n1572 ;
  assign n24312 = ( ~n620 & n17808 ) | ( ~n620 & n24311 ) | ( n17808 & n24311 ) ;
  assign n24313 = ( n6468 & n18270 ) | ( n6468 & n24312 ) | ( n18270 & n24312 ) ;
  assign n24314 = ( n325 & n685 ) | ( n325 & ~n16914 ) | ( n685 & ~n16914 ) ;
  assign n24315 = n14828 ^ n5753 ^ 1'b0 ;
  assign n24316 = ( ~n5616 & n13068 ) | ( ~n5616 & n24315 ) | ( n13068 & n24315 ) ;
  assign n24317 = n5775 & ~n17292 ;
  assign n24318 = n24317 ^ n18773 ^ 1'b0 ;
  assign n24319 = n12266 ^ n7362 ^ 1'b0 ;
  assign n24320 = ( n4755 & ~n24318 ) | ( n4755 & n24319 ) | ( ~n24318 & n24319 ) ;
  assign n24321 = n24320 ^ n11467 ^ n474 ;
  assign n24322 = ( n4538 & n7878 ) | ( n4538 & ~n15653 ) | ( n7878 & ~n15653 ) ;
  assign n24323 = ~n12725 & n24322 ;
  assign n24324 = n24323 ^ n12663 ^ 1'b0 ;
  assign n24325 = n24324 ^ n12341 ^ n7372 ;
  assign n24326 = n448 ^ x164 ^ 1'b0 ;
  assign n24327 = n6774 ^ n5823 ^ 1'b0 ;
  assign n24328 = n10876 & n24327 ;
  assign n24329 = n10743 ^ n8838 ^ 1'b0 ;
  assign n24330 = n21853 ^ n4975 ^ 1'b0 ;
  assign n24331 = ~n6145 & n24330 ;
  assign n24338 = ( n3141 & ~n6992 ) | ( n3141 & n13576 ) | ( ~n6992 & n13576 ) ;
  assign n24332 = n6032 ^ n5404 ^ 1'b0 ;
  assign n24333 = n3004 & ~n24332 ;
  assign n24334 = ~n17246 & n24333 ;
  assign n24335 = n24334 ^ n9067 ^ 1'b0 ;
  assign n24336 = n394 & n6810 ;
  assign n24337 = ( n2365 & ~n24335 ) | ( n2365 & n24336 ) | ( ~n24335 & n24336 ) ;
  assign n24339 = n24338 ^ n24337 ^ n17566 ;
  assign n24340 = n21519 ^ n7187 ^ 1'b0 ;
  assign n24341 = n3347 & n3490 ;
  assign n24342 = n24341 ^ n14131 ^ 1'b0 ;
  assign n24343 = n24342 ^ n23228 ^ n1623 ;
  assign n24344 = n20948 ^ n15910 ^ 1'b0 ;
  assign n24345 = n24343 | n24344 ;
  assign n24346 = ~n14481 & n21638 ;
  assign n24347 = n7187 & n24346 ;
  assign n24348 = n6786 ^ n2727 ^ 1'b0 ;
  assign n24349 = n22353 ^ n22198 ^ n21743 ;
  assign n24350 = n7060 ^ n6027 ^ 1'b0 ;
  assign n24351 = n9946 & n24350 ;
  assign n24352 = n21864 ^ n564 ^ 1'b0 ;
  assign n24353 = ( n3142 & n24351 ) | ( n3142 & ~n24352 ) | ( n24351 & ~n24352 ) ;
  assign n24354 = ( ~n2017 & n24349 ) | ( ~n2017 & n24353 ) | ( n24349 & n24353 ) ;
  assign n24355 = n1064 & n23463 ;
  assign n24356 = n2310 & ~n10412 ;
  assign n24357 = n24356 ^ n13888 ^ 1'b0 ;
  assign n24358 = ~n8103 & n24357 ;
  assign n24359 = n24358 ^ n21867 ^ n18320 ;
  assign n24360 = ( ~n11364 & n13879 ) | ( ~n11364 & n14287 ) | ( n13879 & n14287 ) ;
  assign n24361 = n9492 ^ n4603 ^ 1'b0 ;
  assign n24362 = n2292 & n20424 ;
  assign n24363 = n20645 ^ n14787 ^ n4808 ;
  assign n24364 = n8021 ^ n4925 ^ x127 ;
  assign n24365 = ( ~n2008 & n20096 ) | ( ~n2008 & n24364 ) | ( n20096 & n24364 ) ;
  assign n24366 = ~n3643 & n9595 ;
  assign n24367 = n24366 ^ n2580 ^ 1'b0 ;
  assign n24368 = n24109 ^ n15313 ^ 1'b0 ;
  assign n24369 = n20026 & n24368 ;
  assign n24370 = n4724 & ~n6374 ;
  assign n24371 = ~n9544 & n24370 ;
  assign n24372 = n24371 ^ n21863 ^ n10210 ;
  assign n24373 = n3427 ^ n3254 ^ n1701 ;
  assign n24374 = n24373 ^ n4379 ^ 1'b0 ;
  assign n24375 = ( n3705 & ~n5840 ) | ( n3705 & n10052 ) | ( ~n5840 & n10052 ) ;
  assign n24376 = n24375 ^ n16521 ^ x57 ;
  assign n24377 = ( n14493 & ~n24374 ) | ( n14493 & n24376 ) | ( ~n24374 & n24376 ) ;
  assign n24378 = n5961 | n12563 ;
  assign n24379 = ( ~n2064 & n5981 ) | ( ~n2064 & n24378 ) | ( n5981 & n24378 ) ;
  assign n24380 = n24379 ^ n12544 ^ 1'b0 ;
  assign n24381 = ~n3509 & n4768 ;
  assign n24382 = n24381 ^ n15182 ^ 1'b0 ;
  assign n24383 = n6485 ^ n3549 ^ 1'b0 ;
  assign n24384 = ~n24382 & n24383 ;
  assign n24385 = n13372 ^ n12260 ^ n6586 ;
  assign n24386 = n24385 ^ n11659 ^ n2396 ;
  assign n24387 = ( ~n5812 & n24384 ) | ( ~n5812 & n24386 ) | ( n24384 & n24386 ) ;
  assign n24388 = n1054 & ~n18192 ;
  assign n24389 = ( n14875 & ~n18593 ) | ( n14875 & n24388 ) | ( ~n18593 & n24388 ) ;
  assign n24391 = n16013 ^ n10244 ^ n6616 ;
  assign n24390 = n10831 & n18157 ;
  assign n24392 = n24391 ^ n24390 ^ 1'b0 ;
  assign n24393 = n7355 | n13888 ;
  assign n24394 = ~n3798 & n7621 ;
  assign n24395 = ( n5328 & ~n14671 ) | ( n5328 & n24394 ) | ( ~n14671 & n24394 ) ;
  assign n24396 = n24395 ^ n18885 ^ 1'b0 ;
  assign n24397 = n2390 | n14754 ;
  assign n24398 = ( ~n5110 & n13027 ) | ( ~n5110 & n24397 ) | ( n13027 & n24397 ) ;
  assign n24399 = n9879 ^ n8820 ^ n258 ;
  assign n24400 = n1886 & ~n24399 ;
  assign n24401 = n24400 ^ n9103 ^ 1'b0 ;
  assign n24402 = n15374 & n24401 ;
  assign n24403 = n17855 ^ n4864 ^ n2325 ;
  assign n24404 = n22970 ^ n4819 ^ 1'b0 ;
  assign n24405 = ~n2021 & n24404 ;
  assign n24406 = ( n9538 & n17004 ) | ( n9538 & ~n24008 ) | ( n17004 & ~n24008 ) ;
  assign n24408 = n6753 | n7718 ;
  assign n24409 = n24408 ^ n14419 ^ 1'b0 ;
  assign n24410 = n24409 ^ n5440 ^ n4759 ;
  assign n24411 = n24410 ^ n7568 ^ 1'b0 ;
  assign n24407 = n5186 | n12290 ;
  assign n24412 = n24411 ^ n24407 ^ 1'b0 ;
  assign n24413 = n4063 & ~n5613 ;
  assign n24414 = n5264 & ~n19654 ;
  assign n24415 = ~n6338 & n24414 ;
  assign n24416 = ( n5251 & ~n22827 ) | ( n5251 & n24415 ) | ( ~n22827 & n24415 ) ;
  assign n24417 = n24413 | n24416 ;
  assign n24418 = n11120 ^ n3366 ^ n1632 ;
  assign n24419 = n22119 & n24418 ;
  assign n24420 = n4228 & n20816 ;
  assign n24423 = ( n5041 & n11175 ) | ( n5041 & n16021 ) | ( n11175 & n16021 ) ;
  assign n24422 = n16824 ^ n7700 ^ n1064 ;
  assign n24421 = n23250 ^ n11044 ^ n9508 ;
  assign n24424 = n24423 ^ n24422 ^ n24421 ;
  assign n24425 = n23169 ^ n15105 ^ 1'b0 ;
  assign n24426 = ( ~n8028 & n10653 ) | ( ~n8028 & n24013 ) | ( n10653 & n24013 ) ;
  assign n24427 = n4045 | n14787 ;
  assign n24428 = ( n15526 & n24426 ) | ( n15526 & n24427 ) | ( n24426 & n24427 ) ;
  assign n24429 = n24428 ^ n7498 ^ 1'b0 ;
  assign n24430 = n24425 & n24429 ;
  assign n24431 = n10098 | n12624 ;
  assign n24432 = n24431 ^ n12990 ^ 1'b0 ;
  assign n24433 = n18780 ^ n8803 ^ n3349 ;
  assign n24434 = n24433 ^ n23442 ^ 1'b0 ;
  assign n24435 = n8821 ^ n3771 ^ 1'b0 ;
  assign n24436 = ( n572 & ~n909 ) | ( n572 & n1398 ) | ( ~n909 & n1398 ) ;
  assign n24437 = n22479 & ~n24436 ;
  assign n24438 = n24437 ^ n9607 ^ 1'b0 ;
  assign n24439 = ( n1849 & ~n24435 ) | ( n1849 & n24438 ) | ( ~n24435 & n24438 ) ;
  assign n24440 = ~n1519 & n2992 ;
  assign n24441 = n24440 ^ n7757 ^ 1'b0 ;
  assign n24442 = n24441 ^ n2487 ^ n821 ;
  assign n24443 = n19850 & n24442 ;
  assign n24444 = ~n4738 & n24443 ;
  assign n24445 = n13229 ^ n9892 ^ 1'b0 ;
  assign n24446 = ( ~n3172 & n6161 ) | ( ~n3172 & n24445 ) | ( n6161 & n24445 ) ;
  assign n24447 = n24446 ^ n8297 ^ 1'b0 ;
  assign n24448 = n8157 & n9535 ;
  assign n24449 = n5717 & n24448 ;
  assign n24450 = n24447 & n24449 ;
  assign n24451 = ( ~n2255 & n21670 ) | ( ~n2255 & n24450 ) | ( n21670 & n24450 ) ;
  assign n24452 = n12296 ^ n2526 ^ 1'b0 ;
  assign n24453 = n999 & n24452 ;
  assign n24454 = n1823 & n3253 ;
  assign n24455 = ( ~n18612 & n23007 ) | ( ~n18612 & n24454 ) | ( n23007 & n24454 ) ;
  assign n24456 = n7638 ^ n2931 ^ 1'b0 ;
  assign n24457 = n23258 & n24456 ;
  assign n24458 = n24457 ^ n8958 ^ n1790 ;
  assign n24459 = n24455 & n24458 ;
  assign n24460 = ~n24453 & n24459 ;
  assign n24461 = ( n7352 & ~n8774 ) | ( n7352 & n21844 ) | ( ~n8774 & n21844 ) ;
  assign n24462 = n24461 ^ n15729 ^ n2671 ;
  assign n24463 = n21236 ^ n12881 ^ 1'b0 ;
  assign n24464 = n19823 ^ n5015 ^ n1665 ;
  assign n24465 = n9835 | n24464 ;
  assign n24466 = n23302 ^ n13028 ^ 1'b0 ;
  assign n24467 = n24465 | n24466 ;
  assign n24470 = ( n416 & ~n4965 ) | ( n416 & n8743 ) | ( ~n4965 & n8743 ) ;
  assign n24469 = n10574 | n19064 ;
  assign n24471 = n24470 ^ n24469 ^ 1'b0 ;
  assign n24468 = n1131 | n4927 ;
  assign n24472 = n24471 ^ n24468 ^ 1'b0 ;
  assign n24473 = n11248 & n24472 ;
  assign n24474 = n24473 ^ n8862 ^ n4902 ;
  assign n24475 = ~n16922 & n20849 ;
  assign n24476 = ~n12442 & n24475 ;
  assign n24477 = n1558 & ~n22011 ;
  assign n24478 = n24476 & n24477 ;
  assign n24482 = ~n5548 & n8393 ;
  assign n24479 = n5997 & n9815 ;
  assign n24480 = n9575 & n24479 ;
  assign n24481 = n589 | n24480 ;
  assign n24483 = n24482 ^ n24481 ^ 1'b0 ;
  assign n24484 = n8836 & ~n20663 ;
  assign n24485 = n12311 & n24484 ;
  assign n24486 = n9942 & n12568 ;
  assign n24487 = ~n12568 & n24486 ;
  assign n24488 = ( n4650 & n5754 ) | ( n4650 & n19806 ) | ( n5754 & n19806 ) ;
  assign n24489 = n24488 ^ n19517 ^ n3016 ;
  assign n24490 = n17338 ^ n16350 ^ 1'b0 ;
  assign n24491 = n8241 | n24490 ;
  assign n24492 = ( ~n8458 & n10038 ) | ( ~n8458 & n16061 ) | ( n10038 & n16061 ) ;
  assign n24493 = n24492 ^ n943 ^ 1'b0 ;
  assign n24494 = n24493 ^ n12053 ^ n6479 ;
  assign n24495 = n4402 ^ n2748 ^ 1'b0 ;
  assign n24496 = ~n5188 & n5194 ;
  assign n24497 = n23029 | n24496 ;
  assign n24498 = ( n1806 & ~n19346 ) | ( n1806 & n24497 ) | ( ~n19346 & n24497 ) ;
  assign n24499 = n10516 & n15034 ;
  assign n24500 = n1208 & n24499 ;
  assign n24512 = n4499 & n6157 ;
  assign n24501 = n4829 ^ n2413 ^ 1'b0 ;
  assign n24502 = ~n642 & n24501 ;
  assign n24503 = n11789 & n24502 ;
  assign n24508 = n7568 ^ n2822 ^ n1138 ;
  assign n24509 = ( n2402 & n7778 ) | ( n2402 & n24508 ) | ( n7778 & n24508 ) ;
  assign n24506 = n17081 ^ n8506 ^ 1'b0 ;
  assign n24504 = ( n7588 & n11324 ) | ( n7588 & ~n11998 ) | ( n11324 & ~n11998 ) ;
  assign n24505 = ( n13543 & n23104 ) | ( n13543 & n24504 ) | ( n23104 & n24504 ) ;
  assign n24507 = n24506 ^ n24505 ^ 1'b0 ;
  assign n24510 = n24509 ^ n24507 ^ n13863 ;
  assign n24511 = ( n3999 & ~n24503 ) | ( n3999 & n24510 ) | ( ~n24503 & n24510 ) ;
  assign n24513 = n24512 ^ n24511 ^ 1'b0 ;
  assign n24514 = ( n10163 & n18188 ) | ( n10163 & ~n18504 ) | ( n18188 & ~n18504 ) ;
  assign n24515 = n24514 ^ n6374 ^ 1'b0 ;
  assign n24516 = n10033 ^ n9565 ^ n4983 ;
  assign n24521 = n12495 ^ n2333 ^ 1'b0 ;
  assign n24517 = ( n6100 & n10832 ) | ( n6100 & ~n24290 ) | ( n10832 & ~n24290 ) ;
  assign n24518 = ( n984 & n21254 ) | ( n984 & ~n24517 ) | ( n21254 & ~n24517 ) ;
  assign n24519 = n24518 ^ n8492 ^ n511 ;
  assign n24520 = ( n9601 & n9672 ) | ( n9601 & ~n24519 ) | ( n9672 & ~n24519 ) ;
  assign n24522 = n24521 ^ n24520 ^ n12914 ;
  assign n24523 = ( n14060 & n19791 ) | ( n14060 & ~n24522 ) | ( n19791 & ~n24522 ) ;
  assign n24524 = ( n24515 & n24516 ) | ( n24515 & n24523 ) | ( n24516 & n24523 ) ;
  assign n24525 = n12945 ^ n12510 ^ 1'b0 ;
  assign n24526 = n5269 & n24525 ;
  assign n24527 = n24526 ^ n16800 ^ n9200 ;
  assign n24528 = ( n2605 & ~n6872 ) | ( n2605 & n21607 ) | ( ~n6872 & n21607 ) ;
  assign n24529 = ~n5345 & n17836 ;
  assign n24530 = n19065 | n22325 ;
  assign n24531 = n24529 & ~n24530 ;
  assign n24532 = n541 | n11935 ;
  assign n24533 = n18560 & ~n24532 ;
  assign n24534 = ( n3465 & n24531 ) | ( n3465 & ~n24533 ) | ( n24531 & ~n24533 ) ;
  assign n24535 = n2051 & ~n8160 ;
  assign n24536 = n24535 ^ n23736 ^ 1'b0 ;
  assign n24539 = n5060 ^ n988 ^ n683 ;
  assign n24537 = n1045 | n15930 ;
  assign n24538 = ( n6742 & n24067 ) | ( n6742 & ~n24537 ) | ( n24067 & ~n24537 ) ;
  assign n24540 = n24539 ^ n24538 ^ 1'b0 ;
  assign n24541 = n17713 | n24540 ;
  assign n24542 = n18827 ^ n1838 ^ 1'b0 ;
  assign n24543 = n11956 | n24542 ;
  assign n24544 = n24543 ^ n16691 ^ n2875 ;
  assign n24545 = ~n1772 & n6901 ;
  assign n24546 = ~x81 & n18270 ;
  assign n24547 = n24546 ^ n11526 ^ 1'b0 ;
  assign n24548 = n10824 ^ n3229 ^ 1'b0 ;
  assign n24549 = ~n8954 & n24548 ;
  assign n24550 = n5354 & n24549 ;
  assign n24551 = ~n3162 & n10376 ;
  assign n24552 = ~n2001 & n5399 ;
  assign n24553 = n24552 ^ n7709 ^ 1'b0 ;
  assign n24554 = ( n3917 & n22925 ) | ( n3917 & ~n24553 ) | ( n22925 & ~n24553 ) ;
  assign n24555 = ( ~n7597 & n14274 ) | ( ~n7597 & n16071 ) | ( n14274 & n16071 ) ;
  assign n24556 = ( n3629 & n23495 ) | ( n3629 & ~n24555 ) | ( n23495 & ~n24555 ) ;
  assign n24557 = n12292 | n24556 ;
  assign n24558 = n3704 & n9205 ;
  assign n24559 = n24558 ^ n24080 ^ 1'b0 ;
  assign n24560 = n13905 | n24559 ;
  assign n24561 = n24560 ^ n3363 ^ 1'b0 ;
  assign n24572 = n4591 & n11440 ;
  assign n24573 = n24572 ^ n11857 ^ 1'b0 ;
  assign n24570 = n10574 ^ n3666 ^ n2356 ;
  assign n24569 = n9763 | n11876 ;
  assign n24571 = n24570 ^ n24569 ^ 1'b0 ;
  assign n24574 = n24573 ^ n24571 ^ n19913 ;
  assign n24562 = n2924 & n6529 ;
  assign n24563 = ( ~n5856 & n17091 ) | ( ~n5856 & n24562 ) | ( n17091 & n24562 ) ;
  assign n24564 = n9491 | n24563 ;
  assign n24565 = n22470 & ~n24564 ;
  assign n24566 = n12923 ^ n1629 ^ n606 ;
  assign n24567 = n24566 ^ n4791 ^ 1'b0 ;
  assign n24568 = ~n24565 & n24567 ;
  assign n24575 = n24574 ^ n24568 ^ n7920 ;
  assign n24576 = n4045 | n5133 ;
  assign n24577 = ~n729 & n18445 ;
  assign n24578 = n24577 ^ n556 ^ 1'b0 ;
  assign n24579 = ( x227 & n24576 ) | ( x227 & n24578 ) | ( n24576 & n24578 ) ;
  assign n24580 = ( n3298 & n21272 ) | ( n3298 & ~n24579 ) | ( n21272 & ~n24579 ) ;
  assign n24581 = n3326 & n6416 ;
  assign n24582 = n10294 ^ n8319 ^ 1'b0 ;
  assign n24583 = n10042 ^ n5930 ^ 1'b0 ;
  assign n24584 = ~n4068 & n24583 ;
  assign n24585 = ( ~n24581 & n24582 ) | ( ~n24581 & n24584 ) | ( n24582 & n24584 ) ;
  assign n24586 = n20339 & ~n24585 ;
  assign n24587 = n8319 | n24586 ;
  assign n24588 = n24587 ^ n1447 ^ 1'b0 ;
  assign n24589 = ( n22863 & ~n24580 ) | ( n22863 & n24588 ) | ( ~n24580 & n24588 ) ;
  assign n24590 = n23815 ^ n6797 ^ n6579 ;
  assign n24591 = n1227 & n9252 ;
  assign n24592 = n24591 ^ n16924 ^ n1545 ;
  assign n24593 = n1365 & n12476 ;
  assign n24594 = n24593 ^ n11658 ^ n6489 ;
  assign n24595 = n18377 ^ n3523 ^ n3379 ;
  assign n24596 = n7844 & ~n9989 ;
  assign n24597 = n3016 & n11642 ;
  assign n24598 = n24597 ^ n10518 ^ 1'b0 ;
  assign n24599 = n24596 & ~n24598 ;
  assign n24600 = ~n17301 & n18539 ;
  assign n24601 = n24600 ^ n21444 ^ 1'b0 ;
  assign n24604 = ~n9205 & n11120 ;
  assign n24605 = ( n2018 & n6002 ) | ( n2018 & n24604 ) | ( n6002 & n24604 ) ;
  assign n24606 = n21870 | n24605 ;
  assign n24602 = n19823 ^ n18334 ^ n6355 ;
  assign n24603 = n24602 ^ n22091 ^ n9292 ;
  assign n24607 = n24606 ^ n24603 ^ n14976 ;
  assign n24608 = n20421 ^ n10917 ^ n5350 ;
  assign n24609 = n9852 & ~n13030 ;
  assign n24610 = ( ~n2137 & n24608 ) | ( ~n2137 & n24609 ) | ( n24608 & n24609 ) ;
  assign n24611 = n10639 ^ n8400 ^ 1'b0 ;
  assign n24612 = ( x250 & n5192 ) | ( x250 & ~n14950 ) | ( n5192 & ~n14950 ) ;
  assign n24613 = ~n5966 & n24612 ;
  assign n24614 = n7862 ^ x134 ^ 1'b0 ;
  assign n24615 = ~n5587 & n24614 ;
  assign n24616 = n7926 ^ n2208 ^ n792 ;
  assign n24621 = n1775 & n6887 ;
  assign n24622 = n24621 ^ n4071 ^ n883 ;
  assign n24619 = n20987 ^ n11378 ^ 1'b0 ;
  assign n24617 = n16647 ^ n557 ^ 1'b0 ;
  assign n24618 = n6762 | n24617 ;
  assign n24620 = n24619 ^ n24618 ^ n5400 ;
  assign n24623 = n24622 ^ n24620 ^ n24051 ;
  assign n24624 = n1685 | n3705 ;
  assign n24625 = n3059 | n24624 ;
  assign n24626 = n24625 ^ n17403 ^ 1'b0 ;
  assign n24627 = ~n2791 & n17799 ;
  assign n24628 = n10075 ^ n4348 ^ 1'b0 ;
  assign n24629 = n24627 | n24628 ;
  assign n24630 = n13075 ^ n11579 ^ n697 ;
  assign n24631 = n18868 ^ n9956 ^ n3331 ;
  assign n24632 = ~n24630 & n24631 ;
  assign n24633 = n24386 ^ n8714 ^ n4692 ;
  assign n24634 = n19667 | n24001 ;
  assign n24635 = n7892 & ~n24634 ;
  assign n24636 = n474 & ~n19007 ;
  assign n24637 = n22256 & ~n24636 ;
  assign n24638 = n24332 ^ n8224 ^ 1'b0 ;
  assign n24639 = ~n20206 & n24638 ;
  assign n24642 = ( n4454 & n8331 ) | ( n4454 & n17017 ) | ( n8331 & n17017 ) ;
  assign n24640 = n11944 ^ n5036 ^ n3718 ;
  assign n24641 = ( ~n6932 & n16199 ) | ( ~n6932 & n24640 ) | ( n16199 & n24640 ) ;
  assign n24643 = n24642 ^ n24641 ^ n13272 ;
  assign n24644 = n12520 | n14752 ;
  assign n24645 = n3910 & ~n24644 ;
  assign n24646 = ( ~n6630 & n24643 ) | ( ~n6630 & n24645 ) | ( n24643 & n24645 ) ;
  assign n24649 = n8487 | n10364 ;
  assign n24650 = n24649 ^ n16907 ^ 1'b0 ;
  assign n24651 = n2013 & ~n24650 ;
  assign n24647 = n20599 ^ n3608 ^ 1'b0 ;
  assign n24648 = n7732 | n24647 ;
  assign n24652 = n24651 ^ n24648 ^ n8304 ;
  assign n24658 = n8152 & ~n9560 ;
  assign n24659 = ~n2427 & n24658 ;
  assign n24653 = n5443 | n19552 ;
  assign n24654 = n9664 | n24653 ;
  assign n24655 = ~n10294 & n10362 ;
  assign n24656 = ( ~n730 & n8492 ) | ( ~n730 & n24655 ) | ( n8492 & n24655 ) ;
  assign n24657 = n24654 & ~n24656 ;
  assign n24660 = n24659 ^ n24657 ^ 1'b0 ;
  assign n24661 = n4182 & ~n9153 ;
  assign n24662 = n24661 ^ n22133 ^ n6997 ;
  assign n24663 = n24662 ^ n20053 ^ n8499 ;
  assign n24664 = n20587 ^ n7739 ^ n7521 ;
  assign n24668 = n7070 | n22472 ;
  assign n24669 = n24668 ^ n8527 ^ 1'b0 ;
  assign n24665 = n16530 ^ n500 ^ 1'b0 ;
  assign n24666 = ~n6645 & n24665 ;
  assign n24667 = n24666 ^ n13261 ^ 1'b0 ;
  assign n24670 = n24669 ^ n24667 ^ 1'b0 ;
  assign n24671 = n18876 & ~n24670 ;
  assign n24672 = n24671 ^ n20311 ^ n3436 ;
  assign n24673 = ( n20330 & n23931 ) | ( n20330 & n24672 ) | ( n23931 & n24672 ) ;
  assign n24674 = ( n3823 & ~n11742 ) | ( n3823 & n14481 ) | ( ~n11742 & n14481 ) ;
  assign n24675 = n2672 & ~n5744 ;
  assign n24676 = n24675 ^ n14892 ^ n9081 ;
  assign n24677 = n24676 ^ n5227 ^ 1'b0 ;
  assign n24680 = ( n10516 & n12119 ) | ( n10516 & n24342 ) | ( n12119 & n24342 ) ;
  assign n24678 = n5885 | n21741 ;
  assign n24679 = n10241 & ~n24678 ;
  assign n24681 = n24680 ^ n24679 ^ 1'b0 ;
  assign n24682 = n13974 ^ n5348 ^ n3293 ;
  assign n24683 = n21661 ^ n11459 ^ n8200 ;
  assign n24684 = ( n2680 & n24682 ) | ( n2680 & ~n24683 ) | ( n24682 & ~n24683 ) ;
  assign n24685 = n11944 ^ n6304 ^ 1'b0 ;
  assign n24686 = n4611 ^ n2427 ^ n2255 ;
  assign n24687 = n8703 ^ n5502 ^ 1'b0 ;
  assign n24688 = n24687 ^ n4819 ^ 1'b0 ;
  assign n24689 = ~n1912 & n24688 ;
  assign n24690 = n520 & n24689 ;
  assign n24693 = n9151 ^ n1340 ^ 1'b0 ;
  assign n24691 = n5465 ^ n3904 ^ 1'b0 ;
  assign n24692 = n460 & ~n24691 ;
  assign n24694 = n24693 ^ n24692 ^ n12062 ;
  assign n24695 = n2959 & ~n3899 ;
  assign n24696 = n24695 ^ n12170 ^ 1'b0 ;
  assign n24697 = ~n8854 & n24696 ;
  assign n24698 = ( ~n10799 & n18670 ) | ( ~n10799 & n20742 ) | ( n18670 & n20742 ) ;
  assign n24699 = n874 ^ n264 ^ 1'b0 ;
  assign n24700 = ~n10438 & n24699 ;
  assign n24701 = n24698 & n24700 ;
  assign n24704 = ~n3495 & n4802 ;
  assign n24705 = n24704 ^ n2722 ^ 1'b0 ;
  assign n24702 = ( ~n8667 & n10010 ) | ( ~n8667 & n12431 ) | ( n10010 & n12431 ) ;
  assign n24703 = ( n10835 & n21518 ) | ( n10835 & n24702 ) | ( n21518 & n24702 ) ;
  assign n24706 = n24705 ^ n24703 ^ n20295 ;
  assign n24708 = ~n14956 & n21914 ;
  assign n24709 = n24708 ^ n7917 ^ 1'b0 ;
  assign n24707 = n17811 & ~n23564 ;
  assign n24710 = n24709 ^ n24707 ^ 1'b0 ;
  assign n24711 = n17539 ^ n13665 ^ 1'b0 ;
  assign n24712 = n17246 & n24711 ;
  assign n24713 = ( n17600 & n20162 ) | ( n17600 & ~n24712 ) | ( n20162 & ~n24712 ) ;
  assign n24714 = ( n7013 & ~n8821 ) | ( n7013 & n11723 ) | ( ~n8821 & n11723 ) ;
  assign n24715 = n8498 | n15612 ;
  assign n24716 = n5284 | n24715 ;
  assign n24719 = n4359 & ~n5739 ;
  assign n24717 = ~n2561 & n10907 ;
  assign n24718 = n24717 ^ n17658 ^ 1'b0 ;
  assign n24720 = n24719 ^ n24718 ^ 1'b0 ;
  assign n24721 = n24716 & ~n24720 ;
  assign n24722 = ~n2560 & n4884 ;
  assign n24723 = ( n7434 & n10021 ) | ( n7434 & ~n17061 ) | ( n10021 & ~n17061 ) ;
  assign n24724 = ( n16642 & n24103 ) | ( n16642 & n24723 ) | ( n24103 & n24723 ) ;
  assign n24725 = ( n3101 & ~n24722 ) | ( n3101 & n24724 ) | ( ~n24722 & n24724 ) ;
  assign n24726 = n24721 & n24725 ;
  assign n24727 = n7259 ^ n4726 ^ 1'b0 ;
  assign n24728 = n16971 & n24727 ;
  assign n24730 = n20189 ^ n3954 ^ n2440 ;
  assign n24729 = x53 & n2123 ;
  assign n24731 = n24730 ^ n24729 ^ 1'b0 ;
  assign n24732 = ( n11609 & n23424 ) | ( n11609 & n24449 ) | ( n23424 & n24449 ) ;
  assign n24733 = n19580 ^ n19128 ^ n15787 ;
  assign n24734 = ( n13594 & n18521 ) | ( n13594 & n19945 ) | ( n18521 & n19945 ) ;
  assign n24735 = n9045 | n24734 ;
  assign n24736 = n24735 ^ n6859 ^ 1'b0 ;
  assign n24737 = ( n20531 & n23207 ) | ( n20531 & n23250 ) | ( n23207 & n23250 ) ;
  assign n24738 = ( n464 & ~n6484 ) | ( n464 & n13913 ) | ( ~n6484 & n13913 ) ;
  assign n24739 = n20432 & n24738 ;
  assign n24740 = n14933 | n24739 ;
  assign n24741 = n23136 ^ n1217 ^ 1'b0 ;
  assign n24742 = n15135 & ~n18755 ;
  assign n24743 = n24742 ^ n20942 ^ 1'b0 ;
  assign n24744 = n22609 ^ n8447 ^ 1'b0 ;
  assign n24745 = n10610 ^ n8955 ^ 1'b0 ;
  assign n24746 = n24745 ^ n7259 ^ n7062 ;
  assign n24747 = n1886 & ~n14188 ;
  assign n24748 = n24747 ^ n23885 ^ 1'b0 ;
  assign n24749 = ( ~n24744 & n24746 ) | ( ~n24744 & n24748 ) | ( n24746 & n24748 ) ;
  assign n24750 = ( n3472 & n6326 ) | ( n3472 & n15856 ) | ( n6326 & n15856 ) ;
  assign n24751 = ~n13188 & n24750 ;
  assign n24752 = ( ~n2451 & n5409 ) | ( ~n2451 & n15084 ) | ( n5409 & n15084 ) ;
  assign n24755 = n13515 ^ n12922 ^ 1'b0 ;
  assign n24756 = n7783 & n24755 ;
  assign n24753 = ~n15737 & n22245 ;
  assign n24754 = ~n3780 & n24753 ;
  assign n24757 = n24756 ^ n24754 ^ 1'b0 ;
  assign n24758 = n9871 | n12677 ;
  assign n24759 = n17455 ^ n3645 ^ 1'b0 ;
  assign n24760 = n10014 | n24759 ;
  assign n24761 = n20816 ^ n15185 ^ n9257 ;
  assign n24762 = n22698 ^ n18339 ^ 1'b0 ;
  assign n24763 = n19265 ^ n6610 ^ 1'b0 ;
  assign n24764 = n18593 & n24763 ;
  assign n24765 = n12315 & ~n17566 ;
  assign n24766 = ( n602 & ~n5427 ) | ( n602 & n8652 ) | ( ~n5427 & n8652 ) ;
  assign n24767 = n16604 ^ n3425 ^ n1274 ;
  assign n24768 = ( n719 & n6971 ) | ( n719 & ~n24767 ) | ( n6971 & ~n24767 ) ;
  assign n24769 = n19529 ^ n8301 ^ 1'b0 ;
  assign n24770 = n7122 & n24769 ;
  assign n24771 = ( n24336 & n24768 ) | ( n24336 & n24770 ) | ( n24768 & n24770 ) ;
  assign n24772 = n24771 ^ n15616 ^ n1236 ;
  assign n24773 = ( n13703 & n24766 ) | ( n13703 & ~n24772 ) | ( n24766 & ~n24772 ) ;
  assign n24774 = n6767 ^ n2891 ^ 1'b0 ;
  assign n24775 = n8085 & n24774 ;
  assign n24776 = ( n529 & ~n1671 ) | ( n529 & n24775 ) | ( ~n1671 & n24775 ) ;
  assign n24777 = n24776 ^ n16475 ^ 1'b0 ;
  assign n24778 = n6865 & ~n24777 ;
  assign n24779 = n24044 ^ n19106 ^ n12607 ;
  assign n24780 = n12238 | n18028 ;
  assign n24781 = n24779 & ~n24780 ;
  assign n24782 = ( n630 & n5569 ) | ( n630 & ~n16029 ) | ( n5569 & ~n16029 ) ;
  assign n24783 = n8036 & ~n23388 ;
  assign n24784 = ~n24782 & n24783 ;
  assign n24785 = n24784 ^ n9629 ^ n4776 ;
  assign n24786 = n5730 & ~n24785 ;
  assign n24787 = n24786 ^ n1866 ^ 1'b0 ;
  assign n24788 = n3485 ^ n2638 ^ n1598 ;
  assign n24789 = n21574 ^ n11584 ^ n5229 ;
  assign n24790 = ~n20397 & n24789 ;
  assign n24791 = n24790 ^ n22781 ^ 1'b0 ;
  assign n24792 = n10468 & n16529 ;
  assign n24793 = n7817 ^ n2634 ^ 1'b0 ;
  assign n24794 = ~n13377 & n24793 ;
  assign n24795 = n24792 & n24794 ;
  assign n24796 = n5392 & ~n12109 ;
  assign n24797 = ( ~n2020 & n3029 ) | ( ~n2020 & n5230 ) | ( n3029 & n5230 ) ;
  assign n24798 = n23888 ^ n23557 ^ n2470 ;
  assign n24799 = n24798 ^ n10871 ^ n8083 ;
  assign n24801 = n7070 ^ n3764 ^ 1'b0 ;
  assign n24800 = n3454 | n13025 ;
  assign n24802 = n24801 ^ n24800 ^ n14462 ;
  assign n24803 = n24802 ^ n19584 ^ n3781 ;
  assign n24804 = n24803 ^ n7578 ^ n2904 ;
  assign n24805 = n21518 ^ n8870 ^ 1'b0 ;
  assign n24806 = ~n4572 & n24805 ;
  assign n24807 = n16544 ^ n1365 ^ 1'b0 ;
  assign n24808 = n24806 & ~n24807 ;
  assign n24811 = n7928 & ~n13181 ;
  assign n24809 = n4466 & n9861 ;
  assign n24810 = n13667 | n24809 ;
  assign n24812 = n24811 ^ n24810 ^ n11608 ;
  assign n24813 = n17424 & ~n21668 ;
  assign n24814 = n24812 & ~n24813 ;
  assign n24815 = n16879 & n24814 ;
  assign n24821 = n1686 & n9340 ;
  assign n24822 = n5696 & n24821 ;
  assign n24816 = ( ~n805 & n3732 ) | ( ~n805 & n7842 ) | ( n3732 & n7842 ) ;
  assign n24817 = n22234 ^ n11205 ^ n8011 ;
  assign n24818 = ( n352 & n24816 ) | ( n352 & n24817 ) | ( n24816 & n24817 ) ;
  assign n24819 = ( n13713 & ~n22399 ) | ( n13713 & n24818 ) | ( ~n22399 & n24818 ) ;
  assign n24820 = n24819 ^ n12351 ^ 1'b0 ;
  assign n24823 = n24822 ^ n24820 ^ n7203 ;
  assign n24824 = n7489 ^ n1793 ^ 1'b0 ;
  assign n24825 = ~n24823 & n24824 ;
  assign n24826 = ( ~n1648 & n10927 ) | ( ~n1648 & n15612 ) | ( n10927 & n15612 ) ;
  assign n24827 = ( n12455 & n14260 ) | ( n12455 & ~n24826 ) | ( n14260 & ~n24826 ) ;
  assign n24837 = ( n3279 & ~n7235 ) | ( n3279 & n16016 ) | ( ~n7235 & n16016 ) ;
  assign n24838 = ~n17079 & n24837 ;
  assign n24835 = n3731 & ~n11824 ;
  assign n24836 = ~n11674 & n24835 ;
  assign n24828 = n19151 ^ n9230 ^ n4939 ;
  assign n24829 = ( ~n1452 & n17534 ) | ( ~n1452 & n24828 ) | ( n17534 & n24828 ) ;
  assign n24830 = n24829 ^ n14281 ^ n2048 ;
  assign n24831 = n1020 | n24830 ;
  assign n24832 = n24831 ^ n8983 ^ 1'b0 ;
  assign n24833 = n258 & ~n24832 ;
  assign n24834 = n24833 ^ n7254 ^ 1'b0 ;
  assign n24839 = n24838 ^ n24836 ^ n24834 ;
  assign n24840 = n6356 ^ n500 ^ 1'b0 ;
  assign n24841 = ( n1302 & n7629 ) | ( n1302 & ~n20670 ) | ( n7629 & ~n20670 ) ;
  assign n24842 = n21567 & n24841 ;
  assign n24843 = n24842 ^ n15420 ^ 1'b0 ;
  assign n24844 = n24843 ^ n23630 ^ n7563 ;
  assign n24845 = n7078 & n19798 ;
  assign n24846 = ( n1721 & ~n13712 ) | ( n1721 & n24845 ) | ( ~n13712 & n24845 ) ;
  assign n24847 = n5281 & ~n6762 ;
  assign n24848 = n24847 ^ n9010 ^ 1'b0 ;
  assign n24849 = ( n4356 & n24846 ) | ( n4356 & n24848 ) | ( n24846 & n24848 ) ;
  assign n24850 = n9116 | n24225 ;
  assign n24851 = n8609 | n24850 ;
  assign n24852 = n24851 ^ n22110 ^ 1'b0 ;
  assign n24853 = n2357 | n23867 ;
  assign n24854 = n3097 | n24853 ;
  assign n24855 = n4180 & ~n6398 ;
  assign n24856 = n7431 & n24855 ;
  assign n24857 = n5361 & n24856 ;
  assign n24858 = ( ~n7964 & n24854 ) | ( ~n7964 & n24857 ) | ( n24854 & n24857 ) ;
  assign n24859 = ( n2844 & n5773 ) | ( n2844 & n9438 ) | ( n5773 & n9438 ) ;
  assign n24860 = ~n4564 & n24553 ;
  assign n24861 = n7198 & n8066 ;
  assign n24862 = n24040 & n24861 ;
  assign n24863 = n24862 ^ n17905 ^ n11933 ;
  assign n24864 = ~n24860 & n24863 ;
  assign n24865 = n24864 ^ n18664 ^ 1'b0 ;
  assign n24866 = n24859 & ~n24865 ;
  assign n24867 = ( ~n7448 & n23979 ) | ( ~n7448 & n24508 ) | ( n23979 & n24508 ) ;
  assign n24868 = n19049 ^ n17908 ^ 1'b0 ;
  assign n24869 = n1910 & ~n24868 ;
  assign n24870 = n24869 ^ n16075 ^ 1'b0 ;
  assign n24871 = ~n2497 & n12585 ;
  assign n24872 = ~n5498 & n24871 ;
  assign n24873 = n18999 & ~n24872 ;
  assign n24874 = x96 & n1866 ;
  assign n24875 = n24874 ^ n17526 ^ n12116 ;
  assign n24876 = n24875 ^ n9606 ^ n5047 ;
  assign n24877 = ~n24873 & n24876 ;
  assign n24878 = ( n8210 & ~n11467 ) | ( n8210 & n13458 ) | ( ~n11467 & n13458 ) ;
  assign n24879 = ( n2874 & ~n12220 ) | ( n2874 & n24878 ) | ( ~n12220 & n24878 ) ;
  assign n24880 = n9739 & ~n24879 ;
  assign n24881 = n24880 ^ n6076 ^ 1'b0 ;
  assign n24882 = n6511 | n14215 ;
  assign n24883 = n24882 ^ n24129 ^ 1'b0 ;
  assign n24884 = n14657 & n22371 ;
  assign n24885 = n24884 ^ n18184 ^ 1'b0 ;
  assign n24886 = n18241 ^ n6323 ^ n5809 ;
  assign n24887 = n16924 ^ n6806 ^ 1'b0 ;
  assign n24888 = ( n10849 & ~n24886 ) | ( n10849 & n24887 ) | ( ~n24886 & n24887 ) ;
  assign n24889 = n23257 ^ n7700 ^ n2513 ;
  assign n24890 = ( n10240 & n15531 ) | ( n10240 & n21054 ) | ( n15531 & n21054 ) ;
  assign n24891 = n24890 ^ n17924 ^ 1'b0 ;
  assign n24893 = ( n7167 & n12487 ) | ( n7167 & ~n18710 ) | ( n12487 & ~n18710 ) ;
  assign n24892 = x184 & n14560 ;
  assign n24894 = n24893 ^ n24892 ^ 1'b0 ;
  assign n24895 = n18070 ^ n10207 ^ 1'b0 ;
  assign n24896 = ~n8213 & n24895 ;
  assign n24897 = n24896 ^ n8533 ^ 1'b0 ;
  assign n24898 = n6602 & n24897 ;
  assign n24899 = ~n24894 & n24898 ;
  assign n24900 = n24899 ^ n18704 ^ 1'b0 ;
  assign n24901 = n2348 | n8239 ;
  assign n24902 = n24901 ^ n23950 ^ n2391 ;
  assign n24903 = n12080 & ~n21741 ;
  assign n24904 = n23827 ^ n14996 ^ 1'b0 ;
  assign n24905 = ~n514 & n24904 ;
  assign n24906 = n9221 & ~n22158 ;
  assign n24907 = ( n18362 & ~n24905 ) | ( n18362 & n24906 ) | ( ~n24905 & n24906 ) ;
  assign n24908 = n8595 & n10921 ;
  assign n24909 = ~n24602 & n24908 ;
  assign n24910 = n19398 | n24909 ;
  assign n24911 = n24910 ^ n4046 ^ 1'b0 ;
  assign n24912 = n24911 ^ n21660 ^ n9637 ;
  assign n24915 = n18325 ^ n12562 ^ n9926 ;
  assign n24913 = n11724 ^ n8400 ^ n4024 ;
  assign n24914 = n24913 ^ n711 ^ 1'b0 ;
  assign n24916 = n24915 ^ n24914 ^ 1'b0 ;
  assign n24919 = ( ~n12190 & n17767 ) | ( ~n12190 & n19276 ) | ( n17767 & n19276 ) ;
  assign n24917 = ( n4552 & n7007 ) | ( n4552 & n18970 ) | ( n7007 & n18970 ) ;
  assign n24918 = n2891 & n24917 ;
  assign n24920 = n24919 ^ n24918 ^ 1'b0 ;
  assign n24921 = n17667 ^ n15981 ^ 1'b0 ;
  assign n24922 = n9916 & ~n13250 ;
  assign n24923 = ~n5905 & n8400 ;
  assign n24926 = n9684 ^ n812 ^ 1'b0 ;
  assign n24924 = n960 & ~n2793 ;
  assign n24925 = n24924 ^ n1049 ^ 1'b0 ;
  assign n24927 = n24926 ^ n24925 ^ n1408 ;
  assign n24928 = n13240 ^ n6483 ^ n5994 ;
  assign n24929 = ( ~n7627 & n8213 ) | ( ~n7627 & n24928 ) | ( n8213 & n24928 ) ;
  assign n24930 = ~n24927 & n24929 ;
  assign n24931 = n4857 & n17049 ;
  assign n24935 = n12177 & ~n20360 ;
  assign n24932 = ( n412 & n5827 ) | ( n412 & ~n11010 ) | ( n5827 & ~n11010 ) ;
  assign n24933 = ( ~n1994 & n2619 ) | ( ~n1994 & n24932 ) | ( n2619 & n24932 ) ;
  assign n24934 = n24933 ^ n9844 ^ 1'b0 ;
  assign n24936 = n24935 ^ n24934 ^ 1'b0 ;
  assign n24937 = ( n8889 & n13756 ) | ( n8889 & ~n16471 ) | ( n13756 & ~n16471 ) ;
  assign n24938 = n24045 & ~n24937 ;
  assign n24939 = n15406 ^ n7795 ^ n315 ;
  assign n24940 = n9606 ^ n2711 ^ 1'b0 ;
  assign n24941 = n16050 & n24940 ;
  assign n24942 = ( n793 & n8396 ) | ( n793 & ~n9265 ) | ( n8396 & ~n9265 ) ;
  assign n24943 = ( n8047 & ~n9739 ) | ( n8047 & n24942 ) | ( ~n9739 & n24942 ) ;
  assign n24944 = ( n9075 & ~n10010 ) | ( n9075 & n24943 ) | ( ~n10010 & n24943 ) ;
  assign n24945 = ( ~n10314 & n24941 ) | ( ~n10314 & n24944 ) | ( n24941 & n24944 ) ;
  assign n24946 = n24945 ^ n21344 ^ n7139 ;
  assign n24947 = n24946 ^ n6086 ^ n1306 ;
  assign n24949 = n1450 | n10941 ;
  assign n24950 = n19552 ^ n7136 ^ n1793 ;
  assign n24951 = ( n9665 & ~n24949 ) | ( n9665 & n24950 ) | ( ~n24949 & n24950 ) ;
  assign n24948 = n6544 ^ n3157 ^ 1'b0 ;
  assign n24952 = n24951 ^ n24948 ^ 1'b0 ;
  assign n24953 = n1415 & n24952 ;
  assign n24954 = n24953 ^ n11615 ^ n2398 ;
  assign n24955 = n15055 ^ n664 ^ 1'b0 ;
  assign n24956 = n376 | n24955 ;
  assign n24957 = ( ~n6916 & n8580 ) | ( ~n6916 & n14060 ) | ( n8580 & n14060 ) ;
  assign n24958 = ( ~n10052 & n14479 ) | ( ~n10052 & n24957 ) | ( n14479 & n24957 ) ;
  assign n24959 = ( ~n3080 & n9512 ) | ( ~n3080 & n12756 ) | ( n9512 & n12756 ) ;
  assign n24960 = n5278 ^ n1706 ^ 1'b0 ;
  assign n24961 = n7676 | n24960 ;
  assign n24962 = n20238 & ~n24961 ;
  assign n24963 = ~n24959 & n24962 ;
  assign n24967 = n8705 ^ n7506 ^ n7397 ;
  assign n24964 = n4239 & ~n17698 ;
  assign n24965 = n17530 & n24964 ;
  assign n24966 = n17144 | n24965 ;
  assign n24968 = n24967 ^ n24966 ^ 1'b0 ;
  assign n24969 = n20404 & ~n24968 ;
  assign n24970 = n19284 ^ n10545 ^ 1'b0 ;
  assign n24971 = n17863 ^ n15439 ^ 1'b0 ;
  assign n24972 = n24970 & ~n24971 ;
  assign n24973 = n24972 ^ n21101 ^ 1'b0 ;
  assign n24974 = n10497 ^ n9990 ^ 1'b0 ;
  assign n24975 = n22010 | n24974 ;
  assign n24976 = n24409 ^ n15744 ^ n9085 ;
  assign n24977 = n24976 ^ n6564 ^ 1'b0 ;
  assign n24978 = n7716 & n13077 ;
  assign n24979 = ~n2934 & n24978 ;
  assign n24980 = ( n16813 & n23239 ) | ( n16813 & n24979 ) | ( n23239 & n24979 ) ;
  assign n24981 = n24980 ^ n22919 ^ n10574 ;
  assign n24982 = ( n3515 & n16920 ) | ( n3515 & ~n24981 ) | ( n16920 & ~n24981 ) ;
  assign n24983 = n16307 ^ n15737 ^ n11331 ;
  assign n24984 = ~n293 & n4365 ;
  assign n24985 = n24984 ^ n1813 ^ 1'b0 ;
  assign n24986 = ( n5825 & ~n14967 ) | ( n5825 & n24985 ) | ( ~n14967 & n24985 ) ;
  assign n24987 = n24986 ^ n1881 ^ 1'b0 ;
  assign n24988 = n15276 ^ n15134 ^ n8274 ;
  assign n24989 = n24988 ^ n4169 ^ 1'b0 ;
  assign n24990 = ( n3884 & n13405 ) | ( n3884 & n24989 ) | ( n13405 & n24989 ) ;
  assign n24991 = n10854 ^ n6951 ^ 1'b0 ;
  assign n24992 = ~n5404 & n24991 ;
  assign n24993 = n24992 ^ n23440 ^ 1'b0 ;
  assign n24994 = n4475 & ~n15334 ;
  assign n24995 = n18605 | n24994 ;
  assign n24999 = n17440 ^ n13977 ^ n5624 ;
  assign n24996 = n17973 ^ n665 ^ n549 ;
  assign n24997 = n20653 & n24996 ;
  assign n24998 = n24997 ^ n4943 ^ 1'b0 ;
  assign n25000 = n24999 ^ n24998 ^ n9698 ;
  assign n25001 = ( n5328 & n7469 ) | ( n5328 & n17650 ) | ( n7469 & n17650 ) ;
  assign n25002 = ( n5217 & n13986 ) | ( n5217 & n25001 ) | ( n13986 & n25001 ) ;
  assign n25003 = ( n3500 & n3840 ) | ( n3500 & n11560 ) | ( n3840 & n11560 ) ;
  assign n25004 = ( n493 & n17410 ) | ( n493 & ~n25003 ) | ( n17410 & ~n25003 ) ;
  assign n25005 = ( n1894 & ~n2217 ) | ( n1894 & n25004 ) | ( ~n2217 & n25004 ) ;
  assign n25006 = n24130 ^ n8997 ^ 1'b0 ;
  assign n25007 = n20880 ^ n5587 ^ 1'b0 ;
  assign n25008 = n7789 & ~n9542 ;
  assign n25009 = n25008 ^ n10350 ^ 1'b0 ;
  assign n25010 = ( n3664 & ~n8770 ) | ( n3664 & n21410 ) | ( ~n8770 & n21410 ) ;
  assign n25011 = n19228 ^ n16480 ^ n8859 ;
  assign n25012 = ~n1133 & n13364 ;
  assign n25013 = n25012 ^ n1677 ^ 1'b0 ;
  assign n25014 = n25013 ^ n6120 ^ 1'b0 ;
  assign n25015 = n25014 ^ n22073 ^ n16297 ;
  assign n25016 = n20994 ^ n575 ^ 1'b0 ;
  assign n25017 = n25016 ^ n6365 ^ 1'b0 ;
  assign n25018 = ~n12589 & n25017 ;
  assign n25019 = n19843 ^ n19299 ^ 1'b0 ;
  assign n25020 = n25018 & n25019 ;
  assign n25021 = n8892 ^ n8380 ^ 1'b0 ;
  assign n25022 = n2797 & ~n25021 ;
  assign n25023 = n20339 ^ n10661 ^ 1'b0 ;
  assign n25024 = ( n16695 & n18822 ) | ( n16695 & ~n25023 ) | ( n18822 & ~n25023 ) ;
  assign n25025 = n8114 & ~n23545 ;
  assign n25026 = n25025 ^ x145 ^ 1'b0 ;
  assign n25027 = n2763 ^ n1736 ^ n1236 ;
  assign n25028 = n25027 ^ n13702 ^ n6625 ;
  assign n25029 = n25028 ^ n11220 ^ 1'b0 ;
  assign n25030 = ( n1284 & n4547 ) | ( n1284 & ~n13290 ) | ( n4547 & ~n13290 ) ;
  assign n25031 = n7091 & n19945 ;
  assign n25032 = n5762 & n25031 ;
  assign n25033 = n7985 & ~n25032 ;
  assign n25034 = ( n7680 & n25030 ) | ( n7680 & ~n25033 ) | ( n25030 & ~n25033 ) ;
  assign n25036 = ~n2810 & n8152 ;
  assign n25037 = n15250 & n25036 ;
  assign n25038 = n25037 ^ n10717 ^ n7157 ;
  assign n25035 = n14032 & n14394 ;
  assign n25039 = n25038 ^ n25035 ^ 1'b0 ;
  assign n25040 = n25039 ^ n3495 ^ 1'b0 ;
  assign n25044 = ( n7334 & ~n8983 ) | ( n7334 & n20405 ) | ( ~n8983 & n20405 ) ;
  assign n25041 = n6255 & n19535 ;
  assign n25042 = n25041 ^ n1474 ^ 1'b0 ;
  assign n25043 = ( n2353 & ~n9850 ) | ( n2353 & n25042 ) | ( ~n9850 & n25042 ) ;
  assign n25045 = n25044 ^ n25043 ^ n4897 ;
  assign n25048 = n15981 ^ n10804 ^ n5309 ;
  assign n25046 = ( n3217 & ~n5598 ) | ( n3217 & n23192 ) | ( ~n5598 & n23192 ) ;
  assign n25047 = n2222 & n25046 ;
  assign n25049 = n25048 ^ n25047 ^ n17264 ;
  assign n25050 = n15078 ^ n14583 ^ n3357 ;
  assign n25051 = n11705 & ~n25050 ;
  assign n25052 = n25051 ^ n3654 ^ 1'b0 ;
  assign n25053 = ( n11647 & ~n18992 ) | ( n11647 & n25052 ) | ( ~n18992 & n25052 ) ;
  assign n25054 = ~n1010 & n11226 ;
  assign n25055 = n25053 & n25054 ;
  assign n25056 = n4853 ^ n3557 ^ 1'b0 ;
  assign n25057 = x79 & ~n25056 ;
  assign n25058 = ( n3472 & n11343 ) | ( n3472 & ~n25057 ) | ( n11343 & ~n25057 ) ;
  assign n25059 = ( n17206 & n18508 ) | ( n17206 & ~n25058 ) | ( n18508 & ~n25058 ) ;
  assign n25060 = n3402 | n6236 ;
  assign n25061 = n25060 ^ n1148 ^ 1'b0 ;
  assign n25062 = n25061 ^ n5708 ^ 1'b0 ;
  assign n25063 = n25062 ^ n13888 ^ n10549 ;
  assign n25064 = n25059 & ~n25063 ;
  assign n25065 = n16084 & n25064 ;
  assign n25066 = n4210 ^ n2332 ^ 1'b0 ;
  assign n25067 = ~n8457 & n25066 ;
  assign n25068 = n25067 ^ n13436 ^ n364 ;
  assign n25069 = n992 & ~n4784 ;
  assign n25070 = ( n23301 & ~n25068 ) | ( n23301 & n25069 ) | ( ~n25068 & n25069 ) ;
  assign n25071 = ( n1304 & n5559 ) | ( n1304 & ~n12238 ) | ( n5559 & ~n12238 ) ;
  assign n25072 = n13123 ^ n10355 ^ 1'b0 ;
  assign n25073 = n18087 & ~n25072 ;
  assign n25074 = ( n10728 & ~n15443 ) | ( n10728 & n25073 ) | ( ~n15443 & n25073 ) ;
  assign n25075 = n21281 & n25074 ;
  assign n25076 = n25075 ^ n24441 ^ 1'b0 ;
  assign n25077 = n10907 & ~n16778 ;
  assign n25078 = ~n11217 & n25077 ;
  assign n25080 = n10045 ^ n8468 ^ 1'b0 ;
  assign n25081 = n7150 & ~n25080 ;
  assign n25079 = ( ~n5835 & n7674 ) | ( ~n5835 & n9417 ) | ( n7674 & n9417 ) ;
  assign n25082 = n25081 ^ n25079 ^ n9007 ;
  assign n25083 = ( ~n4782 & n6037 ) | ( ~n4782 & n12857 ) | ( n6037 & n12857 ) ;
  assign n25084 = ~n4128 & n17557 ;
  assign n25085 = n25084 ^ n3746 ^ 1'b0 ;
  assign n25086 = n20779 & n25085 ;
  assign n25087 = n14311 & n16228 ;
  assign n25088 = n12198 & n25087 ;
  assign n25089 = n679 ^ x221 ^ 1'b0 ;
  assign n25090 = n25088 | n25089 ;
  assign n25091 = n21409 ^ n14100 ^ n11972 ;
  assign n25092 = n9945 ^ n3397 ^ 1'b0 ;
  assign n25095 = ( n5723 & ~n11529 ) | ( n5723 & n11727 ) | ( ~n11529 & n11727 ) ;
  assign n25096 = ( n2061 & n7900 ) | ( n2061 & n25095 ) | ( n7900 & n25095 ) ;
  assign n25093 = ~n8442 & n18257 ;
  assign n25094 = n25093 ^ n20395 ^ n10267 ;
  assign n25097 = n25096 ^ n25094 ^ n15659 ;
  assign n25098 = ( n320 & n18235 ) | ( n320 & n25097 ) | ( n18235 & n25097 ) ;
  assign n25099 = ~n11905 & n19318 ;
  assign n25100 = n18929 & n25099 ;
  assign n25101 = n1278 | n1466 ;
  assign n25104 = n16386 ^ n1495 ^ 1'b0 ;
  assign n25102 = n20804 ^ n6247 ^ 1'b0 ;
  assign n25103 = n15411 | n25102 ;
  assign n25105 = n25104 ^ n25103 ^ n23381 ;
  assign n25106 = n24817 ^ n15994 ^ 1'b0 ;
  assign n25107 = n23797 ^ n8669 ^ n5976 ;
  assign n25108 = ( n3621 & n19954 ) | ( n3621 & n25107 ) | ( n19954 & n25107 ) ;
  assign n25109 = n25108 ^ n19378 ^ n10939 ;
  assign n25110 = ( n4265 & n8168 ) | ( n4265 & ~n25109 ) | ( n8168 & ~n25109 ) ;
  assign n25111 = ~n14577 & n16361 ;
  assign n25112 = ( x80 & n14710 ) | ( x80 & ~n25111 ) | ( n14710 & ~n25111 ) ;
  assign n25113 = n10777 ^ n9499 ^ 1'b0 ;
  assign n25114 = ~n4325 & n25113 ;
  assign n25115 = n25114 ^ n8595 ^ n5997 ;
  assign n25116 = ( n3169 & ~n7346 ) | ( n3169 & n20163 ) | ( ~n7346 & n20163 ) ;
  assign n25117 = n3037 | n12753 ;
  assign n25118 = n25117 ^ n2282 ^ 1'b0 ;
  assign n25119 = n7870 ^ n3784 ^ n1271 ;
  assign n25120 = n25119 ^ n18058 ^ n14418 ;
  assign n25121 = n12234 ^ n6789 ^ n2349 ;
  assign n25122 = ( ~n5227 & n15389 ) | ( ~n5227 & n22055 ) | ( n15389 & n22055 ) ;
  assign n25123 = ( n11794 & ~n16599 ) | ( n11794 & n25122 ) | ( ~n16599 & n25122 ) ;
  assign n25124 = ( n9134 & n10884 ) | ( n9134 & n25123 ) | ( n10884 & n25123 ) ;
  assign n25126 = n12042 ^ n11754 ^ 1'b0 ;
  assign n25127 = ~n17377 & n25126 ;
  assign n25125 = ~n4945 & n22613 ;
  assign n25128 = n25127 ^ n25125 ^ 1'b0 ;
  assign n25129 = n18410 ^ n5253 ^ 1'b0 ;
  assign n25130 = n25128 | n25129 ;
  assign n25133 = n7544 ^ n6585 ^ 1'b0 ;
  assign n25134 = ~n4244 & n25133 ;
  assign n25131 = n16570 ^ n13505 ^ n4480 ;
  assign n25132 = ( ~n8290 & n11954 ) | ( ~n8290 & n25131 ) | ( n11954 & n25131 ) ;
  assign n25135 = n25134 ^ n25132 ^ 1'b0 ;
  assign n25136 = n13132 & n25135 ;
  assign n25137 = ~n13807 & n25136 ;
  assign n25138 = n11286 & n25137 ;
  assign n25139 = n477 & ~n2272 ;
  assign n25140 = ( n12714 & n18242 ) | ( n12714 & n19984 ) | ( n18242 & n19984 ) ;
  assign n25141 = n4895 & n25140 ;
  assign n25142 = ~n2381 & n25141 ;
  assign n25145 = n19111 ^ n4437 ^ n3632 ;
  assign n25143 = n7442 & ~n9074 ;
  assign n25144 = n13408 | n25143 ;
  assign n25146 = n25145 ^ n25144 ^ 1'b0 ;
  assign n25147 = n9325 | n25146 ;
  assign n25148 = n19794 & ~n25147 ;
  assign n25149 = n3838 | n21794 ;
  assign n25150 = n4284 ^ n509 ^ 1'b0 ;
  assign n25151 = n5362 & ~n25150 ;
  assign n25152 = ~n25149 & n25151 ;
  assign n25153 = x138 & ~n11171 ;
  assign n25154 = ( n17811 & ~n20066 ) | ( n17811 & n25153 ) | ( ~n20066 & n25153 ) ;
  assign n25155 = n13990 & n14518 ;
  assign n25156 = n9604 & n19945 ;
  assign n25157 = n626 & n25156 ;
  assign n25158 = n12359 & ~n25157 ;
  assign n25159 = ( ~n10196 & n16587 ) | ( ~n10196 & n25158 ) | ( n16587 & n25158 ) ;
  assign n25164 = n21058 ^ n13627 ^ 1'b0 ;
  assign n25165 = ~n1803 & n25164 ;
  assign n25166 = ( ~n2623 & n14976 ) | ( ~n2623 & n25165 ) | ( n14976 & n25165 ) ;
  assign n25160 = n3754 ^ n2463 ^ 1'b0 ;
  assign n25161 = n25160 ^ n1046 ^ 1'b0 ;
  assign n25162 = n11488 | n25161 ;
  assign n25163 = ( n10361 & n22616 ) | ( n10361 & ~n25162 ) | ( n22616 & ~n25162 ) ;
  assign n25167 = n25166 ^ n25163 ^ n5896 ;
  assign n25168 = n20902 ^ n10695 ^ n1445 ;
  assign n25169 = n10645 ^ n9614 ^ 1'b0 ;
  assign n25170 = n18981 ^ n13330 ^ 1'b0 ;
  assign n25171 = n13436 | n25170 ;
  assign n25172 = ( n2086 & n5065 ) | ( n2086 & ~n10668 ) | ( n5065 & ~n10668 ) ;
  assign n25173 = n2276 | n10294 ;
  assign n25174 = n25173 ^ n8661 ^ 1'b0 ;
  assign n25175 = n19420 ^ n6458 ^ 1'b0 ;
  assign n25176 = n25174 & ~n25175 ;
  assign n25177 = n8025 & n25176 ;
  assign n25178 = n25172 & n25177 ;
  assign n25179 = ( n1821 & n2152 ) | ( n1821 & ~n20467 ) | ( n2152 & ~n20467 ) ;
  assign n25180 = ( ~n1419 & n8896 ) | ( ~n1419 & n25179 ) | ( n8896 & n25179 ) ;
  assign n25181 = n18707 | n19944 ;
  assign n25182 = n25181 ^ n3210 ^ 1'b0 ;
  assign n25183 = n5407 | n6536 ;
  assign n25184 = x114 | n25183 ;
  assign n25185 = n8163 ^ n3953 ^ n433 ;
  assign n25186 = n14873 & ~n25185 ;
  assign n25187 = n24553 ^ n10570 ^ 1'b0 ;
  assign n25188 = ( n1378 & n6926 ) | ( n1378 & ~n25187 ) | ( n6926 & ~n25187 ) ;
  assign n25189 = ( ~n10589 & n25186 ) | ( ~n10589 & n25188 ) | ( n25186 & n25188 ) ;
  assign n25190 = n372 & n20348 ;
  assign n25191 = n25190 ^ n20772 ^ 1'b0 ;
  assign n25192 = n16452 ^ n9938 ^ n5357 ;
  assign n25193 = n25192 ^ n15851 ^ n13385 ;
  assign n25194 = n25193 ^ n20382 ^ n3982 ;
  assign n25195 = n15330 & ~n25194 ;
  assign n25196 = ( n3910 & n5156 ) | ( n3910 & ~n5353 ) | ( n5156 & ~n5353 ) ;
  assign n25197 = n25196 ^ n17198 ^ n4450 ;
  assign n25198 = ( ~n1686 & n2967 ) | ( ~n1686 & n20976 ) | ( n2967 & n20976 ) ;
  assign n25199 = n25198 ^ n23054 ^ n12418 ;
  assign n25200 = ( n6883 & n25197 ) | ( n6883 & ~n25199 ) | ( n25197 & ~n25199 ) ;
  assign n25201 = n18428 & ~n25200 ;
  assign n25202 = n1928 & ~n13241 ;
  assign n25212 = ( x62 & n1236 ) | ( x62 & ~n8838 ) | ( n1236 & ~n8838 ) ;
  assign n25203 = n11634 & n15112 ;
  assign n25204 = ( ~n18863 & n21409 ) | ( ~n18863 & n25203 ) | ( n21409 & n25203 ) ;
  assign n25205 = n2080 | n10626 ;
  assign n25206 = n25205 ^ n810 ^ 1'b0 ;
  assign n25207 = n10124 ^ n4830 ^ 1'b0 ;
  assign n25208 = n5905 & ~n25207 ;
  assign n25209 = ( n569 & n25206 ) | ( n569 & n25208 ) | ( n25206 & n25208 ) ;
  assign n25210 = ( n5507 & n25204 ) | ( n5507 & ~n25209 ) | ( n25204 & ~n25209 ) ;
  assign n25211 = n22580 & n25210 ;
  assign n25213 = n25212 ^ n25211 ^ 1'b0 ;
  assign n25214 = n14303 ^ n5786 ^ 1'b0 ;
  assign n25215 = n25214 ^ n24915 ^ 1'b0 ;
  assign n25216 = n3339 & ~n25215 ;
  assign n25217 = n15491 & ~n17453 ;
  assign n25218 = n14586 ^ n13305 ^ n10979 ;
  assign n25219 = ( ~n13493 & n15169 ) | ( ~n13493 & n25218 ) | ( n15169 & n25218 ) ;
  assign n25220 = n25219 ^ n23537 ^ n10201 ;
  assign n25221 = ( n1220 & n1403 ) | ( n1220 & ~n6960 ) | ( n1403 & ~n6960 ) ;
  assign n25222 = n17297 & n25221 ;
  assign n25223 = n10724 & n13099 ;
  assign n25224 = n7991 & ~n10531 ;
  assign n25225 = n4772 | n16414 ;
  assign n25226 = n25224 & ~n25225 ;
  assign n25227 = n13429 ^ n7247 ^ n4050 ;
  assign n25228 = ~n4301 & n22381 ;
  assign n25229 = ( n4664 & ~n19121 ) | ( n4664 & n25228 ) | ( ~n19121 & n25228 ) ;
  assign n25230 = ( n9044 & n25227 ) | ( n9044 & ~n25229 ) | ( n25227 & ~n25229 ) ;
  assign n25231 = n25230 ^ n16935 ^ n550 ;
  assign n25232 = ( n979 & n22332 ) | ( n979 & n23852 ) | ( n22332 & n23852 ) ;
  assign n25233 = n25231 | n25232 ;
  assign n25234 = n11900 ^ n6923 ^ 1'b0 ;
  assign n25235 = n11633 & ~n25234 ;
  assign n25236 = n1189 | n15502 ;
  assign n25237 = n11513 & ~n18489 ;
  assign n25238 = ~n16965 & n25237 ;
  assign n25239 = ( ~n21642 & n22711 ) | ( ~n21642 & n25238 ) | ( n22711 & n25238 ) ;
  assign n25240 = n25239 ^ n11952 ^ n3518 ;
  assign n25242 = ( ~n17480 & n18169 ) | ( ~n17480 & n18696 ) | ( n18169 & n18696 ) ;
  assign n25241 = n21036 ^ n13277 ^ 1'b0 ;
  assign n25243 = n25242 ^ n25241 ^ 1'b0 ;
  assign n25244 = n17963 ^ n17169 ^ n10706 ;
  assign n25245 = n16462 ^ n12046 ^ n8215 ;
  assign n25246 = n25245 ^ n8241 ^ 1'b0 ;
  assign n25247 = n25246 ^ n14611 ^ n7836 ;
  assign n25248 = ( ~n4229 & n5369 ) | ( ~n4229 & n5881 ) | ( n5369 & n5881 ) ;
  assign n25249 = n4618 & n25248 ;
  assign n25250 = ( x123 & n1076 ) | ( x123 & n8266 ) | ( n1076 & n8266 ) ;
  assign n25251 = n11618 & n25250 ;
  assign n25252 = ( n8416 & n25249 ) | ( n8416 & ~n25251 ) | ( n25249 & ~n25251 ) ;
  assign n25253 = n4005 & ~n18174 ;
  assign n25254 = n25253 ^ n5924 ^ n5740 ;
  assign n25255 = n8309 & n10089 ;
  assign n25256 = n13070 ^ n8371 ^ 1'b0 ;
  assign n25257 = n15683 | n25256 ;
  assign n25258 = n24605 & ~n25257 ;
  assign n25259 = n289 & ~n25258 ;
  assign n25260 = n7746 ^ n6785 ^ n2538 ;
  assign n25261 = n3848 & n8157 ;
  assign n25262 = n25261 ^ n350 ^ 1'b0 ;
  assign n25263 = n11473 & ~n25262 ;
  assign n25264 = n25263 ^ n4263 ^ 1'b0 ;
  assign n25265 = n8032 & ~n25264 ;
  assign n25266 = n17557 & ~n23144 ;
  assign n25267 = ~n22829 & n25266 ;
  assign n25268 = n18713 & n25267 ;
  assign n25273 = n17905 ^ n4157 ^ n419 ;
  assign n25272 = ( ~n1101 & n9984 ) | ( ~n1101 & n14956 ) | ( n9984 & n14956 ) ;
  assign n25270 = n18421 ^ n11946 ^ n11310 ;
  assign n25269 = ~n15044 & n18062 ;
  assign n25271 = n25270 ^ n25269 ^ 1'b0 ;
  assign n25274 = n25273 ^ n25272 ^ n25271 ;
  assign n25275 = n10332 ^ n1419 ^ 1'b0 ;
  assign n25276 = ( n4351 & n24450 ) | ( n4351 & n25275 ) | ( n24450 & n25275 ) ;
  assign n25277 = ( ~n12761 & n15822 ) | ( ~n12761 & n23875 ) | ( n15822 & n23875 ) ;
  assign n25278 = n25276 | n25277 ;
  assign n25279 = x228 & n6758 ;
  assign n25280 = n25279 ^ n12927 ^ 1'b0 ;
  assign n25281 = n19080 ^ n5180 ^ 1'b0 ;
  assign n25282 = ( n8780 & n25280 ) | ( n8780 & n25281 ) | ( n25280 & n25281 ) ;
  assign n25283 = n16550 ^ n13208 ^ 1'b0 ;
  assign n25284 = n17739 ^ n14108 ^ n7601 ;
  assign n25285 = ( n13440 & ~n18736 ) | ( n13440 & n19517 ) | ( ~n18736 & n19517 ) ;
  assign n25286 = n5522 ^ n5268 ^ 1'b0 ;
  assign n25287 = n25286 ^ n16236 ^ n4358 ;
  assign n25288 = ( x156 & n1400 ) | ( x156 & n16870 ) | ( n1400 & n16870 ) ;
  assign n25289 = n24356 ^ n9252 ^ 1'b0 ;
  assign n25290 = n25042 & ~n25289 ;
  assign n25291 = n25290 ^ n24411 ^ 1'b0 ;
  assign n25292 = n9231 | n25291 ;
  assign n25294 = n24199 ^ n20246 ^ n12766 ;
  assign n25293 = ~n2782 & n3961 ;
  assign n25295 = n25294 ^ n25293 ^ 1'b0 ;
  assign n25296 = n7199 ^ n1507 ^ x19 ;
  assign n25297 = n5290 & ~n25296 ;
  assign n25298 = n19580 ^ n8972 ^ 1'b0 ;
  assign n25299 = ( ~n5710 & n7912 ) | ( ~n5710 & n25298 ) | ( n7912 & n25298 ) ;
  assign n25300 = ( n8658 & n12609 ) | ( n8658 & n25299 ) | ( n12609 & n25299 ) ;
  assign n25301 = n12870 & n25300 ;
  assign n25302 = ~n21982 & n23455 ;
  assign n25305 = n5700 ^ n4367 ^ 1'b0 ;
  assign n25306 = ( ~n15661 & n17439 ) | ( ~n15661 & n25305 ) | ( n17439 & n25305 ) ;
  assign n25307 = ~n21251 & n25306 ;
  assign n25303 = ( n10667 & ~n11044 ) | ( n10667 & n16435 ) | ( ~n11044 & n16435 ) ;
  assign n25304 = ( n8038 & ~n13272 ) | ( n8038 & n25303 ) | ( ~n13272 & n25303 ) ;
  assign n25308 = n25307 ^ n25304 ^ n21795 ;
  assign n25309 = ( n8297 & n10139 ) | ( n8297 & n23038 ) | ( n10139 & n23038 ) ;
  assign n25310 = n18955 ^ n17855 ^ 1'b0 ;
  assign n25311 = n11570 & ~n25310 ;
  assign n25312 = n14471 ^ n4403 ^ 1'b0 ;
  assign n25313 = n11552 & ~n25312 ;
  assign n25314 = n17042 ^ n15876 ^ 1'b0 ;
  assign n25315 = n8262 & n25314 ;
  assign n25316 = n25315 ^ n16354 ^ n1974 ;
  assign n25317 = n25313 & ~n25316 ;
  assign n25318 = ( n10770 & ~n17417 ) | ( n10770 & n20807 ) | ( ~n17417 & n20807 ) ;
  assign n25319 = ( ~n1606 & n17589 ) | ( ~n1606 & n23466 ) | ( n17589 & n23466 ) ;
  assign n25320 = n25318 & ~n25319 ;
  assign n25322 = ( ~n638 & n4696 ) | ( ~n638 & n13002 ) | ( n4696 & n13002 ) ;
  assign n25323 = n25322 ^ n679 ^ 1'b0 ;
  assign n25324 = ~n15230 & n25323 ;
  assign n25321 = n1297 | n11516 ;
  assign n25325 = n25324 ^ n25321 ^ 1'b0 ;
  assign n25326 = n2470 | n10827 ;
  assign n25327 = ( n5242 & ~n25325 ) | ( n5242 & n25326 ) | ( ~n25325 & n25326 ) ;
  assign n25328 = n10441 ^ n5533 ^ 1'b0 ;
  assign n25329 = ~n15812 & n25328 ;
  assign n25330 = ~n23416 & n25329 ;
  assign n25331 = n7721 & n25330 ;
  assign n25332 = ( ~n11415 & n11924 ) | ( ~n11415 & n25331 ) | ( n11924 & n25331 ) ;
  assign n25333 = ( ~n15378 & n25271 ) | ( ~n15378 & n25332 ) | ( n25271 & n25332 ) ;
  assign n25334 = ( n7195 & n8893 ) | ( n7195 & n14416 ) | ( n8893 & n14416 ) ;
  assign n25335 = ~n8290 & n24012 ;
  assign n25336 = n21676 ^ n4855 ^ n4224 ;
  assign n25337 = ( n10219 & ~n25335 ) | ( n10219 & n25336 ) | ( ~n25335 & n25336 ) ;
  assign n25338 = ~n25334 & n25337 ;
  assign n25339 = n25338 ^ n24518 ^ 1'b0 ;
  assign n25340 = n6236 | n25339 ;
  assign n25341 = n9534 ^ n8564 ^ 1'b0 ;
  assign n25342 = n17489 | n25341 ;
  assign n25343 = n11677 & ~n19175 ;
  assign n25344 = n25342 & n25343 ;
  assign n25345 = n8616 ^ n7836 ^ 1'b0 ;
  assign n25346 = ( n13990 & n14683 ) | ( n13990 & n25345 ) | ( n14683 & n25345 ) ;
  assign n25347 = ( n1894 & ~n17462 ) | ( n1894 & n25346 ) | ( ~n17462 & n25346 ) ;
  assign n25351 = n23758 ^ n6668 ^ 1'b0 ;
  assign n25348 = ( n792 & n6884 ) | ( n792 & ~n7214 ) | ( n6884 & ~n7214 ) ;
  assign n25349 = n849 & ~n6574 ;
  assign n25350 = n25348 & n25349 ;
  assign n25352 = n25351 ^ n25350 ^ 1'b0 ;
  assign n25353 = ~n2908 & n25352 ;
  assign n25354 = ( n12078 & n16654 ) | ( n12078 & n25353 ) | ( n16654 & n25353 ) ;
  assign n25355 = n25354 ^ n20177 ^ n2155 ;
  assign n25362 = n332 & n11258 ;
  assign n25363 = ~n8680 & n25362 ;
  assign n25364 = ( n957 & ~n22368 ) | ( n957 & n25363 ) | ( ~n22368 & n25363 ) ;
  assign n25356 = ( n3420 & n6014 ) | ( n3420 & n11663 ) | ( n6014 & n11663 ) ;
  assign n25357 = n3449 & ~n5150 ;
  assign n25358 = n1582 & n25357 ;
  assign n25359 = n25358 ^ n8644 ^ 1'b0 ;
  assign n25360 = n25359 ^ n23446 ^ n12744 ;
  assign n25361 = ( n4906 & ~n25356 ) | ( n4906 & n25360 ) | ( ~n25356 & n25360 ) ;
  assign n25365 = n25364 ^ n25361 ^ n2176 ;
  assign n25366 = ( n717 & ~n10707 ) | ( n717 & n13361 ) | ( ~n10707 & n13361 ) ;
  assign n25367 = n25365 & ~n25366 ;
  assign n25369 = n10533 ^ n8996 ^ n6174 ;
  assign n25370 = ( ~n5519 & n10408 ) | ( ~n5519 & n25369 ) | ( n10408 & n25369 ) ;
  assign n25368 = n2282 | n20802 ;
  assign n25371 = n25370 ^ n25368 ^ n24382 ;
  assign n25372 = n2803 | n25371 ;
  assign n25373 = ~n652 & n7705 ;
  assign n25374 = ~n22583 & n25373 ;
  assign n25375 = ( n5648 & n6369 ) | ( n5648 & ~n19001 ) | ( n6369 & ~n19001 ) ;
  assign n25376 = n949 | n6829 ;
  assign n25377 = n6471 | n25376 ;
  assign n25378 = n25377 ^ n16314 ^ 1'b0 ;
  assign n25379 = n25378 ^ n21638 ^ 1'b0 ;
  assign n25380 = n25379 ^ n12518 ^ 1'b0 ;
  assign n25381 = ~n6768 & n25380 ;
  assign n25382 = ~n25375 & n25381 ;
  assign n25383 = n25382 ^ n725 ^ 1'b0 ;
  assign n25384 = ( n5450 & n9175 ) | ( n5450 & n11296 ) | ( n9175 & n11296 ) ;
  assign n25385 = ( n1791 & n3649 ) | ( n1791 & ~n4601 ) | ( n3649 & ~n4601 ) ;
  assign n25386 = n6181 & ~n25385 ;
  assign n25387 = n25384 & n25386 ;
  assign n25388 = n19742 ^ n12705 ^ 1'b0 ;
  assign n25389 = n9464 | n25388 ;
  assign n25390 = x127 & ~n4006 ;
  assign n25391 = n25390 ^ n13795 ^ 1'b0 ;
  assign n25392 = n25391 ^ n12315 ^ n7201 ;
  assign n25393 = ( n11452 & ~n15785 ) | ( n11452 & n25392 ) | ( ~n15785 & n25392 ) ;
  assign n25394 = ~n2187 & n4464 ;
  assign n25395 = n25394 ^ n14757 ^ n11258 ;
  assign n25396 = n5190 ^ n2632 ^ n1572 ;
  assign n25397 = n25396 ^ n19111 ^ n10288 ;
  assign n25398 = n25397 ^ n585 ^ 1'b0 ;
  assign n25399 = ( n15990 & n24640 ) | ( n15990 & n24879 ) | ( n24640 & n24879 ) ;
  assign n25400 = n25399 ^ n17515 ^ n735 ;
  assign n25401 = n15139 & n18575 ;
  assign n25402 = n16789 & n25401 ;
  assign n25403 = ~n12977 & n15305 ;
  assign n25404 = n8807 ^ n7895 ^ n2288 ;
  assign n25405 = n25404 ^ n21386 ^ n2187 ;
  assign n25406 = n8725 ^ n6737 ^ 1'b0 ;
  assign n25407 = n6477 & ~n21694 ;
  assign n25408 = n12729 ^ n3449 ^ 1'b0 ;
  assign n25409 = ( n3525 & n12562 ) | ( n3525 & ~n25408 ) | ( n12562 & ~n25408 ) ;
  assign n25410 = n962 & n25176 ;
  assign n25412 = ( n4418 & ~n6622 ) | ( n4418 & n25196 ) | ( ~n6622 & n25196 ) ;
  assign n25411 = n18386 ^ n16577 ^ n8110 ;
  assign n25413 = n25412 ^ n25411 ^ 1'b0 ;
  assign n25414 = ( n3981 & n5142 ) | ( n3981 & n14462 ) | ( n5142 & n14462 ) ;
  assign n25415 = n25414 ^ n24182 ^ 1'b0 ;
  assign n25416 = ( n3635 & n5484 ) | ( n3635 & n21562 ) | ( n5484 & n21562 ) ;
  assign n25417 = n18970 & ~n25416 ;
  assign n25418 = n25417 ^ n24812 ^ 1'b0 ;
  assign n25419 = n10116 ^ n6039 ^ 1'b0 ;
  assign n25420 = n17678 ^ n1803 ^ 1'b0 ;
  assign n25421 = ~n3918 & n5328 ;
  assign n25422 = n25421 ^ n17658 ^ n12227 ;
  assign n25423 = ~n8897 & n25422 ;
  assign n25424 = ~n4583 & n25423 ;
  assign n25425 = ( ~n6456 & n25420 ) | ( ~n6456 & n25424 ) | ( n25420 & n25424 ) ;
  assign n25426 = ( n256 & n25419 ) | ( n256 & ~n25425 ) | ( n25419 & ~n25425 ) ;
  assign n25427 = n6403 & ~n8112 ;
  assign n25428 = ( n10801 & ~n12670 ) | ( n10801 & n25427 ) | ( ~n12670 & n25427 ) ;
  assign n25429 = n25428 ^ n16753 ^ n12236 ;
  assign n25432 = n5616 & n6934 ;
  assign n25433 = n23228 & n25432 ;
  assign n25430 = n1067 | n14972 ;
  assign n25431 = n10256 & ~n25430 ;
  assign n25434 = n25433 ^ n25431 ^ n8444 ;
  assign n25435 = n6983 & n25434 ;
  assign n25436 = n864 | n10769 ;
  assign n25437 = n8473 & ~n25436 ;
  assign n25438 = n9101 & ~n25437 ;
  assign n25439 = n12750 ^ n8799 ^ 1'b0 ;
  assign n25440 = n25438 & n25439 ;
  assign n25441 = ( n16960 & n23052 ) | ( n16960 & n25440 ) | ( n23052 & n25440 ) ;
  assign n25442 = n12247 ^ n4216 ^ n990 ;
  assign n25443 = n25442 ^ n9296 ^ 1'b0 ;
  assign n25444 = n25443 ^ n5472 ^ 1'b0 ;
  assign n25445 = n25444 ^ n1460 ^ 1'b0 ;
  assign n25446 = ( ~n4123 & n10210 ) | ( ~n4123 & n15576 ) | ( n10210 & n15576 ) ;
  assign n25447 = ( n7719 & ~n11538 ) | ( n7719 & n25446 ) | ( ~n11538 & n25446 ) ;
  assign n25448 = ( n751 & n2365 ) | ( n751 & n6815 ) | ( n2365 & n6815 ) ;
  assign n25449 = n25448 ^ x137 ^ 1'b0 ;
  assign n25450 = n10254 & n25449 ;
  assign n25451 = ~n7072 & n25450 ;
  assign n25452 = n13502 & n25451 ;
  assign n25453 = n25452 ^ n12275 ^ n1455 ;
  assign n25454 = n14619 & n15782 ;
  assign n25455 = ~n17690 & n25454 ;
  assign n25456 = n21487 ^ n16942 ^ n2498 ;
  assign n25457 = ( n9739 & n9814 ) | ( n9739 & ~n25456 ) | ( n9814 & ~n25456 ) ;
  assign n25458 = n1044 & n16457 ;
  assign n25459 = n25458 ^ n5891 ^ 1'b0 ;
  assign n25460 = ~n15644 & n19745 ;
  assign n25461 = n25460 ^ n21001 ^ 1'b0 ;
  assign n25462 = ( n8173 & n25459 ) | ( n8173 & ~n25461 ) | ( n25459 & ~n25461 ) ;
  assign n25463 = n12057 ^ n3743 ^ n2179 ;
  assign n25464 = ( ~x212 & n7277 ) | ( ~x212 & n16873 ) | ( n7277 & n16873 ) ;
  assign n25465 = n7196 ^ n3863 ^ 1'b0 ;
  assign n25466 = ( n9059 & n17150 ) | ( n9059 & n19877 ) | ( n17150 & n19877 ) ;
  assign n25467 = n12998 ^ n12485 ^ n7931 ;
  assign n25468 = n25467 ^ n20325 ^ 1'b0 ;
  assign n25469 = ( n8209 & n8744 ) | ( n8209 & ~n18865 ) | ( n8744 & ~n18865 ) ;
  assign n25470 = n13235 & ~n24888 ;
  assign n25471 = n10740 ^ n9983 ^ 1'b0 ;
  assign n25472 = n25471 ^ n25364 ^ n5670 ;
  assign n25473 = ( n8323 & n13004 ) | ( n8323 & n15261 ) | ( n13004 & n15261 ) ;
  assign n25474 = n3625 & n25473 ;
  assign n25475 = ( n20989 & n22171 ) | ( n20989 & n25474 ) | ( n22171 & n25474 ) ;
  assign n25476 = n10293 & n15883 ;
  assign n25477 = n25476 ^ n8484 ^ 1'b0 ;
  assign n25478 = n4985 | n11903 ;
  assign n25479 = n25478 ^ n12483 ^ 1'b0 ;
  assign n25480 = n3468 & ~n25479 ;
  assign n25481 = n419 & ~n8468 ;
  assign n25482 = n25481 ^ n11663 ^ n4298 ;
  assign n25483 = ( n4348 & ~n11827 ) | ( n4348 & n16230 ) | ( ~n11827 & n16230 ) ;
  assign n25484 = n25483 ^ n22267 ^ n20161 ;
  assign n25485 = n25484 ^ n22256 ^ 1'b0 ;
  assign n25486 = n9499 ^ n2428 ^ n469 ;
  assign n25487 = n10939 & n25486 ;
  assign n25488 = n15250 & n25487 ;
  assign n25489 = n1644 & ~n25488 ;
  assign n25490 = ~n3647 & n24905 ;
  assign n25491 = n24979 ^ n24241 ^ n2333 ;
  assign n25492 = n25491 ^ n6505 ^ 1'b0 ;
  assign n25493 = n25490 & ~n25492 ;
  assign n25501 = n14516 ^ n10475 ^ n1482 ;
  assign n25499 = ( n3078 & n5701 ) | ( n3078 & n6995 ) | ( n5701 & n6995 ) ;
  assign n25494 = n8621 ^ n6229 ^ n2952 ;
  assign n25495 = ( n5042 & n10991 ) | ( n5042 & n25494 ) | ( n10991 & n25494 ) ;
  assign n25496 = n7136 ^ n4003 ^ n2062 ;
  assign n25497 = ( ~n13626 & n17611 ) | ( ~n13626 & n25496 ) | ( n17611 & n25496 ) ;
  assign n25498 = n25495 & ~n25497 ;
  assign n25500 = n25499 ^ n25498 ^ 1'b0 ;
  assign n25502 = n25501 ^ n25500 ^ n8224 ;
  assign n25503 = n21258 ^ n7018 ^ n4884 ;
  assign n25504 = n25503 ^ n23549 ^ n16557 ;
  assign n25505 = n13528 & ~n14745 ;
  assign n25506 = ~n6938 & n25505 ;
  assign n25507 = n6314 | n25506 ;
  assign n25508 = n23112 ^ n16352 ^ 1'b0 ;
  assign n25509 = n16649 ^ n3430 ^ 1'b0 ;
  assign n25510 = ( n9652 & n9739 ) | ( n9652 & n18905 ) | ( n9739 & n18905 ) ;
  assign n25511 = n11875 ^ n9451 ^ 1'b0 ;
  assign n25512 = n1846 & ~n25511 ;
  assign n25513 = ~n8463 & n25512 ;
  assign n25518 = n13989 ^ n6948 ^ 1'b0 ;
  assign n25519 = n10862 & ~n25518 ;
  assign n25514 = ( ~n13634 & n18818 ) | ( ~n13634 & n25404 ) | ( n18818 & n25404 ) ;
  assign n25515 = n16034 ^ n10482 ^ n9731 ;
  assign n25516 = n25515 ^ n18887 ^ 1'b0 ;
  assign n25517 = ( n17275 & n25514 ) | ( n17275 & n25516 ) | ( n25514 & n25516 ) ;
  assign n25520 = n25519 ^ n25517 ^ n2313 ;
  assign n25523 = n6209 & ~n11666 ;
  assign n25524 = ( n5266 & n5646 ) | ( n5266 & ~n25523 ) | ( n5646 & ~n25523 ) ;
  assign n25521 = n12239 ^ n11083 ^ n7905 ;
  assign n25522 = ( n1977 & n13069 ) | ( n1977 & n25521 ) | ( n13069 & n25521 ) ;
  assign n25525 = n25524 ^ n25522 ^ 1'b0 ;
  assign n25526 = n25520 & ~n25525 ;
  assign n25527 = n3257 & n16586 ;
  assign n25528 = ~n19945 & n25527 ;
  assign n25529 = n25016 ^ n7629 ^ 1'b0 ;
  assign n25530 = n25528 | n25529 ;
  assign n25531 = n13200 ^ n7780 ^ 1'b0 ;
  assign n25532 = n21263 ^ n1504 ^ 1'b0 ;
  assign n25537 = n23090 ^ n11355 ^ n10244 ;
  assign n25533 = n4117 | n4622 ;
  assign n25534 = n25533 ^ n4063 ^ 1'b0 ;
  assign n25535 = n9969 & n25534 ;
  assign n25536 = n18665 & n25535 ;
  assign n25538 = n25537 ^ n25536 ^ n11727 ;
  assign n25541 = n1449 | n20976 ;
  assign n25539 = n7293 & n8105 ;
  assign n25540 = n25539 ^ n10281 ^ 1'b0 ;
  assign n25542 = n25541 ^ n25540 ^ 1'b0 ;
  assign n25543 = n25542 ^ n15975 ^ 1'b0 ;
  assign n25544 = n14821 | n25543 ;
  assign n25545 = ( n7259 & n7574 ) | ( n7259 & n17036 ) | ( n7574 & n17036 ) ;
  assign n25546 = n3267 ^ n604 ^ 1'b0 ;
  assign n25547 = n18156 & n25546 ;
  assign n25548 = n16251 ^ n7133 ^ n4458 ;
  assign n25549 = n25548 ^ n18647 ^ n7870 ;
  assign n25550 = n20273 & ~n25549 ;
  assign n25551 = n25550 ^ n17190 ^ 1'b0 ;
  assign n25552 = n20557 ^ n20262 ^ 1'b0 ;
  assign n25553 = n8816 | n22251 ;
  assign n25554 = n18647 & ~n25553 ;
  assign n25555 = n25554 ^ n12897 ^ 1'b0 ;
  assign n25556 = n5944 & ~n25555 ;
  assign n25557 = n10361 ^ n3705 ^ n2273 ;
  assign n25558 = ( n2426 & n11229 ) | ( n2426 & ~n25557 ) | ( n11229 & ~n25557 ) ;
  assign n25559 = n15825 ^ n13888 ^ n13171 ;
  assign n25565 = ~n652 & n12062 ;
  assign n25560 = n14781 ^ n8935 ^ 1'b0 ;
  assign n25561 = ~n11658 & n25560 ;
  assign n25562 = n25561 ^ n19905 ^ 1'b0 ;
  assign n25563 = n7449 & n25562 ;
  assign n25564 = n25563 ^ n4638 ^ n500 ;
  assign n25566 = n25565 ^ n25564 ^ n7139 ;
  assign n25567 = ( n773 & ~n1703 ) | ( n773 & n19515 ) | ( ~n1703 & n19515 ) ;
  assign n25568 = n20619 & ~n25567 ;
  assign n25569 = n25568 ^ n12464 ^ 1'b0 ;
  assign n25570 = n14622 & ~n25569 ;
  assign n25571 = n5281 | n25570 ;
  assign n25572 = ~n4922 & n13678 ;
  assign n25573 = n13218 ^ n6437 ^ n5832 ;
  assign n25574 = n18328 ^ n7926 ^ n4491 ;
  assign n25575 = n25573 | n25574 ;
  assign n25576 = n25575 ^ n19615 ^ 1'b0 ;
  assign n25577 = ~n2059 & n25576 ;
  assign n25581 = n18543 ^ n2734 ^ n1326 ;
  assign n25578 = ( ~n4884 & n10200 ) | ( ~n4884 & n17179 ) | ( n10200 & n17179 ) ;
  assign n25579 = ( n690 & ~n20095 ) | ( n690 & n25578 ) | ( ~n20095 & n25578 ) ;
  assign n25580 = n25579 ^ n506 ^ 1'b0 ;
  assign n25582 = n25581 ^ n25580 ^ n23077 ;
  assign n25583 = n13450 | n15022 ;
  assign n25589 = n9693 ^ n8313 ^ 1'b0 ;
  assign n25587 = ( ~n4376 & n19792 ) | ( ~n4376 & n22616 ) | ( n19792 & n22616 ) ;
  assign n25584 = ( ~n456 & n7822 ) | ( ~n456 & n8169 ) | ( n7822 & n8169 ) ;
  assign n25585 = ~n447 & n892 ;
  assign n25586 = n25584 & n25585 ;
  assign n25588 = n25587 ^ n25586 ^ 1'b0 ;
  assign n25590 = n25589 ^ n25588 ^ n2271 ;
  assign n25591 = n6522 & n19581 ;
  assign n25592 = n25591 ^ n15654 ^ 1'b0 ;
  assign n25593 = n21023 ^ n19713 ^ n15608 ;
  assign n25594 = n14278 ^ n13041 ^ x186 ;
  assign n25595 = n25594 ^ n4975 ^ 1'b0 ;
  assign n25596 = ( ~n8480 & n14219 ) | ( ~n8480 & n22253 ) | ( n14219 & n22253 ) ;
  assign n25597 = ( n5416 & n20516 ) | ( n5416 & ~n25596 ) | ( n20516 & ~n25596 ) ;
  assign n25598 = n25597 ^ n16138 ^ 1'b0 ;
  assign n25599 = n12983 ^ n6957 ^ n6322 ;
  assign n25600 = n6698 & n7492 ;
  assign n25601 = n1131 & n25600 ;
  assign n25602 = ( n17361 & n25599 ) | ( n17361 & n25601 ) | ( n25599 & n25601 ) ;
  assign n25603 = ( n5820 & ~n7834 ) | ( n5820 & n8257 ) | ( ~n7834 & n8257 ) ;
  assign n25604 = n15496 ^ n14193 ^ n10125 ;
  assign n25605 = ( n8980 & n25603 ) | ( n8980 & ~n25604 ) | ( n25603 & ~n25604 ) ;
  assign n25606 = n25605 ^ n19681 ^ 1'b0 ;
  assign n25607 = n18084 ^ n3309 ^ n1766 ;
  assign n25608 = n8857 ^ n3490 ^ 1'b0 ;
  assign n25609 = ~n5368 & n25608 ;
  assign n25610 = n1734 | n25609 ;
  assign n25611 = ( n11393 & n19748 ) | ( n11393 & n25392 ) | ( n19748 & n25392 ) ;
  assign n25612 = ( n25607 & ~n25610 ) | ( n25607 & n25611 ) | ( ~n25610 & n25611 ) ;
  assign n25613 = ( n5202 & n20053 ) | ( n5202 & ~n23238 ) | ( n20053 & ~n23238 ) ;
  assign n25614 = n19450 & ~n25613 ;
  assign n25615 = ~n25612 & n25614 ;
  assign n25619 = n13314 ^ n9455 ^ 1'b0 ;
  assign n25616 = n15542 ^ n14868 ^ n6563 ;
  assign n25617 = ( n1485 & n10131 ) | ( n1485 & n12509 ) | ( n10131 & n12509 ) ;
  assign n25618 = ( ~n15245 & n25616 ) | ( ~n15245 & n25617 ) | ( n25616 & n25617 ) ;
  assign n25620 = n25619 ^ n25618 ^ n19398 ;
  assign n25622 = n10356 & n23959 ;
  assign n25623 = n25622 ^ n8725 ^ n6411 ;
  assign n25621 = ( n4119 & n12394 ) | ( n4119 & ~n16137 ) | ( n12394 & ~n16137 ) ;
  assign n25624 = n25623 ^ n25621 ^ n2327 ;
  assign n25625 = n19555 ^ n13738 ^ 1'b0 ;
  assign n25626 = n16475 ^ n3820 ^ 1'b0 ;
  assign n25627 = ~n9263 & n25626 ;
  assign n25628 = n25627 ^ n491 ^ 1'b0 ;
  assign n25629 = n1887 & ~n5305 ;
  assign n25630 = n25629 ^ n3333 ^ 1'b0 ;
  assign n25631 = n7985 | n25630 ;
  assign n25632 = n11927 & n25631 ;
  assign n25633 = n25632 ^ n3139 ^ 1'b0 ;
  assign n25634 = ( n1510 & n25628 ) | ( n1510 & ~n25633 ) | ( n25628 & ~n25633 ) ;
  assign n25635 = n22289 ^ n14827 ^ 1'b0 ;
  assign n25636 = n824 & ~n25635 ;
  assign n25637 = ( n8026 & n25634 ) | ( n8026 & n25636 ) | ( n25634 & n25636 ) ;
  assign n25643 = ( n2729 & ~n13372 ) | ( n2729 & n19762 ) | ( ~n13372 & n19762 ) ;
  assign n25644 = n15449 & n25643 ;
  assign n25645 = ~n9869 & n25644 ;
  assign n25638 = ( n10751 & ~n11472 ) | ( n10751 & n12872 ) | ( ~n11472 & n12872 ) ;
  assign n25639 = n23486 ^ n3142 ^ 1'b0 ;
  assign n25640 = n25638 & n25639 ;
  assign n25641 = n9875 & n25640 ;
  assign n25642 = n16970 & n25641 ;
  assign n25646 = n25645 ^ n25642 ^ n15569 ;
  assign n25647 = n10327 ^ n397 ^ 1'b0 ;
  assign n25648 = n4652 & n22223 ;
  assign n25649 = n25648 ^ n9305 ^ 1'b0 ;
  assign n25650 = n4449 & ~n10627 ;
  assign n25651 = n11867 & ~n25650 ;
  assign n25652 = n25651 ^ n2317 ^ x66 ;
  assign n25653 = ( n11645 & ~n17661 ) | ( n11645 & n22216 ) | ( ~n17661 & n22216 ) ;
  assign n25654 = ( n22220 & ~n23101 ) | ( n22220 & n25653 ) | ( ~n23101 & n25653 ) ;
  assign n25655 = n25654 ^ n21843 ^ n1164 ;
  assign n25656 = ~n2050 & n9655 ;
  assign n25657 = n2357 & n25656 ;
  assign n25658 = ( n13495 & ~n18775 ) | ( n13495 & n25657 ) | ( ~n18775 & n25657 ) ;
  assign n25659 = n25658 ^ n10049 ^ 1'b0 ;
  assign n25660 = n2605 | n19818 ;
  assign n25661 = n20953 & ~n25660 ;
  assign n25662 = n25661 ^ n13804 ^ n10546 ;
  assign n25663 = ~n12244 & n20508 ;
  assign n25664 = n23015 & ~n25663 ;
  assign n25665 = n17120 & n25664 ;
  assign n25666 = ( n6567 & ~n10843 ) | ( n6567 & n18129 ) | ( ~n10843 & n18129 ) ;
  assign n25667 = n25666 ^ n20386 ^ n7556 ;
  assign n25668 = n7878 & n25667 ;
  assign n25669 = ~n3340 & n25668 ;
  assign n25670 = ( ~n16160 & n19051 ) | ( ~n16160 & n25534 ) | ( n19051 & n25534 ) ;
  assign n25671 = ~n8402 & n15836 ;
  assign n25672 = n25670 & n25671 ;
  assign n25673 = ( n697 & n18318 ) | ( n697 & ~n25672 ) | ( n18318 & ~n25672 ) ;
  assign n25674 = n3643 | n4764 ;
  assign n25675 = n25674 ^ n22079 ^ n1643 ;
  assign n25676 = ~n13041 & n17327 ;
  assign n25677 = ~n12759 & n25676 ;
  assign n25678 = n23888 ^ n8733 ^ 1'b0 ;
  assign n25679 = ~n25677 & n25678 ;
  assign n25680 = ~n1025 & n19423 ;
  assign n25681 = n25680 ^ n1760 ^ 1'b0 ;
  assign n25682 = n9669 ^ n943 ^ 1'b0 ;
  assign n25683 = n25681 & ~n25682 ;
  assign n25684 = n25456 ^ n18020 ^ n10785 ;
  assign n25685 = n3367 & ~n4884 ;
  assign n25686 = n9697 & n25685 ;
  assign n25687 = n25686 ^ n10955 ^ 1'b0 ;
  assign n25688 = ( n2250 & ~n25684 ) | ( n2250 & n25687 ) | ( ~n25684 & n25687 ) ;
  assign n25691 = n13778 ^ n5323 ^ n3860 ;
  assign n25692 = n7743 & ~n23137 ;
  assign n25693 = n25691 & n25692 ;
  assign n25689 = n18752 ^ n2404 ^ 1'b0 ;
  assign n25690 = ( n9985 & ~n21820 ) | ( n9985 & n25689 ) | ( ~n21820 & n25689 ) ;
  assign n25694 = n25693 ^ n25690 ^ n4717 ;
  assign n25695 = n7405 & ~n25694 ;
  assign n25696 = n17143 ^ n2992 ^ 1'b0 ;
  assign n25697 = n12594 ^ n8423 ^ 1'b0 ;
  assign n25698 = n3985 | n25697 ;
  assign n25699 = n25698 ^ n7471 ^ n381 ;
  assign n25700 = n25699 ^ n12860 ^ 1'b0 ;
  assign n25701 = ( n12377 & n17340 ) | ( n12377 & ~n25700 ) | ( n17340 & ~n25700 ) ;
  assign n25702 = n7780 ^ n5014 ^ n833 ;
  assign n25703 = ~n23653 & n25702 ;
  assign n25704 = n25703 ^ x126 ^ 1'b0 ;
  assign n25711 = n17283 & ~n17539 ;
  assign n25712 = n24270 ^ n15941 ^ 1'b0 ;
  assign n25713 = n25711 & n25712 ;
  assign n25705 = n15676 ^ n13274 ^ n10010 ;
  assign n25706 = n3182 | n3421 ;
  assign n25707 = n25706 ^ n9221 ^ 1'b0 ;
  assign n25708 = n16071 | n25707 ;
  assign n25709 = n25705 | n25708 ;
  assign n25710 = n20882 & n25709 ;
  assign n25714 = n25713 ^ n25710 ^ 1'b0 ;
  assign n25715 = n15413 ^ n4759 ^ n1279 ;
  assign n25716 = n25715 ^ n5804 ^ 1'b0 ;
  assign n25717 = n1419 & ~n25716 ;
  assign n25718 = ~n2291 & n25717 ;
  assign n25719 = n25718 ^ n24852 ^ n20488 ;
  assign n25720 = ( n4493 & ~n17889 ) | ( n4493 & n18008 ) | ( ~n17889 & n18008 ) ;
  assign n25721 = n15326 & ~n16024 ;
  assign n25722 = n25721 ^ n3203 ^ 1'b0 ;
  assign n25725 = n19599 ^ n9758 ^ n6709 ;
  assign n25726 = n17540 | n18239 ;
  assign n25727 = n25725 | n25726 ;
  assign n25723 = ( n3583 & n13974 ) | ( n3583 & n17468 ) | ( n13974 & n17468 ) ;
  assign n25724 = ~n13623 & n25723 ;
  assign n25728 = n25727 ^ n25724 ^ 1'b0 ;
  assign n25729 = n11215 | n18098 ;
  assign n25730 = n13962 ^ n1827 ^ 1'b0 ;
  assign n25731 = ( n3962 & n9723 ) | ( n3962 & ~n22368 ) | ( n9723 & ~n22368 ) ;
  assign n25732 = n18180 ^ n5354 ^ n2298 ;
  assign n25733 = n25732 ^ n20816 ^ 1'b0 ;
  assign n25734 = n16430 ^ x78 ^ 1'b0 ;
  assign n25735 = n887 & n25734 ;
  assign n25736 = n25735 ^ n6661 ^ 1'b0 ;
  assign n25737 = n6961 | n23297 ;
  assign n25738 = n3357 & n3545 ;
  assign n25739 = n2809 | n13006 ;
  assign n25740 = n13249 | n25739 ;
  assign n25741 = ( n3090 & n25738 ) | ( n3090 & n25740 ) | ( n25738 & n25740 ) ;
  assign n25742 = n25741 ^ n12083 ^ n4965 ;
  assign n25743 = n25742 ^ n21712 ^ n4990 ;
  assign n25744 = ~n25737 & n25743 ;
  assign n25745 = n21930 & n25744 ;
  assign n25749 = ~n2937 & n19051 ;
  assign n25746 = ( n3798 & ~n12156 ) | ( n3798 & n14220 ) | ( ~n12156 & n14220 ) ;
  assign n25747 = ~n6074 & n25746 ;
  assign n25748 = n25747 ^ n24258 ^ 1'b0 ;
  assign n25750 = n25749 ^ n25748 ^ n401 ;
  assign n25753 = n8836 & ~n12198 ;
  assign n25754 = n25753 ^ n15546 ^ 1'b0 ;
  assign n25751 = n14393 ^ n8060 ^ 1'b0 ;
  assign n25752 = ( n17216 & n19511 ) | ( n17216 & n25751 ) | ( n19511 & n25751 ) ;
  assign n25755 = n25754 ^ n25752 ^ n10751 ;
  assign n25756 = n22859 ^ n7294 ^ 1'b0 ;
  assign n25757 = n10510 ^ n4312 ^ 1'b0 ;
  assign n25758 = n20369 ^ n16066 ^ n9108 ;
  assign n25763 = n2113 | n6198 ;
  assign n25760 = n8536 & ~n14823 ;
  assign n25761 = n25760 ^ n5231 ^ 1'b0 ;
  assign n25759 = ( ~n5875 & n7128 ) | ( ~n5875 & n11828 ) | ( n7128 & n11828 ) ;
  assign n25762 = n25761 ^ n25759 ^ n7464 ;
  assign n25764 = n25763 ^ n25762 ^ n5333 ;
  assign n25765 = ( n1182 & n9064 ) | ( n1182 & n25764 ) | ( n9064 & n25764 ) ;
  assign n25766 = x127 & n22268 ;
  assign n25767 = n14431 & ~n20670 ;
  assign n25768 = ~n25766 & n25767 ;
  assign n25772 = n8886 ^ n5685 ^ n1899 ;
  assign n25773 = n25772 ^ n24785 ^ 1'b0 ;
  assign n25774 = n4160 | n25773 ;
  assign n25769 = ( n6216 & n7464 ) | ( n6216 & ~n18653 ) | ( n7464 & ~n18653 ) ;
  assign n25770 = n8128 ^ n6048 ^ n1771 ;
  assign n25771 = n25769 | n25770 ;
  assign n25775 = n25774 ^ n25771 ^ 1'b0 ;
  assign n25776 = ( n10382 & n25768 ) | ( n10382 & n25775 ) | ( n25768 & n25775 ) ;
  assign n25777 = n9973 ^ x37 ^ 1'b0 ;
  assign n25778 = n25777 ^ n9556 ^ n6336 ;
  assign n25779 = n23064 ^ n15973 ^ 1'b0 ;
  assign n25780 = ( n5809 & ~n19058 ) | ( n5809 & n24942 ) | ( ~n19058 & n24942 ) ;
  assign n25781 = n14593 ^ n1476 ^ n432 ;
  assign n25782 = x168 & n25781 ;
  assign n25783 = n25780 & ~n25782 ;
  assign n25784 = n25779 & n25783 ;
  assign n25785 = ~n4045 & n11099 ;
  assign n25786 = n2652 & n25785 ;
  assign n25787 = ( n6083 & ~n24576 ) | ( n6083 & n25786 ) | ( ~n24576 & n25786 ) ;
  assign n25788 = n697 & n23730 ;
  assign n25789 = ( n2470 & n4924 ) | ( n2470 & ~n4958 ) | ( n4924 & ~n4958 ) ;
  assign n25790 = n19067 ^ n781 ^ 1'b0 ;
  assign n25791 = n9084 & n25790 ;
  assign n25792 = ( n14648 & n22408 ) | ( n14648 & ~n25791 ) | ( n22408 & ~n25791 ) ;
  assign n25793 = ( ~n1160 & n25789 ) | ( ~n1160 & n25792 ) | ( n25789 & n25792 ) ;
  assign n25796 = n4929 ^ n4136 ^ n2652 ;
  assign n25797 = ( n2575 & n6408 ) | ( n2575 & ~n25796 ) | ( n6408 & ~n25796 ) ;
  assign n25794 = n6971 & ~n22632 ;
  assign n25795 = ( n5589 & n12291 ) | ( n5589 & n25794 ) | ( n12291 & n25794 ) ;
  assign n25798 = n25797 ^ n25795 ^ n4441 ;
  assign n25799 = n7410 ^ n6553 ^ n332 ;
  assign n25800 = n25799 ^ n25104 ^ n23010 ;
  assign n25801 = n25800 ^ n25517 ^ n16064 ;
  assign n25802 = n1887 & n11534 ;
  assign n25803 = ( n4277 & ~n10535 ) | ( n4277 & n11198 ) | ( ~n10535 & n11198 ) ;
  assign n25804 = ( ~n9788 & n19886 ) | ( ~n9788 & n25803 ) | ( n19886 & n25803 ) ;
  assign n25805 = ( n3103 & ~n24594 ) | ( n3103 & n25804 ) | ( ~n24594 & n25804 ) ;
  assign n25806 = n10920 ^ n8599 ^ 1'b0 ;
  assign n25807 = n9159 | n25806 ;
  assign n25808 = n13738 ^ n4310 ^ 1'b0 ;
  assign n25809 = n25807 | n25808 ;
  assign n25810 = n25805 & ~n25809 ;
  assign n25811 = n14967 & n19765 ;
  assign n25812 = n25811 ^ n11083 ^ 1'b0 ;
  assign n25813 = n8384 & n8619 ;
  assign n25814 = n513 & ~n6168 ;
  assign n25815 = ~n24338 & n25814 ;
  assign n25816 = n3549 & ~n4552 ;
  assign n25817 = n25816 ^ n23035 ^ n9281 ;
  assign n25818 = n3075 | n24605 ;
  assign n25819 = n25818 ^ n11370 ^ n10260 ;
  assign n25820 = n15345 | n25819 ;
  assign n25821 = n25820 ^ n20442 ^ 1'b0 ;
  assign n25822 = n6611 ^ n530 ^ 1'b0 ;
  assign n25823 = n1748 & ~n25822 ;
  assign n25824 = n25823 ^ x218 ^ 1'b0 ;
  assign n25825 = n25824 ^ n13527 ^ n2637 ;
  assign n25826 = n3113 ^ n739 ^ 1'b0 ;
  assign n25827 = n20398 ^ n17150 ^ n3348 ;
  assign n25828 = ~n4227 & n25827 ;
  assign n25829 = n2340 & ~n9415 ;
  assign n25830 = ( ~n1884 & n21522 ) | ( ~n1884 & n25829 ) | ( n21522 & n25829 ) ;
  assign n25831 = n18686 ^ n14023 ^ n11229 ;
  assign n25832 = n21373 ^ n5184 ^ 1'b0 ;
  assign n25833 = n15086 ^ n1228 ^ 1'b0 ;
  assign n25834 = n25833 ^ n17767 ^ n17225 ;
  assign n25835 = n25834 ^ n19601 ^ n4896 ;
  assign n25836 = n6662 | n14178 ;
  assign n25837 = n25836 ^ n560 ^ 1'b0 ;
  assign n25845 = n18421 ^ n7702 ^ n2914 ;
  assign n25839 = n11892 ^ n4082 ^ n1455 ;
  assign n25838 = n1455 | n15863 ;
  assign n25840 = n25839 ^ n25838 ^ 1'b0 ;
  assign n25841 = ~n6056 & n9025 ;
  assign n25842 = n8753 & n25841 ;
  assign n25843 = n25840 & n25842 ;
  assign n25844 = n15027 | n25843 ;
  assign n25846 = n25845 ^ n25844 ^ 1'b0 ;
  assign n25847 = n17574 ^ n7449 ^ 1'b0 ;
  assign n25849 = ( n7106 & n7390 ) | ( n7106 & n23598 ) | ( n7390 & n23598 ) ;
  assign n25850 = n12373 ^ n7622 ^ 1'b0 ;
  assign n25851 = n14859 | n25850 ;
  assign n25852 = n25849 & ~n25851 ;
  assign n25853 = n1785 & n25852 ;
  assign n25848 = n6007 & n23324 ;
  assign n25854 = n25853 ^ n25848 ^ n13157 ;
  assign n25855 = ( n2009 & n3182 ) | ( n2009 & n9993 ) | ( n3182 & n9993 ) ;
  assign n25856 = n25855 ^ n1895 ^ 1'b0 ;
  assign n25857 = ~n19441 & n25856 ;
  assign n25858 = n2832 & n3073 ;
  assign n25859 = ~n3073 & n25858 ;
  assign n25860 = n591 & ~n25859 ;
  assign n25861 = ~n591 & n25860 ;
  assign n25862 = n5294 | n25861 ;
  assign n25863 = n18893 & ~n25862 ;
  assign n25864 = n2402 & ~n25863 ;
  assign n25865 = n2591 & n25864 ;
  assign n25866 = n6961 ^ n6917 ^ 1'b0 ;
  assign n25867 = n1197 & n25866 ;
  assign n25868 = ( n20284 & ~n24129 ) | ( n20284 & n25867 ) | ( ~n24129 & n25867 ) ;
  assign n25869 = ~n6581 & n7844 ;
  assign n25870 = n10722 & n25869 ;
  assign n25871 = ( n4015 & n18782 ) | ( n4015 & n25870 ) | ( n18782 & n25870 ) ;
  assign n25872 = n9856 | n17494 ;
  assign n25873 = n25872 ^ n20126 ^ 1'b0 ;
  assign n25874 = ( n671 & n8015 ) | ( n671 & n11343 ) | ( n8015 & n11343 ) ;
  assign n25876 = n3374 & n4595 ;
  assign n25877 = ~n5018 & n25876 ;
  assign n25875 = ( n1499 & n9450 ) | ( n1499 & n14127 ) | ( n9450 & n14127 ) ;
  assign n25878 = n25877 ^ n25875 ^ 1'b0 ;
  assign n25879 = n17083 ^ n16907 ^ 1'b0 ;
  assign n25880 = ~n21211 & n23239 ;
  assign n25881 = ( n9496 & ~n11532 ) | ( n9496 & n17657 ) | ( ~n11532 & n17657 ) ;
  assign n25882 = n25881 ^ n23308 ^ 1'b0 ;
  assign n25883 = n5378 | n25882 ;
  assign n25884 = ( ~n2669 & n4837 ) | ( ~n2669 & n6379 ) | ( n4837 & n6379 ) ;
  assign n25885 = n13220 | n25884 ;
  assign n25886 = n4991 & n10015 ;
  assign n25897 = ( n1733 & n11824 ) | ( n1733 & ~n11985 ) | ( n11824 & ~n11985 ) ;
  assign n25896 = ~n2671 & n6846 ;
  assign n25898 = n25897 ^ n25896 ^ 1'b0 ;
  assign n25899 = ( n2371 & n9126 ) | ( n2371 & n13289 ) | ( n9126 & n13289 ) ;
  assign n25900 = n19473 & ~n25899 ;
  assign n25901 = ~n25898 & n25900 ;
  assign n25888 = ( n2172 & ~n8011 ) | ( n2172 & n14188 ) | ( ~n8011 & n14188 ) ;
  assign n25889 = n1395 | n25888 ;
  assign n25890 = n25889 ^ n23144 ^ 1'b0 ;
  assign n25891 = n19139 ^ n10104 ^ 1'b0 ;
  assign n25892 = n4756 ^ n2690 ^ 1'b0 ;
  assign n25893 = n9512 & n25892 ;
  assign n25894 = n25891 & n25893 ;
  assign n25895 = ~n25890 & n25894 ;
  assign n25887 = n22209 ^ n21086 ^ n982 ;
  assign n25902 = n25901 ^ n25895 ^ n25887 ;
  assign n25903 = ~n1561 & n5707 ;
  assign n25904 = n25903 ^ n16841 ^ 1'b0 ;
  assign n25905 = n6808 & ~n9449 ;
  assign n25906 = n25905 ^ n17482 ^ 1'b0 ;
  assign n25907 = n5183 & n6376 ;
  assign n25908 = n25907 ^ n5634 ^ 1'b0 ;
  assign n25909 = n6896 | n25908 ;
  assign n25910 = n25909 ^ n2684 ^ 1'b0 ;
  assign n25911 = n17936 & ~n25910 ;
  assign n25912 = ~n4173 & n7988 ;
  assign n25913 = n25912 ^ n16271 ^ x50 ;
  assign n25914 = ( n8719 & n10206 ) | ( n8719 & n25913 ) | ( n10206 & n25913 ) ;
  assign n25915 = n4395 & ~n4409 ;
  assign n25916 = ~n25914 & n25915 ;
  assign n25917 = n25916 ^ n15778 ^ 1'b0 ;
  assign n25919 = n16216 ^ n11791 ^ n6213 ;
  assign n25918 = ( ~n10203 & n17520 ) | ( ~n10203 & n21789 ) | ( n17520 & n21789 ) ;
  assign n25920 = n25919 ^ n25918 ^ n21978 ;
  assign n25921 = ( ~n1532 & n15843 ) | ( ~n1532 & n21785 ) | ( n15843 & n21785 ) ;
  assign n25922 = n14452 & ~n25200 ;
  assign n25923 = n25452 ^ n3218 ^ 1'b0 ;
  assign n25924 = ~n14980 & n25923 ;
  assign n25925 = ( n8803 & ~n24999 ) | ( n8803 & n25924 ) | ( ~n24999 & n25924 ) ;
  assign n25926 = n16348 & ~n24915 ;
  assign n25927 = n10195 & n25926 ;
  assign n25928 = ( n10004 & n14951 ) | ( n10004 & ~n17971 ) | ( n14951 & ~n17971 ) ;
  assign n25929 = n25928 ^ n14283 ^ 1'b0 ;
  assign n25930 = ~n13870 & n25929 ;
  assign n25931 = n8986 ^ n8063 ^ n2908 ;
  assign n25932 = n16971 & ~n25931 ;
  assign n25933 = n25932 ^ n19370 ^ 1'b0 ;
  assign n25934 = n6440 & ~n25933 ;
  assign n25935 = n1930 & n25934 ;
  assign n25936 = ( ~n14093 & n23003 ) | ( ~n14093 & n25935 ) | ( n23003 & n25935 ) ;
  assign n25942 = n6120 & ~n7272 ;
  assign n25943 = n25942 ^ n6268 ^ 1'b0 ;
  assign n25939 = ( ~x239 & n1113 ) | ( ~x239 & n2306 ) | ( n1113 & n2306 ) ;
  assign n25940 = n25939 ^ n805 ^ 1'b0 ;
  assign n25941 = ~n8575 & n25940 ;
  assign n25937 = n25131 ^ n16503 ^ n11428 ;
  assign n25938 = ( n9022 & n11147 ) | ( n9022 & n25937 ) | ( n11147 & n25937 ) ;
  assign n25944 = n25943 ^ n25941 ^ n25938 ;
  assign n25945 = n19713 ^ n18851 ^ n12584 ;
  assign n25952 = n5467 & ~n15807 ;
  assign n25947 = n6481 ^ n2684 ^ 1'b0 ;
  assign n25946 = n8686 | n13020 ;
  assign n25948 = n25947 ^ n25946 ^ n11852 ;
  assign n25949 = n477 & ~n25948 ;
  assign n25950 = n25949 ^ n3407 ^ 1'b0 ;
  assign n25951 = n10837 | n25950 ;
  assign n25953 = n25952 ^ n25951 ^ 1'b0 ;
  assign n25954 = n22396 ^ n16161 ^ n7987 ;
  assign n25955 = n25954 ^ n24651 ^ n6130 ;
  assign n25956 = ~n3692 & n18410 ;
  assign n25957 = ( ~n9552 & n21731 ) | ( ~n9552 & n25956 ) | ( n21731 & n25956 ) ;
  assign n25958 = ( n4621 & n22842 ) | ( n4621 & n25957 ) | ( n22842 & n25957 ) ;
  assign n25959 = n7174 ^ n6097 ^ 1'b0 ;
  assign n25960 = n25959 ^ n1569 ^ 1'b0 ;
  assign n25961 = ( n4240 & n15488 ) | ( n4240 & n25960 ) | ( n15488 & n25960 ) ;
  assign n25962 = n13047 & n25961 ;
  assign n25963 = ~n19850 & n25962 ;
  assign n25964 = ( ~n4566 & n18779 ) | ( ~n4566 & n25963 ) | ( n18779 & n25963 ) ;
  assign n25965 = n7268 & n12204 ;
  assign n25966 = ~n10534 & n25965 ;
  assign n25967 = ( n2631 & n10337 ) | ( n2631 & ~n25966 ) | ( n10337 & ~n25966 ) ;
  assign n25968 = n25967 ^ n15934 ^ n8790 ;
  assign n25969 = ( n8894 & n9324 ) | ( n8894 & n18709 ) | ( n9324 & n18709 ) ;
  assign n25970 = ~n10005 & n15908 ;
  assign n25971 = n16032 ^ n5256 ^ n2316 ;
  assign n25972 = n5486 & n25971 ;
  assign n25973 = ~n25970 & n25972 ;
  assign n25974 = n20814 ^ n3503 ^ n2250 ;
  assign n25975 = n20430 ^ n13603 ^ n1313 ;
  assign n25976 = ( ~n25973 & n25974 ) | ( ~n25973 & n25975 ) | ( n25974 & n25975 ) ;
  assign n25977 = ~n3015 & n23091 ;
  assign n25978 = n25977 ^ n7009 ^ 1'b0 ;
  assign n25979 = n9767 ^ n6257 ^ n4378 ;
  assign n25980 = n25979 ^ n16131 ^ n5587 ;
  assign n25981 = n25978 & ~n25980 ;
  assign n25982 = n16619 | n25981 ;
  assign n25983 = n22313 | n25982 ;
  assign n25984 = n6628 ^ n4425 ^ n2353 ;
  assign n25985 = n16057 ^ n8716 ^ 1'b0 ;
  assign n25986 = n23951 & ~n25985 ;
  assign n25987 = n25986 ^ n18858 ^ n14093 ;
  assign n25988 = ( ~n2909 & n25984 ) | ( ~n2909 & n25987 ) | ( n25984 & n25987 ) ;
  assign n25989 = n20611 ^ n4568 ^ 1'b0 ;
  assign n25990 = n25988 & ~n25989 ;
  assign n25991 = n17603 ^ n3494 ^ 1'b0 ;
  assign n25992 = n25991 ^ n11609 ^ 1'b0 ;
  assign n25993 = n14909 | n25992 ;
  assign n25999 = n1068 ^ n1058 ^ 1'b0 ;
  assign n26000 = n7224 | n25999 ;
  assign n25996 = n2050 | n19913 ;
  assign n25997 = n25996 ^ n11935 ^ 1'b0 ;
  assign n25998 = n25997 ^ n18215 ^ 1'b0 ;
  assign n25994 = n12232 | n22236 ;
  assign n25995 = n25702 | n25994 ;
  assign n26001 = n26000 ^ n25998 ^ n25995 ;
  assign n26002 = n4498 & ~n5748 ;
  assign n26003 = ~n2387 & n26002 ;
  assign n26004 = n25294 & ~n26003 ;
  assign n26005 = n11387 | n11555 ;
  assign n26006 = n26005 ^ x49 ^ 1'b0 ;
  assign n26019 = n6211 ^ n4386 ^ 1'b0 ;
  assign n26020 = n4286 & ~n26019 ;
  assign n26014 = ( n9121 & ~n10243 ) | ( n9121 & n16645 ) | ( ~n10243 & n16645 ) ;
  assign n26015 = n26014 ^ n5051 ^ n2495 ;
  assign n26016 = n26015 ^ n24464 ^ n4857 ;
  assign n26017 = n19520 ^ n3976 ^ 1'b0 ;
  assign n26018 = ~n26016 & n26017 ;
  assign n26021 = n26020 ^ n26018 ^ n21799 ;
  assign n26007 = n423 | n22927 ;
  assign n26008 = n26007 ^ n8913 ^ n4680 ;
  assign n26009 = ( ~n19439 & n22711 ) | ( ~n19439 & n26008 ) | ( n22711 & n26008 ) ;
  assign n26010 = n26009 ^ n4319 ^ 1'b0 ;
  assign n26011 = n11638 & ~n26010 ;
  assign n26012 = ~n3526 & n26011 ;
  assign n26013 = n26012 ^ n15409 ^ 1'b0 ;
  assign n26022 = n26021 ^ n26013 ^ n15008 ;
  assign n26023 = n7579 | n25013 ;
  assign n26024 = n26023 ^ n6755 ^ 1'b0 ;
  assign n26025 = n21292 | n26024 ;
  assign n26026 = n15779 | n26025 ;
  assign n26027 = ( n1721 & n4100 ) | ( n1721 & n26026 ) | ( n4100 & n26026 ) ;
  assign n26028 = n8299 ^ n2928 ^ 1'b0 ;
  assign n26029 = n21876 ^ n5753 ^ 1'b0 ;
  assign n26030 = ( n5129 & n6749 ) | ( n5129 & n17279 ) | ( n6749 & n17279 ) ;
  assign n26031 = n26030 ^ n15319 ^ 1'b0 ;
  assign n26032 = x174 & n26031 ;
  assign n26033 = ( n12769 & n26029 ) | ( n12769 & n26032 ) | ( n26029 & n26032 ) ;
  assign n26034 = n17619 & n18644 ;
  assign n26035 = ~n26033 & n26034 ;
  assign n26036 = n10687 ^ n9597 ^ 1'b0 ;
  assign n26037 = n1840 & n26036 ;
  assign n26038 = n10685 ^ n9042 ^ n8798 ;
  assign n26039 = n10046 & n26038 ;
  assign n26040 = ( n3365 & ~n7741 ) | ( n3365 & n23690 ) | ( ~n7741 & n23690 ) ;
  assign n26041 = ~n601 & n759 ;
  assign n26042 = n20339 & n26041 ;
  assign n26043 = ~n13627 & n26042 ;
  assign n26044 = n1414 | n9516 ;
  assign n26045 = n1114 & ~n26044 ;
  assign n26046 = n11595 & ~n14455 ;
  assign n26047 = x156 & n26046 ;
  assign n26048 = n26045 & n26047 ;
  assign n26049 = n13167 & ~n26048 ;
  assign n26050 = n25421 ^ n5402 ^ n4268 ;
  assign n26051 = n566 | n1784 ;
  assign n26052 = n5346 ^ x49 ^ 1'b0 ;
  assign n26053 = n4626 ^ x19 ^ 1'b0 ;
  assign n26054 = x102 & ~n26053 ;
  assign n26055 = n4630 & n6827 ;
  assign n26056 = ~n26054 & n26055 ;
  assign n26057 = n3587 ^ n1990 ^ n1376 ;
  assign n26058 = x134 & n26057 ;
  assign n26059 = n26056 & n26058 ;
  assign n26060 = n386 & n24602 ;
  assign n26061 = n26060 ^ n2466 ^ 1'b0 ;
  assign n26063 = n9727 ^ n2850 ^ 1'b0 ;
  assign n26064 = n1442 | n26063 ;
  assign n26062 = n9365 & n15943 ;
  assign n26065 = n26064 ^ n26062 ^ n2633 ;
  assign n26066 = n21338 ^ n18620 ^ n893 ;
  assign n26067 = n11062 ^ n10308 ^ n2708 ;
  assign n26068 = n8130 ^ n4109 ^ 1'b0 ;
  assign n26069 = n10873 | n26068 ;
  assign n26070 = ~n8376 & n13977 ;
  assign n26071 = ( n25939 & n26069 ) | ( n25939 & n26070 ) | ( n26069 & n26070 ) ;
  assign n26072 = n26071 ^ n21098 ^ n6639 ;
  assign n26083 = ~n17654 & n19535 ;
  assign n26084 = n26083 ^ n1351 ^ 1'b0 ;
  assign n26073 = n8032 ^ x55 ^ 1'b0 ;
  assign n26074 = n26073 ^ n12478 ^ n2903 ;
  assign n26075 = ( n6973 & n8900 ) | ( n6973 & ~n16179 ) | ( n8900 & ~n16179 ) ;
  assign n26076 = n15033 & ~n26075 ;
  assign n26077 = ( n2193 & n8113 ) | ( n2193 & ~n26076 ) | ( n8113 & ~n26076 ) ;
  assign n26079 = n25377 ^ n3997 ^ n1940 ;
  assign n26078 = ~n1293 & n12830 ;
  assign n26080 = n26079 ^ n26078 ^ 1'b0 ;
  assign n26081 = ( n589 & n26077 ) | ( n589 & n26080 ) | ( n26077 & n26080 ) ;
  assign n26082 = ~n26074 & n26081 ;
  assign n26085 = n26084 ^ n26082 ^ 1'b0 ;
  assign n26086 = x95 & ~n14995 ;
  assign n26087 = n26086 ^ n5572 ^ 1'b0 ;
  assign n26088 = n25286 ^ n19079 ^ n6086 ;
  assign n26089 = ~n10198 & n14223 ;
  assign n26090 = n13475 & n26089 ;
  assign n26091 = ( ~n6037 & n16209 ) | ( ~n6037 & n26090 ) | ( n16209 & n26090 ) ;
  assign n26092 = ( n20146 & n23331 ) | ( n20146 & ~n24924 ) | ( n23331 & ~n24924 ) ;
  assign n26093 = ( n3498 & ~n4902 ) | ( n3498 & n21696 ) | ( ~n4902 & n21696 ) ;
  assign n26094 = ( n12179 & ~n19600 ) | ( n12179 & n26093 ) | ( ~n19600 & n26093 ) ;
  assign n26095 = ( n5730 & n15518 ) | ( n5730 & n17614 ) | ( n15518 & n17614 ) ;
  assign n26096 = n6200 | n11949 ;
  assign n26097 = n19382 | n26096 ;
  assign n26098 = ~n8493 & n26097 ;
  assign n26099 = n26095 & n26098 ;
  assign n26100 = ( ~n947 & n22293 ) | ( ~n947 & n24650 ) | ( n22293 & n24650 ) ;
  assign n26101 = n9524 & ~n21650 ;
  assign n26102 = n2582 & n11092 ;
  assign n26103 = n26101 & n26102 ;
  assign n26104 = ( n23127 & n26100 ) | ( n23127 & n26103 ) | ( n26100 & n26103 ) ;
  assign n26105 = n12112 | n17569 ;
  assign n26106 = n26105 ^ n2791 ^ 1'b0 ;
  assign n26107 = n26106 ^ n11588 ^ n4507 ;
  assign n26108 = ( n3430 & ~n21669 ) | ( n3430 & n26107 ) | ( ~n21669 & n26107 ) ;
  assign n26109 = ( n8436 & n10578 ) | ( n8436 & n23932 ) | ( n10578 & n23932 ) ;
  assign n26110 = n17654 | n24418 ;
  assign n26111 = ( n2955 & n8836 ) | ( n2955 & ~n20824 ) | ( n8836 & ~n20824 ) ;
  assign n26112 = n799 | n19004 ;
  assign n26113 = n26112 ^ n4394 ^ 1'b0 ;
  assign n26114 = ~n22729 & n26113 ;
  assign n26115 = n26114 ^ n14284 ^ 1'b0 ;
  assign n26116 = n14500 ^ n11050 ^ 1'b0 ;
  assign n26117 = n1940 & ~n26116 ;
  assign n26118 = ( n327 & n17076 ) | ( n327 & ~n17696 ) | ( n17076 & ~n17696 ) ;
  assign n26119 = ( ~n4847 & n26117 ) | ( ~n4847 & n26118 ) | ( n26117 & n26118 ) ;
  assign n26120 = n26115 & n26119 ;
  assign n26121 = n26120 ^ n12116 ^ 1'b0 ;
  assign n26122 = ( n8587 & n26111 ) | ( n8587 & ~n26121 ) | ( n26111 & ~n26121 ) ;
  assign n26124 = n1410 | n11578 ;
  assign n26123 = n2470 | n3145 ;
  assign n26125 = n26124 ^ n26123 ^ 1'b0 ;
  assign n26126 = n17426 & ~n18088 ;
  assign n26127 = ( ~n504 & n3768 ) | ( ~n504 & n7377 ) | ( n3768 & n7377 ) ;
  assign n26128 = ( n22225 & n26126 ) | ( n22225 & ~n26127 ) | ( n26126 & ~n26127 ) ;
  assign n26129 = n1239 ^ n1113 ^ 1'b0 ;
  assign n26130 = n23125 & ~n26129 ;
  assign n26131 = n14908 ^ n9148 ^ 1'b0 ;
  assign n26132 = n7641 ^ n5110 ^ 1'b0 ;
  assign n26133 = n26131 & n26132 ;
  assign n26134 = n4049 & ~n8333 ;
  assign n26135 = ( n542 & ~n8623 ) | ( n542 & n26134 ) | ( ~n8623 & n26134 ) ;
  assign n26136 = n26135 ^ n13859 ^ n1555 ;
  assign n26137 = n18455 ^ n14560 ^ n360 ;
  assign n26138 = n5435 ^ n3335 ^ 1'b0 ;
  assign n26139 = ( ~n6195 & n18697 ) | ( ~n6195 & n26138 ) | ( n18697 & n26138 ) ;
  assign n26142 = x2 & n18297 ;
  assign n26143 = n26142 ^ n9499 ^ 1'b0 ;
  assign n26144 = x164 & n26143 ;
  assign n26145 = n26144 ^ n21458 ^ 1'b0 ;
  assign n26140 = ( n1225 & ~n4478 ) | ( n1225 & n12746 ) | ( ~n4478 & n12746 ) ;
  assign n26141 = ( n11604 & n12358 ) | ( n11604 & ~n26140 ) | ( n12358 & ~n26140 ) ;
  assign n26146 = n26145 ^ n26141 ^ 1'b0 ;
  assign n26147 = n26139 | n26146 ;
  assign n26148 = ( n14981 & ~n19727 ) | ( n14981 & n24976 ) | ( ~n19727 & n24976 ) ;
  assign n26149 = n2337 & ~n4153 ;
  assign n26150 = n10309 ^ n811 ^ 1'b0 ;
  assign n26151 = n830 & ~n26150 ;
  assign n26152 = ~n20687 & n26151 ;
  assign n26153 = n26152 ^ n19329 ^ 1'b0 ;
  assign n26154 = ~n329 & n7297 ;
  assign n26155 = n20887 ^ n12478 ^ n2343 ;
  assign n26156 = n26154 & n26155 ;
  assign n26157 = ~n2590 & n26156 ;
  assign n26158 = ( n2187 & ~n4544 ) | ( n2187 & n5430 ) | ( ~n4544 & n5430 ) ;
  assign n26159 = n24164 | n26158 ;
  assign n26160 = n26157 & ~n26159 ;
  assign n26164 = n717 & ~n9327 ;
  assign n26161 = n7286 & n8763 ;
  assign n26162 = ~n6211 & n26161 ;
  assign n26163 = ( n8311 & ~n11492 ) | ( n8311 & n26162 ) | ( ~n11492 & n26162 ) ;
  assign n26165 = n26164 ^ n26163 ^ n2413 ;
  assign n26166 = n26165 ^ n9390 ^ 1'b0 ;
  assign n26167 = ~n950 & n26166 ;
  assign n26168 = n3956 | n9876 ;
  assign n26169 = n10088 | n26168 ;
  assign n26170 = n26169 ^ n23899 ^ 1'b0 ;
  assign n26171 = n718 | n10895 ;
  assign n26172 = n26171 ^ n7698 ^ n5809 ;
  assign n26173 = ( n9076 & n15851 ) | ( n9076 & n22130 ) | ( n15851 & n22130 ) ;
  assign n26174 = n19270 ^ n10278 ^ n5853 ;
  assign n26175 = n26174 ^ n25818 ^ n21318 ;
  assign n26176 = n25913 ^ n10676 ^ 1'b0 ;
  assign n26177 = n2469 & n26176 ;
  assign n26178 = n13548 ^ n9381 ^ 1'b0 ;
  assign n26179 = n17597 | n18466 ;
  assign n26180 = n26179 ^ n24139 ^ 1'b0 ;
  assign n26181 = n3377 & ~n10563 ;
  assign n26182 = n26181 ^ n9250 ^ 1'b0 ;
  assign n26186 = n902 & ~n22747 ;
  assign n26187 = n26186 ^ n10408 ^ 1'b0 ;
  assign n26188 = n26187 ^ n7592 ^ 1'b0 ;
  assign n26189 = n26188 ^ n4271 ^ 1'b0 ;
  assign n26190 = ( n4506 & n8723 ) | ( n4506 & n26189 ) | ( n8723 & n26189 ) ;
  assign n26183 = n25984 ^ n3176 ^ 1'b0 ;
  assign n26184 = n26183 ^ n19230 ^ 1'b0 ;
  assign n26185 = n2291 & ~n26184 ;
  assign n26191 = n26190 ^ n26185 ^ n11008 ;
  assign n26192 = n20920 ^ n11172 ^ n6233 ;
  assign n26193 = n2610 | n11353 ;
  assign n26194 = n26193 ^ n23091 ^ 1'b0 ;
  assign n26195 = n26194 ^ n701 ^ 1'b0 ;
  assign n26196 = ~n26192 & n26195 ;
  assign n26197 = n26196 ^ n22600 ^ n5477 ;
  assign n26198 = n3590 ^ n1899 ^ 1'b0 ;
  assign n26199 = n12138 | n20007 ;
  assign n26200 = n26198 | n26199 ;
  assign n26201 = n3184 ^ n896 ^ 1'b0 ;
  assign n26202 = n564 | n26201 ;
  assign n26203 = ~n7334 & n26202 ;
  assign n26204 = ( n5156 & ~n8376 ) | ( n5156 & n17727 ) | ( ~n8376 & n17727 ) ;
  assign n26205 = n26204 ^ n12120 ^ 1'b0 ;
  assign n26206 = ~n740 & n26205 ;
  assign n26207 = n26206 ^ n11416 ^ n2681 ;
  assign n26208 = ( ~n2234 & n12104 ) | ( ~n2234 & n23007 ) | ( n12104 & n23007 ) ;
  assign n26209 = ( n2076 & n10945 ) | ( n2076 & n26208 ) | ( n10945 & n26208 ) ;
  assign n26210 = n16395 ^ n12601 ^ n3491 ;
  assign n26211 = n26210 ^ n4514 ^ 1'b0 ;
  assign n26212 = ~n1712 & n26211 ;
  assign n26213 = n23430 ^ n15856 ^ n6135 ;
  assign n26214 = n22396 ^ n21958 ^ 1'b0 ;
  assign n26215 = n26213 | n26214 ;
  assign n26216 = n6239 & ~n9403 ;
  assign n26217 = n26216 ^ n11896 ^ 1'b0 ;
  assign n26218 = n5092 & ~n26217 ;
  assign n26219 = n26218 ^ n21936 ^ 1'b0 ;
  assign n26220 = n4966 ^ n508 ^ 1'b0 ;
  assign n26221 = n26220 ^ n8109 ^ 1'b0 ;
  assign n26222 = n18950 & ~n26221 ;
  assign n26223 = n4046 ^ n1575 ^ n932 ;
  assign n26224 = ~n6134 & n7345 ;
  assign n26227 = n25107 ^ n2105 ^ 1'b0 ;
  assign n26225 = n16602 ^ n10406 ^ 1'b0 ;
  assign n26226 = n1442 | n26225 ;
  assign n26228 = n26227 ^ n26226 ^ n14956 ;
  assign n26229 = n3704 & n10319 ;
  assign n26230 = n26228 & n26229 ;
  assign n26231 = n12030 ^ n8820 ^ n7759 ;
  assign n26232 = ~n11456 & n14351 ;
  assign n26233 = n26232 ^ n8774 ^ 1'b0 ;
  assign n26234 = n4780 & n26233 ;
  assign n26235 = n12663 | n23441 ;
  assign n26236 = ( ~n9613 & n12688 ) | ( ~n9613 & n17943 ) | ( n12688 & n17943 ) ;
  assign n26237 = n14188 ^ n12729 ^ n9437 ;
  assign n26238 = n26237 ^ n3018 ^ 1'b0 ;
  assign n26240 = n11984 | n18080 ;
  assign n26241 = n26240 ^ n1216 ^ 1'b0 ;
  assign n26239 = n1465 & ~n5283 ;
  assign n26242 = n26241 ^ n26239 ^ 1'b0 ;
  assign n26243 = n17940 ^ n1166 ^ 1'b0 ;
  assign n26244 = n26243 ^ n18413 ^ n8548 ;
  assign n26245 = ( n4100 & n25305 ) | ( n4100 & n26244 ) | ( n25305 & n26244 ) ;
  assign n26246 = n20352 ^ n5775 ^ n2111 ;
  assign n26247 = n23221 ^ n6476 ^ 1'b0 ;
  assign n26248 = ( ~n19868 & n20139 ) | ( ~n19868 & n25549 ) | ( n20139 & n25549 ) ;
  assign n26249 = ( n3931 & n14980 ) | ( n3931 & ~n23174 ) | ( n14980 & ~n23174 ) ;
  assign n26250 = n26249 ^ n22251 ^ 1'b0 ;
  assign n26251 = n16433 ^ n9067 ^ n3263 ;
  assign n26252 = ~n6127 & n26251 ;
  assign n26253 = n21549 | n26252 ;
  assign n26254 = n22876 ^ n9094 ^ n317 ;
  assign n26257 = ( n3123 & ~n4837 ) | ( n3123 & n21628 ) | ( ~n4837 & n21628 ) ;
  assign n26258 = n15785 | n26257 ;
  assign n26259 = n13504 | n26258 ;
  assign n26255 = n15132 & ~n18246 ;
  assign n26256 = n26255 ^ n25725 ^ n7337 ;
  assign n26260 = n26259 ^ n26256 ^ n7763 ;
  assign n26261 = n9688 | n26260 ;
  assign n26262 = n26261 ^ n4128 ^ 1'b0 ;
  assign n26263 = ~n2481 & n15521 ;
  assign n26264 = n8473 & n9456 ;
  assign n26265 = n12167 & ~n26264 ;
  assign n26266 = n26263 & ~n26265 ;
  assign n26267 = ~n8281 & n12576 ;
  assign n26268 = n10802 & n26267 ;
  assign n26269 = n26268 ^ n2878 ^ n2517 ;
  assign n26270 = n26269 ^ n17356 ^ n928 ;
  assign n26271 = ( n609 & n1260 ) | ( n609 & ~n4646 ) | ( n1260 & ~n4646 ) ;
  assign n26272 = n22613 ^ n4994 ^ 1'b0 ;
  assign n26273 = n26271 | n26272 ;
  assign n26274 = n10258 ^ x132 ^ 1'b0 ;
  assign n26275 = n13528 & n26274 ;
  assign n26276 = ( n9908 & n9954 ) | ( n9908 & n26275 ) | ( n9954 & n26275 ) ;
  assign n26277 = n26276 ^ n2670 ^ 1'b0 ;
  assign n26278 = n6904 & n26277 ;
  assign n26279 = ( ~n3069 & n26273 ) | ( ~n3069 & n26278 ) | ( n26273 & n26278 ) ;
  assign n26280 = ( n766 & n2043 ) | ( n766 & n11809 ) | ( n2043 & n11809 ) ;
  assign n26281 = n26280 ^ n22505 ^ n13368 ;
  assign n26282 = ( n13961 & n22064 ) | ( n13961 & ~n25777 ) | ( n22064 & ~n25777 ) ;
  assign n26283 = n5110 ^ n2898 ^ 1'b0 ;
  assign n26284 = ( ~n8813 & n26032 ) | ( ~n8813 & n26283 ) | ( n26032 & n26283 ) ;
  assign n26285 = ( n4576 & n17461 ) | ( n4576 & n26284 ) | ( n17461 & n26284 ) ;
  assign n26286 = n26285 ^ n17554 ^ n16855 ;
  assign n26287 = n5051 ^ n1411 ^ 1'b0 ;
  assign n26288 = ( n5170 & ~n12211 ) | ( n5170 & n26287 ) | ( ~n12211 & n26287 ) ;
  assign n26289 = n13976 ^ n5595 ^ 1'b0 ;
  assign n26290 = n6549 & n26289 ;
  assign n26291 = n26290 ^ n16317 ^ 1'b0 ;
  assign n26292 = n9122 & n12382 ;
  assign n26293 = n20162 & n26292 ;
  assign n26294 = n26293 ^ n6006 ^ n5578 ;
  assign n26295 = ( n8286 & n19322 ) | ( n8286 & n20282 ) | ( n19322 & n20282 ) ;
  assign n26296 = n26295 ^ n16410 ^ n6566 ;
  assign n26297 = n26296 ^ n9138 ^ 1'b0 ;
  assign n26298 = n5937 & n26297 ;
  assign n26299 = n16679 ^ n3615 ^ 1'b0 ;
  assign n26300 = n18536 & ~n26299 ;
  assign n26301 = ~n529 & n1161 ;
  assign n26302 = ~n11729 & n26301 ;
  assign n26303 = ( ~x103 & n620 ) | ( ~x103 & n9567 ) | ( n620 & n9567 ) ;
  assign n26304 = n22779 ^ n19689 ^ n9938 ;
  assign n26305 = n26304 ^ n6573 ^ 1'b0 ;
  assign n26306 = n15933 & n24426 ;
  assign n26307 = n26306 ^ n18246 ^ 1'b0 ;
  assign n26308 = n13814 ^ n10792 ^ 1'b0 ;
  assign n26309 = n22370 ^ x154 ^ 1'b0 ;
  assign n26310 = n26309 ^ n6769 ^ n3505 ;
  assign n26311 = ( n9314 & n9385 ) | ( n9314 & n26310 ) | ( n9385 & n26310 ) ;
  assign n26312 = n14142 ^ n2676 ^ 1'b0 ;
  assign n26313 = ( ~n4552 & n8947 ) | ( ~n4552 & n26312 ) | ( n8947 & n26312 ) ;
  assign n26314 = ( n679 & n1632 ) | ( n679 & ~n3794 ) | ( n1632 & ~n3794 ) ;
  assign n26315 = n26314 ^ n3501 ^ 1'b0 ;
  assign n26316 = n26315 ^ n8973 ^ n1676 ;
  assign n26317 = n24395 ^ n11601 ^ n7016 ;
  assign n26318 = n4549 | n14593 ;
  assign n26319 = n6925 & ~n26318 ;
  assign n26320 = n26319 ^ n18052 ^ n13275 ;
  assign n26321 = n15487 ^ n13992 ^ n3011 ;
  assign n26322 = n16561 ^ n8495 ^ n4345 ;
  assign n26323 = n3329 & ~n14970 ;
  assign n26324 = ~n26322 & n26323 ;
  assign n26325 = n26321 | n26324 ;
  assign n26326 = ( n3253 & n3453 ) | ( n3253 & ~n7585 ) | ( n3453 & ~n7585 ) ;
  assign n26327 = ( ~n3917 & n7748 ) | ( ~n3917 & n8480 ) | ( n7748 & n8480 ) ;
  assign n26328 = ( n3224 & n21754 ) | ( n3224 & ~n25971 ) | ( n21754 & ~n25971 ) ;
  assign n26329 = n21245 ^ n7618 ^ 1'b0 ;
  assign n26330 = n26328 & ~n26329 ;
  assign n26331 = n26327 | n26330 ;
  assign n26332 = n13817 & ~n18252 ;
  assign n26333 = n6768 | n21359 ;
  assign n26334 = n13651 & n21137 ;
  assign n26335 = ~n9610 & n11634 ;
  assign n26336 = n26335 ^ n11292 ^ n3052 ;
  assign n26337 = n26334 & ~n26336 ;
  assign n26338 = n25221 ^ n9972 ^ 1'b0 ;
  assign n26339 = ~n15115 & n26338 ;
  assign n26340 = n26339 ^ n20747 ^ n18776 ;
  assign n26342 = n6009 ^ n1600 ^ 1'b0 ;
  assign n26343 = ( n6565 & n19635 ) | ( n6565 & ~n26342 ) | ( n19635 & ~n26342 ) ;
  assign n26341 = ( n6236 & n11863 ) | ( n6236 & n13321 ) | ( n11863 & n13321 ) ;
  assign n26344 = n26343 ^ n26341 ^ n1492 ;
  assign n26345 = n16960 & n26344 ;
  assign n26346 = n26345 ^ n12106 ^ 1'b0 ;
  assign n26347 = n15779 ^ n2128 ^ 1'b0 ;
  assign n26348 = n26346 | n26347 ;
  assign n26349 = n24310 ^ n21014 ^ n690 ;
  assign n26350 = n26349 ^ n24046 ^ n4809 ;
  assign n26351 = n6376 | n9306 ;
  assign n26352 = ( n1814 & ~n6466 ) | ( n1814 & n26351 ) | ( ~n6466 & n26351 ) ;
  assign n26353 = n26352 ^ n5723 ^ n977 ;
  assign n26354 = n3655 & n25276 ;
  assign n26355 = n1494 | n5653 ;
  assign n26356 = n9052 ^ n7249 ^ 1'b0 ;
  assign n26357 = n26355 & ~n26356 ;
  assign n26358 = n19338 ^ n3233 ^ 1'b0 ;
  assign n26359 = n26357 & ~n26358 ;
  assign n26362 = n8538 ^ n5004 ^ 1'b0 ;
  assign n26366 = n1648 ^ n296 ^ 1'b0 ;
  assign n26363 = n3886 | n4950 ;
  assign n26364 = n8562 ^ n1164 ^ 1'b0 ;
  assign n26365 = n26363 & n26364 ;
  assign n26367 = n26366 ^ n26365 ^ n12329 ;
  assign n26368 = ~n11503 & n12172 ;
  assign n26369 = n26368 ^ n1761 ^ 1'b0 ;
  assign n26370 = n10861 & ~n23039 ;
  assign n26371 = ~n26369 & n26370 ;
  assign n26372 = ( n26362 & ~n26367 ) | ( n26362 & n26371 ) | ( ~n26367 & n26371 ) ;
  assign n26360 = ( n603 & ~n2628 ) | ( n603 & n3202 ) | ( ~n2628 & n3202 ) ;
  assign n26361 = n17718 & ~n26360 ;
  assign n26373 = n26372 ^ n26361 ^ 1'b0 ;
  assign n26374 = n23356 ^ n13884 ^ n5921 ;
  assign n26375 = n8112 ^ n5339 ^ 1'b0 ;
  assign n26376 = n26041 ^ n7531 ^ n3436 ;
  assign n26377 = ( ~n407 & n1908 ) | ( ~n407 & n26376 ) | ( n1908 & n26376 ) ;
  assign n26378 = ( ~n6840 & n23308 ) | ( ~n6840 & n26377 ) | ( n23308 & n26377 ) ;
  assign n26379 = n26378 ^ n15912 ^ 1'b0 ;
  assign n26380 = n26375 & ~n26379 ;
  assign n26381 = ~n18411 & n26380 ;
  assign n26382 = n26374 & n26381 ;
  assign n26383 = n25693 ^ n8917 ^ 1'b0 ;
  assign n26384 = n1319 & ~n26383 ;
  assign n26385 = n21227 ^ n13862 ^ n9931 ;
  assign n26386 = n19098 ^ n10492 ^ 1'b0 ;
  assign n26387 = n26385 & ~n26386 ;
  assign n26388 = ( n13802 & n26384 ) | ( n13802 & n26387 ) | ( n26384 & n26387 ) ;
  assign n26396 = n18455 ^ n16625 ^ n14319 ;
  assign n26394 = n19006 ^ n7536 ^ n5761 ;
  assign n26390 = n3941 & ~n9063 ;
  assign n26391 = n4743 ^ n593 ^ 1'b0 ;
  assign n26392 = n3689 & ~n26391 ;
  assign n26393 = ( n14404 & ~n26390 ) | ( n14404 & n26392 ) | ( ~n26390 & n26392 ) ;
  assign n26395 = n26394 ^ n26393 ^ n21251 ;
  assign n26389 = n8475 ^ n4051 ^ 1'b0 ;
  assign n26397 = n26396 ^ n26395 ^ n26389 ;
  assign n26398 = ~n7964 & n14311 ;
  assign n26399 = ~n25766 & n26398 ;
  assign n26400 = n18505 & ~n26399 ;
  assign n26401 = n6351 & n26400 ;
  assign n26402 = ( ~n1422 & n5416 ) | ( ~n1422 & n21013 ) | ( n5416 & n21013 ) ;
  assign n26403 = ( ~n16440 & n23804 ) | ( ~n16440 & n26402 ) | ( n23804 & n26402 ) ;
  assign n26404 = ( n3661 & n20135 ) | ( n3661 & n22627 ) | ( n20135 & n22627 ) ;
  assign n26405 = n9674 ^ n1408 ^ 1'b0 ;
  assign n26406 = n26405 ^ n21695 ^ 1'b0 ;
  assign n26407 = n12198 ^ n3684 ^ 1'b0 ;
  assign n26408 = n6807 & n13675 ;
  assign n26409 = n26408 ^ x89 ^ 1'b0 ;
  assign n26410 = n6951 | n19101 ;
  assign n26411 = n26410 ^ n20813 ^ 1'b0 ;
  assign n26412 = n26411 ^ n15262 ^ x14 ;
  assign n26413 = n26409 | n26412 ;
  assign n26414 = n14281 ^ n6829 ^ n1524 ;
  assign n26415 = ( n4492 & ~n9527 ) | ( n4492 & n12441 ) | ( ~n9527 & n12441 ) ;
  assign n26416 = ( ~n1645 & n17468 ) | ( ~n1645 & n26415 ) | ( n17468 & n26415 ) ;
  assign n26417 = ~n26414 & n26416 ;
  assign n26418 = n2677 & n26417 ;
  assign n26419 = ~n26413 & n26418 ;
  assign n26420 = n20424 ^ n2043 ^ 1'b0 ;
  assign n26421 = ~n11809 & n26420 ;
  assign n26422 = n11056 ^ n9893 ^ n829 ;
  assign n26423 = ~n5760 & n15201 ;
  assign n26424 = n26423 ^ n3000 ^ 1'b0 ;
  assign n26425 = n16927 ^ n4554 ^ 1'b0 ;
  assign n26426 = ( ~n26422 & n26424 ) | ( ~n26422 & n26425 ) | ( n26424 & n26425 ) ;
  assign n26427 = n1419 & n1468 ;
  assign n26428 = n2172 & n26427 ;
  assign n26429 = ( n644 & n8355 ) | ( n644 & ~n11192 ) | ( n8355 & ~n11192 ) ;
  assign n26430 = n24675 & ~n26429 ;
  assign n26431 = ( n7622 & ~n11771 ) | ( n7622 & n26430 ) | ( ~n11771 & n26430 ) ;
  assign n26432 = n7772 & n26431 ;
  assign n26433 = n26432 ^ n8077 ^ 1'b0 ;
  assign n26434 = ~n14568 & n26433 ;
  assign n26435 = n3458 & ~n5395 ;
  assign n26436 = n23269 & n26435 ;
  assign n26437 = n26436 ^ n8406 ^ 1'b0 ;
  assign n26438 = n23166 & n24246 ;
  assign n26439 = ~n1784 & n5386 ;
  assign n26441 = n6625 ^ n5812 ^ n4490 ;
  assign n26440 = ~n6395 & n17132 ;
  assign n26442 = n26441 ^ n26440 ^ 1'b0 ;
  assign n26443 = n8400 & n26442 ;
  assign n26444 = n734 & n26443 ;
  assign n26445 = n26439 & n26444 ;
  assign n26448 = n7685 ^ n3608 ^ 1'b0 ;
  assign n26446 = n20528 ^ n20085 ^ n8468 ;
  assign n26447 = ~n13719 & n26446 ;
  assign n26449 = n26448 ^ n26447 ^ 1'b0 ;
  assign n26450 = n13728 ^ n10132 ^ n4167 ;
  assign n26451 = n26450 ^ n13006 ^ 1'b0 ;
  assign n26452 = n10294 ^ n7310 ^ 1'b0 ;
  assign n26453 = n6037 | n26452 ;
  assign n26454 = n26453 ^ n16172 ^ n8701 ;
  assign n26455 = ( n7625 & n20001 ) | ( n7625 & n25563 ) | ( n20001 & n25563 ) ;
  assign n26456 = ( ~n26231 & n26454 ) | ( ~n26231 & n26455 ) | ( n26454 & n26455 ) ;
  assign n26457 = n25696 ^ n11737 ^ 1'b0 ;
  assign n26458 = ~n12979 & n26457 ;
  assign n26459 = n19101 ^ n6944 ^ 1'b0 ;
  assign n26466 = x186 & n8085 ;
  assign n26467 = n26466 ^ n4678 ^ 1'b0 ;
  assign n26465 = n8208 & ~n17880 ;
  assign n26468 = n26467 ^ n26465 ^ 1'b0 ;
  assign n26461 = ( n3942 & n6023 ) | ( n3942 & n17562 ) | ( n6023 & n17562 ) ;
  assign n26462 = n11932 ^ n917 ^ 1'b0 ;
  assign n26463 = ~n2928 & n26462 ;
  assign n26464 = ( n19818 & ~n26461 ) | ( n19818 & n26463 ) | ( ~n26461 & n26463 ) ;
  assign n26460 = ~n6090 & n11425 ;
  assign n26469 = n26468 ^ n26464 ^ n26460 ;
  assign n26470 = n20975 ^ n17937 ^ n11635 ;
  assign n26471 = n20276 | n23333 ;
  assign n26472 = ( n5651 & n19991 ) | ( n5651 & ~n20471 ) | ( n19991 & ~n20471 ) ;
  assign n26473 = n9662 | n12371 ;
  assign n26474 = n25224 ^ n10905 ^ 1'b0 ;
  assign n26475 = n26473 & ~n26474 ;
  assign n26476 = ~n26472 & n26475 ;
  assign n26477 = n23570 | n25956 ;
  assign n26478 = ~n1449 & n26477 ;
  assign n26479 = n26476 & n26478 ;
  assign n26480 = n24044 & n25419 ;
  assign n26481 = n16741 ^ n4265 ^ n3914 ;
  assign n26482 = ( n1295 & ~n9617 ) | ( n1295 & n14151 ) | ( ~n9617 & n14151 ) ;
  assign n26483 = n26481 & ~n26482 ;
  assign n26484 = n10138 ^ n8902 ^ n6455 ;
  assign n26485 = n8730 ^ n5733 ^ n4594 ;
  assign n26486 = n18312 ^ n10438 ^ n6299 ;
  assign n26487 = ~n2743 & n12821 ;
  assign n26488 = n18487 & n26487 ;
  assign n26489 = ( ~n9191 & n26486 ) | ( ~n9191 & n26488 ) | ( n26486 & n26488 ) ;
  assign n26490 = ( n12766 & n26485 ) | ( n12766 & ~n26489 ) | ( n26485 & ~n26489 ) ;
  assign n26491 = ~n10268 & n22845 ;
  assign n26492 = ( n5373 & ~n6608 ) | ( n5373 & n9131 ) | ( ~n6608 & n9131 ) ;
  assign n26493 = n26492 ^ n12207 ^ n3635 ;
  assign n26494 = n9887 | n26493 ;
  assign n26495 = n25076 ^ n5158 ^ 1'b0 ;
  assign n26496 = n1927 & n26495 ;
  assign n26497 = n11863 ^ n1989 ^ n1199 ;
  assign n26498 = ( ~n16577 & n17047 ) | ( ~n16577 & n26497 ) | ( n17047 & n26497 ) ;
  assign n26499 = n3835 & n16885 ;
  assign n26500 = n24553 ^ n2177 ^ 1'b0 ;
  assign n26501 = n23904 & n26500 ;
  assign n26502 = ~n11448 & n26501 ;
  assign n26503 = ( n3083 & n26499 ) | ( n3083 & n26502 ) | ( n26499 & n26502 ) ;
  assign n26504 = n1109 ^ n617 ^ 1'b0 ;
  assign n26505 = ~n6554 & n26504 ;
  assign n26506 = n9468 ^ n7175 ^ 1'b0 ;
  assign n26507 = ~n5312 & n26506 ;
  assign n26508 = n15887 & n26507 ;
  assign n26509 = ( n15659 & n26505 ) | ( n15659 & ~n26508 ) | ( n26505 & ~n26508 ) ;
  assign n26510 = n2152 & n13446 ;
  assign n26511 = n26510 ^ n26424 ^ 1'b0 ;
  assign n26512 = n7899 ^ n4274 ^ 1'b0 ;
  assign n26513 = n6500 & ~n26512 ;
  assign n26514 = ~n2471 & n26513 ;
  assign n26515 = ( n5115 & ~n5265 ) | ( n5115 & n13865 ) | ( ~n5265 & n13865 ) ;
  assign n26516 = n6876 ^ n963 ^ 1'b0 ;
  assign n26517 = n26515 | n26516 ;
  assign n26518 = ~n14116 & n21947 ;
  assign n26519 = n26517 & n26518 ;
  assign n26520 = n18276 ^ n8124 ^ 1'b0 ;
  assign n26521 = n26520 ^ n21892 ^ n5679 ;
  assign n26522 = n26416 ^ n14297 ^ 1'b0 ;
  assign n26523 = n13677 ^ n8801 ^ 1'b0 ;
  assign n26524 = ~n6887 & n26523 ;
  assign n26527 = ~n11025 & n20272 ;
  assign n26526 = n2607 ^ n2039 ^ 1'b0 ;
  assign n26525 = ~n5426 & n11521 ;
  assign n26528 = n26527 ^ n26526 ^ n26525 ;
  assign n26529 = n8973 ^ n3739 ^ 1'b0 ;
  assign n26530 = ( n9420 & n11536 ) | ( n9420 & ~n20321 ) | ( n11536 & ~n20321 ) ;
  assign n26531 = ~n2764 & n7828 ;
  assign n26532 = ~n2096 & n26531 ;
  assign n26533 = ( n26529 & n26530 ) | ( n26529 & n26532 ) | ( n26530 & n26532 ) ;
  assign n26534 = ~n9861 & n17181 ;
  assign n26535 = n26534 ^ n26441 ^ n7382 ;
  assign n26536 = n6607 & n26535 ;
  assign n26537 = n11335 & n26536 ;
  assign n26541 = ~n2166 & n4674 ;
  assign n26538 = ( ~n13038 & n17255 ) | ( ~n13038 & n19038 ) | ( n17255 & n19038 ) ;
  assign n26539 = n2070 & n21607 ;
  assign n26540 = ~n26538 & n26539 ;
  assign n26542 = n26541 ^ n26540 ^ n7686 ;
  assign n26543 = ( n9875 & n16732 ) | ( n9875 & n22588 ) | ( n16732 & n22588 ) ;
  assign n26544 = ( n2292 & n12908 ) | ( n2292 & n13563 ) | ( n12908 & n13563 ) ;
  assign n26545 = n18527 ^ n8684 ^ n1767 ;
  assign n26546 = ~n11885 & n26545 ;
  assign n26547 = n16622 ^ n12870 ^ n9008 ;
  assign n26548 = n5944 & n6995 ;
  assign n26549 = ~n9871 & n13072 ;
  assign n26550 = n26548 & n26549 ;
  assign n26551 = n11948 | n14494 ;
  assign n26552 = n26550 & ~n26551 ;
  assign n26553 = n23486 ^ n18384 ^ 1'b0 ;
  assign n26554 = n6783 ^ n812 ^ 1'b0 ;
  assign n26555 = n13384 & n24719 ;
  assign n26556 = n10536 & n26555 ;
  assign n26557 = n4787 & ~n7906 ;
  assign n26558 = n26557 ^ n289 ^ 1'b0 ;
  assign n26559 = n26558 ^ n3353 ^ 1'b0 ;
  assign n26560 = ~n16732 & n26559 ;
  assign n26562 = ( ~n818 & n1920 ) | ( ~n818 & n6097 ) | ( n1920 & n6097 ) ;
  assign n26563 = n13794 & ~n26562 ;
  assign n26561 = n22710 ^ n18125 ^ n6861 ;
  assign n26564 = n26563 ^ n26561 ^ 1'b0 ;
  assign n26567 = ( n1239 & n5809 ) | ( n1239 & ~n11735 ) | ( n5809 & ~n11735 ) ;
  assign n26568 = n26567 ^ n15313 ^ 1'b0 ;
  assign n26565 = n12244 & ~n14307 ;
  assign n26566 = ~n2940 & n26565 ;
  assign n26569 = n26568 ^ n26566 ^ 1'b0 ;
  assign n26570 = n4465 & n7450 ;
  assign n26571 = n26570 ^ n7683 ^ 1'b0 ;
  assign n26572 = n10680 ^ n4201 ^ 1'b0 ;
  assign n26573 = n26571 & ~n26572 ;
  assign n26574 = ( n5995 & ~n25534 ) | ( n5995 & n26573 ) | ( ~n25534 & n26573 ) ;
  assign n26575 = n22047 ^ n20085 ^ 1'b0 ;
  assign n26576 = n26575 ^ n10418 ^ 1'b0 ;
  assign n26577 = n15479 ^ n9008 ^ 1'b0 ;
  assign n26578 = n10393 & n14210 ;
  assign n26579 = n24539 & n26578 ;
  assign n26580 = n26579 ^ n19481 ^ 1'b0 ;
  assign n26581 = n26577 & n26580 ;
  assign n26582 = ~n1756 & n26500 ;
  assign n26583 = n15012 ^ n2350 ^ 1'b0 ;
  assign n26584 = n14051 ^ n9314 ^ n2958 ;
  assign n26585 = ( n3002 & ~n14459 ) | ( n3002 & n26584 ) | ( ~n14459 & n26584 ) ;
  assign n26586 = ( ~n21449 & n26583 ) | ( ~n21449 & n26585 ) | ( n26583 & n26585 ) ;
  assign n26588 = n2273 & n2879 ;
  assign n26589 = ~n7541 & n26588 ;
  assign n26590 = n26280 & ~n26589 ;
  assign n26591 = n26590 ^ n5230 ^ 1'b0 ;
  assign n26587 = n6387 | n26257 ;
  assign n26592 = n26591 ^ n26587 ^ 1'b0 ;
  assign n26593 = n26592 ^ n12936 ^ n7719 ;
  assign n26594 = n969 & ~n18024 ;
  assign n26595 = n17265 ^ n14126 ^ 1'b0 ;
  assign n26596 = n923 & n14106 ;
  assign n26597 = n22254 ^ n21830 ^ n4618 ;
  assign n26598 = n26597 ^ n13829 ^ 1'b0 ;
  assign n26599 = n12967 & ~n16709 ;
  assign n26600 = n2098 | n11209 ;
  assign n26601 = n26599 & ~n26600 ;
  assign n26603 = ( n1725 & ~n20572 ) | ( n1725 & n26126 ) | ( ~n20572 & n26126 ) ;
  assign n26602 = n4161 & n7827 ;
  assign n26604 = n26603 ^ n26602 ^ 1'b0 ;
  assign n26605 = n3201 ^ n2126 ^ x161 ;
  assign n26606 = n11123 & n20653 ;
  assign n26607 = n26606 ^ n11796 ^ 1'b0 ;
  assign n26608 = ( n13557 & n26605 ) | ( n13557 & n26607 ) | ( n26605 & n26607 ) ;
  assign n26609 = ( n17540 & ~n23147 ) | ( n17540 & n26608 ) | ( ~n23147 & n26608 ) ;
  assign n26611 = ~n8370 & n8979 ;
  assign n26610 = n21642 ^ n19564 ^ n7030 ;
  assign n26612 = n26611 ^ n26610 ^ 1'b0 ;
  assign n26613 = n7906 | n25736 ;
  assign n26614 = n15825 & ~n26613 ;
  assign n26615 = n10724 ^ n803 ^ 1'b0 ;
  assign n26616 = n14055 | n26615 ;
  assign n26617 = n4158 | n10196 ;
  assign n26618 = n6919 | n26617 ;
  assign n26619 = n26618 ^ n2308 ^ 1'b0 ;
  assign n26620 = n15856 ^ n1872 ^ n1102 ;
  assign n26621 = n18767 ^ n10521 ^ n10468 ;
  assign n26622 = n26621 ^ n21802 ^ n17833 ;
  assign n26623 = n16440 ^ n9077 ^ n1111 ;
  assign n26624 = n11476 | n26623 ;
  assign n26625 = n26624 ^ n3464 ^ 1'b0 ;
  assign n26626 = n25853 ^ n17982 ^ x4 ;
  assign n26627 = n14290 ^ n5548 ^ n3415 ;
  assign n26628 = ~n6392 & n26627 ;
  assign n26629 = n26626 | n26628 ;
  assign n26630 = n15714 ^ n5125 ^ 1'b0 ;
  assign n26631 = ~n21742 & n26630 ;
  assign n26632 = n26631 ^ n16266 ^ 1'b0 ;
  assign n26633 = n8104 ^ n7086 ^ n4829 ;
  assign n26634 = n24914 ^ n16184 ^ 1'b0 ;
  assign n26637 = n19628 ^ n7475 ^ x12 ;
  assign n26636 = n8883 ^ n7973 ^ 1'b0 ;
  assign n26638 = n26637 ^ n26636 ^ n24719 ;
  assign n26639 = n26638 ^ n6420 ^ 1'b0 ;
  assign n26635 = ~n1221 & n4716 ;
  assign n26640 = n26639 ^ n26635 ^ 1'b0 ;
  assign n26641 = ( ~n3050 & n7862 ) | ( ~n3050 & n26640 ) | ( n7862 & n26640 ) ;
  assign n26642 = ( x141 & ~n1505 ) | ( x141 & n3660 ) | ( ~n1505 & n3660 ) ;
  assign n26643 = n387 | n26642 ;
  assign n26645 = n10651 & ~n11533 ;
  assign n26644 = n19105 ^ n1250 ^ 1'b0 ;
  assign n26646 = n26645 ^ n26644 ^ n23249 ;
  assign n26647 = n17879 ^ n8224 ^ 1'b0 ;
  assign n26648 = n9261 ^ n5931 ^ n5889 ;
  assign n26649 = n9164 | n26648 ;
  assign n26650 = n26647 & ~n26649 ;
  assign n26651 = ( n4613 & n6773 ) | ( n4613 & ~n26650 ) | ( n6773 & ~n26650 ) ;
  assign n26655 = ( n2004 & ~n3111 ) | ( n2004 & n7410 ) | ( ~n3111 & n7410 ) ;
  assign n26652 = n24427 ^ n3887 ^ 1'b0 ;
  assign n26653 = ~n335 & n26652 ;
  assign n26654 = n18822 & n26653 ;
  assign n26656 = n26655 ^ n26654 ^ 1'b0 ;
  assign n26657 = n20594 ^ n7409 ^ 1'b0 ;
  assign n26658 = n18823 ^ n9998 ^ 1'b0 ;
  assign n26659 = n10574 | n12913 ;
  assign n26660 = n12262 | n26659 ;
  assign n26661 = ( n15316 & ~n26658 ) | ( n15316 & n26660 ) | ( ~n26658 & n26660 ) ;
  assign n26662 = ( ~n25288 & n26657 ) | ( ~n25288 & n26661 ) | ( n26657 & n26661 ) ;
  assign n26663 = n26662 ^ n16623 ^ n9730 ;
  assign n26664 = n11811 ^ n5367 ^ n1286 ;
  assign n26665 = ~n11352 & n26664 ;
  assign n26666 = n9389 & n26665 ;
  assign n26667 = ~n6211 & n10546 ;
  assign n26668 = n21161 | n21346 ;
  assign n26669 = ( n7247 & n19346 ) | ( n7247 & ~n20135 ) | ( n19346 & ~n20135 ) ;
  assign n26670 = n24186 ^ n18620 ^ n2804 ;
  assign n26672 = ~n8657 & n23332 ;
  assign n26673 = ~n9616 & n26672 ;
  assign n26674 = n26673 ^ n13849 ^ n4599 ;
  assign n26671 = ( n8094 & ~n17263 ) | ( n8094 & n18180 ) | ( ~n17263 & n18180 ) ;
  assign n26675 = n26674 ^ n26671 ^ 1'b0 ;
  assign n26680 = n693 & ~n11730 ;
  assign n26677 = n7131 ^ x193 ^ 1'b0 ;
  assign n26678 = ~n2771 & n26677 ;
  assign n26679 = n26678 ^ n10727 ^ 1'b0 ;
  assign n26681 = n26680 ^ n26679 ^ n5897 ;
  assign n26682 = ( n1691 & n4899 ) | ( n1691 & ~n10782 ) | ( n4899 & ~n10782 ) ;
  assign n26683 = n26681 & n26682 ;
  assign n26684 = n26683 ^ n5043 ^ 1'b0 ;
  assign n26676 = ( ~n12300 & n14412 ) | ( ~n12300 & n17807 ) | ( n14412 & n17807 ) ;
  assign n26685 = n26684 ^ n26676 ^ x4 ;
  assign n26689 = ( x28 & ~n5231 ) | ( x28 & n5283 ) | ( ~n5231 & n5283 ) ;
  assign n26686 = n12929 ^ n7169 ^ 1'b0 ;
  assign n26687 = n26686 ^ n15022 ^ n14138 ;
  assign n26688 = ~n6451 & n26687 ;
  assign n26690 = n26689 ^ n26688 ^ 1'b0 ;
  assign n26691 = n16764 & ~n26690 ;
  assign n26692 = ( n23968 & ~n26685 ) | ( n23968 & n26691 ) | ( ~n26685 & n26691 ) ;
  assign n26693 = n17191 ^ n7700 ^ n6593 ;
  assign n26694 = x129 & ~n8657 ;
  assign n26695 = n26694 ^ n15190 ^ 1'b0 ;
  assign n26696 = ( n25520 & n26693 ) | ( n25520 & n26695 ) | ( n26693 & n26695 ) ;
  assign n26697 = n7203 ^ n1431 ^ 1'b0 ;
  assign n26698 = n26697 ^ n11429 ^ 1'b0 ;
  assign n26699 = n10307 ^ n4555 ^ 1'b0 ;
  assign n26700 = ( n7094 & ~n18651 ) | ( n7094 & n25799 ) | ( ~n18651 & n25799 ) ;
  assign n26701 = n1481 & ~n4333 ;
  assign n26702 = n1809 & n26701 ;
  assign n26703 = n26702 ^ n23172 ^ n11217 ;
  assign n26704 = n26703 ^ n7044 ^ n2013 ;
  assign n26705 = n26700 | n26704 ;
  assign n26706 = n11671 | n26705 ;
  assign n26707 = n26706 ^ n6177 ^ 1'b0 ;
  assign n26708 = ~n23144 & n26707 ;
  assign n26709 = n26699 & n26708 ;
  assign n26710 = ( ~n10020 & n10766 ) | ( ~n10020 & n21708 ) | ( n10766 & n21708 ) ;
  assign n26711 = n26710 ^ n12205 ^ n10800 ;
  assign n26712 = n15511 ^ n10086 ^ n2046 ;
  assign n26717 = n9176 ^ n8217 ^ x202 ;
  assign n26715 = n8447 | n10845 ;
  assign n26713 = n6485 & ~n16275 ;
  assign n26714 = n26713 ^ n24602 ^ 1'b0 ;
  assign n26716 = n26715 ^ n26714 ^ n835 ;
  assign n26718 = n26717 ^ n26716 ^ n13451 ;
  assign n26719 = ( n4707 & ~n6557 ) | ( n4707 & n9945 ) | ( ~n6557 & n9945 ) ;
  assign n26720 = n26719 ^ n7330 ^ 1'b0 ;
  assign n26721 = n19182 & n26720 ;
  assign n26722 = n26721 ^ n19323 ^ 1'b0 ;
  assign n26723 = ~n23016 & n26722 ;
  assign n26724 = n26723 ^ n1221 ^ 1'b0 ;
  assign n26725 = n22866 ^ n4785 ^ 1'b0 ;
  assign n26726 = n8893 & ~n26725 ;
  assign n26727 = n5783 | n23099 ;
  assign n26728 = x181 | n26727 ;
  assign n26729 = n26728 ^ n14677 ^ 1'b0 ;
  assign n26730 = n26729 ^ n16156 ^ n5616 ;
  assign n26731 = ( n2217 & ~n8654 ) | ( n2217 & n26730 ) | ( ~n8654 & n26730 ) ;
  assign n26732 = ( ~n2317 & n14165 ) | ( ~n2317 & n19070 ) | ( n14165 & n19070 ) ;
  assign n26733 = n25752 ^ n4732 ^ 1'b0 ;
  assign n26734 = ( n2840 & ~n8233 ) | ( n2840 & n26733 ) | ( ~n8233 & n26733 ) ;
  assign n26738 = n12835 ^ n10027 ^ 1'b0 ;
  assign n26739 = ( n1836 & ~n14065 ) | ( n1836 & n26738 ) | ( ~n14065 & n26738 ) ;
  assign n26735 = n1951 ^ n1891 ^ 1'b0 ;
  assign n26736 = n23156 & n26735 ;
  assign n26737 = n22412 & n26736 ;
  assign n26740 = n26739 ^ n26737 ^ 1'b0 ;
  assign n26741 = ( n10861 & n16202 ) | ( n10861 & ~n17091 ) | ( n16202 & ~n17091 ) ;
  assign n26742 = ( n1416 & n17333 ) | ( n1416 & n26741 ) | ( n17333 & n26741 ) ;
  assign n26743 = n24494 ^ n6630 ^ 1'b0 ;
  assign n26744 = n26742 | n26743 ;
  assign n26745 = n17727 ^ n14952 ^ n8393 ;
  assign n26746 = n26745 ^ n11878 ^ n3117 ;
  assign n26747 = n23730 ^ n19655 ^ n4759 ;
  assign n26748 = n16507 ^ n13560 ^ 1'b0 ;
  assign n26749 = n26748 ^ n2536 ^ 1'b0 ;
  assign n26750 = ~n26747 & n26749 ;
  assign n26751 = ( n4303 & n18074 ) | ( n4303 & ~n26750 ) | ( n18074 & ~n26750 ) ;
  assign n26753 = ( n2014 & ~n4424 ) | ( n2014 & n8398 ) | ( ~n4424 & n8398 ) ;
  assign n26754 = n4596 & ~n26753 ;
  assign n26755 = n26754 ^ n17191 ^ 1'b0 ;
  assign n26752 = ~n6752 & n9282 ;
  assign n26756 = n26755 ^ n26752 ^ 1'b0 ;
  assign n26759 = n8838 & n10862 ;
  assign n26760 = n26759 ^ n5785 ^ 1'b0 ;
  assign n26757 = ( n1708 & n12780 ) | ( n1708 & ~n16399 ) | ( n12780 & ~n16399 ) ;
  assign n26758 = n26757 ^ n9233 ^ 1'b0 ;
  assign n26761 = n26760 ^ n26758 ^ n667 ;
  assign n26762 = n9324 & ~n26761 ;
  assign n26763 = n17607 ^ n13158 ^ n8732 ;
  assign n26764 = n7241 ^ n4771 ^ n2673 ;
  assign n26765 = n26763 | n26764 ;
  assign n26766 = n20671 & ~n21397 ;
  assign n26767 = n2448 & n26766 ;
  assign n26768 = n26767 ^ n3420 ^ 1'b0 ;
  assign n26769 = ~n630 & n12447 ;
  assign n26770 = ~n2538 & n26769 ;
  assign n26771 = n26770 ^ n9135 ^ 1'b0 ;
  assign n26772 = n14795 | n26771 ;
  assign n26773 = n26772 ^ n22223 ^ n11357 ;
  assign n26774 = n26760 ^ n1708 ^ 1'b0 ;
  assign n26775 = n1776 | n26774 ;
  assign n26776 = ( ~n8884 & n12385 ) | ( ~n8884 & n12856 ) | ( n12385 & n12856 ) ;
  assign n26777 = n8984 & n26776 ;
  assign n26782 = ( n8947 & ~n14747 ) | ( n8947 & n17222 ) | ( ~n14747 & n17222 ) ;
  assign n26778 = n990 & ~n24999 ;
  assign n26779 = ~n4234 & n26778 ;
  assign n26780 = n20088 ^ n2632 ^ n969 ;
  assign n26781 = n26779 & ~n26780 ;
  assign n26783 = n26782 ^ n26781 ^ n21079 ;
  assign n26785 = n3972 & ~n9621 ;
  assign n26786 = n26785 ^ n11443 ^ 1'b0 ;
  assign n26784 = ( ~n873 & n6180 ) | ( ~n873 & n11984 ) | ( n6180 & n11984 ) ;
  assign n26787 = n26786 ^ n26784 ^ n8588 ;
  assign n26788 = ~n861 & n10352 ;
  assign n26789 = n8270 & n26788 ;
  assign n26790 = n4156 & ~n26789 ;
  assign n26791 = n13860 & ~n26790 ;
  assign n26792 = n26791 ^ n9579 ^ 1'b0 ;
  assign n26793 = n16596 | n26792 ;
  assign n26794 = ~n13465 & n26793 ;
  assign n26795 = n13509 & ~n19468 ;
  assign n26796 = ~n1785 & n11848 ;
  assign n26797 = ~n13677 & n26796 ;
  assign n26798 = n20854 ^ n6959 ^ n4448 ;
  assign n26799 = x205 & n15312 ;
  assign n26800 = ~n5267 & n26799 ;
  assign n26801 = n5752 ^ n4209 ^ 1'b0 ;
  assign n26802 = ~n26800 & n26801 ;
  assign n26803 = ( ~n24696 & n26798 ) | ( ~n24696 & n26802 ) | ( n26798 & n26802 ) ;
  assign n26804 = n26797 | n26803 ;
  assign n26805 = n20076 ^ n12234 ^ 1'b0 ;
  assign n26806 = n25088 | n26805 ;
  assign n26807 = n7850 ^ n883 ^ 1'b0 ;
  assign n26808 = n6297 | n26807 ;
  assign n26809 = n9267 | n26808 ;
  assign n26810 = n26809 ^ n21391 ^ 1'b0 ;
  assign n26811 = n18229 ^ n9990 ^ 1'b0 ;
  assign n26812 = n1731 & ~n26811 ;
  assign n26813 = n26812 ^ n18722 ^ n10588 ;
  assign n26814 = n26813 ^ n11231 ^ n7452 ;
  assign n26815 = n6017 ^ n2451 ^ 1'b0 ;
  assign n26816 = ~n1306 & n26815 ;
  assign n26817 = n19601 & n26816 ;
  assign n26818 = n1650 | n16141 ;
  assign n26819 = ~n270 & n25095 ;
  assign n26820 = n26819 ^ n23377 ^ 1'b0 ;
  assign n26821 = n8540 ^ n4224 ^ n586 ;
  assign n26822 = ~n3746 & n26821 ;
  assign n26823 = x59 & n868 ;
  assign n26824 = n26823 ^ n11124 ^ 1'b0 ;
  assign n26825 = n26824 ^ n13274 ^ n3060 ;
  assign n26826 = ( x61 & n24571 ) | ( x61 & n26825 ) | ( n24571 & n26825 ) ;
  assign n26827 = ( n2052 & n2947 ) | ( n2052 & n12845 ) | ( n2947 & n12845 ) ;
  assign n26828 = ( ~n8091 & n26826 ) | ( ~n8091 & n26827 ) | ( n26826 & n26827 ) ;
  assign n26829 = ( n6238 & n7376 ) | ( n6238 & n18386 ) | ( n7376 & n18386 ) ;
  assign n26830 = ( ~n12944 & n15120 ) | ( ~n12944 & n15347 ) | ( n15120 & n15347 ) ;
  assign n26831 = n3770 | n6407 ;
  assign n26832 = n26831 ^ n2364 ^ 1'b0 ;
  assign n26833 = ( n2188 & ~n5391 ) | ( n2188 & n15423 ) | ( ~n5391 & n15423 ) ;
  assign n26834 = ( n18169 & n26832 ) | ( n18169 & ~n26833 ) | ( n26832 & ~n26833 ) ;
  assign n26835 = ( n25547 & ~n26830 ) | ( n25547 & n26834 ) | ( ~n26830 & n26834 ) ;
  assign n26836 = x86 & n8184 ;
  assign n26837 = ~n20671 & n26836 ;
  assign n26838 = n22260 & ~n26837 ;
  assign n26839 = n26838 ^ n10916 ^ 1'b0 ;
  assign n26840 = n25650 ^ n16360 ^ n640 ;
  assign n26841 = n4009 & ~n11628 ;
  assign n26842 = ( n11271 & n26840 ) | ( n11271 & ~n26841 ) | ( n26840 & ~n26841 ) ;
  assign n26843 = n26842 ^ n15339 ^ 1'b0 ;
  assign n26844 = n26843 ^ n21822 ^ n12935 ;
  assign n26847 = n9944 ^ n4165 ^ n1440 ;
  assign n26845 = n15886 ^ n7670 ^ 1'b0 ;
  assign n26846 = ( n9108 & n19001 ) | ( n9108 & n26845 ) | ( n19001 & n26845 ) ;
  assign n26848 = n26847 ^ n26846 ^ n1564 ;
  assign n26849 = n26848 ^ n5275 ^ 1'b0 ;
  assign n26850 = n26844 | n26849 ;
  assign n26851 = n8156 & ~n18207 ;
  assign n26852 = ( ~n10538 & n12542 ) | ( ~n10538 & n26851 ) | ( n12542 & n26851 ) ;
  assign n26853 = n26852 ^ n14822 ^ n4221 ;
  assign n26854 = ( ~n761 & n11830 ) | ( ~n761 & n13462 ) | ( n11830 & n13462 ) ;
  assign n26855 = n26854 ^ n9321 ^ 1'b0 ;
  assign n26858 = n16781 ^ n12556 ^ n11379 ;
  assign n26856 = x244 & n6260 ;
  assign n26857 = ~n15831 & n26856 ;
  assign n26859 = n26858 ^ n26857 ^ n2067 ;
  assign n26860 = ( ~n14966 & n25074 ) | ( ~n14966 & n26859 ) | ( n25074 & n26859 ) ;
  assign n26861 = ( n4818 & ~n11180 ) | ( n4818 & n24529 ) | ( ~n11180 & n24529 ) ;
  assign n26862 = n1135 & ~n26861 ;
  assign n26863 = ~n20317 & n20371 ;
  assign n26864 = n26863 ^ n13980 ^ 1'b0 ;
  assign n26865 = ( n3310 & ~n6632 ) | ( n3310 & n16694 ) | ( ~n6632 & n16694 ) ;
  assign n26866 = ( x107 & n2127 ) | ( x107 & n20832 ) | ( n2127 & n20832 ) ;
  assign n26867 = n13181 & ~n18401 ;
  assign n26868 = n26867 ^ n20210 ^ 1'b0 ;
  assign n26869 = n26866 | n26868 ;
  assign n26870 = n26869 ^ n16953 ^ 1'b0 ;
  assign n26871 = n23726 ^ n1897 ^ x231 ;
  assign n26872 = n26871 ^ n14543 ^ n6671 ;
  assign n26873 = n20446 ^ n5547 ^ n5519 ;
  assign n26874 = n1315 | n9542 ;
  assign n26875 = ~n14624 & n26874 ;
  assign n26876 = n26875 ^ n26579 ^ 1'b0 ;
  assign n26877 = n17110 ^ n13271 ^ 1'b0 ;
  assign n26878 = n24687 ^ n6312 ^ 1'b0 ;
  assign n26879 = n26878 ^ n22081 ^ n21908 ;
  assign n26880 = n3635 | n14787 ;
  assign n26881 = ( n3956 & n19621 ) | ( n3956 & ~n26880 ) | ( n19621 & ~n26880 ) ;
  assign n26883 = n1620 & n8902 ;
  assign n26882 = ~n5960 & n23217 ;
  assign n26884 = n26883 ^ n26882 ^ 1'b0 ;
  assign n26886 = ( n2324 & ~n7352 ) | ( n2324 & n7919 ) | ( ~n7352 & n7919 ) ;
  assign n26885 = n9507 ^ n6323 ^ 1'b0 ;
  assign n26887 = n26886 ^ n26885 ^ n20008 ;
  assign n26888 = ( n4371 & n4549 ) | ( n4371 & ~n26887 ) | ( n4549 & ~n26887 ) ;
  assign n26889 = n5484 & ~n26888 ;
  assign n26890 = ( ~n2904 & n8259 ) | ( ~n2904 & n16228 ) | ( n8259 & n16228 ) ;
  assign n26891 = ( ~n7106 & n8158 ) | ( ~n7106 & n16198 ) | ( n8158 & n16198 ) ;
  assign n26894 = n10641 ^ n1652 ^ 1'b0 ;
  assign n26895 = ~n1208 & n26894 ;
  assign n26892 = n3232 & ~n13390 ;
  assign n26893 = n26892 ^ n9257 ^ 1'b0 ;
  assign n26896 = n26895 ^ n26893 ^ n1189 ;
  assign n26897 = ( ~n5707 & n8191 ) | ( ~n5707 & n26896 ) | ( n8191 & n26896 ) ;
  assign n26898 = n26897 ^ n20403 ^ n19995 ;
  assign n26899 = n18382 ^ n15539 ^ n13838 ;
  assign n26900 = ~n1193 & n26899 ;
  assign n26901 = ( n3565 & ~n14818 ) | ( n3565 & n16773 ) | ( ~n14818 & n16773 ) ;
  assign n26902 = n26901 ^ n17135 ^ 1'b0 ;
  assign n26903 = ( n8164 & ~n13333 ) | ( n8164 & n13648 ) | ( ~n13333 & n13648 ) ;
  assign n26904 = n26020 ^ n9271 ^ n4659 ;
  assign n26905 = ( x179 & n23576 ) | ( x179 & ~n26904 ) | ( n23576 & ~n26904 ) ;
  assign n26906 = n20225 ^ n1198 ^ 1'b0 ;
  assign n26907 = n2030 | n26906 ;
  assign n26908 = n26907 ^ n20730 ^ n4917 ;
  assign n26909 = ~n15499 & n26908 ;
  assign n26915 = x207 & ~n20073 ;
  assign n26916 = n26915 ^ n6987 ^ 1'b0 ;
  assign n26910 = n22268 ^ n2470 ^ 1'b0 ;
  assign n26911 = ( n7352 & n15926 ) | ( n7352 & n26910 ) | ( n15926 & n26910 ) ;
  assign n26912 = ~n7703 & n24693 ;
  assign n26913 = n8806 & n26912 ;
  assign n26914 = ( n1680 & n26911 ) | ( n1680 & n26913 ) | ( n26911 & n26913 ) ;
  assign n26917 = n26916 ^ n26914 ^ n12486 ;
  assign n26921 = n4797 & n9132 ;
  assign n26922 = n26921 ^ n4818 ^ 1'b0 ;
  assign n26918 = n13333 ^ n12176 ^ n11653 ;
  assign n26919 = n25377 ^ n14998 ^ 1'b0 ;
  assign n26920 = ~n26918 & n26919 ;
  assign n26923 = n26922 ^ n26920 ^ n9358 ;
  assign n26924 = n17635 ^ n8190 ^ n1346 ;
  assign n26925 = n25305 ^ n11849 ^ 1'b0 ;
  assign n26926 = ( n13515 & n26924 ) | ( n13515 & ~n26925 ) | ( n26924 & ~n26925 ) ;
  assign n26927 = ( ~n1581 & n4883 ) | ( ~n1581 & n13027 ) | ( n4883 & n13027 ) ;
  assign n26928 = n26927 ^ n16049 ^ 1'b0 ;
  assign n26929 = ~n1460 & n14833 ;
  assign n26930 = ~n16239 & n26929 ;
  assign n26931 = n23782 ^ n20720 ^ n858 ;
  assign n26932 = ~n11866 & n13284 ;
  assign n26933 = n26932 ^ n20669 ^ 1'b0 ;
  assign n26934 = ( n11922 & n13306 ) | ( n11922 & ~n26933 ) | ( n13306 & ~n26933 ) ;
  assign n26935 = ( x228 & n15729 ) | ( x228 & n18120 ) | ( n15729 & n18120 ) ;
  assign n26936 = n5014 | n26935 ;
  assign n26937 = n26936 ^ n15796 ^ 1'b0 ;
  assign n26939 = n20354 ^ n14697 ^ n7296 ;
  assign n26938 = n2250 | n7345 ;
  assign n26940 = n26939 ^ n26938 ^ 1'b0 ;
  assign n26941 = n18916 | n26940 ;
  assign n26942 = n16964 ^ n15321 ^ n360 ;
  assign n26943 = n4478 & n16443 ;
  assign n26944 = n5831 | n18352 ;
  assign n26945 = ~n5054 & n26944 ;
  assign n26946 = ( ~n15190 & n26943 ) | ( ~n15190 & n26945 ) | ( n26943 & n26945 ) ;
  assign n26947 = n10904 ^ n5093 ^ 1'b0 ;
  assign n26953 = n6031 & n6390 ;
  assign n26950 = n14873 | n15486 ;
  assign n26951 = n26950 ^ n12829 ^ n11885 ;
  assign n26952 = ( n12263 & ~n22840 ) | ( n12263 & n26951 ) | ( ~n22840 & n26951 ) ;
  assign n26948 = ( n7385 & n10306 ) | ( n7385 & ~n18008 ) | ( n10306 & ~n18008 ) ;
  assign n26949 = n26948 ^ n6825 ^ 1'b0 ;
  assign n26954 = n26953 ^ n26952 ^ n26949 ;
  assign n26955 = n5760 | n7722 ;
  assign n26956 = n26955 ^ n9630 ^ 1'b0 ;
  assign n26957 = ~n8459 & n26956 ;
  assign n26958 = n26957 ^ n8287 ^ 1'b0 ;
  assign n26960 = ~n4656 & n5284 ;
  assign n26961 = n26960 ^ n3339 ^ 1'b0 ;
  assign n26959 = n13874 & n17733 ;
  assign n26962 = n26961 ^ n26959 ^ 1'b0 ;
  assign n26963 = ( n19624 & n26958 ) | ( n19624 & ~n26962 ) | ( n26958 & ~n26962 ) ;
  assign n26964 = n4836 & n14369 ;
  assign n26965 = n26963 & n26964 ;
  assign n26966 = n24817 ^ n11541 ^ n4379 ;
  assign n26967 = ( n3247 & n9437 ) | ( n3247 & ~n11439 ) | ( n9437 & ~n11439 ) ;
  assign n26968 = ~n24555 & n26967 ;
  assign n26969 = n23651 ^ n17333 ^ n7641 ;
  assign n26970 = ( n705 & n18703 ) | ( n705 & n26673 ) | ( n18703 & n26673 ) ;
  assign n26971 = n23667 | n26970 ;
  assign n26972 = ( ~n3172 & n6642 ) | ( ~n3172 & n13109 ) | ( n6642 & n13109 ) ;
  assign n26973 = ( ~n4040 & n15548 ) | ( ~n4040 & n26972 ) | ( n15548 & n26972 ) ;
  assign n26982 = n19370 ^ n17198 ^ 1'b0 ;
  assign n26983 = n8072 & ~n26982 ;
  assign n26979 = ( n4175 & n4431 ) | ( n4175 & n7637 ) | ( n4431 & n7637 ) ;
  assign n26980 = n13265 ^ n6686 ^ 1'b0 ;
  assign n26981 = n26979 & ~n26980 ;
  assign n26974 = n3720 ^ n3106 ^ 1'b0 ;
  assign n26975 = n1271 & ~n26974 ;
  assign n26976 = ~n7536 & n26975 ;
  assign n26977 = ~n7664 & n26976 ;
  assign n26978 = n9131 & n26977 ;
  assign n26984 = n26983 ^ n26981 ^ n26978 ;
  assign n26985 = ~n3898 & n10000 ;
  assign n26986 = n17465 ^ n6584 ^ 1'b0 ;
  assign n26987 = n7144 & n26986 ;
  assign n26988 = n26287 ^ n4544 ^ 1'b0 ;
  assign n26989 = n26987 & n26988 ;
  assign n26990 = n26989 ^ n15402 ^ 1'b0 ;
  assign n26991 = n26990 ^ n2070 ^ 1'b0 ;
  assign n26994 = n24005 ^ n10935 ^ n1685 ;
  assign n26992 = n736 | n3119 ;
  assign n26993 = ~n3159 & n26992 ;
  assign n26995 = n26994 ^ n26993 ^ 1'b0 ;
  assign n26996 = n26995 ^ n20673 ^ n2163 ;
  assign n26997 = ( n22740 & n26991 ) | ( n22740 & n26996 ) | ( n26991 & n26996 ) ;
  assign n26998 = n14985 & ~n15438 ;
  assign n26999 = ~n1301 & n4322 ;
  assign n27000 = n26999 ^ n1644 ^ 1'b0 ;
  assign n27001 = n27000 ^ n16347 ^ 1'b0 ;
  assign n27002 = ~n934 & n27001 ;
  assign n27003 = n20184 ^ n2598 ^ 1'b0 ;
  assign n27007 = n10268 ^ n6218 ^ x240 ;
  assign n27004 = ~n3538 & n21276 ;
  assign n27005 = ( n13082 & ~n21833 ) | ( n13082 & n27004 ) | ( ~n21833 & n27004 ) ;
  assign n27006 = n17815 | n27005 ;
  assign n27008 = n27007 ^ n27006 ^ n6558 ;
  assign n27009 = n24268 & n27008 ;
  assign n27010 = n1656 ^ n550 ^ 1'b0 ;
  assign n27011 = ( ~n9930 & n24514 ) | ( ~n9930 & n27010 ) | ( n24514 & n27010 ) ;
  assign n27012 = n5725 | n6110 ;
  assign n27013 = n12739 & ~n27012 ;
  assign n27014 = n989 & n5195 ;
  assign n27015 = n27013 & n27014 ;
  assign n27016 = n27015 ^ n22154 ^ n13363 ;
  assign n27018 = n10777 ^ n550 ^ 1'b0 ;
  assign n27017 = n18421 ^ n3991 ^ 1'b0 ;
  assign n27019 = n27018 ^ n27017 ^ n15899 ;
  assign n27020 = n10077 & ~n18771 ;
  assign n27021 = n27020 ^ n25987 ^ n4210 ;
  assign n27022 = n23457 ^ n5368 ^ 1'b0 ;
  assign n27023 = n27022 ^ n12219 ^ 1'b0 ;
  assign n27024 = ~n8374 & n27023 ;
  assign n27025 = n9693 | n25807 ;
  assign n27026 = n2592 | n8729 ;
  assign n27027 = n27026 ^ n18894 ^ 1'b0 ;
  assign n27028 = n25921 & n27027 ;
  assign n27033 = n10379 & ~n13670 ;
  assign n27034 = n27033 ^ n5010 ^ n4074 ;
  assign n27035 = ( ~n5183 & n11758 ) | ( ~n5183 & n27034 ) | ( n11758 & n27034 ) ;
  assign n27031 = n8917 & ~n11149 ;
  assign n27032 = n12255 & n27031 ;
  assign n27029 = n12503 ^ n11381 ^ n502 ;
  assign n27030 = n27029 ^ n7391 ^ 1'b0 ;
  assign n27036 = n27035 ^ n27032 ^ n27030 ;
  assign n27037 = ~n7862 & n11588 ;
  assign n27038 = n27037 ^ n14821 ^ n12982 ;
  assign n27039 = n23404 & ~n23736 ;
  assign n27040 = n14552 ^ n9519 ^ n1227 ;
  assign n27041 = n27040 ^ n6382 ^ n4645 ;
  assign n27042 = ( x156 & n7259 ) | ( x156 & n27041 ) | ( n7259 & n27041 ) ;
  assign n27043 = ( n3499 & n13807 ) | ( n3499 & n20707 ) | ( n13807 & n20707 ) ;
  assign n27044 = ~n11265 & n20393 ;
  assign n27045 = n27044 ^ n7125 ^ 1'b0 ;
  assign n27046 = n11151 ^ n6425 ^ n3306 ;
  assign n27047 = n1526 & n3428 ;
  assign n27048 = n27047 ^ n17211 ^ 1'b0 ;
  assign n27049 = n20483 ^ n4991 ^ 1'b0 ;
  assign n27050 = n8203 & n11653 ;
  assign n27051 = n27049 & n27050 ;
  assign n27052 = n27051 ^ n5885 ^ 1'b0 ;
  assign n27053 = ( n27046 & n27048 ) | ( n27046 & n27052 ) | ( n27048 & n27052 ) ;
  assign n27054 = n16813 & ~n20073 ;
  assign n27055 = ( ~n7913 & n11492 ) | ( ~n7913 & n27054 ) | ( n11492 & n27054 ) ;
  assign n27056 = ( n7417 & n18064 ) | ( n7417 & ~n27055 ) | ( n18064 & ~n27055 ) ;
  assign n27057 = ( ~n10594 & n19885 ) | ( ~n10594 & n27056 ) | ( n19885 & n27056 ) ;
  assign n27058 = n2354 & n6873 ;
  assign n27059 = n27058 ^ n10609 ^ 1'b0 ;
  assign n27060 = n27057 & n27059 ;
  assign n27061 = n4295 & n6184 ;
  assign n27062 = n27061 ^ n8184 ^ 1'b0 ;
  assign n27063 = n11749 | n27062 ;
  assign n27064 = n11319 & n27063 ;
  assign n27065 = n22134 ^ n12899 ^ n3860 ;
  assign n27066 = n27065 ^ n10610 ^ 1'b0 ;
  assign n27067 = ~n8741 & n27066 ;
  assign n27068 = ~n3129 & n18560 ;
  assign n27069 = n20766 ^ n12197 ^ n9940 ;
  assign n27070 = n27069 ^ n3028 ^ 1'b0 ;
  assign n27079 = n3991 ^ n2584 ^ n2183 ;
  assign n27080 = n9017 ^ n2850 ^ 1'b0 ;
  assign n27081 = n27079 | n27080 ;
  assign n27071 = ~n451 & n2248 ;
  assign n27072 = n27071 ^ n1291 ^ 1'b0 ;
  assign n27073 = n17530 ^ n10874 ^ 1'b0 ;
  assign n27074 = n9972 & ~n27073 ;
  assign n27075 = n9725 & ~n15548 ;
  assign n27076 = ( ~n27072 & n27074 ) | ( ~n27072 & n27075 ) | ( n27074 & n27075 ) ;
  assign n27077 = n17152 & n27076 ;
  assign n27078 = ~n1264 & n27077 ;
  assign n27082 = n27081 ^ n27078 ^ n6628 ;
  assign n27083 = ( ~n625 & n12213 ) | ( ~n625 & n14605 ) | ( n12213 & n14605 ) ;
  assign n27084 = n17851 ^ n15224 ^ n10021 ;
  assign n27085 = n3765 | n27084 ;
  assign n27086 = ( n833 & ~n9197 ) | ( n833 & n18605 ) | ( ~n9197 & n18605 ) ;
  assign n27087 = ( ~n9984 & n26935 ) | ( ~n9984 & n27086 ) | ( n26935 & n27086 ) ;
  assign n27088 = n21949 ^ n11579 ^ 1'b0 ;
  assign n27089 = n27088 ^ n26033 ^ n3408 ;
  assign n27090 = n461 & n3058 ;
  assign n27091 = n5516 & ~n27090 ;
  assign n27092 = ~x59 & n27091 ;
  assign n27093 = n27092 ^ n10172 ^ n2353 ;
  assign n27094 = n4601 & ~n27093 ;
  assign n27095 = ~n2072 & n27094 ;
  assign n27096 = n5953 | n7137 ;
  assign n27097 = n5821 | n27096 ;
  assign n27100 = ( ~n1536 & n2671 ) | ( ~n1536 & n3863 ) | ( n2671 & n3863 ) ;
  assign n27098 = x178 & n5197 ;
  assign n27099 = ~n14657 & n27098 ;
  assign n27101 = n27100 ^ n27099 ^ n20897 ;
  assign n27102 = ~n14696 & n27101 ;
  assign n27103 = ~n3718 & n26472 ;
  assign n27104 = n27103 ^ x31 ^ 1'b0 ;
  assign n27105 = ( ~n489 & n6325 ) | ( ~n489 & n8539 ) | ( n6325 & n8539 ) ;
  assign n27106 = ( n22889 & n27104 ) | ( n22889 & n27105 ) | ( n27104 & n27105 ) ;
  assign n27107 = n6493 & ~n21188 ;
  assign n27108 = ~n12216 & n27107 ;
  assign n27109 = ( n2536 & n16113 ) | ( n2536 & n27108 ) | ( n16113 & n27108 ) ;
  assign n27110 = n27109 ^ n12515 ^ n6889 ;
  assign n27112 = n10260 ^ x106 ^ 1'b0 ;
  assign n27111 = n12194 & ~n15230 ;
  assign n27113 = n27112 ^ n27111 ^ 1'b0 ;
  assign n27114 = n20787 ^ n11353 ^ 1'b0 ;
  assign n27115 = n21720 & n27114 ;
  assign n27116 = n1651 | n18707 ;
  assign n27117 = n27116 ^ n11906 ^ 1'b0 ;
  assign n27118 = n27117 ^ n23482 ^ n9412 ;
  assign n27119 = n3444 | n23026 ;
  assign n27120 = n27119 ^ n25046 ^ 1'b0 ;
  assign n27121 = n9858 | n9872 ;
  assign n27122 = n8199 & n27121 ;
  assign n27123 = n25250 ^ n24058 ^ 1'b0 ;
  assign n27124 = n27122 | n27123 ;
  assign n27125 = n9096 ^ n6911 ^ n3333 ;
  assign n27126 = n27125 ^ n6661 ^ n4409 ;
  assign n27127 = n10874 ^ n5376 ^ 1'b0 ;
  assign n27128 = n7795 & ~n23041 ;
  assign n27129 = n27127 & ~n27128 ;
  assign n27130 = n1582 & n6389 ;
  assign n27131 = ~x130 & n27130 ;
  assign n27132 = ( n9412 & n24893 ) | ( n9412 & ~n27131 ) | ( n24893 & ~n27131 ) ;
  assign n27133 = ( n15075 & ~n17231 ) | ( n15075 & n24830 ) | ( ~n17231 & n24830 ) ;
  assign n27134 = n821 & ~n27133 ;
  assign n27135 = n21665 ^ n3421 ^ 1'b0 ;
  assign n27136 = ~n7498 & n27135 ;
  assign n27137 = n27136 ^ n23174 ^ 1'b0 ;
  assign n27138 = n5712 ^ n1385 ^ 1'b0 ;
  assign n27139 = n10281 | n27138 ;
  assign n27140 = n1794 | n27139 ;
  assign n27141 = ( n6671 & n27137 ) | ( n6671 & n27140 ) | ( n27137 & n27140 ) ;
  assign n27142 = n27141 ^ n3952 ^ 1'b0 ;
  assign n27143 = n20013 ^ n1777 ^ 1'b0 ;
  assign n27144 = n17136 & ~n27143 ;
  assign n27145 = n20081 ^ n5881 ^ x124 ;
  assign n27146 = n18135 & ~n27145 ;
  assign n27147 = ~n27144 & n27146 ;
  assign n27148 = n27147 ^ n20557 ^ n12814 ;
  assign n27149 = ~n21820 & n27148 ;
  assign n27150 = n12999 & ~n18226 ;
  assign n27151 = ~x84 & n27150 ;
  assign n27152 = ( ~n4297 & n7181 ) | ( ~n4297 & n22706 ) | ( n7181 & n22706 ) ;
  assign n27153 = n3471 & n16075 ;
  assign n27154 = ~n7171 & n27153 ;
  assign n27155 = n27154 ^ n14924 ^ 1'b0 ;
  assign n27156 = n27152 & ~n27155 ;
  assign n27157 = n27156 ^ n12494 ^ 1'b0 ;
  assign n27160 = n13915 ^ n9069 ^ n3132 ;
  assign n27158 = n8944 ^ n5294 ^ 1'b0 ;
  assign n27159 = n4775 | n27158 ;
  assign n27161 = n27160 ^ n27159 ^ 1'b0 ;
  assign n27162 = n27161 ^ n14966 ^ n6173 ;
  assign n27163 = n14811 & n27162 ;
  assign n27164 = n27163 ^ n9524 ^ n620 ;
  assign n27165 = n12692 ^ n2530 ^ n1979 ;
  assign n27166 = n11702 | n27165 ;
  assign n27167 = ~n22609 & n27166 ;
  assign n27171 = n9192 ^ n8903 ^ 1'b0 ;
  assign n27168 = n521 & ~n6989 ;
  assign n27169 = ~n8272 & n27168 ;
  assign n27170 = n26750 & ~n27169 ;
  assign n27172 = n27171 ^ n27170 ^ 1'b0 ;
  assign n27173 = n25378 ^ n21256 ^ n15235 ;
  assign n27174 = ( n13100 & n24565 ) | ( n13100 & n27173 ) | ( n24565 & n27173 ) ;
  assign n27175 = n10081 ^ n8784 ^ n2149 ;
  assign n27176 = n9013 ^ n6186 ^ 1'b0 ;
  assign n27177 = ~n5595 & n27176 ;
  assign n27178 = n16057 & ~n18630 ;
  assign n27179 = ~n21148 & n27178 ;
  assign n27181 = n11158 ^ n8280 ^ n2935 ;
  assign n27182 = ( ~n2547 & n15360 ) | ( ~n2547 & n27181 ) | ( n15360 & n27181 ) ;
  assign n27180 = ~n10788 & n17256 ;
  assign n27183 = n27182 ^ n27180 ^ 1'b0 ;
  assign n27184 = ~n25754 & n27183 ;
  assign n27185 = n20404 ^ n15252 ^ n2552 ;
  assign n27186 = n27185 ^ n2550 ^ 1'b0 ;
  assign n27187 = n22470 ^ n10081 ^ 1'b0 ;
  assign n27188 = ( n7489 & n8897 ) | ( n7489 & n19446 ) | ( n8897 & n19446 ) ;
  assign n27189 = ( n592 & ~n27187 ) | ( n592 & n27188 ) | ( ~n27187 & n27188 ) ;
  assign n27190 = n12833 & ~n12835 ;
  assign n27191 = x77 & n4117 ;
  assign n27192 = n5141 & n27191 ;
  assign n27193 = n11570 ^ n5522 ^ n494 ;
  assign n27194 = ~n6995 & n27193 ;
  assign n27195 = n27192 & n27194 ;
  assign n27196 = n27195 ^ n25717 ^ n14260 ;
  assign n27197 = n27196 ^ n15095 ^ 1'b0 ;
  assign n27198 = ~n7459 & n27197 ;
  assign n27201 = ( n1232 & ~n9087 ) | ( n1232 & n12676 ) | ( ~n9087 & n12676 ) ;
  assign n27202 = n6776 & ~n11908 ;
  assign n27203 = n27202 ^ n13078 ^ 1'b0 ;
  assign n27204 = n27201 & ~n27203 ;
  assign n27205 = ( n3608 & ~n8416 ) | ( n3608 & n27204 ) | ( ~n8416 & n27204 ) ;
  assign n27206 = n27205 ^ n3123 ^ 1'b0 ;
  assign n27199 = n15039 & ~n15968 ;
  assign n27200 = n27199 ^ n844 ^ 1'b0 ;
  assign n27207 = n27206 ^ n27200 ^ 1'b0 ;
  assign n27208 = n5378 & n27207 ;
  assign n27209 = ( n2127 & n20135 ) | ( n2127 & ~n21768 ) | ( n20135 & ~n21768 ) ;
  assign n27210 = ( ~n1148 & n2744 ) | ( ~n1148 & n24699 ) | ( n2744 & n24699 ) ;
  assign n27211 = n27210 ^ n13264 ^ 1'b0 ;
  assign n27212 = n27209 | n27211 ;
  assign n27213 = n687 | n27212 ;
  assign n27214 = n27208 | n27213 ;
  assign n27215 = ~n26348 & n27214 ;
  assign n27216 = n7388 & n26505 ;
  assign n27217 = n13547 ^ n2760 ^ 1'b0 ;
  assign n27218 = ~n2337 & n5050 ;
  assign n27219 = n27218 ^ n23993 ^ n22039 ;
  assign n27220 = n22896 ^ n2359 ^ 1'b0 ;
  assign n27221 = n27219 | n27220 ;
  assign n27222 = n5860 | n12868 ;
  assign n27223 = n9238 ^ n8187 ^ 1'b0 ;
  assign n27224 = n481 & ~n27223 ;
  assign n27225 = n15389 & n27224 ;
  assign n27226 = n27225 ^ n13846 ^ 1'b0 ;
  assign n27227 = n1308 & ~n27226 ;
  assign n27228 = ( n16496 & n27222 ) | ( n16496 & n27227 ) | ( n27222 & n27227 ) ;
  assign n27229 = n14205 ^ n13087 ^ 1'b0 ;
  assign n27230 = ~n11961 & n27229 ;
  assign n27234 = n22150 ^ n19359 ^ n19174 ;
  assign n27231 = ( n2999 & n9642 ) | ( n2999 & n16927 ) | ( n9642 & n16927 ) ;
  assign n27232 = n22665 ^ n17668 ^ 1'b0 ;
  assign n27233 = n27231 | n27232 ;
  assign n27235 = n27234 ^ n27233 ^ n7207 ;
  assign n27236 = n22476 ^ n19912 ^ n19430 ;
  assign n27239 = n13816 ^ n8826 ^ 1'b0 ;
  assign n27237 = ( n3796 & n5604 ) | ( n3796 & ~n25057 ) | ( n5604 & ~n25057 ) ;
  assign n27238 = ~n14051 & n27237 ;
  assign n27240 = n27239 ^ n27238 ^ 1'b0 ;
  assign n27241 = n27240 ^ n24566 ^ n14093 ;
  assign n27242 = n11375 ^ n2956 ^ x137 ;
  assign n27243 = n7535 & n13801 ;
  assign n27244 = n27243 ^ n8721 ^ 1'b0 ;
  assign n27245 = ~n6222 & n11748 ;
  assign n27246 = n9883 & n27245 ;
  assign n27247 = n27246 ^ n16796 ^ n12188 ;
  assign n27248 = ( ~n4841 & n21661 ) | ( ~n4841 & n27247 ) | ( n21661 & n27247 ) ;
  assign n27249 = n27244 | n27248 ;
  assign n27250 = n13707 & n27249 ;
  assign n27251 = ~n12602 & n27250 ;
  assign n27252 = n5708 & ~n8562 ;
  assign n27253 = ~n5125 & n13831 ;
  assign n27258 = n20596 & ~n21289 ;
  assign n27259 = ~n14076 & n27258 ;
  assign n27254 = n20734 ^ n13616 ^ n12238 ;
  assign n27255 = ( n5025 & n12542 ) | ( n5025 & ~n27254 ) | ( n12542 & ~n27254 ) ;
  assign n27256 = n9508 ^ n6797 ^ 1'b0 ;
  assign n27257 = n27255 & n27256 ;
  assign n27260 = n27259 ^ n27257 ^ n21002 ;
  assign n27261 = n5654 ^ n4458 ^ n3905 ;
  assign n27262 = n18570 ^ n13594 ^ 1'b0 ;
  assign n27263 = n2338 & n19760 ;
  assign n27264 = ~n8591 & n27263 ;
  assign n27265 = n9009 & n9246 ;
  assign n27266 = n27265 ^ n13639 ^ 1'b0 ;
  assign n27267 = ~n539 & n27266 ;
  assign n27268 = n27267 ^ n5930 ^ 1'b0 ;
  assign n27269 = ( n9441 & ~n11622 ) | ( n9441 & n13594 ) | ( ~n11622 & n13594 ) ;
  assign n27270 = ( n4460 & n16538 ) | ( n4460 & n27269 ) | ( n16538 & n27269 ) ;
  assign n27271 = n27270 ^ n18091 ^ 1'b0 ;
  assign n27272 = n5495 | n5732 ;
  assign n27273 = ( ~n9083 & n9496 ) | ( ~n9083 & n9804 ) | ( n9496 & n9804 ) ;
  assign n27274 = n27273 ^ n5121 ^ 1'b0 ;
  assign n27275 = n17087 ^ n14219 ^ n467 ;
  assign n27276 = ( n7885 & n14307 ) | ( n7885 & ~n27275 ) | ( n14307 & ~n27275 ) ;
  assign n27277 = n10577 ^ n9016 ^ n2335 ;
  assign n27278 = n27277 ^ n10160 ^ 1'b0 ;
  assign n27279 = n27276 | n27278 ;
  assign n27280 = n22957 ^ n9667 ^ 1'b0 ;
  assign n27281 = n2114 | n27280 ;
  assign n27282 = n27148 | n27281 ;
  assign n27283 = n27282 ^ n18173 ^ 1'b0 ;
  assign n27284 = ( n5387 & n6913 ) | ( n5387 & n6915 ) | ( n6913 & n6915 ) ;
  assign n27285 = n24256 ^ n11697 ^ n10823 ;
  assign n27286 = n10001 & ~n27285 ;
  assign n27287 = n633 & ~n4220 ;
  assign n27288 = ~n7685 & n27287 ;
  assign n27289 = n6368 & ~n27288 ;
  assign n27290 = n27289 ^ n16296 ^ n5311 ;
  assign n27291 = n4056 & ~n5175 ;
  assign n27292 = n10742 & n17498 ;
  assign n27293 = n1434 & n27292 ;
  assign n27294 = ( n23452 & ~n26310 ) | ( n23452 & n27293 ) | ( ~n26310 & n27293 ) ;
  assign n27295 = n15824 & ~n27294 ;
  assign n27296 = n27291 & n27295 ;
  assign n27297 = ~n11022 & n22453 ;
  assign n27298 = ~n6386 & n27297 ;
  assign n27299 = n9342 ^ n4294 ^ n2763 ;
  assign n27300 = ( ~n14813 & n26321 ) | ( ~n14813 & n27299 ) | ( n26321 & n27299 ) ;
  assign n27301 = n5529 & ~n7295 ;
  assign n27304 = n4245 | n6407 ;
  assign n27305 = n4038 | n27304 ;
  assign n27306 = ( ~n1885 & n8749 ) | ( ~n1885 & n27305 ) | ( n8749 & n27305 ) ;
  assign n27307 = n27306 ^ n19344 ^ 1'b0 ;
  assign n27302 = n17678 ^ n6364 ^ x65 ;
  assign n27303 = ( n5726 & n23310 ) | ( n5726 & ~n27302 ) | ( n23310 & ~n27302 ) ;
  assign n27308 = n27307 ^ n27303 ^ n23459 ;
  assign n27309 = n8763 & ~n15812 ;
  assign n27310 = n19486 & n27309 ;
  assign n27311 = ( n17292 & n22194 ) | ( n17292 & ~n27310 ) | ( n22194 & ~n27310 ) ;
  assign n27312 = ( n2184 & ~n6586 ) | ( n2184 & n13082 ) | ( ~n6586 & n13082 ) ;
  assign n27313 = n4063 & ~n27312 ;
  assign n27314 = n5048 & n12931 ;
  assign n27315 = ~n4568 & n27314 ;
  assign n27316 = ~n10641 & n27315 ;
  assign n27317 = n15357 | n27316 ;
  assign n27318 = n27317 ^ n7223 ^ 1'b0 ;
  assign n27319 = ( n10691 & ~n18532 ) | ( n10691 & n23423 ) | ( ~n18532 & n23423 ) ;
  assign n27320 = ( n10432 & n16812 ) | ( n10432 & n27319 ) | ( n16812 & n27319 ) ;
  assign n27324 = n15180 ^ n6849 ^ n3564 ;
  assign n27321 = n23888 ^ n8928 ^ 1'b0 ;
  assign n27322 = n13573 | n27321 ;
  assign n27323 = ( ~n2440 & n7172 ) | ( ~n2440 & n27322 ) | ( n7172 & n27322 ) ;
  assign n27325 = n27324 ^ n27323 ^ n458 ;
  assign n27326 = n23301 ^ n19980 ^ n11099 ;
  assign n27327 = n21132 ^ n3200 ^ 1'b0 ;
  assign n27328 = ( n9802 & ~n21309 ) | ( n9802 & n27327 ) | ( ~n21309 & n27327 ) ;
  assign n27329 = ( n13291 & n15256 ) | ( n13291 & ~n27328 ) | ( n15256 & ~n27328 ) ;
  assign n27330 = n10725 & n13126 ;
  assign n27331 = n27330 ^ n1885 ^ 1'b0 ;
  assign n27332 = n18644 & ~n27331 ;
  assign n27333 = n24581 ^ n16985 ^ 1'b0 ;
  assign n27334 = n21987 ^ n12461 ^ n511 ;
  assign n27335 = n10980 ^ n3206 ^ n477 ;
  assign n27336 = n14516 & n27335 ;
  assign n27337 = n27336 ^ n2558 ^ 1'b0 ;
  assign n27338 = n27337 ^ n14234 ^ 1'b0 ;
  assign n27339 = ~n8064 & n27338 ;
  assign n27340 = n27334 | n27339 ;
  assign n27341 = ~n21891 & n27340 ;
  assign n27342 = ~n27333 & n27341 ;
  assign n27343 = n21847 ^ n7658 ^ n4984 ;
  assign n27344 = n22146 ^ n920 ^ 1'b0 ;
  assign n27345 = ~n6086 & n27344 ;
  assign n27346 = n4814 & n27345 ;
  assign n27347 = ( n3979 & ~n27343 ) | ( n3979 & n27346 ) | ( ~n27343 & n27346 ) ;
  assign n27348 = n3397 & n6591 ;
  assign n27349 = n27348 ^ n10263 ^ 1'b0 ;
  assign n27350 = n25473 & ~n26188 ;
  assign n27351 = n6491 & ~n24454 ;
  assign n27352 = ~n2259 & n11709 ;
  assign n27353 = ~n5403 & n27352 ;
  assign n27354 = ( n5524 & ~n27351 ) | ( n5524 & n27353 ) | ( ~n27351 & n27353 ) ;
  assign n27355 = n27354 ^ n7294 ^ 1'b0 ;
  assign n27356 = ~n7822 & n27355 ;
  assign n27357 = n27356 ^ n13680 ^ 1'b0 ;
  assign n27358 = n27350 & ~n27357 ;
  assign n27359 = n8011 ^ n7089 ^ 1'b0 ;
  assign n27360 = n27359 ^ n11585 ^ 1'b0 ;
  assign n27361 = n6867 & ~n12473 ;
  assign n27362 = n27360 & n27361 ;
  assign n27363 = n15883 ^ n9852 ^ 1'b0 ;
  assign n27364 = n1505 & n27363 ;
  assign n27365 = ~n22286 & n27364 ;
  assign n27366 = n8423 ^ n7637 ^ 1'b0 ;
  assign n27367 = ~n27365 & n27366 ;
  assign n27368 = ( n3764 & n9394 ) | ( n3764 & n13043 ) | ( n9394 & n13043 ) ;
  assign n27369 = ( ~n8338 & n21058 ) | ( ~n8338 & n25142 ) | ( n21058 & n25142 ) ;
  assign n27371 = n7009 ^ n792 ^ 1'b0 ;
  assign n27372 = ( n2338 & n22218 ) | ( n2338 & n27371 ) | ( n22218 & n27371 ) ;
  assign n27370 = ( n10027 & n18484 ) | ( n10027 & n23503 ) | ( n18484 & n23503 ) ;
  assign n27373 = n27372 ^ n27370 ^ n20604 ;
  assign n27376 = ( n4248 & ~n4793 ) | ( n4248 & n20403 ) | ( ~n4793 & n20403 ) ;
  assign n27374 = n18434 | n24891 ;
  assign n27375 = n10602 | n27374 ;
  assign n27377 = n27376 ^ n27375 ^ 1'b0 ;
  assign n27381 = n15304 ^ n4716 ^ n3603 ;
  assign n27380 = ( n4962 & n8160 ) | ( n4962 & n26687 ) | ( n8160 & n26687 ) ;
  assign n27378 = n7136 & n7675 ;
  assign n27379 = n27378 ^ n6503 ^ n3184 ;
  assign n27382 = n27381 ^ n27380 ^ n27379 ;
  assign n27383 = x240 & n3475 ;
  assign n27384 = ~x146 & n27383 ;
  assign n27385 = n27384 ^ n4711 ^ n3117 ;
  assign n27386 = n4768 | n6681 ;
  assign n27387 = ( n2777 & n14756 ) | ( n2777 & n27386 ) | ( n14756 & n27386 ) ;
  assign n27388 = ( ~n6977 & n22529 ) | ( ~n6977 & n25882 ) | ( n22529 & n25882 ) ;
  assign n27389 = n10552 ^ n660 ^ x194 ;
  assign n27390 = n27389 ^ n14923 ^ 1'b0 ;
  assign n27391 = n12297 & n27390 ;
  assign n27392 = n22922 ^ n2883 ^ n1319 ;
  assign n27393 = n27392 ^ n24154 ^ n21377 ;
  assign n27394 = ( n16675 & ~n19374 ) | ( n16675 & n27393 ) | ( ~n19374 & n27393 ) ;
  assign n27395 = n12446 & n26909 ;
  assign n27396 = ~n20729 & n27395 ;
  assign n27397 = n9050 ^ n7479 ^ 1'b0 ;
  assign n27398 = n9438 ^ n258 ^ 1'b0 ;
  assign n27399 = ~n20457 & n27398 ;
  assign n27400 = n14657 ^ n5712 ^ 1'b0 ;
  assign n27401 = n27399 & n27400 ;
  assign n27402 = n27401 ^ n22627 ^ n3126 ;
  assign n27403 = ( n16898 & n17731 ) | ( n16898 & n22674 ) | ( n17731 & n22674 ) ;
  assign n27405 = n14136 ^ n5478 ^ 1'b0 ;
  assign n27406 = ( n4275 & n19423 ) | ( n4275 & ~n27405 ) | ( n19423 & ~n27405 ) ;
  assign n27404 = n26275 ^ n13107 ^ n7934 ;
  assign n27407 = n27406 ^ n27404 ^ n8093 ;
  assign n27408 = n15070 ^ n13345 ^ n11059 ;
  assign n27409 = n14472 ^ n5700 ^ 1'b0 ;
  assign n27410 = ( n2208 & n27408 ) | ( n2208 & ~n27409 ) | ( n27408 & ~n27409 ) ;
  assign n27411 = n27410 ^ n16739 ^ n419 ;
  assign n27412 = n20571 ^ n15589 ^ n9007 ;
  assign n27413 = n22963 ^ n16573 ^ 1'b0 ;
  assign n27414 = n17172 ^ n6567 ^ n6004 ;
  assign n27415 = n2624 & n9007 ;
  assign n27416 = n27415 ^ n12729 ^ 1'b0 ;
  assign n27418 = n17377 ^ n6768 ^ 1'b0 ;
  assign n27419 = n10677 & ~n27418 ;
  assign n27417 = n13791 ^ n4121 ^ 1'b0 ;
  assign n27420 = n27419 ^ n27417 ^ n11440 ;
  assign n27421 = n2120 | n27420 ;
  assign n27422 = n27421 ^ n13652 ^ 1'b0 ;
  assign n27426 = n12703 ^ n10864 ^ n4085 ;
  assign n27424 = n13240 ^ n4448 ^ 1'b0 ;
  assign n27423 = ( n10048 & n12080 ) | ( n10048 & ~n15522 ) | ( n12080 & ~n15522 ) ;
  assign n27425 = n27424 ^ n27423 ^ 1'b0 ;
  assign n27427 = n27426 ^ n27425 ^ n7480 ;
  assign n27428 = ( n3834 & n25421 ) | ( n3834 & n27427 ) | ( n25421 & n27427 ) ;
  assign n27429 = ( n1479 & ~n12113 ) | ( n1479 & n16255 ) | ( ~n12113 & n16255 ) ;
  assign n27430 = n664 | n23446 ;
  assign n27431 = n27430 ^ n7958 ^ 1'b0 ;
  assign n27432 = n25500 & n27431 ;
  assign n27433 = n11966 ^ n7922 ^ n1643 ;
  assign n27434 = n17169 ^ n5919 ^ n4942 ;
  assign n27435 = ( n6313 & n25694 ) | ( n6313 & n27434 ) | ( n25694 & n27434 ) ;
  assign n27436 = ( n979 & n23583 ) | ( n979 & n23868 ) | ( n23583 & n23868 ) ;
  assign n27442 = ( n6153 & n6345 ) | ( n6153 & n6558 ) | ( n6345 & n6558 ) ;
  assign n27443 = n27442 ^ n21840 ^ n12332 ;
  assign n27437 = ( n2707 & n6251 ) | ( n2707 & ~n17678 ) | ( n6251 & ~n17678 ) ;
  assign n27438 = n14435 ^ n11991 ^ n4660 ;
  assign n27439 = n27437 & ~n27438 ;
  assign n27440 = n27439 ^ n18604 ^ 1'b0 ;
  assign n27441 = ( n11850 & ~n19252 ) | ( n11850 & n27440 ) | ( ~n19252 & n27440 ) ;
  assign n27444 = n27443 ^ n27441 ^ 1'b0 ;
  assign n27445 = n27436 & ~n27444 ;
  assign n27446 = n4011 | n12106 ;
  assign n27447 = n19948 ^ n9490 ^ n6190 ;
  assign n27448 = n18441 ^ n13430 ^ 1'b0 ;
  assign n27449 = n10229 & ~n27448 ;
  assign n27450 = ( ~n8164 & n8199 ) | ( ~n8164 & n27449 ) | ( n8199 & n27449 ) ;
  assign n27451 = ( ~n8595 & n16720 ) | ( ~n8595 & n25187 ) | ( n16720 & n25187 ) ;
  assign n27452 = n7391 & ~n24277 ;
  assign n27453 = ~n6616 & n27452 ;
  assign n27454 = n1984 & ~n27453 ;
  assign n27455 = n27454 ^ n9007 ^ 1'b0 ;
  assign n27456 = n15591 ^ n13479 ^ n3479 ;
  assign n27457 = n22800 ^ n4980 ^ 1'b0 ;
  assign n27458 = n12163 & n27457 ;
  assign n27459 = ~n14013 & n27458 ;
  assign n27460 = ( n18803 & ~n27456 ) | ( n18803 & n27459 ) | ( ~n27456 & n27459 ) ;
  assign n27461 = n13692 & ~n27259 ;
  assign n27462 = n25845 & n27461 ;
  assign n27463 = n27462 ^ n12161 ^ 1'b0 ;
  assign n27464 = n9923 ^ n3254 ^ 1'b0 ;
  assign n27465 = n6561 | n27464 ;
  assign n27466 = ( n1544 & n14967 ) | ( n1544 & n27465 ) | ( n14967 & n27465 ) ;
  assign n27467 = n27466 ^ n395 ^ 1'b0 ;
  assign n27468 = n3468 | n12293 ;
  assign n27469 = n27468 ^ n9720 ^ 1'b0 ;
  assign n27470 = ( n8291 & n15076 ) | ( n8291 & n27469 ) | ( n15076 & n27469 ) ;
  assign n27471 = ( n7576 & n8446 ) | ( n7576 & ~n8987 ) | ( n8446 & ~n8987 ) ;
  assign n27472 = n27471 ^ n11055 ^ 1'b0 ;
  assign n27473 = n5213 & ~n27472 ;
  assign n27474 = n23092 & n27473 ;
  assign n27475 = n4300 & n9361 ;
  assign n27476 = n2877 & ~n27475 ;
  assign n27477 = n27476 ^ x186 ^ 1'b0 ;
  assign n27478 = n1853 | n27477 ;
  assign n27479 = n27474 | n27478 ;
  assign n27480 = ~n4015 & n12557 ;
  assign n27481 = n27480 ^ n1746 ^ 1'b0 ;
  assign n27482 = n27481 ^ n547 ^ 1'b0 ;
  assign n27483 = n3516 | n18488 ;
  assign n27484 = n27482 & ~n27483 ;
  assign n27488 = n16905 & n20611 ;
  assign n27489 = n27488 ^ n16029 ^ 1'b0 ;
  assign n27485 = n8413 & ~n14605 ;
  assign n27486 = n27485 ^ n9094 ^ 1'b0 ;
  assign n27487 = ( n11472 & n24970 ) | ( n11472 & ~n27486 ) | ( n24970 & ~n27486 ) ;
  assign n27490 = n27489 ^ n27487 ^ n8157 ;
  assign n27491 = ( ~n1220 & n14695 ) | ( ~n1220 & n24873 ) | ( n14695 & n24873 ) ;
  assign n27492 = ~n23692 & n27491 ;
  assign n27493 = n23586 ^ n9932 ^ n429 ;
  assign n27494 = n5809 | n22304 ;
  assign n27495 = n11574 | n27494 ;
  assign n27496 = n12965 ^ n8148 ^ 1'b0 ;
  assign n27497 = n27495 & n27496 ;
  assign n27498 = n4633 ^ n4441 ^ n2498 ;
  assign n27499 = n14552 ^ n6484 ^ 1'b0 ;
  assign n27500 = n27498 & ~n27499 ;
  assign n27501 = ~n14525 & n27500 ;
  assign n27502 = ( ~n4311 & n22854 ) | ( ~n4311 & n27501 ) | ( n22854 & n27501 ) ;
  assign n27503 = ( n9623 & n27497 ) | ( n9623 & n27502 ) | ( n27497 & n27502 ) ;
  assign n27504 = n20301 ^ n3410 ^ n1323 ;
  assign n27505 = n27504 ^ n10353 ^ n857 ;
  assign n27506 = n7197 & n27505 ;
  assign n27507 = ~n27503 & n27506 ;
  assign n27508 = ~n8408 & n27115 ;
  assign n27509 = n23451 & n27508 ;
  assign n27510 = n22604 ^ n8209 ^ 1'b0 ;
  assign n27511 = n27510 ^ n7817 ^ 1'b0 ;
  assign n27515 = n11366 ^ n603 ^ 1'b0 ;
  assign n27514 = n7129 ^ n6029 ^ n547 ;
  assign n27516 = n27515 ^ n27514 ^ 1'b0 ;
  assign n27517 = n24064 & ~n27516 ;
  assign n27512 = n13754 ^ n10833 ^ 1'b0 ;
  assign n27513 = n20311 & ~n27512 ;
  assign n27518 = n27517 ^ n27513 ^ 1'b0 ;
  assign n27519 = ~n9131 & n10651 ;
  assign n27520 = n12700 & n27519 ;
  assign n27521 = n25248 & ~n27520 ;
  assign n27522 = ~n8003 & n27521 ;
  assign n27523 = n15207 | n27522 ;
  assign n27524 = n27523 ^ n10836 ^ 1'b0 ;
  assign n27525 = n7442 & ~n25686 ;
  assign n27526 = ( n798 & ~n19271 ) | ( n798 & n27525 ) | ( ~n19271 & n27525 ) ;
  assign n27527 = n24504 ^ n4747 ^ 1'b0 ;
  assign n27529 = ~n2194 & n3582 ;
  assign n27528 = ( ~n19428 & n22980 ) | ( ~n19428 & n25185 ) | ( n22980 & n25185 ) ;
  assign n27530 = n27529 ^ n27528 ^ n6878 ;
  assign n27531 = n27530 ^ n18644 ^ 1'b0 ;
  assign n27532 = ( n2632 & ~n18588 ) | ( n2632 & n24518 ) | ( ~n18588 & n24518 ) ;
  assign n27533 = ( n3651 & ~n11143 ) | ( n3651 & n17043 ) | ( ~n11143 & n17043 ) ;
  assign n27534 = n1914 & n7794 ;
  assign n27535 = n19715 ^ n5705 ^ n2094 ;
  assign n27536 = n2944 | n5052 ;
  assign n27537 = ( n6510 & n9349 ) | ( n6510 & ~n10195 ) | ( n9349 & ~n10195 ) ;
  assign n27538 = ( n21047 & n27536 ) | ( n21047 & n27537 ) | ( n27536 & n27537 ) ;
  assign n27539 = ( n10669 & n10792 ) | ( n10669 & ~n17219 ) | ( n10792 & ~n17219 ) ;
  assign n27540 = n27539 ^ n18057 ^ n6181 ;
  assign n27541 = n20135 | n27540 ;
  assign n27542 = n5234 | n26394 ;
  assign n27550 = ~n1921 & n24570 ;
  assign n27551 = n2502 ^ n1798 ^ 1'b0 ;
  assign n27552 = ~n27550 & n27551 ;
  assign n27546 = ~n712 & n18100 ;
  assign n27547 = n27546 ^ n8987 ^ 1'b0 ;
  assign n27548 = n27547 ^ n19961 ^ n14328 ;
  assign n27543 = n6883 | n13616 ;
  assign n27544 = n27543 ^ n2558 ^ 1'b0 ;
  assign n27545 = n12525 & ~n27544 ;
  assign n27549 = n27548 ^ n27545 ^ 1'b0 ;
  assign n27553 = n27552 ^ n27549 ^ 1'b0 ;
  assign n27554 = n27542 | n27553 ;
  assign n27555 = n26816 ^ n16732 ^ 1'b0 ;
  assign n27556 = n27555 ^ n12664 ^ 1'b0 ;
  assign n27557 = n27556 ^ n6709 ^ 1'b0 ;
  assign n27558 = n1822 & n22884 ;
  assign n27559 = ( n2021 & ~n12116 ) | ( n2021 & n16045 ) | ( ~n12116 & n16045 ) ;
  assign n27560 = ( n572 & ~n11018 ) | ( n572 & n27559 ) | ( ~n11018 & n27559 ) ;
  assign n27561 = n1108 & ~n18277 ;
  assign n27562 = n27561 ^ n12087 ^ 1'b0 ;
  assign n27563 = ( n2110 & ~n11470 ) | ( n2110 & n27562 ) | ( ~n11470 & n27562 ) ;
  assign n27564 = n4471 ^ n2152 ^ 1'b0 ;
  assign n27565 = n27564 ^ n12661 ^ 1'b0 ;
  assign n27566 = n11090 & n14633 ;
  assign n27567 = n27566 ^ n15028 ^ 1'b0 ;
  assign n27568 = n27567 ^ n6631 ^ n1810 ;
  assign n27569 = n7086 | n12275 ;
  assign n27570 = n13914 | n27569 ;
  assign n27574 = n7073 ^ n5285 ^ n722 ;
  assign n27575 = ( n2370 & ~n21599 ) | ( n2370 & n27574 ) | ( ~n21599 & n27574 ) ;
  assign n27571 = n21791 & ~n25617 ;
  assign n27572 = n27571 ^ n17351 ^ 1'b0 ;
  assign n27573 = n18522 & n27572 ;
  assign n27576 = n27575 ^ n27573 ^ 1'b0 ;
  assign n27579 = n4134 ^ n3258 ^ 1'b0 ;
  assign n27577 = n17570 ^ n13221 ^ 1'b0 ;
  assign n27578 = n5042 & ~n27577 ;
  assign n27580 = n27579 ^ n27578 ^ n5723 ;
  assign n27581 = n27580 ^ n22513 ^ 1'b0 ;
  assign n27582 = n6666 ^ n3173 ^ n2300 ;
  assign n27583 = n20797 ^ n13869 ^ n7608 ;
  assign n27584 = n1921 | n27583 ;
  assign n27585 = n27584 ^ n13801 ^ 1'b0 ;
  assign n27586 = n935 | n1584 ;
  assign n27587 = n15277 ^ n10777 ^ n7407 ;
  assign n27588 = n7774 ^ n2775 ^ 1'b0 ;
  assign n27589 = ( n7541 & n27587 ) | ( n7541 & n27588 ) | ( n27587 & n27588 ) ;
  assign n27590 = n19463 ^ n16943 ^ n1703 ;
  assign n27591 = n6902 & ~n27590 ;
  assign n27592 = n9136 & n26020 ;
  assign n27593 = n4638 & n27592 ;
  assign n27594 = ( ~n10501 & n26366 ) | ( ~n10501 & n27392 ) | ( n26366 & n27392 ) ;
  assign n27595 = n27594 ^ n13574 ^ 1'b0 ;
  assign n27596 = n20031 ^ n5713 ^ 1'b0 ;
  assign n27597 = ( n2099 & n5702 ) | ( n2099 & ~n13127 ) | ( n5702 & ~n13127 ) ;
  assign n27598 = n1368 & n18075 ;
  assign n27599 = n27598 ^ n4892 ^ 1'b0 ;
  assign n27600 = ( ~n2522 & n27597 ) | ( ~n2522 & n27599 ) | ( n27597 & n27599 ) ;
  assign n27601 = n4053 & n14096 ;
  assign n27602 = n17614 & n27601 ;
  assign n27603 = ~n4208 & n14515 ;
  assign n27605 = n19905 ^ n16497 ^ n1524 ;
  assign n27604 = ( ~n7671 & n12887 ) | ( ~n7671 & n15694 ) | ( n12887 & n15694 ) ;
  assign n27606 = n27605 ^ n27604 ^ 1'b0 ;
  assign n27607 = n27603 | n27606 ;
  assign n27608 = ( n2076 & ~n27602 ) | ( n2076 & n27607 ) | ( ~n27602 & n27607 ) ;
  assign n27609 = n27608 ^ n20622 ^ n9436 ;
  assign n27610 = n21577 ^ n9643 ^ n6320 ;
  assign n27611 = n9375 | n25769 ;
  assign n27612 = n27610 & ~n27611 ;
  assign n27613 = n25519 ^ n8124 ^ n5455 ;
  assign n27614 = n4458 & ~n4480 ;
  assign n27615 = n27614 ^ n5980 ^ 1'b0 ;
  assign n27616 = n27615 ^ n14980 ^ n6446 ;
  assign n27617 = n6968 ^ n6484 ^ n4494 ;
  assign n27618 = n27617 ^ n15202 ^ 1'b0 ;
  assign n27619 = ( n11103 & ~n25088 ) | ( n11103 & n27618 ) | ( ~n25088 & n27618 ) ;
  assign n27620 = n5015 ^ n1945 ^ n569 ;
  assign n27621 = ( n4807 & n14614 ) | ( n4807 & n27620 ) | ( n14614 & n27620 ) ;
  assign n27622 = n17304 | n27621 ;
  assign n27623 = n27622 ^ n19436 ^ n12048 ;
  assign n27624 = ~n14729 & n27623 ;
  assign n27625 = n21339 & n27624 ;
  assign n27626 = n26369 ^ n5337 ^ 1'b0 ;
  assign n27627 = n1732 & n9044 ;
  assign n27628 = n7970 & n27627 ;
  assign n27630 = n2494 & ~n22034 ;
  assign n27631 = n8382 & n27630 ;
  assign n27629 = ~n304 & n7638 ;
  assign n27632 = n27631 ^ n27629 ^ 1'b0 ;
  assign n27633 = ( ~n24199 & n27628 ) | ( ~n24199 & n27632 ) | ( n27628 & n27632 ) ;
  assign n27634 = n15591 ^ n3764 ^ x20 ;
  assign n27635 = n4365 & n27634 ;
  assign n27636 = n27635 ^ n12302 ^ 1'b0 ;
  assign n27637 = n27636 ^ n6889 ^ n4084 ;
  assign n27638 = n27637 ^ n24636 ^ n16029 ;
  assign n27639 = ~n3765 & n17803 ;
  assign n27640 = ~n17024 & n27639 ;
  assign n27641 = n27640 ^ n15145 ^ n13891 ;
  assign n27643 = n18187 ^ n13327 ^ n11971 ;
  assign n27644 = n27643 ^ n18390 ^ 1'b0 ;
  assign n27642 = n25094 ^ n17129 ^ n7247 ;
  assign n27645 = n27644 ^ n27642 ^ 1'b0 ;
  assign n27646 = ~n23627 & n27645 ;
  assign n27647 = ( n3005 & n7187 ) | ( n3005 & ~n8745 ) | ( n7187 & ~n8745 ) ;
  assign n27648 = n27647 ^ n5355 ^ 1'b0 ;
  assign n27649 = n17611 | n27648 ;
  assign n27650 = n27649 ^ n20686 ^ n3870 ;
  assign n27651 = n14013 & n24518 ;
  assign n27652 = n20162 ^ n1647 ^ 1'b0 ;
  assign n27653 = ~n21873 & n27652 ;
  assign n27654 = ~n5693 & n12927 ;
  assign n27655 = n3196 & n27654 ;
  assign n27656 = ( ~n8494 & n27653 ) | ( ~n8494 & n27655 ) | ( n27653 & n27655 ) ;
  assign n27657 = ( ~n6179 & n7604 ) | ( ~n6179 & n10815 ) | ( n7604 & n10815 ) ;
  assign n27658 = n7754 ^ n2002 ^ n261 ;
  assign n27659 = n8614 & n14284 ;
  assign n27660 = ( ~n824 & n27658 ) | ( ~n824 & n27659 ) | ( n27658 & n27659 ) ;
  assign n27661 = n24299 ^ n3661 ^ 1'b0 ;
  assign n27662 = n27660 | n27661 ;
  assign n27663 = n8435 & ~n11730 ;
  assign n27664 = n11099 ^ n9045 ^ n8032 ;
  assign n27665 = n27663 & n27664 ;
  assign n27666 = ( n4173 & n4408 ) | ( n4173 & n7827 ) | ( n4408 & n7827 ) ;
  assign n27667 = n8214 ^ n5265 ^ 1'b0 ;
  assign n27668 = ~n2114 & n27667 ;
  assign n27669 = n27668 ^ n14891 ^ n6944 ;
  assign n27670 = n11147 ^ n9824 ^ 1'b0 ;
  assign n27671 = ( ~n1609 & n6718 ) | ( ~n1609 & n27670 ) | ( n6718 & n27670 ) ;
  assign n27672 = n27671 ^ n21869 ^ n2967 ;
  assign n27673 = n862 & ~n8604 ;
  assign n27674 = n27673 ^ n2863 ^ 1'b0 ;
  assign n27675 = n12473 | n15079 ;
  assign n27676 = n27675 ^ n4298 ^ 1'b0 ;
  assign n27677 = n27676 ^ n10023 ^ n9403 ;
  assign n27678 = n1966 | n27677 ;
  assign n27679 = n18129 ^ n7563 ^ n387 ;
  assign n27680 = n4149 | n27679 ;
  assign n27681 = ( n2344 & ~n5773 ) | ( n2344 & n7878 ) | ( ~n5773 & n7878 ) ;
  assign n27682 = n8813 & n27681 ;
  assign n27683 = n27682 ^ n10926 ^ 1'b0 ;
  assign n27684 = ( n1200 & n27680 ) | ( n1200 & n27683 ) | ( n27680 & n27683 ) ;
  assign n27685 = ( n6177 & ~n13527 ) | ( n6177 & n16726 ) | ( ~n13527 & n16726 ) ;
  assign n27686 = n14859 ^ n7573 ^ n6628 ;
  assign n27687 = ( n1650 & n1993 ) | ( n1650 & n21442 ) | ( n1993 & n21442 ) ;
  assign n27688 = n27687 ^ n1469 ^ 1'b0 ;
  assign n27689 = n27686 | n27688 ;
  assign n27690 = n27689 ^ n15934 ^ 1'b0 ;
  assign n27691 = n27685 & n27690 ;
  assign n27694 = n8755 ^ n5278 ^ n3841 ;
  assign n27692 = n18752 ^ n7257 ^ 1'b0 ;
  assign n27693 = ~n23078 & n27692 ;
  assign n27695 = n27694 ^ n27693 ^ 1'b0 ;
  assign n27700 = ( ~n1952 & n2020 ) | ( ~n1952 & n15389 ) | ( n2020 & n15389 ) ;
  assign n27701 = n27700 ^ n16968 ^ n9720 ;
  assign n27696 = n20872 ^ n20301 ^ 1'b0 ;
  assign n27697 = n11728 & ~n27696 ;
  assign n27698 = n27697 ^ n25153 ^ 1'b0 ;
  assign n27699 = n725 & n27698 ;
  assign n27702 = n27701 ^ n27699 ^ 1'b0 ;
  assign n27703 = n27519 ^ n19291 ^ n16121 ;
  assign n27704 = n13407 & ~n13442 ;
  assign n27705 = n5587 ^ n2272 ^ 1'b0 ;
  assign n27706 = ( n16176 & n21554 ) | ( n16176 & n27705 ) | ( n21554 & n27705 ) ;
  assign n27707 = n27704 | n27706 ;
  assign n27708 = n13366 | n22972 ;
  assign n27709 = n3228 & ~n11841 ;
  assign n27710 = n27709 ^ x165 ^ 1'b0 ;
  assign n27711 = n9754 & n12630 ;
  assign n27712 = n2293 & n13802 ;
  assign n27713 = n8213 ^ n5880 ^ 1'b0 ;
  assign n27714 = n17319 & n27713 ;
  assign n27715 = n24157 ^ n7093 ^ 1'b0 ;
  assign n27716 = n1968 & n27715 ;
  assign n27717 = n27716 ^ n10520 ^ 1'b0 ;
  assign n27718 = n4635 | n6161 ;
  assign n27719 = n27718 ^ n13298 ^ 1'b0 ;
  assign n27720 = n9926 & ~n27719 ;
  assign n27721 = n22254 ^ n838 ^ 1'b0 ;
  assign n27722 = ( n26267 & n27720 ) | ( n26267 & n27721 ) | ( n27720 & n27721 ) ;
  assign n27723 = n6938 & ~n19151 ;
  assign n27724 = n27723 ^ n24896 ^ 1'b0 ;
  assign n27725 = n20669 ^ n18747 ^ n11010 ;
  assign n27726 = n7961 & ~n20677 ;
  assign n27727 = n27726 ^ n4254 ^ 1'b0 ;
  assign n27728 = x63 & n27727 ;
  assign n27729 = ( ~n21112 & n27725 ) | ( ~n21112 & n27728 ) | ( n27725 & n27728 ) ;
  assign n27730 = x25 & ~n4078 ;
  assign n27731 = n27730 ^ n4529 ^ 1'b0 ;
  assign n27732 = n27731 ^ n3262 ^ 1'b0 ;
  assign n27733 = n5846 & ~n27732 ;
  assign n27734 = ( n18745 & ~n19191 ) | ( n18745 & n27733 ) | ( ~n19191 & n27733 ) ;
  assign n27735 = ( n6302 & n8052 ) | ( n6302 & ~n27734 ) | ( n8052 & ~n27734 ) ;
  assign n27736 = n4484 & ~n7698 ;
  assign n27737 = ( x53 & ~n4240 ) | ( x53 & n7922 ) | ( ~n4240 & n7922 ) ;
  assign n27738 = ( n26674 & n27736 ) | ( n26674 & n27737 ) | ( n27736 & n27737 ) ;
  assign n27739 = n485 & n6148 ;
  assign n27740 = ~n2332 & n27739 ;
  assign n27741 = n27740 ^ n18093 ^ n1548 ;
  assign n27742 = n7167 & n8996 ;
  assign n27743 = ~n6783 & n27742 ;
  assign n27744 = n27741 & ~n27743 ;
  assign n27745 = n16277 | n27744 ;
  assign n27746 = n27745 ^ n11615 ^ 1'b0 ;
  assign n27747 = n27746 ^ n10588 ^ 1'b0 ;
  assign n27748 = ~n27738 & n27747 ;
  assign n27749 = n15820 ^ n5441 ^ x48 ;
  assign n27750 = ( n4501 & n4994 ) | ( n4501 & ~n6884 ) | ( n4994 & ~n6884 ) ;
  assign n27751 = n27750 ^ n24425 ^ n11546 ;
  assign n27752 = n11015 & n27751 ;
  assign n27753 = ~n27749 & n27752 ;
  assign n27754 = ~n10350 & n17641 ;
  assign n27755 = n21139 ^ n7984 ^ 1'b0 ;
  assign n27756 = n27754 | n27755 ;
  assign n27757 = ( ~n282 & n9437 ) | ( ~n282 & n15200 ) | ( n9437 & n15200 ) ;
  assign n27758 = n27757 ^ n3648 ^ n1969 ;
  assign n27759 = n11314 ^ n10829 ^ n10465 ;
  assign n27760 = n638 & ~n18031 ;
  assign n27761 = n27759 & n27760 ;
  assign n27763 = n16874 ^ n6015 ^ n632 ;
  assign n27762 = ~n3785 & n4371 ;
  assign n27764 = n27763 ^ n27762 ^ n26812 ;
  assign n27765 = n7788 | n8914 ;
  assign n27766 = n27765 ^ n6027 ^ n1447 ;
  assign n27767 = n2494 & n27766 ;
  assign n27768 = ( n3144 & n11088 ) | ( n3144 & n14998 ) | ( n11088 & n14998 ) ;
  assign n27769 = ( n10388 & ~n21013 ) | ( n10388 & n27768 ) | ( ~n21013 & n27768 ) ;
  assign n27770 = n10076 & n13759 ;
  assign n27771 = ~n16361 & n27770 ;
  assign n27772 = n27771 ^ n1072 ^ 1'b0 ;
  assign n27773 = ~n27769 & n27772 ;
  assign n27774 = n20863 ^ n12323 ^ 1'b0 ;
  assign n27775 = n19698 & ~n20123 ;
  assign n27776 = ~n27774 & n27775 ;
  assign n27777 = n27776 ^ n18434 ^ n2576 ;
  assign n27778 = n14844 | n15616 ;
  assign n27779 = n10277 | n27778 ;
  assign n27780 = n12578 ^ n7790 ^ n2364 ;
  assign n27781 = n27780 ^ n13702 ^ n12032 ;
  assign n27782 = ( ~n11022 & n27779 ) | ( ~n11022 & n27781 ) | ( n27779 & n27781 ) ;
  assign n27783 = ( n8413 & ~n10491 ) | ( n8413 & n22004 ) | ( ~n10491 & n22004 ) ;
  assign n27784 = ~n16084 & n27783 ;
  assign n27785 = n24441 & n27784 ;
  assign n27786 = ( n11034 & ~n18884 ) | ( n11034 & n27206 ) | ( ~n18884 & n27206 ) ;
  assign n27787 = n27786 ^ n17917 ^ n1502 ;
  assign n27789 = n1303 & n18083 ;
  assign n27790 = ~n1553 & n27789 ;
  assign n27788 = n21143 ^ n15978 ^ 1'b0 ;
  assign n27791 = n27790 ^ n27788 ^ n14927 ;
  assign n27792 = n9700 & n12606 ;
  assign n27793 = n27792 ^ x180 ^ 1'b0 ;
  assign n27794 = ( ~n6450 & n6466 ) | ( ~n6450 & n12499 ) | ( n6466 & n12499 ) ;
  assign n27795 = ( n16052 & n27793 ) | ( n16052 & n27794 ) | ( n27793 & n27794 ) ;
  assign n27796 = ( ~n5220 & n12024 ) | ( ~n5220 & n22245 ) | ( n12024 & n22245 ) ;
  assign n27797 = n17612 & n27796 ;
  assign n27798 = ( n3997 & ~n19245 ) | ( n3997 & n27797 ) | ( ~n19245 & n27797 ) ;
  assign n27799 = ( n701 & n27795 ) | ( n701 & n27798 ) | ( n27795 & n27798 ) ;
  assign n27800 = n26919 ^ n20601 ^ n1924 ;
  assign n27803 = n6933 ^ n6002 ^ n2694 ;
  assign n27801 = n8137 ^ n3737 ^ 1'b0 ;
  assign n27802 = n15880 | n27801 ;
  assign n27804 = n27803 ^ n27802 ^ 1'b0 ;
  assign n27805 = n3159 ^ n271 ^ 1'b0 ;
  assign n27806 = n6944 ^ n3403 ^ n2157 ;
  assign n27807 = n6476 & ~n27806 ;
  assign n27808 = ~x227 & n27807 ;
  assign n27809 = n27805 | n27808 ;
  assign n27810 = n7401 | n27809 ;
  assign n27811 = n27810 ^ n10902 ^ x88 ;
  assign n27812 = n23700 ^ n13642 ^ n2382 ;
  assign n27813 = n17851 ^ n2596 ^ 1'b0 ;
  assign n27814 = n14942 & n27813 ;
  assign n27815 = ~n7667 & n27814 ;
  assign n27816 = ~n4396 & n27815 ;
  assign n27817 = n4227 | n10397 ;
  assign n27818 = n27816 & ~n27817 ;
  assign n27819 = n18868 ^ n7824 ^ n3661 ;
  assign n27820 = n27819 ^ n16659 ^ n15454 ;
  assign n27821 = ~n6122 & n10049 ;
  assign n27822 = n27821 ^ n1803 ^ 1'b0 ;
  assign n27823 = n27822 ^ n19589 ^ n3987 ;
  assign n27824 = ( ~n2434 & n19991 ) | ( ~n2434 & n26710 ) | ( n19991 & n26710 ) ;
  assign n27825 = n18093 ^ n2874 ^ 1'b0 ;
  assign n27826 = n15274 ^ n11991 ^ n6165 ;
  assign n27827 = n18132 & ~n27826 ;
  assign n27828 = n20742 & ~n27827 ;
  assign n27829 = n27825 & n27828 ;
  assign n27831 = n26994 ^ n3747 ^ 1'b0 ;
  assign n27830 = n397 & ~n10720 ;
  assign n27832 = n27831 ^ n27830 ^ 1'b0 ;
  assign n27833 = ( n4313 & ~n6230 ) | ( n4313 & n25940 ) | ( ~n6230 & n25940 ) ;
  assign n27834 = ( n4295 & n7899 ) | ( n4295 & ~n27544 ) | ( n7899 & ~n27544 ) ;
  assign n27835 = n3889 ^ n2381 ^ n1993 ;
  assign n27836 = n27835 ^ n17184 ^ 1'b0 ;
  assign n27837 = n12157 & n27836 ;
  assign n27838 = n26032 & n27837 ;
  assign n27839 = ~n27834 & n27838 ;
  assign n27840 = n27833 | n27839 ;
  assign n27841 = n18795 & ~n27840 ;
  assign n27842 = n530 & ~n7833 ;
  assign n27843 = n19905 & ~n27842 ;
  assign n27844 = ( n500 & n6235 ) | ( n500 & ~n9728 ) | ( n6235 & ~n9728 ) ;
  assign n27845 = n27844 ^ n17132 ^ n12775 ;
  assign n27846 = n27843 | n27845 ;
  assign n27847 = n16812 ^ n7421 ^ n5097 ;
  assign n27848 = n14695 ^ n5685 ^ n5417 ;
  assign n27849 = n12537 ^ n2433 ^ 1'b0 ;
  assign n27850 = n16410 & n27849 ;
  assign n27851 = n27850 ^ n8056 ^ 1'b0 ;
  assign n27852 = ( n5939 & ~n11065 ) | ( n5939 & n27851 ) | ( ~n11065 & n27851 ) ;
  assign n27854 = n15288 ^ n3254 ^ n2086 ;
  assign n27853 = n3974 & ~n26308 ;
  assign n27855 = n27854 ^ n27853 ^ 1'b0 ;
  assign n27856 = n17571 ^ n17356 ^ n3618 ;
  assign n27857 = n17602 ^ n6118 ^ 1'b0 ;
  assign n27858 = n3095 & ~n27857 ;
  assign n27860 = n25127 ^ n23125 ^ n18778 ;
  assign n27859 = ~n10162 & n24996 ;
  assign n27861 = n27860 ^ n27859 ^ 1'b0 ;
  assign n27862 = ( ~n2662 & n16983 ) | ( ~n2662 & n26955 ) | ( n16983 & n26955 ) ;
  assign n27863 = n26208 ^ n23145 ^ 1'b0 ;
  assign n27864 = ( n21609 & n27862 ) | ( n21609 & n27863 ) | ( n27862 & n27863 ) ;
  assign n27865 = n664 | n2012 ;
  assign n27866 = ~n1157 & n3843 ;
  assign n27867 = ~n16856 & n27866 ;
  assign n27868 = n27865 & ~n27867 ;
  assign n27869 = n8333 ^ n7280 ^ n5051 ;
  assign n27870 = n14168 & ~n27869 ;
  assign n27871 = n20408 & n27870 ;
  assign n27872 = ( n1491 & n6929 ) | ( n1491 & ~n16743 ) | ( n6929 & ~n16743 ) ;
  assign n27873 = n27871 & ~n27872 ;
  assign n27874 = n9055 ^ n5522 ^ n2131 ;
  assign n27875 = ( n5218 & n12852 ) | ( n5218 & n27874 ) | ( n12852 & n27874 ) ;
  assign n27876 = n1136 & ~n27875 ;
  assign n27877 = n27876 ^ n16023 ^ 1'b0 ;
  assign n27878 = ~n1173 & n27877 ;
  assign n27879 = n4526 & n27878 ;
  assign n27880 = n3898 | n10953 ;
  assign n27881 = n27880 ^ n12508 ^ 1'b0 ;
  assign n27882 = ~n24546 & n27881 ;
  assign n27884 = n4760 & ~n5441 ;
  assign n27885 = ~n3925 & n27884 ;
  assign n27886 = n27885 ^ n9772 ^ n4906 ;
  assign n27883 = n10444 | n25672 ;
  assign n27887 = n27886 ^ n27883 ^ 1'b0 ;
  assign n27888 = n2475 & ~n5901 ;
  assign n27889 = n13025 ^ n2240 ^ n355 ;
  assign n27890 = n16697 & n22260 ;
  assign n27891 = ~n27889 & n27890 ;
  assign n27892 = ( n9062 & n22228 ) | ( n9062 & ~n27891 ) | ( n22228 & ~n27891 ) ;
  assign n27893 = n27144 & n27892 ;
  assign n27894 = n27893 ^ n23586 ^ 1'b0 ;
  assign n27895 = ( ~n27887 & n27888 ) | ( ~n27887 & n27894 ) | ( n27888 & n27894 ) ;
  assign n27896 = n27895 ^ n20464 ^ 1'b0 ;
  assign n27897 = ~n912 & n27896 ;
  assign n27898 = n27897 ^ n2962 ^ 1'b0 ;
  assign n27899 = ( n3520 & n4563 ) | ( n3520 & n10917 ) | ( n4563 & n10917 ) ;
  assign n27900 = ( ~n3586 & n10589 ) | ( ~n3586 & n27899 ) | ( n10589 & n27899 ) ;
  assign n27901 = ( ~n14527 & n17967 ) | ( ~n14527 & n27900 ) | ( n17967 & n27900 ) ;
  assign n27902 = ( n2812 & n12563 ) | ( n2812 & n27901 ) | ( n12563 & n27901 ) ;
  assign n27903 = ( n2184 & ~n11450 ) | ( n2184 & n27902 ) | ( ~n11450 & n27902 ) ;
  assign n27904 = n23636 ^ n12977 ^ n8272 ;
  assign n27905 = ( n2360 & ~n11819 ) | ( n2360 & n27904 ) | ( ~n11819 & n27904 ) ;
  assign n27906 = n13024 ^ n7689 ^ n6072 ;
  assign n27907 = n7438 & n24092 ;
  assign n27908 = n13038 & n27907 ;
  assign n27909 = n20894 & n21917 ;
  assign n27910 = n16385 | n19692 ;
  assign n27911 = ~n8848 & n17657 ;
  assign n27912 = n1352 & n27911 ;
  assign n27913 = n27912 ^ n27694 ^ n14818 ;
  assign n27914 = n27913 ^ n1758 ^ 1'b0 ;
  assign n27915 = n3499 & n19697 ;
  assign n27916 = ( n20409 & ~n21999 ) | ( n20409 & n27915 ) | ( ~n21999 & n27915 ) ;
  assign n27917 = n14553 ^ n9713 ^ n6919 ;
  assign n27918 = ( ~n2279 & n4075 ) | ( ~n2279 & n25246 ) | ( n4075 & n25246 ) ;
  assign n27919 = ( ~n9244 & n27917 ) | ( ~n9244 & n27918 ) | ( n27917 & n27918 ) ;
  assign n27920 = n9917 & ~n27919 ;
  assign n27923 = n21327 ^ n15181 ^ n4375 ;
  assign n27921 = n3456 & ~n8643 ;
  assign n27922 = n7116 | n27921 ;
  assign n27924 = n27923 ^ n27922 ^ n9895 ;
  assign n27925 = n18328 ^ n14863 ^ n11231 ;
  assign n27926 = n4070 & n12321 ;
  assign n27927 = n27926 ^ n3335 ^ 1'b0 ;
  assign n27928 = ( n12769 & n14818 ) | ( n12769 & n27927 ) | ( n14818 & n27927 ) ;
  assign n27929 = n21296 ^ n2097 ^ 1'b0 ;
  assign n27930 = ~n11003 & n27929 ;
  assign n27931 = n5376 ^ n3739 ^ 1'b0 ;
  assign n27932 = ~n1662 & n6424 ;
  assign n27933 = ~n6660 & n27932 ;
  assign n27934 = n595 & n19780 ;
  assign n27935 = ~n14233 & n27934 ;
  assign n27936 = ( ~n19824 & n27933 ) | ( ~n19824 & n27935 ) | ( n27933 & n27935 ) ;
  assign n27938 = ( ~n7354 & n11108 ) | ( ~n7354 & n21326 ) | ( n11108 & n21326 ) ;
  assign n27939 = n5101 | n27938 ;
  assign n27940 = n14100 | n27939 ;
  assign n27941 = n3815 & ~n26763 ;
  assign n27942 = n2000 & n27941 ;
  assign n27943 = n27942 ^ n8336 ^ n7591 ;
  assign n27944 = n2422 | n27943 ;
  assign n27945 = n27944 ^ n7989 ^ 1'b0 ;
  assign n27946 = n27940 & ~n27945 ;
  assign n27947 = n27946 ^ n8644 ^ 1'b0 ;
  assign n27937 = n15973 | n18039 ;
  assign n27948 = n27947 ^ n27937 ^ 1'b0 ;
  assign n27949 = n8303 & ~n8583 ;
  assign n27950 = n27949 ^ n4017 ^ 1'b0 ;
  assign n27951 = n8945 | n27950 ;
  assign n27952 = n689 & ~n27951 ;
  assign n27955 = n17292 ^ n14074 ^ n9564 ;
  assign n27956 = n3681 | n27955 ;
  assign n27957 = n10218 | n27956 ;
  assign n27953 = ( n1445 & n5449 ) | ( n1445 & ~n11784 ) | ( n5449 & ~n11784 ) ;
  assign n27954 = n27953 ^ n2819 ^ 1'b0 ;
  assign n27958 = n27957 ^ n27954 ^ 1'b0 ;
  assign n27959 = n2560 & ~n15595 ;
  assign n27960 = n17829 & ~n19568 ;
  assign n27961 = n27960 ^ n358 ^ 1'b0 ;
  assign n27962 = x194 & ~n12205 ;
  assign n27963 = n18198 ^ n5752 ^ n5566 ;
  assign n27964 = ~n27962 & n27963 ;
  assign n27965 = ( n5146 & n25890 ) | ( n5146 & ~n27964 ) | ( n25890 & ~n27964 ) ;
  assign n27966 = ( n5478 & n23932 ) | ( n5478 & n27965 ) | ( n23932 & n27965 ) ;
  assign n27967 = n27966 ^ n18753 ^ n8745 ;
  assign n27968 = n16974 ^ n8180 ^ n7009 ;
  assign n27969 = n7316 ^ n4981 ^ 1'b0 ;
  assign n27970 = n16080 | n27969 ;
  assign n27971 = ( n304 & ~n27968 ) | ( n304 & n27970 ) | ( ~n27968 & n27970 ) ;
  assign n27976 = ( n2866 & n5928 ) | ( n2866 & ~n15266 ) | ( n5928 & ~n15266 ) ;
  assign n27973 = ~n5282 & n7201 ;
  assign n27974 = ~n9957 & n27973 ;
  assign n27972 = n11896 & n19470 ;
  assign n27975 = n27974 ^ n27972 ^ 1'b0 ;
  assign n27977 = n27976 ^ n27975 ^ n12938 ;
  assign n27978 = n27977 ^ n27314 ^ n3951 ;
  assign n27979 = n7677 & ~n22097 ;
  assign n27980 = ( n11467 & ~n20497 ) | ( n11467 & n25384 ) | ( ~n20497 & n25384 ) ;
  assign n27981 = n27980 ^ n26833 ^ 1'b0 ;
  assign n27982 = n18679 ^ n11663 ^ 1'b0 ;
  assign n27983 = ( n6995 & n26399 ) | ( n6995 & n27982 ) | ( n26399 & n27982 ) ;
  assign n27984 = ( ~n14768 & n18155 ) | ( ~n14768 & n27983 ) | ( n18155 & n27983 ) ;
  assign n27985 = ( n4082 & n9062 ) | ( n4082 & ~n19084 ) | ( n9062 & ~n19084 ) ;
  assign n27986 = n27985 ^ n10196 ^ n1294 ;
  assign n27987 = n7387 ^ n2909 ^ 1'b0 ;
  assign n27988 = n12096 & n27987 ;
  assign n27989 = ( ~n4652 & n6398 ) | ( ~n4652 & n7640 ) | ( n6398 & n7640 ) ;
  assign n27990 = n5362 & ~n27989 ;
  assign n27991 = n23867 & n27990 ;
  assign n27992 = n27991 ^ n11771 ^ 1'b0 ;
  assign n27993 = n27988 & n27992 ;
  assign n27994 = ~n21432 & n24913 ;
  assign n27995 = n27994 ^ n280 ^ 1'b0 ;
  assign n27996 = ~n10314 & n27995 ;
  assign n27997 = ~n27993 & n27996 ;
  assign n28002 = ( n1508 & n2353 ) | ( n1508 & ~n3347 ) | ( n2353 & ~n3347 ) ;
  assign n27998 = n6793 & ~n12131 ;
  assign n27999 = n27998 ^ n20001 ^ n446 ;
  assign n28000 = n5595 & n27999 ;
  assign n28001 = n16838 & n28000 ;
  assign n28003 = n28002 ^ n28001 ^ 1'b0 ;
  assign n28004 = n8943 ^ n5288 ^ n423 ;
  assign n28005 = ( n24845 & n25918 ) | ( n24845 & ~n28004 ) | ( n25918 & ~n28004 ) ;
  assign n28006 = ( ~n2177 & n22632 ) | ( ~n2177 & n28005 ) | ( n22632 & n28005 ) ;
  assign n28007 = n12218 & n22010 ;
  assign n28008 = n28007 ^ n10967 ^ 1'b0 ;
  assign n28009 = n28008 ^ n23578 ^ n1486 ;
  assign n28011 = ( ~n1900 & n11538 ) | ( ~n1900 & n12823 ) | ( n11538 & n12823 ) ;
  assign n28010 = ( n5998 & ~n11242 ) | ( n5998 & n21549 ) | ( ~n11242 & n21549 ) ;
  assign n28012 = n28011 ^ n28010 ^ n17147 ;
  assign n28013 = n9098 & n12682 ;
  assign n28014 = n28013 ^ n5232 ^ 1'b0 ;
  assign n28015 = n4224 | n14017 ;
  assign n28016 = n28015 ^ n24702 ^ 1'b0 ;
  assign n28017 = n28016 ^ n4057 ^ 1'b0 ;
  assign n28018 = n6304 & n13312 ;
  assign n28019 = n1276 & ~n17307 ;
  assign n28020 = n11286 | n28019 ;
  assign n28021 = n28020 ^ n9279 ^ 1'b0 ;
  assign n28022 = n5190 & n28021 ;
  assign n28023 = n28022 ^ n7296 ^ 1'b0 ;
  assign n28024 = ~n14801 & n28023 ;
  assign n28025 = ( n10961 & n25805 ) | ( n10961 & ~n28024 ) | ( n25805 & ~n28024 ) ;
  assign n28026 = ~n1245 & n22286 ;
  assign n28027 = ~n13590 & n28026 ;
  assign n28028 = ( ~n22250 & n24854 ) | ( ~n22250 & n28027 ) | ( n24854 & n28027 ) ;
  assign n28029 = n23015 & ~n23249 ;
  assign n28030 = n3969 & n28029 ;
  assign n28032 = n7995 ^ n1684 ^ 1'b0 ;
  assign n28033 = ~n2329 & n28032 ;
  assign n28031 = ( ~n10292 & n18193 ) | ( ~n10292 & n19515 ) | ( n18193 & n19515 ) ;
  assign n28034 = n28033 ^ n28031 ^ 1'b0 ;
  assign n28035 = ~n7269 & n10671 ;
  assign n28036 = ~n8802 & n28035 ;
  assign n28037 = ( n9120 & ~n15659 ) | ( n9120 & n28036 ) | ( ~n15659 & n28036 ) ;
  assign n28038 = n22346 ^ n12779 ^ 1'b0 ;
  assign n28039 = n28038 ^ n2755 ^ n2382 ;
  assign n28040 = ( x215 & n24231 ) | ( x215 & ~n25849 ) | ( n24231 & ~n25849 ) ;
  assign n28041 = n28040 ^ n14257 ^ n11577 ;
  assign n28042 = n6621 | n14279 ;
  assign n28043 = n28042 ^ n15716 ^ n298 ;
  assign n28044 = n16069 ^ n11216 ^ 1'b0 ;
  assign n28045 = n28044 ^ n22791 ^ 1'b0 ;
  assign n28046 = ( n1839 & n18093 ) | ( n1839 & n22532 ) | ( n18093 & n22532 ) ;
  assign n28047 = n28046 ^ n23929 ^ n1041 ;
  assign n28048 = ( n2442 & n9670 ) | ( n2442 & ~n28047 ) | ( n9670 & ~n28047 ) ;
  assign n28049 = n23736 ^ n22107 ^ n4584 ;
  assign n28051 = n23856 ^ n6032 ^ n554 ;
  assign n28050 = n16749 ^ n6106 ^ 1'b0 ;
  assign n28052 = n28051 ^ n28050 ^ n10733 ;
  assign n28053 = ( ~n12746 & n13892 ) | ( ~n12746 & n18579 ) | ( n13892 & n18579 ) ;
  assign n28054 = n22996 ^ n10380 ^ 1'b0 ;
  assign n28055 = n3355 & n9452 ;
  assign n28056 = ( n8678 & n15692 ) | ( n8678 & ~n28055 ) | ( n15692 & ~n28055 ) ;
  assign n28057 = ( n910 & n12455 ) | ( n910 & n21962 ) | ( n12455 & n21962 ) ;
  assign n28058 = ( n4462 & ~n28056 ) | ( n4462 & n28057 ) | ( ~n28056 & n28057 ) ;
  assign n28059 = n4683 & ~n4729 ;
  assign n28060 = n28059 ^ n11503 ^ 1'b0 ;
  assign n28061 = n28060 ^ n7796 ^ 1'b0 ;
  assign n28062 = n28061 ^ n8233 ^ 1'b0 ;
  assign n28063 = ~n6077 & n28062 ;
  assign n28064 = n8360 | n28063 ;
  assign n28068 = n1458 & n9262 ;
  assign n28066 = n1191 & ~n6345 ;
  assign n28067 = n4387 & n28066 ;
  assign n28065 = ( n1444 & ~n6391 ) | ( n1444 & n8334 ) | ( ~n6391 & n8334 ) ;
  assign n28069 = n28068 ^ n28067 ^ n28065 ;
  assign n28070 = n15334 ^ n2247 ^ 1'b0 ;
  assign n28071 = n24775 ^ n4394 ^ 1'b0 ;
  assign n28072 = n20014 ^ n16511 ^ n3632 ;
  assign n28073 = ( ~n5722 & n14255 ) | ( ~n5722 & n15234 ) | ( n14255 & n15234 ) ;
  assign n28074 = n18968 ^ n7662 ^ 1'b0 ;
  assign n28075 = n5344 & ~n28074 ;
  assign n28076 = n24687 ^ n7401 ^ 1'b0 ;
  assign n28077 = n10281 | n26929 ;
  assign n28078 = n28077 ^ n11477 ^ 1'b0 ;
  assign n28079 = n28076 & ~n28078 ;
  assign n28080 = n1429 & ~n1492 ;
  assign n28081 = n19295 ^ n15142 ^ n7750 ;
  assign n28082 = n16893 & n28081 ;
  assign n28083 = n28080 & n28082 ;
  assign n28084 = n639 | n22241 ;
  assign n28085 = n1848 & ~n28084 ;
  assign n28086 = n28085 ^ n13195 ^ 1'b0 ;
  assign n28087 = n20726 & n28086 ;
  assign n28088 = n28087 ^ n5417 ^ 1'b0 ;
  assign n28089 = n14592 & n28088 ;
  assign n28090 = n28089 ^ n18940 ^ 1'b0 ;
  assign n28091 = ( n8018 & ~n8810 ) | ( n8018 & n11172 ) | ( ~n8810 & n11172 ) ;
  assign n28092 = n12583 & ~n17218 ;
  assign n28093 = ( n5410 & n10631 ) | ( n5410 & n16857 ) | ( n10631 & n16857 ) ;
  assign n28095 = n22875 ^ n16654 ^ 1'b0 ;
  assign n28096 = n19766 & ~n28095 ;
  assign n28094 = n17638 ^ n13088 ^ n11105 ;
  assign n28097 = n28096 ^ n28094 ^ 1'b0 ;
  assign n28098 = n28097 ^ n1475 ^ 1'b0 ;
  assign n28099 = n28093 & n28098 ;
  assign n28100 = ( n758 & ~n24753 ) | ( n758 & n28099 ) | ( ~n24753 & n28099 ) ;
  assign n28104 = ( n3216 & n6650 ) | ( n3216 & ~n8732 ) | ( n6650 & ~n8732 ) ;
  assign n28105 = x78 & ~n28104 ;
  assign n28106 = n28105 ^ n22807 ^ 1'b0 ;
  assign n28103 = ( ~n11338 & n11580 ) | ( ~n11338 & n20305 ) | ( n11580 & n20305 ) ;
  assign n28101 = n2121 | n12826 ;
  assign n28102 = n1940 | n28101 ;
  assign n28107 = n28106 ^ n28103 ^ n28102 ;
  assign n28108 = n18286 & ~n19583 ;
  assign n28109 = n28108 ^ n2857 ^ 1'b0 ;
  assign n28110 = n10086 ^ n7313 ^ 1'b0 ;
  assign n28111 = ( x244 & n21572 ) | ( x244 & ~n28110 ) | ( n21572 & ~n28110 ) ;
  assign n28112 = ~n4192 & n28111 ;
  assign n28113 = n12619 ^ n10121 ^ 1'b0 ;
  assign n28114 = ( ~n9361 & n24515 ) | ( ~n9361 & n25604 ) | ( n24515 & n25604 ) ;
  assign n28115 = n14146 | n17997 ;
  assign n28116 = n28115 ^ n17435 ^ 1'b0 ;
  assign n28117 = n14596 ^ n12414 ^ 1'b0 ;
  assign n28118 = n5237 & n28117 ;
  assign n28119 = n8198 ^ n4582 ^ n595 ;
  assign n28120 = n1685 & n8475 ;
  assign n28121 = ( n7369 & n23074 ) | ( n7369 & ~n23653 ) | ( n23074 & ~n23653 ) ;
  assign n28122 = n28121 ^ n7950 ^ 1'b0 ;
  assign n28123 = n3028 | n27456 ;
  assign n28124 = n28123 ^ n3408 ^ 1'b0 ;
  assign n28125 = n13408 ^ n7741 ^ 1'b0 ;
  assign n28126 = ~n4950 & n16250 ;
  assign n28127 = ( n16596 & ~n28125 ) | ( n16596 & n28126 ) | ( ~n28125 & n28126 ) ;
  assign n28130 = ( n3959 & n7902 ) | ( n3959 & ~n17030 ) | ( n7902 & ~n17030 ) ;
  assign n28128 = n27885 ^ n15127 ^ 1'b0 ;
  assign n28129 = n13018 & n28128 ;
  assign n28131 = n28130 ^ n28129 ^ n7627 ;
  assign n28132 = n15930 ^ n15478 ^ n6718 ;
  assign n28133 = n28132 ^ n16129 ^ 1'b0 ;
  assign n28134 = n4290 ^ n1543 ^ 1'b0 ;
  assign n28135 = n6193 | n13183 ;
  assign n28136 = n12244 & ~n28135 ;
  assign n28137 = n2859 & ~n28136 ;
  assign n28138 = ~n28134 & n28137 ;
  assign n28139 = n9222 ^ n3587 ^ n1019 ;
  assign n28140 = n5340 | n14104 ;
  assign n28141 = n28139 | n28140 ;
  assign n28142 = ~n13361 & n28141 ;
  assign n28143 = n11435 ^ n2356 ^ 1'b0 ;
  assign n28145 = n23882 ^ n15335 ^ n9857 ;
  assign n28144 = n6741 ^ n3377 ^ n1630 ;
  assign n28146 = n28145 ^ n28144 ^ n13456 ;
  assign n28147 = x196 & n13305 ;
  assign n28148 = n21609 ^ n19107 ^ n8465 ;
  assign n28154 = ( n447 & ~n5110 ) | ( n447 & n8179 ) | ( ~n5110 & n8179 ) ;
  assign n28149 = n20186 ^ n17414 ^ n13002 ;
  assign n28150 = n12843 & n16546 ;
  assign n28151 = n28149 & n28150 ;
  assign n28152 = n7879 & n10139 ;
  assign n28153 = ~n28151 & n28152 ;
  assign n28155 = n28154 ^ n28153 ^ n12884 ;
  assign n28156 = ( ~n16328 & n28148 ) | ( ~n16328 & n28155 ) | ( n28148 & n28155 ) ;
  assign n28157 = n10665 & n13586 ;
  assign n28158 = ( n23760 & n27281 ) | ( n23760 & ~n28157 ) | ( n27281 & ~n28157 ) ;
  assign n28159 = n5386 & n16016 ;
  assign n28160 = ( n10019 & n12996 ) | ( n10019 & n15924 ) | ( n12996 & n15924 ) ;
  assign n28161 = n12442 & ~n28160 ;
  assign n28162 = n16393 & n28161 ;
  assign n28163 = n21442 & n28162 ;
  assign n28164 = n25673 ^ x46 ^ 1'b0 ;
  assign n28165 = ~n5673 & n28164 ;
  assign n28166 = n11138 ^ n10593 ^ n5142 ;
  assign n28167 = n12070 ^ n9531 ^ n4902 ;
  assign n28168 = ( n12461 & n15338 ) | ( n12461 & ~n28167 ) | ( n15338 & ~n28167 ) ;
  assign n28169 = n12220 ^ n9402 ^ n2035 ;
  assign n28170 = n20246 ^ n12525 ^ 1'b0 ;
  assign n28171 = ~n17987 & n28170 ;
  assign n28180 = n1169 ^ n822 ^ 1'b0 ;
  assign n28181 = ~n19569 & n28180 ;
  assign n28182 = ( n15447 & ~n15791 ) | ( n15447 & n28181 ) | ( ~n15791 & n28181 ) ;
  assign n28178 = n13535 ^ n5285 ^ 1'b0 ;
  assign n28179 = ( n1123 & ~n3195 ) | ( n1123 & n28178 ) | ( ~n3195 & n28178 ) ;
  assign n28172 = n8094 ^ n1484 ^ 1'b0 ;
  assign n28173 = n10115 & n28172 ;
  assign n28174 = ( n14235 & ~n14576 ) | ( n14235 & n28173 ) | ( ~n14576 & n28173 ) ;
  assign n28175 = ( n2633 & ~n6987 ) | ( n2633 & n15834 ) | ( ~n6987 & n15834 ) ;
  assign n28176 = ( n13737 & ~n28174 ) | ( n13737 & n28175 ) | ( ~n28174 & n28175 ) ;
  assign n28177 = ( n13510 & n16974 ) | ( n13510 & n28176 ) | ( n16974 & n28176 ) ;
  assign n28183 = n28182 ^ n28179 ^ n28177 ;
  assign n28184 = ~n11643 & n15568 ;
  assign n28185 = n10596 & ~n18727 ;
  assign n28186 = ( n8843 & ~n15393 ) | ( n8843 & n28185 ) | ( ~n15393 & n28185 ) ;
  assign n28187 = ( ~n12272 & n28184 ) | ( ~n12272 & n28186 ) | ( n28184 & n28186 ) ;
  assign n28188 = n1710 & n9468 ;
  assign n28189 = n28188 ^ n1271 ^ 1'b0 ;
  assign n28190 = n4601 & n21160 ;
  assign n28191 = n2200 & n28190 ;
  assign n28192 = n28191 ^ n12431 ^ n7402 ;
  assign n28193 = ( n10185 & n24702 ) | ( n10185 & n28192 ) | ( n24702 & n28192 ) ;
  assign n28194 = ( n9519 & ~n28189 ) | ( n9519 & n28193 ) | ( ~n28189 & n28193 ) ;
  assign n28195 = n20311 ^ n17724 ^ n1206 ;
  assign n28196 = n23015 ^ n6332 ^ 1'b0 ;
  assign n28197 = n28196 ^ n6165 ^ 1'b0 ;
  assign n28198 = ( n10232 & n17867 ) | ( n10232 & n28130 ) | ( n17867 & n28130 ) ;
  assign n28199 = n28198 ^ n16262 ^ n6305 ;
  assign n28200 = ~n21959 & n28199 ;
  assign n28201 = ( n5257 & n6032 ) | ( n5257 & n12621 ) | ( n6032 & n12621 ) ;
  assign n28202 = ( ~n5004 & n6646 ) | ( ~n5004 & n9374 ) | ( n6646 & n9374 ) ;
  assign n28203 = n4063 & n28202 ;
  assign n28204 = ~n28201 & n28203 ;
  assign n28205 = n3092 ^ n2837 ^ n1679 ;
  assign n28206 = ( ~n815 & n7125 ) | ( ~n815 & n28205 ) | ( n7125 & n28205 ) ;
  assign n28207 = n12190 | n12263 ;
  assign n28208 = ( n14921 & ~n17360 ) | ( n14921 & n28207 ) | ( ~n17360 & n28207 ) ;
  assign n28209 = n15441 & n20556 ;
  assign n28210 = n15546 ^ n14456 ^ 1'b0 ;
  assign n28212 = n3149 & n7053 ;
  assign n28213 = n22108 & n28212 ;
  assign n28214 = n28213 ^ n873 ^ 1'b0 ;
  assign n28211 = n11771 | n25970 ;
  assign n28215 = n28214 ^ n28211 ^ n1461 ;
  assign n28216 = ~n17982 & n27548 ;
  assign n28217 = n28216 ^ n25954 ^ 1'b0 ;
  assign n28218 = n23549 ^ n15071 ^ n8461 ;
  assign n28219 = n18540 ^ n4983 ^ 1'b0 ;
  assign n28220 = ~n16134 & n28219 ;
  assign n28221 = ~n1400 & n28220 ;
  assign n28222 = n3268 & ~n10372 ;
  assign n28223 = ( n2237 & ~n17475 ) | ( n2237 & n22896 ) | ( ~n17475 & n22896 ) ;
  assign n28224 = n2301 & ~n3847 ;
  assign n28225 = n28224 ^ n10411 ^ n9496 ;
  assign n28226 = n28225 ^ n4999 ^ 1'b0 ;
  assign n28227 = n16021 ^ n12759 ^ 1'b0 ;
  assign n28228 = n19220 & ~n25931 ;
  assign n28229 = ( n10590 & n23398 ) | ( n10590 & n28228 ) | ( n23398 & n28228 ) ;
  assign n28230 = ~n14061 & n16329 ;
  assign n28231 = n22521 & n28230 ;
  assign n28232 = ( n2386 & n2527 ) | ( n2386 & n28231 ) | ( n2527 & n28231 ) ;
  assign n28233 = ( n15002 & n15319 ) | ( n15002 & ~n15685 ) | ( n15319 & ~n15685 ) ;
  assign n28234 = n28232 | n28233 ;
  assign n28235 = ( n8538 & ~n13788 ) | ( n8538 & n28234 ) | ( ~n13788 & n28234 ) ;
  assign n28236 = n9046 | n10342 ;
  assign n28237 = n8898 | n17603 ;
  assign n28238 = ( ~n900 & n1567 ) | ( ~n900 & n28237 ) | ( n1567 & n28237 ) ;
  assign n28239 = n24328 & ~n28238 ;
  assign n28240 = n2077 & n28239 ;
  assign n28241 = n5620 ^ n1789 ^ 1'b0 ;
  assign n28242 = ( n2711 & ~n4339 ) | ( n2711 & n28241 ) | ( ~n4339 & n28241 ) ;
  assign n28243 = n16442 & n28242 ;
  assign n28244 = ( n7514 & n9650 ) | ( n7514 & ~n11509 ) | ( n9650 & ~n11509 ) ;
  assign n28245 = n2594 & ~n8369 ;
  assign n28246 = ~n18237 & n28245 ;
  assign n28247 = n11164 | n16539 ;
  assign n28248 = n28247 ^ n15890 ^ 1'b0 ;
  assign n28249 = n23797 & ~n24714 ;
  assign n28250 = n14659 & n28249 ;
  assign n28251 = ( ~n6157 & n15226 ) | ( ~n6157 & n28250 ) | ( n15226 & n28250 ) ;
  assign n28252 = n2776 | n4068 ;
  assign n28253 = n21034 ^ n5544 ^ n2752 ;
  assign n28254 = n17430 & ~n28253 ;
  assign n28255 = n28254 ^ n11828 ^ 1'b0 ;
  assign n28256 = n28252 | n28255 ;
  assign n28257 = n23829 | n28256 ;
  assign n28259 = n8791 ^ n8751 ^ n6927 ;
  assign n28260 = n10534 & ~n28259 ;
  assign n28261 = n22793 & ~n28260 ;
  assign n28262 = n28261 ^ n24549 ^ 1'b0 ;
  assign n28258 = ( n4316 & n12735 ) | ( n4316 & ~n18345 ) | ( n12735 & ~n18345 ) ;
  assign n28263 = n28262 ^ n28258 ^ n4331 ;
  assign n28264 = ( n1011 & n6800 ) | ( n1011 & ~n7403 ) | ( n6800 & ~n7403 ) ;
  assign n28265 = n28264 ^ n19010 ^ n6534 ;
  assign n28267 = n15066 ^ n5202 ^ 1'b0 ;
  assign n28268 = n4230 | n28267 ;
  assign n28266 = ( n8481 & ~n8983 ) | ( n8481 & n13085 ) | ( ~n8983 & n13085 ) ;
  assign n28269 = n28268 ^ n28266 ^ 1'b0 ;
  assign n28270 = n5013 & ~n20535 ;
  assign n28271 = ( x35 & n4650 ) | ( x35 & n4990 ) | ( n4650 & n4990 ) ;
  assign n28272 = n16284 | n28271 ;
  assign n28273 = ~n21525 & n26696 ;
  assign n28274 = n28272 & n28273 ;
  assign n28275 = n10228 & n15153 ;
  assign n28276 = n28275 ^ n21509 ^ 1'b0 ;
  assign n28277 = n25618 ^ n25085 ^ n20135 ;
  assign n28278 = n9191 & n10060 ;
  assign n28279 = ( n5799 & ~n9627 ) | ( n5799 & n28278 ) | ( ~n9627 & n28278 ) ;
  assign n28280 = n11914 ^ n3844 ^ 1'b0 ;
  assign n28281 = n10565 & ~n28280 ;
  assign n28282 = ~n19608 & n28281 ;
  assign n28283 = n28282 ^ n4577 ^ 1'b0 ;
  assign n28284 = ( n3475 & n3586 ) | ( n3475 & n14542 ) | ( n3586 & n14542 ) ;
  assign n28285 = n16808 & n28284 ;
  assign n28286 = ~n28283 & n28285 ;
  assign n28287 = ( n3593 & ~n25316 ) | ( n3593 & n28286 ) | ( ~n25316 & n28286 ) ;
  assign n28288 = ( ~n4963 & n8943 ) | ( ~n4963 & n9872 ) | ( n8943 & n9872 ) ;
  assign n28289 = ( n2585 & n11760 ) | ( n2585 & ~n28288 ) | ( n11760 & ~n28288 ) ;
  assign n28290 = n3642 & n13904 ;
  assign n28291 = ~n6414 & n28290 ;
  assign n28292 = n28291 ^ n8461 ^ n1156 ;
  assign n28293 = ( n8914 & n12479 ) | ( n8914 & ~n28292 ) | ( n12479 & ~n28292 ) ;
  assign n28294 = n9066 | n22406 ;
  assign n28295 = n28294 ^ n19038 ^ 1'b0 ;
  assign n28296 = ~n28293 & n28295 ;
  assign n28297 = ( n10140 & n28289 ) | ( n10140 & n28296 ) | ( n28289 & n28296 ) ;
  assign n28298 = n5992 ^ n5475 ^ 1'b0 ;
  assign n28299 = n6634 ^ n3765 ^ n640 ;
  assign n28300 = n28299 ^ n24157 ^ 1'b0 ;
  assign n28302 = ( n745 & n1806 ) | ( n745 & n3643 ) | ( n1806 & n3643 ) ;
  assign n28303 = ( n4844 & n16341 ) | ( n4844 & ~n28302 ) | ( n16341 & ~n28302 ) ;
  assign n28301 = n4487 ^ n4155 ^ 1'b0 ;
  assign n28304 = n28303 ^ n28301 ^ n18542 ;
  assign n28305 = n18143 & ~n28304 ;
  assign n28306 = n27063 & n28305 ;
  assign n28307 = n8174 ^ n704 ^ n688 ;
  assign n28308 = ( n3011 & n8777 ) | ( n3011 & n28307 ) | ( n8777 & n28307 ) ;
  assign n28309 = ~n10864 & n13652 ;
  assign n28310 = n5288 ^ n4373 ^ n3200 ;
  assign n28311 = ~n13318 & n28051 ;
  assign n28312 = ~n28310 & n28311 ;
  assign n28313 = ~n12546 & n14466 ;
  assign n28314 = n28313 ^ n25548 ^ 1'b0 ;
  assign n28315 = n27854 ^ n20334 ^ n5017 ;
  assign n28316 = n28315 ^ n15735 ^ 1'b0 ;
  assign n28317 = ( n1188 & n4222 ) | ( n1188 & ~n8389 ) | ( n4222 & ~n8389 ) ;
  assign n28318 = n23722 ^ n10222 ^ 1'b0 ;
  assign n28319 = n16677 | n28318 ;
  assign n28320 = n22100 ^ n12036 ^ n10807 ;
  assign n28321 = n23007 ^ n10921 ^ n9286 ;
  assign n28322 = n28321 ^ n13943 ^ n13318 ;
  assign n28323 = n28322 ^ n4045 ^ 1'b0 ;
  assign n28324 = n28320 & n28323 ;
  assign n28325 = n28324 ^ n26914 ^ n26827 ;
  assign n28326 = ( n9074 & ~n18939 ) | ( n9074 & n28202 ) | ( ~n18939 & n28202 ) ;
  assign n28327 = n10911 | n15829 ;
  assign n28328 = n6631 | n20295 ;
  assign n28329 = n28327 & ~n28328 ;
  assign n28330 = ( ~n2809 & n7452 ) | ( ~n2809 & n28329 ) | ( n7452 & n28329 ) ;
  assign n28331 = n28330 ^ n21582 ^ 1'b0 ;
  assign n28332 = n18850 & ~n28331 ;
  assign n28333 = ( n7215 & n21649 ) | ( n7215 & n23913 ) | ( n21649 & n23913 ) ;
  assign n28334 = n520 | n28333 ;
  assign n28335 = n22218 & ~n28334 ;
  assign n28336 = n18835 ^ n11071 ^ n7723 ;
  assign n28337 = ( n516 & ~n14721 ) | ( n516 & n28336 ) | ( ~n14721 & n28336 ) ;
  assign n28338 = n28337 ^ n25537 ^ n7946 ;
  assign n28339 = ( n8979 & ~n14036 ) | ( n8979 & n23544 ) | ( ~n14036 & n23544 ) ;
  assign n28345 = ( ~n15521 & n15663 ) | ( ~n15521 & n16877 ) | ( n15663 & n16877 ) ;
  assign n28344 = n19774 ^ n17098 ^ n14690 ;
  assign n28346 = n28345 ^ n28344 ^ n6242 ;
  assign n28340 = n20413 ^ n18447 ^ 1'b0 ;
  assign n28341 = n25303 | n28340 ;
  assign n28342 = n3446 & ~n28341 ;
  assign n28343 = ~n11025 & n28342 ;
  assign n28347 = n28346 ^ n28343 ^ 1'b0 ;
  assign n28348 = ( n3894 & ~n6427 ) | ( n3894 & n7722 ) | ( ~n6427 & n7722 ) ;
  assign n28349 = n13851 ^ n8413 ^ 1'b0 ;
  assign n28350 = n7459 | n28349 ;
  assign n28351 = n10641 & ~n28350 ;
  assign n28352 = n28351 ^ n22638 ^ 1'b0 ;
  assign n28353 = ( ~n4195 & n28348 ) | ( ~n4195 & n28352 ) | ( n28348 & n28352 ) ;
  assign n28354 = n28353 ^ n6587 ^ 1'b0 ;
  assign n28357 = ~n6565 & n13664 ;
  assign n28358 = n28357 ^ n26972 ^ 1'b0 ;
  assign n28359 = n1351 & ~n28358 ;
  assign n28355 = n775 & n18751 ;
  assign n28356 = n6253 & n28355 ;
  assign n28360 = n28359 ^ n28356 ^ n24373 ;
  assign n28361 = n28360 ^ n20051 ^ 1'b0 ;
  assign n28362 = n8531 & ~n14956 ;
  assign n28363 = n28362 ^ n20662 ^ 1'b0 ;
  assign n28364 = ( n1790 & n2234 ) | ( n1790 & n5512 ) | ( n2234 & n5512 ) ;
  assign n28365 = ( n1940 & ~n3026 ) | ( n1940 & n6919 ) | ( ~n3026 & n6919 ) ;
  assign n28366 = ~n26135 & n28365 ;
  assign n28367 = ( n18851 & ~n28364 ) | ( n18851 & n28366 ) | ( ~n28364 & n28366 ) ;
  assign n28368 = n2733 | n7670 ;
  assign n28369 = n23579 & n28368 ;
  assign n28370 = n6851 & n28369 ;
  assign n28371 = n28370 ^ n10781 ^ n6887 ;
  assign n28372 = n28371 ^ n14572 ^ n6753 ;
  assign n28373 = ( n6973 & n10844 ) | ( n6973 & ~n23516 ) | ( n10844 & ~n23516 ) ;
  assign n28374 = ~n27328 & n28373 ;
  assign n28375 = n28372 & n28374 ;
  assign n28376 = n28367 & ~n28375 ;
  assign n28377 = ~n8649 & n18188 ;
  assign n28378 = ~n1052 & n28377 ;
  assign n28379 = ( n16297 & n26355 ) | ( n16297 & n28378 ) | ( n26355 & n28378 ) ;
  assign n28380 = n25334 ^ n20898 ^ 1'b0 ;
  assign n28381 = ( n17240 & n20184 ) | ( n17240 & ~n26697 ) | ( n20184 & ~n26697 ) ;
  assign n28382 = n7576 | n19275 ;
  assign n28383 = ( ~n10596 & n12260 ) | ( ~n10596 & n18461 ) | ( n12260 & n18461 ) ;
  assign n28384 = ( n10678 & n12446 ) | ( n10678 & ~n28383 ) | ( n12446 & ~n28383 ) ;
  assign n28385 = ~n28382 & n28384 ;
  assign n28386 = n28385 ^ n24488 ^ 1'b0 ;
  assign n28390 = ( n10169 & n14840 ) | ( n10169 & ~n21713 ) | ( n14840 & ~n21713 ) ;
  assign n28391 = n28390 ^ n13888 ^ n6656 ;
  assign n28387 = ( n3115 & ~n4850 ) | ( n3115 & n8127 ) | ( ~n4850 & n8127 ) ;
  assign n28388 = n19792 ^ n9582 ^ n1652 ;
  assign n28389 = n28387 | n28388 ;
  assign n28392 = n28391 ^ n28389 ^ 1'b0 ;
  assign n28393 = x37 & n4650 ;
  assign n28394 = n20807 ^ n19972 ^ n8026 ;
  assign n28395 = n13747 ^ n3997 ^ 1'b0 ;
  assign n28396 = n1039 | n28395 ;
  assign n28397 = n10749 | n28396 ;
  assign n28398 = n28397 ^ n17361 ^ 1'b0 ;
  assign n28399 = n10001 & n28398 ;
  assign n28400 = ( n16540 & ~n24626 ) | ( n16540 & n28399 ) | ( ~n24626 & n28399 ) ;
  assign n28401 = n3109 & n11033 ;
  assign n28402 = n28401 ^ n4199 ^ 1'b0 ;
  assign n28403 = ( n17038 & n27112 ) | ( n17038 & n28402 ) | ( n27112 & n28402 ) ;
  assign n28404 = ~n7904 & n28403 ;
  assign n28405 = n28404 ^ n12756 ^ 1'b0 ;
  assign n28406 = n469 & n9820 ;
  assign n28407 = n28406 ^ n18853 ^ 1'b0 ;
  assign n28408 = n16634 ^ n8937 ^ x113 ;
  assign n28409 = ( x106 & n7957 ) | ( x106 & ~n9482 ) | ( n7957 & ~n9482 ) ;
  assign n28410 = n19077 ^ n3861 ^ 1'b0 ;
  assign n28411 = n28409 & n28410 ;
  assign n28412 = ( n14479 & n28408 ) | ( n14479 & n28411 ) | ( n28408 & n28411 ) ;
  assign n28416 = n11504 ^ n7378 ^ n5545 ;
  assign n28417 = n28416 ^ n7753 ^ 1'b0 ;
  assign n28414 = n25214 ^ n16158 ^ 1'b0 ;
  assign n28415 = n27572 & ~n28414 ;
  assign n28418 = n28417 ^ n28415 ^ n4560 ;
  assign n28413 = n25014 ^ n21958 ^ n10872 ;
  assign n28419 = n28418 ^ n28413 ^ n22766 ;
  assign n28420 = n25067 ^ n9280 ^ x69 ;
  assign n28421 = ( n2171 & n14474 ) | ( n2171 & n19393 ) | ( n14474 & n19393 ) ;
  assign n28422 = n15772 ^ n14382 ^ n13739 ;
  assign n28423 = n27048 ^ n13744 ^ n6769 ;
  assign n28424 = ~n28422 & n28423 ;
  assign n28425 = n28424 ^ n2769 ^ 1'b0 ;
  assign n28430 = n1155 & ~n20305 ;
  assign n28429 = n4064 & ~n16918 ;
  assign n28431 = n28430 ^ n28429 ^ 1'b0 ;
  assign n28426 = n16252 ^ n2556 ^ 1'b0 ;
  assign n28427 = n28426 ^ n13486 ^ n874 ;
  assign n28428 = ~n15490 & n28427 ;
  assign n28432 = n28431 ^ n28428 ^ n20215 ;
  assign n28433 = ~n12668 & n28212 ;
  assign n28434 = n24514 ^ n688 ^ 1'b0 ;
  assign n28435 = n20387 | n28434 ;
  assign n28436 = n6431 & n7479 ;
  assign n28441 = n28152 ^ n11245 ^ n4785 ;
  assign n28442 = n28441 ^ n1362 ^ 1'b0 ;
  assign n28439 = n26686 ^ n10615 ^ 1'b0 ;
  assign n28437 = n17693 ^ n11346 ^ 1'b0 ;
  assign n28438 = n8996 & ~n28437 ;
  assign n28440 = n28439 ^ n28438 ^ n17865 ;
  assign n28443 = n28442 ^ n28440 ^ n1296 ;
  assign n28446 = n7881 & ~n15210 ;
  assign n28444 = n10134 ^ n5165 ^ n1034 ;
  assign n28445 = n18360 & ~n28444 ;
  assign n28447 = n28446 ^ n28445 ^ 1'b0 ;
  assign n28448 = ~n24818 & n28447 ;
  assign n28449 = n10451 ^ n6701 ^ 1'b0 ;
  assign n28453 = n10556 ^ n9076 ^ n2765 ;
  assign n28450 = ( ~n971 & n4044 ) | ( ~n971 & n19477 ) | ( n4044 & n19477 ) ;
  assign n28451 = ( x94 & n349 ) | ( x94 & n25419 ) | ( n349 & n25419 ) ;
  assign n28452 = ( n23825 & ~n28450 ) | ( n23825 & n28451 ) | ( ~n28450 & n28451 ) ;
  assign n28454 = n28453 ^ n28452 ^ 1'b0 ;
  assign n28455 = n17821 | n27689 ;
  assign n28456 = n23947 | n28455 ;
  assign n28457 = n4649 & n28456 ;
  assign n28458 = n25379 | n28457 ;
  assign n28459 = ( n4440 & n12172 ) | ( n4440 & n14923 ) | ( n12172 & n14923 ) ;
  assign n28460 = n7879 ^ n588 ^ 1'b0 ;
  assign n28461 = x150 | n28460 ;
  assign n28462 = n28461 ^ n22037 ^ n3504 ;
  assign n28463 = n8024 | n9146 ;
  assign n28464 = n7419 | n28463 ;
  assign n28465 = ~n9279 & n28464 ;
  assign n28466 = n28462 & n28465 ;
  assign n28467 = ( n10556 & ~n28459 ) | ( n10556 & n28466 ) | ( ~n28459 & n28466 ) ;
  assign n28468 = ~n4134 & n5826 ;
  assign n28469 = n18455 ^ n7859 ^ 1'b0 ;
  assign n28470 = ( n8184 & ~n9401 ) | ( n8184 & n28469 ) | ( ~n9401 & n28469 ) ;
  assign n28471 = ~n2790 & n28470 ;
  assign n28472 = n8403 | n10364 ;
  assign n28473 = n2976 & ~n28472 ;
  assign n28474 = n20448 & n28473 ;
  assign n28475 = n3215 ^ n2340 ^ 1'b0 ;
  assign n28476 = ~n19794 & n28475 ;
  assign n28477 = n14854 ^ n4735 ^ 1'b0 ;
  assign n28478 = ( n14121 & ~n16903 ) | ( n14121 & n28477 ) | ( ~n16903 & n28477 ) ;
  assign n28479 = n14294 | n20778 ;
  assign n28480 = n28479 ^ n26075 ^ n21333 ;
  assign n28481 = n28478 | n28480 ;
  assign n28482 = n24232 | n28481 ;
  assign n28483 = n13634 & ~n24816 ;
  assign n28484 = n28483 ^ n4004 ^ 1'b0 ;
  assign n28485 = n28484 ^ n7322 ^ x81 ;
  assign n28486 = n26640 ^ x73 ^ 1'b0 ;
  assign n28490 = n24231 ^ n1454 ^ 1'b0 ;
  assign n28487 = ~n1581 & n24625 ;
  assign n28488 = ~n7977 & n28487 ;
  assign n28489 = ( n7723 & ~n15618 ) | ( n7723 & n28488 ) | ( ~n15618 & n28488 ) ;
  assign n28491 = n28490 ^ n28489 ^ 1'b0 ;
  assign n28494 = ( n2611 & n4937 ) | ( n2611 & n12803 ) | ( n4937 & n12803 ) ;
  assign n28495 = n12948 | n23951 ;
  assign n28496 = ( n24157 & n28494 ) | ( n24157 & ~n28495 ) | ( n28494 & ~n28495 ) ;
  assign n28493 = n9575 & n22153 ;
  assign n28492 = n24612 ^ n15653 ^ 1'b0 ;
  assign n28497 = n28496 ^ n28493 ^ n28492 ;
  assign n28503 = ( n8057 & n10854 ) | ( n8057 & n24585 ) | ( n10854 & n24585 ) ;
  assign n28504 = ( n7086 & ~n13337 ) | ( n7086 & n28503 ) | ( ~n13337 & n28503 ) ;
  assign n28498 = n9951 ^ n5873 ^ 1'b0 ;
  assign n28499 = ( ~n1130 & n4591 ) | ( ~n1130 & n28498 ) | ( n4591 & n28498 ) ;
  assign n28500 = n939 | n16307 ;
  assign n28501 = n28500 ^ n6905 ^ 1'b0 ;
  assign n28502 = n28499 & ~n28501 ;
  assign n28505 = n28504 ^ n28502 ^ n4492 ;
  assign n28506 = n7417 ^ n6927 ^ n4342 ;
  assign n28507 = n21478 ^ n3148 ^ 1'b0 ;
  assign n28508 = n28506 & ~n28507 ;
  assign n28510 = ( ~n8538 & n19948 ) | ( ~n8538 & n20863 ) | ( n19948 & n20863 ) ;
  assign n28509 = ~n8734 & n9617 ;
  assign n28511 = n28510 ^ n28509 ^ n5860 ;
  assign n28512 = n4951 ^ n2459 ^ x149 ;
  assign n28513 = n1592 & ~n28512 ;
  assign n28514 = n6731 & ~n28513 ;
  assign n28515 = n28514 ^ n6459 ^ 1'b0 ;
  assign n28518 = ( n8999 & n14883 ) | ( n8999 & ~n25296 ) | ( n14883 & ~n25296 ) ;
  assign n28516 = n16483 ^ n10984 ^ n5685 ;
  assign n28517 = n26573 & ~n28516 ;
  assign n28519 = n28518 ^ n28517 ^ 1'b0 ;
  assign n28520 = n18157 ^ n12874 ^ 1'b0 ;
  assign n28522 = n28148 ^ n6068 ^ 1'b0 ;
  assign n28521 = n2884 & ~n13737 ;
  assign n28523 = n28522 ^ n28521 ^ 1'b0 ;
  assign n28524 = ~n20531 & n28523 ;
  assign n28525 = n4478 ^ n2936 ^ 1'b0 ;
  assign n28526 = n18500 ^ n6678 ^ n4466 ;
  assign n28527 = n7333 | n17417 ;
  assign n28528 = n7704 | n28527 ;
  assign n28529 = ~n2053 & n6283 ;
  assign n28530 = n10886 & ~n20127 ;
  assign n28531 = ( n5784 & n16676 ) | ( n5784 & n20669 ) | ( n16676 & n20669 ) ;
  assign n28532 = ( x14 & n8134 ) | ( x14 & ~n11301 ) | ( n8134 & ~n11301 ) ;
  assign n28533 = n28531 & ~n28532 ;
  assign n28534 = n5793 & n19035 ;
  assign n28535 = n10709 & n28534 ;
  assign n28536 = n28535 ^ n6350 ^ n1793 ;
  assign n28537 = n28536 ^ n1564 ^ x107 ;
  assign n28538 = ( n19931 & n28241 ) | ( n19931 & n28537 ) | ( n28241 & n28537 ) ;
  assign n28539 = ( n1558 & n2086 ) | ( n1558 & n22054 ) | ( n2086 & n22054 ) ;
  assign n28540 = n15566 ^ n13052 ^ n332 ;
  assign n28541 = n21376 ^ n2513 ^ n2426 ;
  assign n28542 = n28541 ^ n27869 ^ n1236 ;
  assign n28543 = n16887 ^ n5407 ^ n1896 ;
  assign n28544 = n28543 ^ n7672 ^ n662 ;
  assign n28545 = ( n555 & ~n1816 ) | ( n555 & n3032 ) | ( ~n1816 & n3032 ) ;
  assign n28546 = n28545 ^ n23432 ^ n3904 ;
  assign n28547 = n20592 ^ n2207 ^ 1'b0 ;
  assign n28548 = n17642 & ~n28547 ;
  assign n28549 = n2007 | n20277 ;
  assign n28550 = n1319 | n28549 ;
  assign n28551 = n9085 ^ n6308 ^ 1'b0 ;
  assign n28552 = ~n8616 & n28551 ;
  assign n28553 = n24911 ^ n19598 ^ 1'b0 ;
  assign n28554 = n28552 & n28553 ;
  assign n28557 = n18153 ^ n741 ^ 1'b0 ;
  assign n28558 = n7630 | n28557 ;
  assign n28559 = n28558 ^ n16093 ^ n13070 ;
  assign n28555 = ~n1384 & n11257 ;
  assign n28556 = ~n261 & n28555 ;
  assign n28560 = n28559 ^ n28556 ^ n25280 ;
  assign n28563 = n4354 & n6591 ;
  assign n28564 = n28563 ^ n5672 ^ 1'b0 ;
  assign n28561 = n15998 ^ n4638 ^ n4101 ;
  assign n28562 = n16684 | n28561 ;
  assign n28565 = n28564 ^ n28562 ^ n2964 ;
  assign n28566 = n6962 & n15004 ;
  assign n28568 = ~n9294 & n12980 ;
  assign n28567 = n3092 & n6092 ;
  assign n28569 = n28568 ^ n28567 ^ 1'b0 ;
  assign n28570 = n28569 ^ n18061 ^ 1'b0 ;
  assign n28571 = ~n609 & n28570 ;
  assign n28572 = n1173 | n1289 ;
  assign n28573 = n28572 ^ n12060 ^ 1'b0 ;
  assign n28574 = ( ~n1004 & n25067 ) | ( ~n1004 & n28573 ) | ( n25067 & n28573 ) ;
  assign n28575 = n11321 & ~n11849 ;
  assign n28576 = n28575 ^ n1424 ^ 1'b0 ;
  assign n28577 = n8849 & ~n28576 ;
  assign n28578 = n2455 ^ n1592 ^ 1'b0 ;
  assign n28579 = n9401 & ~n28578 ;
  assign n28580 = n9804 ^ n3689 ^ 1'b0 ;
  assign n28581 = ~n7608 & n28580 ;
  assign n28582 = n28581 ^ n15561 ^ 1'b0 ;
  assign n28583 = n25691 ^ n4263 ^ 1'b0 ;
  assign n28584 = n28582 | n28583 ;
  assign n28585 = ( ~n25231 & n28579 ) | ( ~n25231 & n28584 ) | ( n28579 & n28584 ) ;
  assign n28589 = n4586 ^ n2640 ^ 1'b0 ;
  assign n28590 = n3499 & n28589 ;
  assign n28591 = ~n271 & n28590 ;
  assign n28586 = ~n8094 & n11492 ;
  assign n28587 = n28586 ^ n2000 ^ 1'b0 ;
  assign n28588 = n28587 ^ n28201 ^ n1863 ;
  assign n28592 = n28591 ^ n28588 ^ n12089 ;
  assign n28593 = n18944 ^ n12442 ^ n10521 ;
  assign n28594 = n10247 & n20694 ;
  assign n28595 = ~n843 & n28594 ;
  assign n28596 = ( n5545 & n28593 ) | ( n5545 & n28595 ) | ( n28593 & n28595 ) ;
  assign n28597 = n28592 & ~n28596 ;
  assign n28598 = n28597 ^ n19267 ^ 1'b0 ;
  assign n28599 = ( ~n13907 & n15321 ) | ( ~n13907 & n28598 ) | ( n15321 & n28598 ) ;
  assign n28600 = n289 & n28599 ;
  assign n28601 = n28600 ^ n9905 ^ 1'b0 ;
  assign n28602 = n26502 ^ n323 ^ 1'b0 ;
  assign n28603 = n28602 ^ n21039 ^ n13238 ;
  assign n28604 = n25378 ^ n1845 ^ 1'b0 ;
  assign n28605 = n2348 & ~n14992 ;
  assign n28606 = ( n4623 & ~n21380 ) | ( n4623 & n28605 ) | ( ~n21380 & n28605 ) ;
  assign n28607 = ( n1634 & ~n3546 ) | ( n1634 & n11881 ) | ( ~n3546 & n11881 ) ;
  assign n28608 = n2960 & ~n11567 ;
  assign n28609 = n28608 ^ n21058 ^ 1'b0 ;
  assign n28610 = n28609 ^ n14813 ^ 1'b0 ;
  assign n28611 = ( n19363 & ~n28607 ) | ( n19363 & n28610 ) | ( ~n28607 & n28610 ) ;
  assign n28612 = n10450 & ~n28611 ;
  assign n28613 = ~n28606 & n28612 ;
  assign n28614 = n10086 ^ n7947 ^ 1'b0 ;
  assign n28615 = n28614 ^ n18792 ^ n17736 ;
  assign n28618 = n11009 ^ n10744 ^ n2679 ;
  assign n28616 = ~n5514 & n6977 ;
  assign n28617 = n28616 ^ n5609 ^ 1'b0 ;
  assign n28619 = n28618 ^ n28617 ^ n10609 ;
  assign n28620 = ( n10240 & n16195 ) | ( n10240 & n24232 ) | ( n16195 & n24232 ) ;
  assign n28621 = ~n1187 & n4733 ;
  assign n28622 = ( ~n5720 & n28620 ) | ( ~n5720 & n28621 ) | ( n28620 & n28621 ) ;
  assign n28623 = n11079 | n22919 ;
  assign n28624 = n10620 | n28623 ;
  assign n28625 = n683 | n14613 ;
  assign n28626 = n28625 ^ n20799 ^ 1'b0 ;
  assign n28628 = n1378 | n4527 ;
  assign n28629 = n1447 & ~n28628 ;
  assign n28627 = ( n7362 & n9728 ) | ( n7362 & ~n19510 ) | ( n9728 & ~n19510 ) ;
  assign n28630 = n28629 ^ n28627 ^ n8566 ;
  assign n28632 = n14561 ^ n5270 ^ 1'b0 ;
  assign n28633 = n19084 | n28632 ;
  assign n28631 = n12170 | n17237 ;
  assign n28634 = n28633 ^ n28631 ^ 1'b0 ;
  assign n28635 = ( ~n2538 & n6749 ) | ( ~n2538 & n28634 ) | ( n6749 & n28634 ) ;
  assign n28636 = n28635 ^ n4781 ^ 1'b0 ;
  assign n28637 = n19392 ^ n15676 ^ 1'b0 ;
  assign n28638 = ( n1317 & n13801 ) | ( n1317 & ~n28637 ) | ( n13801 & ~n28637 ) ;
  assign n28639 = n10895 ^ n8407 ^ 1'b0 ;
  assign n28640 = n10676 ^ n6129 ^ n1644 ;
  assign n28641 = ~n5057 & n28640 ;
  assign n28642 = n8820 ^ n8523 ^ n4291 ;
  assign n28643 = n265 & n28642 ;
  assign n28644 = ~n1980 & n10073 ;
  assign n28645 = n28644 ^ n4438 ^ 1'b0 ;
  assign n28646 = n25530 | n28645 ;
  assign n28647 = n3355 | n28646 ;
  assign n28648 = n19489 ^ n12169 ^ 1'b0 ;
  assign n28649 = n28648 ^ n16119 ^ n16073 ;
  assign n28651 = ( n7350 & n7482 ) | ( n7350 & ~n13218 ) | ( n7482 & ~n13218 ) ;
  assign n28650 = n15941 ^ n11906 ^ n6791 ;
  assign n28652 = n28651 ^ n28650 ^ n5098 ;
  assign n28653 = n950 | n8762 ;
  assign n28654 = n7306 & ~n28653 ;
  assign n28655 = n22479 & ~n27482 ;
  assign n28656 = n28655 ^ n26273 ^ 1'b0 ;
  assign n28659 = ~n5361 & n8463 ;
  assign n28660 = ~n4971 & n28659 ;
  assign n28657 = n20457 ^ n5935 ^ 1'b0 ;
  assign n28658 = n16179 & n28657 ;
  assign n28661 = n28660 ^ n28658 ^ n22061 ;
  assign n28662 = ~n3126 & n28661 ;
  assign n28667 = n12005 | n15641 ;
  assign n28668 = n7795 | n28667 ;
  assign n28665 = n1634 & n3530 ;
  assign n28666 = ( ~n5074 & n10216 ) | ( ~n5074 & n28665 ) | ( n10216 & n28665 ) ;
  assign n28669 = n28668 ^ n28666 ^ n11740 ;
  assign n28663 = n25296 ^ n12289 ^ n6337 ;
  assign n28664 = ( ~n2373 & n4053 ) | ( ~n2373 & n28663 ) | ( n4053 & n28663 ) ;
  assign n28670 = n28669 ^ n28664 ^ n23402 ;
  assign n28671 = n18402 ^ n6033 ^ 1'b0 ;
  assign n28672 = n1479 | n4733 ;
  assign n28674 = n16824 ^ n10782 ^ 1'b0 ;
  assign n28673 = n11261 | n12291 ;
  assign n28675 = n28674 ^ n28673 ^ 1'b0 ;
  assign n28676 = n638 | n17232 ;
  assign n28677 = ( n10310 & ~n19787 ) | ( n10310 & n28676 ) | ( ~n19787 & n28676 ) ;
  assign n28678 = n6947 ^ n2684 ^ 1'b0 ;
  assign n28679 = ( n22049 & n28677 ) | ( n22049 & ~n28678 ) | ( n28677 & ~n28678 ) ;
  assign n28680 = n28679 ^ n9697 ^ 1'b0 ;
  assign n28681 = n15814 ^ n10092 ^ 1'b0 ;
  assign n28684 = n13117 ^ n6246 ^ n2143 ;
  assign n28682 = ( n608 & n723 ) | ( n608 & ~n3704 ) | ( n723 & ~n3704 ) ;
  assign n28683 = n17671 | n28682 ;
  assign n28685 = n28684 ^ n28683 ^ n10582 ;
  assign n28686 = ~n24836 & n28685 ;
  assign n28687 = n28686 ^ n12267 ^ 1'b0 ;
  assign n28688 = ( ~n15544 & n28681 ) | ( ~n15544 & n28687 ) | ( n28681 & n28687 ) ;
  assign n28689 = n6904 & ~n17114 ;
  assign n28690 = n28689 ^ x55 ^ 1'b0 ;
  assign n28691 = n28690 ^ n10174 ^ n3363 ;
  assign n28692 = ( n473 & n6360 ) | ( n473 & n10952 ) | ( n6360 & n10952 ) ;
  assign n28693 = n28692 ^ n20840 ^ 1'b0 ;
  assign n28694 = ~n13969 & n28693 ;
  assign n28695 = n28694 ^ n12603 ^ 1'b0 ;
  assign n28696 = ( n480 & ~n28691 ) | ( n480 & n28695 ) | ( ~n28691 & n28695 ) ;
  assign n28697 = n9447 & n28696 ;
  assign n28698 = n2118 | n12638 ;
  assign n28699 = n27482 ^ n15852 ^ 1'b0 ;
  assign n28700 = ~n4307 & n17330 ;
  assign n28701 = ( n1304 & n14149 ) | ( n1304 & ~n23574 ) | ( n14149 & ~n23574 ) ;
  assign n28702 = n25725 ^ n22455 ^ n9031 ;
  assign n28703 = ( n7899 & n18715 ) | ( n7899 & n28702 ) | ( n18715 & n28702 ) ;
  assign n28704 = ~n13356 & n21519 ;
  assign n28705 = n8017 & n28704 ;
  assign n28710 = n10533 ^ n6188 ^ 1'b0 ;
  assign n28711 = n666 & n28710 ;
  assign n28712 = n9576 & n28711 ;
  assign n28713 = n7069 & n28712 ;
  assign n28706 = n8881 & n9932 ;
  assign n28707 = n28706 ^ n7561 ^ 1'b0 ;
  assign n28708 = n19408 ^ n14219 ^ 1'b0 ;
  assign n28709 = ( n18548 & n28707 ) | ( n18548 & n28708 ) | ( n28707 & n28708 ) ;
  assign n28714 = n28713 ^ n28709 ^ 1'b0 ;
  assign n28715 = n28705 | n28714 ;
  assign n28716 = n9696 ^ n7365 ^ n1118 ;
  assign n28717 = n1385 | n11685 ;
  assign n28718 = n28717 ^ n491 ^ 1'b0 ;
  assign n28719 = ( n1861 & n2083 ) | ( n1861 & n28718 ) | ( n2083 & n28718 ) ;
  assign n28720 = n4067 | n28719 ;
  assign n28721 = n11303 ^ n916 ^ n343 ;
  assign n28722 = n28721 ^ n25306 ^ n786 ;
  assign n28723 = ( n15062 & ~n28720 ) | ( n15062 & n28722 ) | ( ~n28720 & n28722 ) ;
  assign n28724 = ( n4995 & n5160 ) | ( n4995 & ~n12399 ) | ( n5160 & ~n12399 ) ;
  assign n28725 = ( ~n20730 & n25524 ) | ( ~n20730 & n28724 ) | ( n25524 & n28724 ) ;
  assign n28726 = n3248 | n17033 ;
  assign n28727 = n18779 ^ n2998 ^ 1'b0 ;
  assign n28728 = n28464 ^ n11068 ^ n1458 ;
  assign n28729 = n15104 | n28728 ;
  assign n28730 = n28729 ^ n7914 ^ 1'b0 ;
  assign n28731 = n25369 ^ n18690 ^ 1'b0 ;
  assign n28732 = ~n22747 & n28731 ;
  assign n28733 = ~n14663 & n28732 ;
  assign n28734 = n28730 & n28733 ;
  assign n28735 = n18586 ^ n13816 ^ n12591 ;
  assign n28736 = ~n20086 & n28735 ;
  assign n28744 = n9227 ^ n6582 ^ 1'b0 ;
  assign n28745 = x239 & ~n28744 ;
  assign n28739 = x55 & ~n2510 ;
  assign n28740 = n28739 ^ n1967 ^ 1'b0 ;
  assign n28737 = ~n847 & n2621 ;
  assign n28738 = n28737 ^ n21853 ^ 1'b0 ;
  assign n28741 = n28740 ^ n28738 ^ n19174 ;
  assign n28742 = n28741 ^ n11810 ^ n2480 ;
  assign n28743 = ( ~n3878 & n7415 ) | ( ~n3878 & n28742 ) | ( n7415 & n28742 ) ;
  assign n28746 = n28745 ^ n28743 ^ 1'b0 ;
  assign n28747 = n25059 & ~n28746 ;
  assign n28749 = ( n2265 & ~n2508 ) | ( n2265 & n12338 ) | ( ~n2508 & n12338 ) ;
  assign n28750 = n28749 ^ n17166 ^ 1'b0 ;
  assign n28748 = n13720 & n20240 ;
  assign n28751 = n28750 ^ n28748 ^ 1'b0 ;
  assign n28752 = ~n5226 & n14585 ;
  assign n28753 = n15092 | n28752 ;
  assign n28754 = ( n19528 & n22840 ) | ( n19528 & ~n28753 ) | ( n22840 & ~n28753 ) ;
  assign n28755 = ( n8019 & n16503 ) | ( n8019 & ~n23121 ) | ( n16503 & ~n23121 ) ;
  assign n28756 = n28755 ^ n19753 ^ n17397 ;
  assign n28757 = n5946 & n13569 ;
  assign n28760 = n485 & n8324 ;
  assign n28761 = n28760 ^ n20596 ^ 1'b0 ;
  assign n28758 = n5471 ^ n1838 ^ 1'b0 ;
  assign n28759 = n13128 & n28758 ;
  assign n28762 = n28761 ^ n28759 ^ 1'b0 ;
  assign n28763 = n16123 & n22884 ;
  assign n28765 = n9664 & ~n17732 ;
  assign n28766 = n28765 ^ n7766 ^ 1'b0 ;
  assign n28764 = n5031 & n5424 ;
  assign n28767 = n28766 ^ n28764 ^ 1'b0 ;
  assign n28768 = ~n28763 & n28767 ;
  assign n28769 = ~n5260 & n28768 ;
  assign n28770 = n3993 ^ n1790 ^ n1656 ;
  assign n28771 = n28770 ^ n21453 ^ n917 ;
  assign n28772 = n28771 ^ n21965 ^ n13043 ;
  assign n28774 = n13647 & ~n17671 ;
  assign n28775 = n28774 ^ n14788 ^ n9353 ;
  assign n28773 = ( n9685 & n18645 ) | ( n9685 & ~n26626 ) | ( n18645 & ~n26626 ) ;
  assign n28776 = n28775 ^ n28773 ^ n26263 ;
  assign n28777 = ( n4839 & n8888 ) | ( n4839 & ~n16602 ) | ( n8888 & ~n16602 ) ;
  assign n28778 = n6860 & n28777 ;
  assign n28779 = n28778 ^ n6323 ^ n1734 ;
  assign n28780 = n3019 | n16395 ;
  assign n28781 = n28780 ^ n18711 ^ n17924 ;
  assign n28782 = n16205 & ~n19335 ;
  assign n28783 = ~n4609 & n28782 ;
  assign n28784 = n17646 ^ n9067 ^ 1'b0 ;
  assign n28785 = n28784 ^ n24174 ^ 1'b0 ;
  assign n28786 = n18751 & n28785 ;
  assign n28788 = n1839 & ~n2595 ;
  assign n28787 = ( n13519 & n15249 ) | ( n13519 & ~n17472 ) | ( n15249 & ~n17472 ) ;
  assign n28789 = n28788 ^ n28787 ^ n16917 ;
  assign n28790 = n18819 & ~n19828 ;
  assign n28791 = n28084 ^ n4189 ^ 1'b0 ;
  assign n28792 = n11996 & ~n28791 ;
  assign n28793 = ( n4983 & n7531 ) | ( n4983 & ~n9798 ) | ( n7531 & ~n9798 ) ;
  assign n28794 = n28793 ^ n10377 ^ 1'b0 ;
  assign n28795 = n28794 ^ n20343 ^ 1'b0 ;
  assign n28796 = ( n28790 & n28792 ) | ( n28790 & ~n28795 ) | ( n28792 & ~n28795 ) ;
  assign n28797 = n15027 ^ n12370 ^ 1'b0 ;
  assign n28798 = n15490 | n28797 ;
  assign n28799 = ( ~n8986 & n9810 ) | ( ~n8986 & n28798 ) | ( n9810 & n28798 ) ;
  assign n28800 = ~n1381 & n26618 ;
  assign n28801 = n1020 | n2445 ;
  assign n28802 = ~n4325 & n28801 ;
  assign n28803 = ~n9967 & n28802 ;
  assign n28804 = n28803 ^ n1697 ^ 1'b0 ;
  assign n28805 = n28800 & n28804 ;
  assign n28806 = n19990 ^ n15229 ^ 1'b0 ;
  assign n28807 = n20135 ^ n19400 ^ 1'b0 ;
  assign n28808 = n26044 ^ n24858 ^ 1'b0 ;
  assign n28809 = n26243 ^ n17875 ^ 1'b0 ;
  assign n28810 = n26140 ^ n2097 ^ 1'b0 ;
  assign n28811 = n15552 ^ n1938 ^ 1'b0 ;
  assign n28812 = n5768 | n28811 ;
  assign n28813 = n2976 | n6182 ;
  assign n28814 = n20073 ^ n17416 ^ 1'b0 ;
  assign n28815 = ( ~n5337 & n28813 ) | ( ~n5337 & n28814 ) | ( n28813 & n28814 ) ;
  assign n28816 = ( ~n9944 & n11729 ) | ( ~n9944 & n20207 ) | ( n11729 & n20207 ) ;
  assign n28817 = ( n28812 & n28815 ) | ( n28812 & ~n28816 ) | ( n28815 & ~n28816 ) ;
  assign n28818 = ( ~n2138 & n9656 ) | ( ~n2138 & n28817 ) | ( n9656 & n28817 ) ;
  assign n28819 = ~n12402 & n16855 ;
  assign n28820 = n2931 & n28819 ;
  assign n28821 = n13233 ^ n6411 ^ 1'b0 ;
  assign n28822 = n14271 | n28821 ;
  assign n28823 = n8549 & ~n13913 ;
  assign n28824 = n28823 ^ n16367 ^ n2421 ;
  assign n28826 = ( ~n638 & n8052 ) | ( ~n638 & n13164 ) | ( n8052 & n13164 ) ;
  assign n28825 = ~n10683 & n20092 ;
  assign n28827 = n28826 ^ n28825 ^ 1'b0 ;
  assign n28828 = ~n19181 & n28827 ;
  assign n28829 = ~n28824 & n28828 ;
  assign n28831 = ~n2728 & n14977 ;
  assign n28832 = n28831 ^ n19503 ^ 1'b0 ;
  assign n28833 = ~n12808 & n17435 ;
  assign n28834 = n28832 & n28833 ;
  assign n28830 = n19652 & n21161 ;
  assign n28835 = n28834 ^ n28830 ^ 1'b0 ;
  assign n28836 = n3605 & ~n15522 ;
  assign n28837 = n28836 ^ n18940 ^ 1'b0 ;
  assign n28839 = ( ~n1034 & n8127 ) | ( ~n1034 & n11916 ) | ( n8127 & n11916 ) ;
  assign n28838 = n9363 | n12446 ;
  assign n28840 = n28839 ^ n28838 ^ n2274 ;
  assign n28841 = n28840 ^ n15631 ^ n6705 ;
  assign n28842 = n9770 ^ n6548 ^ n5604 ;
  assign n28843 = n12062 & n28842 ;
  assign n28844 = n3755 & n28843 ;
  assign n28845 = ( n17053 & ~n27825 ) | ( n17053 & n28844 ) | ( ~n27825 & n28844 ) ;
  assign n28846 = n13396 ^ n368 ^ 1'b0 ;
  assign n28847 = n28845 & n28846 ;
  assign n28848 = ( n10526 & ~n13319 ) | ( n10526 & n18195 ) | ( ~n13319 & n18195 ) ;
  assign n28849 = ( n3206 & n11218 ) | ( n3206 & ~n28848 ) | ( n11218 & ~n28848 ) ;
  assign n28850 = n27694 ^ n7003 ^ n4213 ;
  assign n28851 = n26771 ^ n25354 ^ n23644 ;
  assign n28852 = ( n22028 & n24545 ) | ( n22028 & n28851 ) | ( n24545 & n28851 ) ;
  assign n28853 = n13400 | n22907 ;
  assign n28854 = n4391 | n28853 ;
  assign n28855 = n17497 ^ n9433 ^ n1838 ;
  assign n28856 = ~n27063 & n28855 ;
  assign n28857 = ~n28854 & n28856 ;
  assign n28858 = n28202 | n28857 ;
  assign n28860 = ( ~n1984 & n6654 ) | ( ~n1984 & n23140 ) | ( n6654 & n23140 ) ;
  assign n28859 = n10751 & ~n12562 ;
  assign n28861 = n28860 ^ n28859 ^ 1'b0 ;
  assign n28862 = n2382 | n16311 ;
  assign n28863 = n1451 & ~n17879 ;
  assign n28864 = n2952 & n28863 ;
  assign n28865 = ( n6903 & n9371 ) | ( n6903 & n17636 ) | ( n9371 & n17636 ) ;
  assign n28866 = ( ~n2092 & n9909 ) | ( ~n2092 & n10046 ) | ( n9909 & n10046 ) ;
  assign n28867 = n28866 ^ n17599 ^ n4367 ;
  assign n28868 = ( ~n28864 & n28865 ) | ( ~n28864 & n28867 ) | ( n28865 & n28867 ) ;
  assign n28869 = n17858 ^ n10207 ^ 1'b0 ;
  assign n28870 = n14108 | n28869 ;
  assign n28871 = ( ~n25374 & n26443 ) | ( ~n25374 & n28870 ) | ( n26443 & n28870 ) ;
  assign n28872 = n16893 ^ n11404 ^ 1'b0 ;
  assign n28873 = ~n10827 & n15597 ;
  assign n28874 = n14593 ^ n6959 ^ 1'b0 ;
  assign n28875 = ~n28873 & n28874 ;
  assign n28876 = ~n6883 & n28875 ;
  assign n28877 = n28872 & n28876 ;
  assign n28878 = ( n313 & ~n17421 ) | ( n313 & n27576 ) | ( ~n17421 & n27576 ) ;
  assign n28880 = n26394 ^ n21143 ^ n14268 ;
  assign n28879 = ~n21665 & n23815 ;
  assign n28881 = n28880 ^ n28879 ^ 1'b0 ;
  assign n28882 = ( ~n7339 & n9964 ) | ( ~n7339 & n28881 ) | ( n9964 & n28881 ) ;
  assign n28883 = n17083 ^ n11545 ^ 1'b0 ;
  assign n28884 = x32 & n28883 ;
  assign n28885 = n17732 ^ n7236 ^ n5670 ;
  assign n28886 = n28885 ^ n13943 ^ 1'b0 ;
  assign n28887 = n14383 | n28886 ;
  assign n28888 = n28887 ^ n15463 ^ 1'b0 ;
  assign n28889 = n17407 ^ n13573 ^ 1'b0 ;
  assign n28890 = ( n2210 & n15976 ) | ( n2210 & n19193 ) | ( n15976 & n19193 ) ;
  assign n28891 = ( ~n4693 & n28333 ) | ( ~n4693 & n28890 ) | ( n28333 & n28890 ) ;
  assign n28892 = n5175 ^ n3276 ^ 1'b0 ;
  assign n28893 = n28892 ^ n9385 ^ 1'b0 ;
  assign n28894 = n21367 & ~n28893 ;
  assign n28895 = n28894 ^ n4551 ^ 1'b0 ;
  assign n28896 = ( n5838 & n12222 ) | ( n5838 & n13423 ) | ( n12222 & n13423 ) ;
  assign n28897 = n2380 | n28896 ;
  assign n28898 = n28897 ^ n15124 ^ n7292 ;
  assign n28904 = n7196 ^ n7124 ^ 1'b0 ;
  assign n28899 = n1595 & n6998 ;
  assign n28900 = n1979 ^ n1421 ^ 1'b0 ;
  assign n28901 = n28900 ^ n25653 ^ 1'b0 ;
  assign n28902 = n15501 | n28901 ;
  assign n28903 = n28899 | n28902 ;
  assign n28905 = n28904 ^ n28903 ^ 1'b0 ;
  assign n28906 = n11051 ^ n1753 ^ 1'b0 ;
  assign n28907 = n6259 & ~n11110 ;
  assign n28908 = n28907 ^ n12005 ^ 1'b0 ;
  assign n28909 = ( x144 & n3208 ) | ( x144 & n28908 ) | ( n3208 & n28908 ) ;
  assign n28910 = n20510 ^ n16143 ^ n5114 ;
  assign n28911 = n16830 | n20733 ;
  assign n28912 = n28911 ^ n21006 ^ 1'b0 ;
  assign n28913 = n28320 | n28912 ;
  assign n28914 = n27046 ^ n14125 ^ 1'b0 ;
  assign n28917 = n9409 ^ n7498 ^ n4693 ;
  assign n28915 = n7633 | n8869 ;
  assign n28916 = n28915 ^ n18074 ^ n4066 ;
  assign n28918 = n28917 ^ n28916 ^ n16668 ;
  assign n28922 = n5498 ^ n325 ^ n289 ;
  assign n28919 = n20053 ^ n7672 ^ n3861 ;
  assign n28920 = n28919 ^ n21348 ^ n934 ;
  assign n28921 = n28920 ^ n14271 ^ n12158 ;
  assign n28923 = n28922 ^ n28921 ^ 1'b0 ;
  assign n28924 = ( x211 & n2096 ) | ( x211 & n17879 ) | ( n2096 & n17879 ) ;
  assign n28925 = n12376 & ~n13879 ;
  assign n28926 = n12026 & ~n16226 ;
  assign n28927 = n11071 & n28926 ;
  assign n28928 = ( n5471 & n18998 ) | ( n5471 & ~n28927 ) | ( n18998 & ~n28927 ) ;
  assign n28929 = n19408 ^ n426 ^ 1'b0 ;
  assign n28930 = ( n5254 & n5874 ) | ( n5254 & ~n7097 ) | ( n5874 & ~n7097 ) ;
  assign n28931 = n10870 | n28582 ;
  assign n28932 = n28930 | n28931 ;
  assign n28933 = ~n12146 & n28932 ;
  assign n28934 = n21706 ^ n624 ^ 1'b0 ;
  assign n28935 = ~n22945 & n28934 ;
  assign n28936 = ~n15064 & n28935 ;
  assign n28937 = n28936 ^ n13446 ^ 1'b0 ;
  assign n28938 = n22766 | n28937 ;
  assign n28939 = ( ~n21436 & n23147 ) | ( ~n21436 & n25725 ) | ( n23147 & n25725 ) ;
  assign n28940 = n3706 | n24608 ;
  assign n28941 = n18469 ^ n658 ^ 1'b0 ;
  assign n28942 = n17573 & ~n28941 ;
  assign n28943 = ( ~n3140 & n28940 ) | ( ~n3140 & n28942 ) | ( n28940 & n28942 ) ;
  assign n28944 = n17448 | n28943 ;
  assign n28945 = ( n8691 & ~n10984 ) | ( n8691 & n28944 ) | ( ~n10984 & n28944 ) ;
  assign n28946 = n16420 ^ n6476 ^ 1'b0 ;
  assign n28947 = n28946 ^ n22083 ^ n20161 ;
  assign n28948 = n19934 ^ n8704 ^ n6255 ;
  assign n28949 = n9730 | n28948 ;
  assign n28950 = n13372 ^ n5456 ^ 1'b0 ;
  assign n28951 = n8109 & n28950 ;
  assign n28952 = n297 & ~n11034 ;
  assign n28953 = n28952 ^ n22613 ^ n12680 ;
  assign n28954 = n28953 ^ n27763 ^ n11285 ;
  assign n28955 = ( ~x130 & n15221 ) | ( ~x130 & n28954 ) | ( n15221 & n28954 ) ;
  assign n28960 = n14365 ^ n7737 ^ n2206 ;
  assign n28961 = n28960 ^ n12542 ^ n1866 ;
  assign n28958 = ~n3861 & n26405 ;
  assign n28959 = n28958 ^ n26375 ^ 1'b0 ;
  assign n28956 = ( n5741 & ~n10260 ) | ( n5741 & n17610 ) | ( ~n10260 & n17610 ) ;
  assign n28957 = n28956 ^ n28301 ^ n10755 ;
  assign n28962 = n28961 ^ n28959 ^ n28957 ;
  assign n28963 = n1390 & n1798 ;
  assign n28964 = n1826 & n28963 ;
  assign n28965 = n2948 & ~n11177 ;
  assign n28966 = ( n7914 & n28964 ) | ( n7914 & ~n28965 ) | ( n28964 & ~n28965 ) ;
  assign n28967 = n15304 ^ n7962 ^ n3675 ;
  assign n28968 = ( n6611 & n28966 ) | ( n6611 & n28967 ) | ( n28966 & n28967 ) ;
  assign n28969 = ( ~n3611 & n14956 ) | ( ~n3611 & n28968 ) | ( n14956 & n28968 ) ;
  assign n28970 = n22244 ^ n21679 ^ 1'b0 ;
  assign n28971 = ~n22379 & n28970 ;
  assign n28972 = n28971 ^ n23954 ^ 1'b0 ;
  assign n28973 = n15912 ^ n8403 ^ 1'b0 ;
  assign n28974 = ( n6091 & ~n7859 ) | ( n6091 & n10266 ) | ( ~n7859 & n10266 ) ;
  assign n28975 = n28974 ^ n25081 ^ 1'b0 ;
  assign n28976 = ( ~n8773 & n20786 ) | ( ~n8773 & n28975 ) | ( n20786 & n28975 ) ;
  assign n28977 = ( n7483 & ~n18920 ) | ( n7483 & n26517 ) | ( ~n18920 & n26517 ) ;
  assign n28978 = ( n5367 & n8260 ) | ( n5367 & ~n11634 ) | ( n8260 & ~n11634 ) ;
  assign n28979 = n23059 | n26897 ;
  assign n28980 = ( n23484 & n28978 ) | ( n23484 & n28979 ) | ( n28978 & n28979 ) ;
  assign n28981 = n4812 ^ x12 ^ 1'b0 ;
  assign n28982 = n23043 ^ n8911 ^ n5754 ;
  assign n28983 = ( n268 & ~n14889 ) | ( n268 & n24756 ) | ( ~n14889 & n24756 ) ;
  assign n28986 = n14465 ^ n10367 ^ n6724 ;
  assign n28984 = n19730 ^ n1072 ^ 1'b0 ;
  assign n28985 = ~n24422 & n28984 ;
  assign n28987 = n28986 ^ n28985 ^ n27559 ;
  assign n28988 = n12244 ^ n2050 ^ 1'b0 ;
  assign n28989 = ( ~n3166 & n7746 ) | ( ~n3166 & n9192 ) | ( n7746 & n9192 ) ;
  assign n28990 = n12476 & n28989 ;
  assign n28991 = n28990 ^ n3941 ^ 1'b0 ;
  assign n28992 = n17245 ^ n9391 ^ 1'b0 ;
  assign n28993 = ( ~n28988 & n28991 ) | ( ~n28988 & n28992 ) | ( n28991 & n28992 ) ;
  assign n28994 = ( n9541 & n28987 ) | ( n9541 & n28993 ) | ( n28987 & n28993 ) ;
  assign n28995 = ( n16066 & ~n28983 ) | ( n16066 & n28994 ) | ( ~n28983 & n28994 ) ;
  assign n28996 = ( n2482 & ~n16513 ) | ( n2482 & n16849 ) | ( ~n16513 & n16849 ) ;
  assign n28997 = n28996 ^ n22337 ^ n12637 ;
  assign n28998 = ( n20135 & n20748 ) | ( n20135 & n28997 ) | ( n20748 & n28997 ) ;
  assign n28999 = ( n8205 & ~n11416 ) | ( n8205 & n22604 ) | ( ~n11416 & n22604 ) ;
  assign n29000 = n14041 ^ n8356 ^ n7595 ;
  assign n29002 = n18619 ^ n6485 ^ n5342 ;
  assign n29003 = ( n466 & n3837 ) | ( n466 & n7162 ) | ( n3837 & n7162 ) ;
  assign n29004 = ( n7853 & ~n13192 ) | ( n7853 & n29003 ) | ( ~n13192 & n29003 ) ;
  assign n29005 = ( n707 & n29002 ) | ( n707 & n29004 ) | ( n29002 & n29004 ) ;
  assign n29001 = n16710 & ~n24087 ;
  assign n29006 = n29005 ^ n29001 ^ 1'b0 ;
  assign n29007 = ( n9530 & ~n12648 ) | ( n9530 & n15154 ) | ( ~n12648 & n15154 ) ;
  assign n29008 = ( n2651 & n19358 ) | ( n2651 & ~n29007 ) | ( n19358 & ~n29007 ) ;
  assign n29009 = n5033 & n9531 ;
  assign n29010 = n29009 ^ n8364 ^ 1'b0 ;
  assign n29011 = n4387 ^ n3712 ^ 1'b0 ;
  assign n29012 = n29011 ^ n15668 ^ n1934 ;
  assign n29013 = n9153 ^ n1289 ^ 1'b0 ;
  assign n29014 = ( n6204 & n6399 ) | ( n6204 & ~n22182 ) | ( n6399 & ~n22182 ) ;
  assign n29015 = ~n16570 & n29014 ;
  assign n29016 = n29015 ^ n4097 ^ 1'b0 ;
  assign n29017 = n6688 | n27989 ;
  assign n29018 = n8346 | n29017 ;
  assign n29019 = n5924 ^ n5260 ^ n5101 ;
  assign n29020 = n29019 ^ n8682 ^ 1'b0 ;
  assign n29023 = n16497 & ~n25145 ;
  assign n29021 = n17388 ^ n3927 ^ 1'b0 ;
  assign n29022 = ~n11264 & n29021 ;
  assign n29024 = n29023 ^ n29022 ^ 1'b0 ;
  assign n29025 = n29020 & n29024 ;
  assign n29026 = n1633 & ~n21809 ;
  assign n29027 = ~n10544 & n29026 ;
  assign n29028 = ( n4052 & n20818 ) | ( n4052 & n29027 ) | ( n20818 & n29027 ) ;
  assign n29029 = n4517 & ~n26687 ;
  assign n29030 = n15429 ^ n2869 ^ 1'b0 ;
  assign n29031 = n2464 | n9624 ;
  assign n29032 = n26648 | n29031 ;
  assign n29033 = ~n15319 & n17273 ;
  assign n29038 = n7182 & n24016 ;
  assign n29039 = n29038 ^ n3427 ^ 1'b0 ;
  assign n29034 = n2046 & ~n4422 ;
  assign n29035 = n29034 ^ n7853 ^ 1'b0 ;
  assign n29036 = n29035 ^ n6100 ^ n5278 ;
  assign n29037 = n16001 | n29036 ;
  assign n29040 = n29039 ^ n29037 ^ 1'b0 ;
  assign n29041 = n29040 ^ n3202 ^ 1'b0 ;
  assign n29042 = n6115 | n20552 ;
  assign n29043 = n29042 ^ n18504 ^ 1'b0 ;
  assign n29044 = n7640 & n29043 ;
  assign n29045 = n24312 ^ n13497 ^ n8900 ;
  assign n29046 = n29045 ^ n19618 ^ n12968 ;
  assign n29047 = n5789 & n23793 ;
  assign n29048 = n15476 ^ n6451 ^ 1'b0 ;
  assign n29049 = ( n2456 & n8907 ) | ( n2456 & ~n19524 ) | ( n8907 & ~n19524 ) ;
  assign n29050 = n29048 | n29049 ;
  assign n29051 = n29050 ^ n7220 ^ n3017 ;
  assign n29054 = n11129 & ~n11668 ;
  assign n29055 = n29054 ^ n20712 ^ 1'b0 ;
  assign n29053 = ( ~n3348 & n5665 ) | ( ~n3348 & n5909 ) | ( n5665 & n5909 ) ;
  assign n29052 = n21048 ^ n12929 ^ n5139 ;
  assign n29056 = n29055 ^ n29053 ^ n29052 ;
  assign n29057 = n29056 ^ n19412 ^ n10833 ;
  assign n29058 = ( n3522 & ~n4866 ) | ( n3522 & n5186 ) | ( ~n4866 & n5186 ) ;
  assign n29059 = ( ~n6488 & n18575 ) | ( ~n6488 & n29058 ) | ( n18575 & n29058 ) ;
  assign n29060 = n29059 ^ n15323 ^ 1'b0 ;
  assign n29061 = n12513 ^ n473 ^ 1'b0 ;
  assign n29062 = n20781 ^ n2212 ^ 1'b0 ;
  assign n29063 = ~n27860 & n29062 ;
  assign n29064 = ~n29061 & n29063 ;
  assign n29065 = n5417 & ~n16211 ;
  assign n29066 = ( n2077 & n7524 ) | ( n2077 & ~n11760 ) | ( n7524 & ~n11760 ) ;
  assign n29067 = n14865 ^ n11976 ^ 1'b0 ;
  assign n29068 = ( n408 & n8561 ) | ( n408 & n29067 ) | ( n8561 & n29067 ) ;
  assign n29069 = n29066 | n29068 ;
  assign n29070 = n7193 | n29069 ;
  assign n29071 = n25939 ^ n8858 ^ n2908 ;
  assign n29072 = n3323 & ~n13820 ;
  assign n29073 = ~n26026 & n29072 ;
  assign n29074 = n6009 | n29073 ;
  assign n29075 = n29071 & ~n29074 ;
  assign n29076 = n24476 ^ n13618 ^ 1'b0 ;
  assign n29077 = n3692 & n29076 ;
  assign n29078 = n29077 ^ n25037 ^ 1'b0 ;
  assign n29080 = n12328 ^ n11966 ^ 1'b0 ;
  assign n29081 = ( ~n3487 & n11218 ) | ( ~n3487 & n29080 ) | ( n11218 & n29080 ) ;
  assign n29079 = n5504 | n5778 ;
  assign n29082 = n29081 ^ n29079 ^ 1'b0 ;
  assign n29083 = n29082 ^ n28936 ^ n9519 ;
  assign n29093 = n392 ^ n265 ^ 1'b0 ;
  assign n29094 = n3459 & ~n29093 ;
  assign n29095 = ( n5086 & n14361 ) | ( n5086 & ~n18159 ) | ( n14361 & ~n18159 ) ;
  assign n29096 = ( n13698 & n29094 ) | ( n13698 & n29095 ) | ( n29094 & n29095 ) ;
  assign n29084 = n4817 ^ n324 ^ n283 ;
  assign n29085 = n20203 ^ n17541 ^ 1'b0 ;
  assign n29086 = ( n17670 & ~n29084 ) | ( n17670 & n29085 ) | ( ~n29084 & n29085 ) ;
  assign n29087 = n6860 & ~n18352 ;
  assign n29088 = n29086 & n29087 ;
  assign n29089 = n1856 | n2944 ;
  assign n29090 = n29088 & ~n29089 ;
  assign n29091 = n29090 ^ n19561 ^ n17605 ;
  assign n29092 = ( n489 & ~n8594 ) | ( n489 & n29091 ) | ( ~n8594 & n29091 ) ;
  assign n29097 = n29096 ^ n29092 ^ n13042 ;
  assign n29099 = ~n10864 & n20511 ;
  assign n29100 = n28479 & n29099 ;
  assign n29098 = ( ~n2608 & n8738 ) | ( ~n2608 & n12032 ) | ( n8738 & n12032 ) ;
  assign n29101 = n29100 ^ n29098 ^ n15326 ;
  assign n29102 = n24079 & ~n29101 ;
  assign n29103 = n3368 ^ n929 ^ n662 ;
  assign n29104 = n29103 ^ n19760 ^ 1'b0 ;
  assign n29105 = ( n10468 & n22957 ) | ( n10468 & n29104 ) | ( n22957 & n29104 ) ;
  assign n29106 = n11108 & ~n16001 ;
  assign n29107 = ~n13564 & n29106 ;
  assign n29108 = n3584 & ~n8082 ;
  assign n29109 = n29108 ^ n26284 ^ 1'b0 ;
  assign n29110 = n29107 | n29109 ;
  assign n29111 = n14146 ^ n8745 ^ 1'b0 ;
  assign n29112 = n4271 & ~n29111 ;
  assign n29113 = ( n3148 & ~n3315 ) | ( n3148 & n14420 ) | ( ~n3315 & n14420 ) ;
  assign n29114 = n12072 ^ n8400 ^ n7244 ;
  assign n29115 = n29113 & ~n29114 ;
  assign n29116 = ( n29110 & n29112 ) | ( n29110 & ~n29115 ) | ( n29112 & ~n29115 ) ;
  assign n29117 = n1555 ^ n1340 ^ 1'b0 ;
  assign n29118 = n12501 ^ n1246 ^ 1'b0 ;
  assign n29119 = n2026 | n29118 ;
  assign n29120 = ( n12722 & n18681 ) | ( n12722 & ~n29119 ) | ( n18681 & ~n29119 ) ;
  assign n29121 = n3225 | n13134 ;
  assign n29122 = n12653 | n20859 ;
  assign n29123 = n26045 & ~n29122 ;
  assign n29124 = n853 & n14183 ;
  assign n29125 = n28103 ^ n15754 ^ n10761 ;
  assign n29126 = ~n17344 & n23579 ;
  assign n29127 = ~n29125 & n29126 ;
  assign n29128 = n29127 ^ n22875 ^ 1'b0 ;
  assign n29129 = n21682 | n29128 ;
  assign n29130 = n28847 ^ n11686 ^ 1'b0 ;
  assign n29131 = n23804 | n29130 ;
  assign n29132 = ( n2769 & n5092 ) | ( n2769 & n26843 ) | ( n5092 & n26843 ) ;
  assign n29133 = n29108 ^ n12746 ^ n3353 ;
  assign n29134 = n29133 ^ n28125 ^ 1'b0 ;
  assign n29135 = x84 & n4247 ;
  assign n29136 = ~n8567 & n29135 ;
  assign n29137 = n9766 & n29136 ;
  assign n29138 = n14710 & ~n28966 ;
  assign n29139 = n23948 & n29138 ;
  assign n29140 = n20035 ^ n14447 ^ n3115 ;
  assign n29141 = n28708 ^ n21473 ^ n2611 ;
  assign n29142 = ( n8838 & ~n9839 ) | ( n8838 & n23963 ) | ( ~n9839 & n23963 ) ;
  assign n29143 = ( ~n4225 & n8601 ) | ( ~n4225 & n22170 ) | ( n8601 & n22170 ) ;
  assign n29144 = ~n1166 & n29143 ;
  assign n29145 = n5991 ^ n3575 ^ 1'b0 ;
  assign n29146 = ~n6795 & n29145 ;
  assign n29147 = n1892 | n27312 ;
  assign n29148 = ~n29146 & n29147 ;
  assign n29149 = n29144 | n29148 ;
  assign n29150 = n29149 ^ n13642 ^ 1'b0 ;
  assign n29151 = n11820 ^ n2979 ^ 1'b0 ;
  assign n29152 = ~n4605 & n5495 ;
  assign n29153 = ~n13142 & n29152 ;
  assign n29154 = n2804 ^ n1806 ^ 1'b0 ;
  assign n29155 = n13693 | n29154 ;
  assign n29156 = ( n6897 & n23403 ) | ( n6897 & n29155 ) | ( n23403 & n29155 ) ;
  assign n29157 = ( n1515 & n22747 ) | ( n1515 & ~n29156 ) | ( n22747 & ~n29156 ) ;
  assign n29158 = ( n10474 & n25486 ) | ( n10474 & n29157 ) | ( n25486 & n29157 ) ;
  assign n29159 = ~n7658 & n16078 ;
  assign n29160 = n29159 ^ n2376 ^ x124 ;
  assign n29161 = ( n4747 & ~n5426 ) | ( n4747 & n29160 ) | ( ~n5426 & n29160 ) ;
  assign n29162 = n28163 ^ n3204 ^ 1'b0 ;
  assign n29163 = ( ~n13400 & n15441 ) | ( ~n13400 & n21887 ) | ( n15441 & n21887 ) ;
  assign n29164 = n29163 ^ n5984 ^ n3476 ;
  assign n29165 = n29164 ^ n16811 ^ 1'b0 ;
  assign n29166 = n13850 ^ x57 ^ 1'b0 ;
  assign n29167 = n17410 & ~n29166 ;
  assign n29168 = n11798 ^ n3452 ^ x247 ;
  assign n29169 = ~n8843 & n29168 ;
  assign n29170 = ( n10290 & n14636 ) | ( n10290 & n29169 ) | ( n14636 & n29169 ) ;
  assign n29171 = ~n510 & n1193 ;
  assign n29172 = n29170 & ~n29171 ;
  assign n29173 = n29172 ^ n18379 ^ 1'b0 ;
  assign n29174 = ( ~n15816 & n28851 ) | ( ~n15816 & n29173 ) | ( n28851 & n29173 ) ;
  assign n29175 = ~n15502 & n16042 ;
  assign n29176 = n21457 & n29175 ;
  assign n29177 = n8862 ^ n2859 ^ 1'b0 ;
  assign n29178 = ~n29176 & n29177 ;
  assign n29179 = n29178 ^ n1916 ^ 1'b0 ;
  assign n29180 = n27310 ^ n15517 ^ 1'b0 ;
  assign n29181 = n3342 & ~n16741 ;
  assign n29182 = n297 & n29181 ;
  assign n29183 = n10676 & n29182 ;
  assign n29184 = ( n6237 & n29180 ) | ( n6237 & ~n29183 ) | ( n29180 & ~n29183 ) ;
  assign n29185 = n4532 | n10011 ;
  assign n29186 = n29185 ^ n8649 ^ 1'b0 ;
  assign n29187 = n29186 ^ n20275 ^ n16724 ;
  assign n29190 = n27766 ^ n3983 ^ 1'b0 ;
  assign n29188 = ( n897 & n18907 ) | ( n897 & ~n28291 ) | ( n18907 & ~n28291 ) ;
  assign n29189 = ~n20469 & n29188 ;
  assign n29191 = n29190 ^ n29189 ^ 1'b0 ;
  assign n29192 = n29191 ^ n20003 ^ 1'b0 ;
  assign n29193 = ~n25514 & n29192 ;
  assign n29194 = n20698 ^ n4584 ^ 1'b0 ;
  assign n29201 = n25514 ^ n475 ^ 1'b0 ;
  assign n29195 = n12578 ^ n7239 ^ 1'b0 ;
  assign n29196 = ~n4061 & n29195 ;
  assign n29197 = n29196 ^ n5679 ^ 1'b0 ;
  assign n29198 = n17879 | n29197 ;
  assign n29199 = n25970 | n29198 ;
  assign n29200 = ~n19533 & n29199 ;
  assign n29202 = n29201 ^ n29200 ^ 1'b0 ;
  assign n29204 = n15453 ^ n6824 ^ 1'b0 ;
  assign n29203 = n18697 | n19322 ;
  assign n29205 = n29204 ^ n29203 ^ 1'b0 ;
  assign n29206 = ( n15913 & ~n19331 ) | ( n15913 & n29205 ) | ( ~n19331 & n29205 ) ;
  assign n29207 = n17898 ^ n8229 ^ x229 ;
  assign n29208 = n29068 ^ n7027 ^ 1'b0 ;
  assign n29209 = ( n3621 & ~n13243 ) | ( n3621 & n29208 ) | ( ~n13243 & n29208 ) ;
  assign n29210 = n6645 ^ n5323 ^ 1'b0 ;
  assign n29211 = ~n25908 & n29210 ;
  assign n29212 = n18958 | n28996 ;
  assign n29213 = n17482 & ~n29212 ;
  assign n29214 = ( n2230 & n2517 ) | ( n2230 & n26832 ) | ( n2517 & n26832 ) ;
  assign n29215 = n29214 ^ n20428 ^ n7709 ;
  assign n29216 = ~n6523 & n21850 ;
  assign n29217 = ~n19438 & n29216 ;
  assign n29218 = n29215 | n29217 ;
  assign n29219 = n29213 & ~n29218 ;
  assign n29220 = n1673 & n6319 ;
  assign n29221 = ( n3860 & n4393 ) | ( n3860 & n5257 ) | ( n4393 & n5257 ) ;
  assign n29222 = ( ~n21379 & n29220 ) | ( ~n21379 & n29221 ) | ( n29220 & n29221 ) ;
  assign n29223 = n6411 & ~n9310 ;
  assign n29224 = n12196 ^ n8274 ^ 1'b0 ;
  assign n29225 = n29060 & ~n29224 ;
  assign n29226 = n9282 ^ n1152 ^ 1'b0 ;
  assign n29227 = n14452 & ~n29226 ;
  assign n29228 = n29227 ^ n26217 ^ n631 ;
  assign n29229 = n29228 ^ n19905 ^ n5435 ;
  assign n29234 = ~n2593 & n21674 ;
  assign n29232 = ( n12659 & n13799 ) | ( n12659 & n26343 ) | ( n13799 & n26343 ) ;
  assign n29233 = ( n18993 & n20464 ) | ( n18993 & n29232 ) | ( n20464 & n29232 ) ;
  assign n29230 = n22904 ^ n2527 ^ 1'b0 ;
  assign n29231 = ~n3029 & n29230 ;
  assign n29235 = n29234 ^ n29233 ^ n29231 ;
  assign n29236 = ~n681 & n23254 ;
  assign n29237 = ~n25709 & n29236 ;
  assign n29238 = n2381 & n10672 ;
  assign n29239 = n29238 ^ n21141 ^ 1'b0 ;
  assign n29240 = n29239 ^ n1595 ^ 1'b0 ;
  assign n29241 = n27140 & n29240 ;
  assign n29242 = ( n2800 & n7546 ) | ( n2800 & n29241 ) | ( n7546 & n29241 ) ;
  assign n29243 = ~n2282 & n9292 ;
  assign n29244 = ( ~n5734 & n8656 ) | ( ~n5734 & n29243 ) | ( n8656 & n29243 ) ;
  assign n29245 = n29244 ^ n26230 ^ n22220 ;
  assign n29246 = ( n1081 & n21839 ) | ( n1081 & ~n29245 ) | ( n21839 & ~n29245 ) ;
  assign n29247 = n18424 ^ n5378 ^ 1'b0 ;
  assign n29248 = ( ~n5962 & n17494 ) | ( ~n5962 & n29247 ) | ( n17494 & n29247 ) ;
  assign n29249 = n6926 & ~n10781 ;
  assign n29250 = n29249 ^ n27849 ^ 1'b0 ;
  assign n29251 = n4837 | n12702 ;
  assign n29252 = n29251 ^ n9508 ^ 1'b0 ;
  assign n29253 = n19523 & n29252 ;
  assign n29254 = n16153 ^ n13033 ^ 1'b0 ;
  assign n29255 = n5193 | n29254 ;
  assign n29256 = n11948 & n16329 ;
  assign n29257 = n29256 ^ n28037 ^ 1'b0 ;
  assign n29258 = n17543 & ~n29257 ;
  assign n29264 = ( n4263 & n12297 ) | ( n4263 & n18744 ) | ( n12297 & n18744 ) ;
  assign n29259 = n5403 ^ n4779 ^ n3325 ;
  assign n29260 = n9221 ^ n5456 ^ 1'b0 ;
  assign n29261 = ~n21136 & n29260 ;
  assign n29262 = n29259 & n29261 ;
  assign n29263 = ~n16077 & n29262 ;
  assign n29265 = n29264 ^ n29263 ^ 1'b0 ;
  assign n29268 = ~n9959 & n16209 ;
  assign n29269 = n29268 ^ n12390 ^ 1'b0 ;
  assign n29270 = n29269 ^ n10464 ^ 1'b0 ;
  assign n29266 = n19316 ^ n9854 ^ n5309 ;
  assign n29267 = n29266 ^ n12018 ^ n7537 ;
  assign n29271 = n29270 ^ n29267 ^ n16188 ;
  assign n29272 = n11115 ^ n4393 ^ n4045 ;
  assign n29273 = n1558 & n29272 ;
  assign n29274 = ~n8191 & n29273 ;
  assign n29275 = n4793 & ~n5147 ;
  assign n29276 = n29275 ^ n12544 ^ 1'b0 ;
  assign n29277 = ( n12012 & n29274 ) | ( n12012 & ~n29276 ) | ( n29274 & ~n29276 ) ;
  assign n29278 = ~n16649 & n20404 ;
  assign n29279 = ~n21446 & n29278 ;
  assign n29280 = ( n1210 & n4317 ) | ( n1210 & n5044 ) | ( n4317 & n5044 ) ;
  assign n29281 = ( n1227 & ~n8127 ) | ( n1227 & n29280 ) | ( ~n8127 & n29280 ) ;
  assign n29282 = n29281 ^ n10823 ^ n9156 ;
  assign n29285 = n15132 ^ n13599 ^ n10190 ;
  assign n29283 = n9491 ^ n4923 ^ 1'b0 ;
  assign n29284 = n8592 | n29283 ;
  assign n29286 = n29285 ^ n29284 ^ n14833 ;
  assign n29290 = n9876 ^ x117 ^ 1'b0 ;
  assign n29287 = n7217 ^ n7082 ^ n352 ;
  assign n29288 = n29287 ^ n9299 ^ n1751 ;
  assign n29289 = n29288 ^ n7686 ^ n5557 ;
  assign n29291 = n29290 ^ n29289 ^ 1'b0 ;
  assign n29292 = n693 & n5415 ;
  assign n29293 = n29292 ^ n1311 ^ 1'b0 ;
  assign n29294 = n11919 | n15796 ;
  assign n29295 = ( n5611 & ~n21264 ) | ( n5611 & n25057 ) | ( ~n21264 & n25057 ) ;
  assign n29296 = n26185 ^ n21542 ^ n5867 ;
  assign n29297 = ( ~n10005 & n12008 ) | ( ~n10005 & n28080 ) | ( n12008 & n28080 ) ;
  assign n29298 = n967 | n16588 ;
  assign n29299 = n19174 | n29298 ;
  assign n29301 = n13564 ^ n1372 ^ 1'b0 ;
  assign n29302 = n3070 | n29301 ;
  assign n29300 = n9349 & ~n21944 ;
  assign n29303 = n29302 ^ n29300 ^ 1'b0 ;
  assign n29304 = n21769 ^ n13181 ^ n4933 ;
  assign n29307 = n5052 | n20559 ;
  assign n29308 = n29307 ^ n4740 ^ 1'b0 ;
  assign n29309 = n18389 | n29308 ;
  assign n29310 = n29309 ^ n13088 ^ 1'b0 ;
  assign n29305 = n20246 ^ n13616 ^ n2378 ;
  assign n29306 = n5263 & ~n29305 ;
  assign n29311 = n29310 ^ n29306 ^ n17693 ;
  assign n29312 = ( ~n17075 & n29304 ) | ( ~n17075 & n29311 ) | ( n29304 & n29311 ) ;
  assign n29314 = n25221 ^ n23210 ^ n11478 ;
  assign n29313 = n8987 ^ n6432 ^ n5456 ;
  assign n29315 = n29314 ^ n29313 ^ n12186 ;
  assign n29317 = n17888 ^ n6036 ^ n5297 ;
  assign n29316 = ( ~n2386 & n4317 ) | ( ~n2386 & n18516 ) | ( n4317 & n18516 ) ;
  assign n29318 = n29317 ^ n29316 ^ 1'b0 ;
  assign n29319 = n20135 ^ n564 ^ 1'b0 ;
  assign n29320 = n25643 & n29319 ;
  assign n29322 = n7835 ^ n6740 ^ 1'b0 ;
  assign n29323 = n23318 & ~n29322 ;
  assign n29321 = ~n657 & n4476 ;
  assign n29324 = n29323 ^ n29321 ^ 1'b0 ;
  assign n29325 = n29320 | n29324 ;
  assign n29326 = ( n1264 & ~n3186 ) | ( n1264 & n27270 ) | ( ~n3186 & n27270 ) ;
  assign n29327 = ~n25142 & n25540 ;
  assign n29328 = n29327 ^ n9673 ^ 1'b0 ;
  assign n29329 = n10124 & ~n26601 ;
  assign n29330 = n29329 ^ n8959 ^ 1'b0 ;
  assign n29334 = n2752 | n4793 ;
  assign n29335 = ( ~n12315 & n26575 ) | ( ~n12315 & n29334 ) | ( n26575 & n29334 ) ;
  assign n29331 = n2084 & n26376 ;
  assign n29332 = n29331 ^ n21825 ^ n7675 ;
  assign n29333 = n17708 & ~n29332 ;
  assign n29336 = n29335 ^ n29333 ^ 1'b0 ;
  assign n29337 = n14838 ^ n767 ^ 1'b0 ;
  assign n29338 = n29336 | n29337 ;
  assign n29339 = n23052 ^ n16543 ^ n2386 ;
  assign n29340 = n1494 & n7577 ;
  assign n29341 = n29340 ^ n5437 ^ 1'b0 ;
  assign n29342 = ( n9582 & ~n16603 ) | ( n9582 & n29341 ) | ( ~n16603 & n29341 ) ;
  assign n29343 = n6448 | n29342 ;
  assign n29344 = n22293 ^ n1652 ^ 1'b0 ;
  assign n29345 = ( n320 & n7732 ) | ( n320 & ~n29344 ) | ( n7732 & ~n29344 ) ;
  assign n29346 = n6253 | n29345 ;
  assign n29347 = n29346 ^ n8648 ^ 1'b0 ;
  assign n29348 = n4340 ^ x173 ^ 1'b0 ;
  assign n29349 = n12772 & ~n27075 ;
  assign n29350 = n29349 ^ n16942 ^ n11461 ;
  assign n29351 = n29348 | n29350 ;
  assign n29352 = n29351 ^ n24533 ^ 1'b0 ;
  assign n29353 = n9617 | n14446 ;
  assign n29354 = n21049 ^ n14645 ^ n4101 ;
  assign n29355 = ( n7931 & n29353 ) | ( n7931 & ~n29354 ) | ( n29353 & ~n29354 ) ;
  assign n29356 = n10532 ^ n1511 ^ 1'b0 ;
  assign n29357 = n29355 & n29356 ;
  assign n29358 = n436 & n15157 ;
  assign n29359 = ( n8320 & ~n15804 ) | ( n8320 & n27160 ) | ( ~n15804 & n27160 ) ;
  assign n29360 = ( ~n6046 & n26294 ) | ( ~n6046 & n29359 ) | ( n26294 & n29359 ) ;
  assign n29361 = n7253 ^ n6484 ^ n5696 ;
  assign n29362 = n29361 ^ n14310 ^ n13069 ;
  assign n29363 = n23663 ^ n2485 ^ 1'b0 ;
  assign n29364 = n7574 | n29363 ;
  assign n29365 = n7759 & ~n29364 ;
  assign n29366 = ~n29362 & n29365 ;
  assign n29367 = n29366 ^ n17132 ^ n12346 ;
  assign n29368 = n5064 | n10019 ;
  assign n29369 = n29368 ^ n23978 ^ 1'b0 ;
  assign n29370 = ~n3636 & n29369 ;
  assign n29371 = n18354 ^ n7786 ^ 1'b0 ;
  assign n29372 = ~n16603 & n29371 ;
  assign n29373 = ( n6448 & ~n10465 ) | ( n6448 & n20052 ) | ( ~n10465 & n20052 ) ;
  assign n29374 = n1733 & ~n5918 ;
  assign n29375 = ~n29373 & n29374 ;
  assign n29376 = n1610 & ~n19689 ;
  assign n29377 = n29376 ^ n28728 ^ 1'b0 ;
  assign n29380 = ( n14544 & n17768 ) | ( n14544 & ~n23976 ) | ( n17768 & ~n23976 ) ;
  assign n29378 = n1953 ^ x184 ^ 1'b0 ;
  assign n29379 = ( ~n1277 & n7234 ) | ( ~n1277 & n29378 ) | ( n7234 & n29378 ) ;
  assign n29381 = n29380 ^ n29379 ^ n11709 ;
  assign n29382 = n29381 ^ n7616 ^ n1668 ;
  assign n29383 = ~n2282 & n29382 ;
  assign n29384 = n25385 ^ n13859 ^ 1'b0 ;
  assign n29385 = ( n4066 & n5831 ) | ( n4066 & ~n9412 ) | ( n5831 & ~n9412 ) ;
  assign n29386 = n29385 ^ n7477 ^ x225 ;
  assign n29387 = ( n9530 & n10950 ) | ( n9530 & ~n28905 ) | ( n10950 & ~n28905 ) ;
  assign n29388 = n18458 ^ n13772 ^ n8007 ;
  assign n29391 = ( n929 & n4261 ) | ( n929 & ~n7007 ) | ( n4261 & ~n7007 ) ;
  assign n29389 = n27765 ^ n14429 ^ n5088 ;
  assign n29390 = ~n10014 & n29389 ;
  assign n29392 = n29391 ^ n29390 ^ 1'b0 ;
  assign n29393 = n24250 & ~n29392 ;
  assign n29394 = n29393 ^ n3369 ^ 1'b0 ;
  assign n29395 = n28563 & ~n29394 ;
  assign n29396 = n20213 & ~n26914 ;
  assign n29397 = n1032 & n29396 ;
  assign n29398 = n28609 ^ n5338 ^ 1'b0 ;
  assign n29399 = n7233 ^ n2257 ^ n2092 ;
  assign n29400 = n29398 & ~n29399 ;
  assign n29401 = n6752 & ~n27805 ;
  assign n29402 = ( n10056 & n10255 ) | ( n10056 & n21755 ) | ( n10255 & n21755 ) ;
  assign n29403 = n23318 ^ n13504 ^ n6044 ;
  assign n29404 = ~n10952 & n18126 ;
  assign n29405 = ( n959 & ~n7393 ) | ( n959 & n28345 ) | ( ~n7393 & n28345 ) ;
  assign n29406 = n20234 ^ n3696 ^ 1'b0 ;
  assign n29407 = n11373 & n29406 ;
  assign n29408 = n29407 ^ n21332 ^ n11788 ;
  assign n29409 = n11808 & ~n18300 ;
  assign n29410 = n29409 ^ n306 ^ 1'b0 ;
  assign n29411 = n23178 & ~n29410 ;
  assign n29412 = ( ~n5551 & n13977 ) | ( ~n5551 & n29411 ) | ( n13977 & n29411 ) ;
  assign n29413 = n23100 ^ n19432 ^ n8867 ;
  assign n29414 = n5846 & n18158 ;
  assign n29415 = n16412 ^ n3637 ^ 1'b0 ;
  assign n29416 = n27862 ^ n14191 ^ n6923 ;
  assign n29417 = ( n16736 & ~n18788 ) | ( n16736 & n29416 ) | ( ~n18788 & n29416 ) ;
  assign n29418 = n21142 & n29417 ;
  assign n29419 = ~n5746 & n8723 ;
  assign n29420 = n29419 ^ n2640 ^ 1'b0 ;
  assign n29421 = n12230 ^ n6862 ^ 1'b0 ;
  assign n29422 = n561 & ~n1343 ;
  assign n29423 = ~n29421 & n29422 ;
  assign n29424 = n29420 & ~n29423 ;
  assign n29425 = ~n4914 & n29424 ;
  assign n29426 = n2948 & ~n24188 ;
  assign n29427 = n17969 ^ n12301 ^ n11812 ;
  assign n29428 = n7118 & n29427 ;
  assign n29434 = n17799 ^ n10565 ^ n1271 ;
  assign n29435 = ( n8739 & ~n25238 ) | ( n8739 & n29434 ) | ( ~n25238 & n29434 ) ;
  assign n29432 = n16082 ^ n12518 ^ n3819 ;
  assign n29429 = n573 | n8205 ;
  assign n29430 = n29429 ^ n7201 ^ 1'b0 ;
  assign n29431 = ( n320 & ~n11395 ) | ( n320 & n29430 ) | ( ~n11395 & n29430 ) ;
  assign n29433 = n29432 ^ n29431 ^ n16103 ;
  assign n29436 = n29435 ^ n29433 ^ 1'b0 ;
  assign n29437 = n7931 ^ n957 ^ n669 ;
  assign n29440 = n9517 ^ n429 ^ 1'b0 ;
  assign n29441 = n8805 | n29440 ;
  assign n29438 = n26030 ^ n13049 ^ n6981 ;
  assign n29439 = n18651 & n29438 ;
  assign n29442 = n29441 ^ n29439 ^ n6682 ;
  assign n29443 = n29442 ^ n20476 ^ n5812 ;
  assign n29444 = n15334 ^ n11168 ^ n1016 ;
  assign n29445 = ~n4568 & n29444 ;
  assign n29446 = n19348 ^ n1810 ^ n1504 ;
  assign n29447 = ~n13075 & n29446 ;
  assign n29448 = n24817 | n29447 ;
  assign n29449 = n23398 & ~n24449 ;
  assign n29450 = n29449 ^ n18481 ^ 1'b0 ;
  assign n29451 = n29450 ^ n7964 ^ 1'b0 ;
  assign n29452 = n29094 ^ n2053 ^ 1'b0 ;
  assign n29453 = n9788 ^ n6381 ^ n2576 ;
  assign n29454 = n14283 ^ n7917 ^ 1'b0 ;
  assign n29455 = ( n9506 & ~n24767 ) | ( n9506 & n29454 ) | ( ~n24767 & n29454 ) ;
  assign n29456 = n16445 & n29455 ;
  assign n29457 = n28442 ^ n1940 ^ 1'b0 ;
  assign n29458 = n28039 | n29457 ;
  assign n29459 = n29457 & ~n29458 ;
  assign n29460 = n1966 ^ n1513 ^ 1'b0 ;
  assign n29461 = n23220 | n29460 ;
  assign n29462 = n6887 | n11873 ;
  assign n29463 = ( n1054 & n5441 ) | ( n1054 & n6325 ) | ( n5441 & n6325 ) ;
  assign n29464 = n29463 ^ n20792 ^ n9233 ;
  assign n29465 = ~n5448 & n6653 ;
  assign n29466 = ( n2639 & n10512 ) | ( n2639 & ~n20692 ) | ( n10512 & ~n20692 ) ;
  assign n29467 = n29466 ^ n2142 ^ 1'b0 ;
  assign n29468 = n21436 | n29276 ;
  assign n29469 = n26375 | n29468 ;
  assign n29470 = n29469 ^ n26603 ^ n16909 ;
  assign n29472 = n22323 ^ n18111 ^ 1'b0 ;
  assign n29471 = n9670 & ~n12795 ;
  assign n29473 = n29472 ^ n29471 ^ n2864 ;
  assign n29474 = ( ~n9449 & n12690 ) | ( ~n9449 & n28691 ) | ( n12690 & n28691 ) ;
  assign n29475 = x153 & n29474 ;
  assign n29476 = ( n2132 & n29473 ) | ( n2132 & n29475 ) | ( n29473 & n29475 ) ;
  assign n29477 = ~n13226 & n20599 ;
  assign n29478 = ~n20599 & n29477 ;
  assign n29479 = n2293 & n8304 ;
  assign n29480 = n29478 & n29479 ;
  assign n29481 = ( n9298 & n27608 ) | ( n9298 & ~n29480 ) | ( n27608 & ~n29480 ) ;
  assign n29482 = n5394 | n28848 ;
  assign n29483 = n12399 | n22747 ;
  assign n29484 = n23578 & ~n29483 ;
  assign n29485 = ~n3987 & n8514 ;
  assign n29486 = n16392 & n29485 ;
  assign n29487 = ( n6820 & ~n24948 ) | ( n6820 & n25607 ) | ( ~n24948 & n25607 ) ;
  assign n29488 = ( n8281 & ~n28345 ) | ( n8281 & n29487 ) | ( ~n28345 & n29487 ) ;
  assign n29489 = n4682 & n29488 ;
  assign n29490 = n29486 & n29489 ;
  assign n29491 = n3898 | n5354 ;
  assign n29493 = n8288 | n8594 ;
  assign n29492 = n2584 & n22089 ;
  assign n29494 = n29493 ^ n29492 ^ 1'b0 ;
  assign n29495 = ( ~n12321 & n29143 ) | ( ~n12321 & n29494 ) | ( n29143 & n29494 ) ;
  assign n29496 = n29495 ^ n23882 ^ n16543 ;
  assign n29497 = n8168 ^ n7362 ^ 1'b0 ;
  assign n29498 = n9144 ^ n7955 ^ n1020 ;
  assign n29499 = n24699 & ~n28231 ;
  assign n29500 = n13537 & n29499 ;
  assign n29501 = n502 | n29500 ;
  assign n29502 = ( n7126 & n14310 ) | ( n7126 & n22337 ) | ( n14310 & n22337 ) ;
  assign n29503 = n343 & n29502 ;
  assign n29504 = ~n20232 & n29503 ;
  assign n29505 = n13971 ^ n2962 ^ 1'b0 ;
  assign n29506 = ( n7611 & n13438 ) | ( n7611 & n14718 ) | ( n13438 & n14718 ) ;
  assign n29507 = n29505 & ~n29506 ;
  assign n29508 = n29507 ^ n14396 ^ n2359 ;
  assign n29509 = n12563 ^ n6493 ^ 1'b0 ;
  assign n29510 = n2988 & ~n29509 ;
  assign n29511 = ( n3600 & ~n17699 ) | ( n3600 & n29510 ) | ( ~n17699 & n29510 ) ;
  assign n29512 = n29511 ^ n16577 ^ 1'b0 ;
  assign n29513 = n2331 & ~n10113 ;
  assign n29514 = n1364 | n15560 ;
  assign n29515 = n988 | n29514 ;
  assign n29516 = n29515 ^ n6162 ^ 1'b0 ;
  assign n29517 = ~n22974 & n29516 ;
  assign n29523 = n18398 ^ n9161 ^ 1'b0 ;
  assign n29524 = n27181 & n29523 ;
  assign n29518 = n7238 & ~n22616 ;
  assign n29519 = n15632 & n22610 ;
  assign n29520 = n26319 & ~n29519 ;
  assign n29521 = n22849 | n29520 ;
  assign n29522 = n29518 | n29521 ;
  assign n29525 = n29524 ^ n29522 ^ n7573 ;
  assign n29529 = n29332 ^ n1653 ^ 1'b0 ;
  assign n29530 = n16800 | n29529 ;
  assign n29526 = n17297 ^ n12638 ^ 1'b0 ;
  assign n29527 = n12774 ^ n4000 ^ 1'b0 ;
  assign n29528 = n29526 & n29527 ;
  assign n29531 = n29530 ^ n29528 ^ 1'b0 ;
  assign n29532 = ~n737 & n27160 ;
  assign n29533 = n8696 & n10146 ;
  assign n29534 = n25088 & n29533 ;
  assign n29535 = n8732 & n11380 ;
  assign n29536 = ( n7045 & ~n15900 ) | ( n7045 & n20503 ) | ( ~n15900 & n20503 ) ;
  assign n29537 = n19467 & n29536 ;
  assign n29538 = ( ~n11686 & n26926 ) | ( ~n11686 & n29290 ) | ( n26926 & n29290 ) ;
  assign n29539 = ( n1352 & ~n5565 ) | ( n1352 & n22521 ) | ( ~n5565 & n22521 ) ;
  assign n29540 = n13556 & ~n29539 ;
  assign n29541 = n5511 | n27193 ;
  assign n29542 = n29541 ^ n22842 ^ 1'b0 ;
  assign n29543 = ~n9912 & n29542 ;
  assign n29548 = n5165 | n28498 ;
  assign n29544 = ( x237 & ~n2242 ) | ( x237 & n2777 ) | ( ~n2242 & n2777 ) ;
  assign n29545 = ~n16917 & n29544 ;
  assign n29546 = ~n3300 & n29545 ;
  assign n29547 = n2944 | n29546 ;
  assign n29549 = n29548 ^ n29547 ^ 1'b0 ;
  assign n29550 = n11607 | n29549 ;
  assign n29551 = n16847 | n29550 ;
  assign n29553 = n27989 ^ n26349 ^ n18281 ;
  assign n29554 = n29553 ^ n17840 ^ 1'b0 ;
  assign n29555 = n4521 & n29554 ;
  assign n29552 = n27927 ^ n27202 ^ n1570 ;
  assign n29556 = n29555 ^ n29552 ^ n24714 ;
  assign n29558 = ~n1768 & n4317 ;
  assign n29559 = n29558 ^ n3314 ^ 1'b0 ;
  assign n29557 = n27520 ^ n16158 ^ n9329 ;
  assign n29560 = n29559 ^ n29557 ^ n16795 ;
  assign n29563 = n13831 ^ n6844 ^ n4402 ;
  assign n29564 = n29563 ^ n17226 ^ n12263 ;
  assign n29561 = n11331 ^ n6596 ^ n1479 ;
  assign n29562 = n15155 & ~n29561 ;
  assign n29565 = n29564 ^ n29562 ^ n15959 ;
  assign n29566 = n6313 & n8644 ;
  assign n29567 = n29566 ^ n21004 ^ n3925 ;
  assign n29568 = n18670 ^ n11643 ^ n9078 ;
  assign n29569 = n5377 ^ n3331 ^ 1'b0 ;
  assign n29570 = ( n539 & n2909 ) | ( n539 & n29569 ) | ( n2909 & n29569 ) ;
  assign n29571 = n20872 & ~n29570 ;
  assign n29572 = n4819 ^ n2604 ^ 1'b0 ;
  assign n29573 = n29571 | n29572 ;
  assign n29574 = ~n13402 & n22845 ;
  assign n29575 = n8015 ^ n7518 ^ 1'b0 ;
  assign n29576 = n258 & n29575 ;
  assign n29577 = n29574 & n29576 ;
  assign n29578 = ~n1800 & n6826 ;
  assign n29579 = n29578 ^ n19078 ^ 1'b0 ;
  assign n29580 = n8130 ^ n3942 ^ 1'b0 ;
  assign n29581 = n2497 | n29580 ;
  assign n29582 = ~n2404 & n29581 ;
  assign n29583 = ~n14353 & n29582 ;
  assign n29584 = ~n19648 & n26077 ;
  assign n29585 = ( n23576 & n27210 ) | ( n23576 & n29584 ) | ( n27210 & n29584 ) ;
  assign n29586 = n1475 | n3548 ;
  assign n29587 = n13272 & ~n29586 ;
  assign n29588 = n29587 ^ n25912 ^ n2845 ;
  assign n29589 = n29061 ^ n18723 ^ 1'b0 ;
  assign n29590 = n27008 & ~n29589 ;
  assign n29591 = n2970 & ~n7994 ;
  assign n29592 = ~n8696 & n29591 ;
  assign n29593 = n29592 ^ n7316 ^ 1'b0 ;
  assign n29594 = n29593 ^ n21761 ^ n13082 ;
  assign n29595 = n9645 & ~n26195 ;
  assign n29596 = ~n29594 & n29595 ;
  assign n29597 = n10080 ^ n4822 ^ n4047 ;
  assign n29600 = n13052 ^ n9892 ^ n8480 ;
  assign n29598 = n17479 ^ n10743 ^ 1'b0 ;
  assign n29599 = n29598 ^ n1030 ^ 1'b0 ;
  assign n29601 = n29600 ^ n29599 ^ n25622 ;
  assign n29602 = n29081 ^ n7558 ^ 1'b0 ;
  assign n29603 = n29602 ^ n13290 ^ n5027 ;
  assign n29604 = n17347 ^ n12143 ^ n1084 ;
  assign n29605 = n14706 | n25616 ;
  assign n29606 = ( n25998 & n29604 ) | ( n25998 & n29605 ) | ( n29604 & n29605 ) ;
  assign n29608 = ( n2155 & n19038 ) | ( n2155 & n24698 ) | ( n19038 & n24698 ) ;
  assign n29607 = ~n2604 & n8308 ;
  assign n29609 = n29608 ^ n29607 ^ 1'b0 ;
  assign n29614 = n3803 & ~n5831 ;
  assign n29610 = n460 & n9200 ;
  assign n29611 = n22133 & n29610 ;
  assign n29612 = n29611 ^ n7214 ^ 1'b0 ;
  assign n29613 = n10668 & ~n29612 ;
  assign n29615 = n29614 ^ n29613 ^ n23138 ;
  assign n29616 = n14300 ^ n2458 ^ 1'b0 ;
  assign n29617 = ( ~n2110 & n11114 ) | ( ~n2110 & n29616 ) | ( n11114 & n29616 ) ;
  assign n29618 = ( n5325 & ~n17569 ) | ( n5325 & n29617 ) | ( ~n17569 & n29617 ) ;
  assign n29619 = n17038 & n29618 ;
  assign n29621 = n2954 & n10340 ;
  assign n29620 = ( n3064 & n7829 ) | ( n3064 & n18870 ) | ( n7829 & n18870 ) ;
  assign n29622 = n29621 ^ n29620 ^ n24426 ;
  assign n29623 = n8903 & n14191 ;
  assign n29624 = n13738 & n29623 ;
  assign n29625 = n8466 | n13722 ;
  assign n29626 = n29625 ^ n2401 ^ 1'b0 ;
  assign n29627 = n23750 ^ n20622 ^ n15601 ;
  assign n29629 = n18088 ^ n6074 ^ n704 ;
  assign n29628 = n20293 ^ n312 ^ 1'b0 ;
  assign n29630 = n29629 ^ n29628 ^ 1'b0 ;
  assign n29631 = ~n29627 & n29630 ;
  assign n29632 = ( n4942 & n14665 ) | ( n4942 & ~n20053 ) | ( n14665 & ~n20053 ) ;
  assign n29633 = n5125 | n29632 ;
  assign n29635 = ~n10383 & n17589 ;
  assign n29636 = n29635 ^ n19411 ^ 1'b0 ;
  assign n29634 = n21648 ^ n21148 ^ n2711 ;
  assign n29637 = n29636 ^ n29634 ^ n10950 ;
  assign n29638 = n8753 ^ n1239 ^ 1'b0 ;
  assign n29639 = ~n13107 & n29638 ;
  assign n29640 = n29639 ^ n29421 ^ 1'b0 ;
  assign n29641 = ( n11297 & n19101 ) | ( n11297 & n29640 ) | ( n19101 & n29640 ) ;
  assign n29642 = ( ~n4872 & n8361 ) | ( ~n4872 & n10579 ) | ( n8361 & n10579 ) ;
  assign n29643 = n20444 ^ n20062 ^ n9438 ;
  assign n29644 = n29643 ^ n6189 ^ 1'b0 ;
  assign n29645 = n29642 & n29644 ;
  assign n29646 = n5336 ^ n4662 ^ 1'b0 ;
  assign n29647 = ~n4984 & n29646 ;
  assign n29648 = ~n1681 & n29647 ;
  assign n29649 = n17670 & n29648 ;
  assign n29650 = n10229 ^ n6832 ^ n287 ;
  assign n29651 = n2380 & ~n29650 ;
  assign n29652 = n2017 | n7125 ;
  assign n29653 = n564 & ~n29652 ;
  assign n29654 = n12845 | n29653 ;
  assign n29655 = n29651 & ~n29654 ;
  assign n29656 = n29655 ^ n18382 ^ n2755 ;
  assign n29657 = n29649 | n29656 ;
  assign n29658 = n10807 | n29657 ;
  assign n29659 = n12742 | n13337 ;
  assign n29660 = n29659 ^ n4493 ^ 1'b0 ;
  assign n29661 = ( ~n4647 & n6177 ) | ( ~n4647 & n22208 ) | ( n6177 & n22208 ) ;
  assign n29662 = ~n15366 & n27335 ;
  assign n29663 = n29662 ^ n12621 ^ 1'b0 ;
  assign n29664 = ~n23871 & n29663 ;
  assign n29665 = n29664 ^ n20297 ^ 1'b0 ;
  assign n29666 = n3939 | n7019 ;
  assign n29667 = ( n9556 & n13472 ) | ( n9556 & n29666 ) | ( n13472 & n29666 ) ;
  assign n29668 = ~n1254 & n12628 ;
  assign n29669 = n29668 ^ n297 ^ 1'b0 ;
  assign n29680 = n13002 | n17790 ;
  assign n29674 = ~x5 & n1940 ;
  assign n29670 = n4360 & ~n8754 ;
  assign n29671 = ~n4710 & n29670 ;
  assign n29672 = ( n3804 & ~n18949 ) | ( n3804 & n29671 ) | ( ~n18949 & n29671 ) ;
  assign n29673 = n6202 & n29672 ;
  assign n29675 = n29674 ^ n29673 ^ 1'b0 ;
  assign n29676 = ( n2959 & ~n27877 ) | ( n2959 & n29675 ) | ( ~n27877 & n29675 ) ;
  assign n29677 = n15226 & n29676 ;
  assign n29678 = n2393 & n29677 ;
  assign n29679 = n10173 & ~n29678 ;
  assign n29681 = n29680 ^ n29679 ^ 1'b0 ;
  assign n29682 = ~n29669 & n29681 ;
  assign n29683 = n29682 ^ n25564 ^ 1'b0 ;
  assign n29684 = n26493 ^ n20130 ^ n7704 ;
  assign n29685 = ( n5737 & ~n21502 ) | ( n5737 & n27706 ) | ( ~n21502 & n27706 ) ;
  assign n29687 = x249 & n19638 ;
  assign n29688 = n29687 ^ n2004 ^ 1'b0 ;
  assign n29686 = n17541 & n25789 ;
  assign n29689 = n29688 ^ n29686 ^ x95 ;
  assign n29690 = n7902 ^ n3264 ^ x126 ;
  assign n29691 = n29690 ^ n394 ^ 1'b0 ;
  assign n29692 = n29691 ^ n13059 ^ 1'b0 ;
  assign n29693 = ~n23212 & n29692 ;
  assign n29694 = n12098 ^ n8091 ^ 1'b0 ;
  assign n29695 = n20720 & ~n29694 ;
  assign n29696 = n18335 ^ n13581 ^ 1'b0 ;
  assign n29697 = n18293 & n29696 ;
  assign n29699 = n3049 & ~n6268 ;
  assign n29700 = ( n2145 & ~n11417 ) | ( n2145 & n29699 ) | ( ~n11417 & n29699 ) ;
  assign n29701 = n29700 ^ n28966 ^ n5989 ;
  assign n29698 = n3280 | n18082 ;
  assign n29702 = n29701 ^ n29698 ^ 1'b0 ;
  assign n29703 = n11775 ^ n4201 ^ 1'b0 ;
  assign n29704 = ~n3208 & n29703 ;
  assign n29705 = n29704 ^ n19464 ^ n10836 ;
  assign n29706 = n22583 ^ n2611 ^ n1846 ;
  assign n29707 = n640 ^ x41 ^ 1'b0 ;
  assign n29708 = n4782 & ~n29707 ;
  assign n29709 = ( n2215 & ~n4582 ) | ( n2215 & n29708 ) | ( ~n4582 & n29708 ) ;
  assign n29710 = ( n10518 & ~n12202 ) | ( n10518 & n29709 ) | ( ~n12202 & n29709 ) ;
  assign n29711 = ( n3439 & n21837 ) | ( n3439 & n29710 ) | ( n21837 & n29710 ) ;
  assign n29712 = ~n6146 & n29711 ;
  assign n29713 = n29712 ^ x244 ^ 1'b0 ;
  assign n29714 = n13969 ^ n8376 ^ n1922 ;
  assign n29715 = n8591 ^ n5500 ^ 1'b0 ;
  assign n29716 = ~n29714 & n29715 ;
  assign n29717 = n26367 ^ n25294 ^ 1'b0 ;
  assign n29718 = n15985 & n22028 ;
  assign n29719 = n20168 & n29718 ;
  assign n29720 = ( n1366 & n4809 ) | ( n1366 & n19915 ) | ( n4809 & n19915 ) ;
  assign n29721 = n29719 & n29720 ;
  assign n29722 = ~n10191 & n15193 ;
  assign n29723 = n29722 ^ n28408 ^ 1'b0 ;
  assign n29724 = n7844 & ~n11893 ;
  assign n29725 = ( ~n1155 & n17220 ) | ( ~n1155 & n27459 ) | ( n17220 & n27459 ) ;
  assign n29726 = x138 & n29725 ;
  assign n29727 = ( ~n8736 & n11288 ) | ( ~n8736 & n12468 ) | ( n11288 & n12468 ) ;
  assign n29728 = ~n2535 & n29727 ;
  assign n29729 = n29728 ^ n24872 ^ 1'b0 ;
  assign n29730 = ( ~n12427 & n18090 ) | ( ~n12427 & n29729 ) | ( n18090 & n29729 ) ;
  assign n29731 = ( ~n8546 & n9195 ) | ( ~n8546 & n27379 ) | ( n9195 & n27379 ) ;
  assign n29732 = n26328 ^ n17880 ^ n5957 ;
  assign n29733 = n705 & n27169 ;
  assign n29734 = ( n24378 & ~n28819 ) | ( n24378 & n29733 ) | ( ~n28819 & n29733 ) ;
  assign n29735 = ~n13025 & n17370 ;
  assign n29736 = n10083 & n29735 ;
  assign n29737 = n28344 ^ n14692 ^ 1'b0 ;
  assign n29738 = n15445 | n29737 ;
  assign n29747 = n25770 | n26913 ;
  assign n29746 = n3460 & n13438 ;
  assign n29740 = n4137 ^ n3410 ^ n2567 ;
  assign n29739 = n3159 | n8700 ;
  assign n29741 = n29740 ^ n29739 ^ 1'b0 ;
  assign n29742 = n26275 & ~n29741 ;
  assign n29743 = n29742 ^ n4410 ^ 1'b0 ;
  assign n29744 = ~n541 & n18684 ;
  assign n29745 = ~n29743 & n29744 ;
  assign n29748 = n29747 ^ n29746 ^ n29745 ;
  assign n29749 = ~n10967 & n21412 ;
  assign n29750 = n15728 & ~n26637 ;
  assign n29751 = n29750 ^ n19036 ^ 1'b0 ;
  assign n29752 = n29751 ^ n24941 ^ n20553 ;
  assign n29753 = ( n7506 & ~n20683 ) | ( n7506 & n29752 ) | ( ~n20683 & n29752 ) ;
  assign n29754 = ~n11643 & n11984 ;
  assign n29755 = ~n5645 & n12628 ;
  assign n29756 = n24139 & n29755 ;
  assign n29757 = n16185 ^ n7037 ^ 1'b0 ;
  assign n29758 = ( n26642 & ~n27002 ) | ( n26642 & n29757 ) | ( ~n27002 & n29757 ) ;
  assign n29759 = n7454 ^ n3157 ^ 1'b0 ;
  assign n29760 = n29758 | n29759 ;
  assign n29761 = n5180 ^ n3620 ^ n2185 ;
  assign n29762 = ~n1502 & n29761 ;
  assign n29763 = n8376 & n29762 ;
  assign n29764 = n14693 | n29763 ;
  assign n29765 = n29764 ^ n5293 ^ 1'b0 ;
  assign n29766 = ( n18502 & n19086 ) | ( n18502 & n29765 ) | ( n19086 & n29765 ) ;
  assign n29767 = n27259 ^ n1023 ^ 1'b0 ;
  assign n29768 = ( n7736 & ~n10505 ) | ( n7736 & n29767 ) | ( ~n10505 & n29767 ) ;
  assign n29769 = ( n2419 & n2764 ) | ( n2419 & n23488 ) | ( n2764 & n23488 ) ;
  assign n29770 = n29769 ^ n6141 ^ 1'b0 ;
  assign n29771 = ~n25298 & n29770 ;
  assign n29772 = ~n16359 & n29771 ;
  assign n29773 = n29772 ^ n17457 ^ 1'b0 ;
  assign n29774 = ( n4596 & n7291 ) | ( n4596 & ~n14798 ) | ( n7291 & ~n14798 ) ;
  assign n29775 = ( n1351 & n4883 ) | ( n1351 & ~n29774 ) | ( n4883 & ~n29774 ) ;
  assign n29776 = n2489 & ~n14465 ;
  assign n29777 = n29776 ^ n21408 ^ 1'b0 ;
  assign n29778 = n29775 & ~n29777 ;
  assign n29779 = n27420 ^ n16011 ^ n4465 ;
  assign n29780 = ( n7076 & n7157 ) | ( n7076 & n25397 ) | ( n7157 & n25397 ) ;
  assign n29781 = n21408 ^ n18584 ^ n9744 ;
  assign n29782 = n29781 ^ n14312 ^ 1'b0 ;
  assign n29783 = x186 & n29782 ;
  assign n29784 = n17319 & ~n23361 ;
  assign n29785 = ~n29783 & n29784 ;
  assign n29786 = n11593 ^ n5715 ^ 1'b0 ;
  assign n29787 = ~n5816 & n29786 ;
  assign n29788 = n29787 ^ n8158 ^ 1'b0 ;
  assign n29789 = n27784 ^ n27375 ^ n24985 ;
  assign n29790 = n22711 ^ n15408 ^ n8375 ;
  assign n29791 = n5955 & n29790 ;
  assign n29792 = n27991 & n29791 ;
  assign n29793 = n29792 ^ n20588 ^ 1'b0 ;
  assign n29794 = ( n1064 & n4145 ) | ( n1064 & ~n9713 ) | ( n4145 & ~n9713 ) ;
  assign n29795 = n29794 ^ n26217 ^ n23220 ;
  assign n29796 = ( n10724 & ~n17940 ) | ( n10724 & n22791 ) | ( ~n17940 & n22791 ) ;
  assign n29797 = n29796 ^ n18920 ^ 1'b0 ;
  assign n29798 = ~n18584 & n29797 ;
  assign n29799 = n3621 | n7799 ;
  assign n29800 = n29799 ^ n27835 ^ n9312 ;
  assign n29801 = ~n15461 & n29800 ;
  assign n29802 = n10116 | n20535 ;
  assign n29803 = n29802 ^ n7810 ^ 1'b0 ;
  assign n29804 = ( n4984 & n24854 ) | ( n4984 & n29803 ) | ( n24854 & n29803 ) ;
  assign n29805 = n12914 & n27814 ;
  assign n29806 = n29804 & n29805 ;
  assign n29808 = n22875 ^ n15264 ^ n1281 ;
  assign n29807 = n11729 ^ n3201 ^ 1'b0 ;
  assign n29809 = n29808 ^ n29807 ^ 1'b0 ;
  assign n29810 = ( n11893 & n14804 ) | ( n11893 & n29809 ) | ( n14804 & n29809 ) ;
  assign n29811 = n24388 ^ n3301 ^ 1'b0 ;
  assign n29812 = ~n2874 & n29811 ;
  assign n29813 = ( ~n7279 & n9820 ) | ( ~n7279 & n13181 ) | ( n9820 & n13181 ) ;
  assign n29814 = n29813 ^ n20948 ^ n11582 ;
  assign n29815 = n29814 ^ n8827 ^ 1'b0 ;
  assign n29816 = ~n1532 & n29815 ;
  assign n29817 = ( n3725 & n8062 ) | ( n3725 & n17202 ) | ( n8062 & n17202 ) ;
  assign n29818 = ( n29812 & ~n29816 ) | ( n29812 & n29817 ) | ( ~n29816 & n29817 ) ;
  assign n29821 = ~n9905 & n22768 ;
  assign n29822 = n29821 ^ x152 ^ 1'b0 ;
  assign n29819 = n20069 ^ n10267 ^ n9103 ;
  assign n29820 = n29819 ^ n4309 ^ x6 ;
  assign n29823 = n29822 ^ n29820 ^ n24170 ;
  assign n29824 = ~n21119 & n29823 ;
  assign n29826 = n540 & n3140 ;
  assign n29827 = n3718 & n29826 ;
  assign n29825 = n21892 & ~n27522 ;
  assign n29828 = n29827 ^ n29825 ^ 1'b0 ;
  assign n29829 = n18822 ^ n5832 ^ 1'b0 ;
  assign n29830 = n969 & n29829 ;
  assign n29831 = n29830 ^ n22485 ^ 1'b0 ;
  assign n29832 = n14085 ^ n10570 ^ 1'b0 ;
  assign n29833 = n7417 & ~n16764 ;
  assign n29834 = n29833 ^ n5330 ^ 1'b0 ;
  assign n29835 = n4407 ^ x229 ^ 1'b0 ;
  assign n29836 = n29834 | n29835 ;
  assign n29837 = n7473 | n18300 ;
  assign n29838 = n5223 ^ n2549 ^ 1'b0 ;
  assign n29839 = n3106 & ~n29838 ;
  assign n29840 = n29839 ^ n28453 ^ n21335 ;
  assign n29841 = n7350 & n18788 ;
  assign n29842 = n6314 & n6539 ;
  assign n29843 = ~n22688 & n29842 ;
  assign n29844 = n9381 ^ n1047 ^ 1'b0 ;
  assign n29845 = n28777 & n29844 ;
  assign n29846 = n29845 ^ n24338 ^ 1'b0 ;
  assign n29847 = n29846 ^ n4405 ^ 1'b0 ;
  assign n29848 = n29843 & ~n29847 ;
  assign n29849 = n29841 & n29848 ;
  assign n29850 = n11760 | n24442 ;
  assign n29851 = ( x192 & n15216 ) | ( x192 & ~n29850 ) | ( n15216 & ~n29850 ) ;
  assign n29852 = ( n1102 & n2463 ) | ( n1102 & n4575 ) | ( n2463 & n4575 ) ;
  assign n29853 = ( ~n788 & n7037 ) | ( ~n788 & n29852 ) | ( n7037 & n29852 ) ;
  assign n29854 = n8801 & n9227 ;
  assign n29855 = n5710 & ~n7065 ;
  assign n29856 = ( ~n2632 & n29854 ) | ( ~n2632 & n29855 ) | ( n29854 & n29855 ) ;
  assign n29857 = ~n17377 & n29856 ;
  assign n29858 = ( n4869 & n5615 ) | ( n4869 & ~n7955 ) | ( n5615 & ~n7955 ) ;
  assign n29859 = n8545 & ~n18791 ;
  assign n29860 = n29858 & ~n29859 ;
  assign n29865 = n9520 | n23104 ;
  assign n29866 = ( n5809 & n7605 ) | ( n5809 & n29865 ) | ( n7605 & n29865 ) ;
  assign n29862 = n4274 ^ n2529 ^ n1515 ;
  assign n29863 = n17237 | n29862 ;
  assign n29861 = n14189 ^ n13634 ^ n8756 ;
  assign n29864 = n29863 ^ n29861 ^ n6413 ;
  assign n29867 = n29866 ^ n29864 ^ n815 ;
  assign n29868 = n22012 ^ n8478 ^ n8205 ;
  assign n29869 = n6279 & n14431 ;
  assign n29870 = ~n19849 & n29869 ;
  assign n29871 = ~n3892 & n6431 ;
  assign n29872 = n11419 ^ n10692 ^ 1'b0 ;
  assign n29873 = n5730 & ~n29872 ;
  assign n29874 = ~n29871 & n29873 ;
  assign n29875 = ( n518 & ~n29870 ) | ( n518 & n29874 ) | ( ~n29870 & n29874 ) ;
  assign n29876 = n11915 ^ n3066 ^ 1'b0 ;
  assign n29877 = n27404 & ~n29876 ;
  assign n29878 = n12089 & n29877 ;
  assign n29879 = n29878 ^ n9460 ^ 1'b0 ;
  assign n29880 = n11546 ^ n4146 ^ 1'b0 ;
  assign n29881 = n15109 ^ n736 ^ 1'b0 ;
  assign n29882 = ( n29879 & n29880 ) | ( n29879 & n29881 ) | ( n29880 & n29881 ) ;
  assign n29886 = n4680 ^ n3728 ^ 1'b0 ;
  assign n29883 = ~n4374 & n13736 ;
  assign n29884 = ~n5404 & n15835 ;
  assign n29885 = n29883 & ~n29884 ;
  assign n29887 = n29886 ^ n29885 ^ 1'b0 ;
  assign n29888 = ( n5225 & n12668 ) | ( n5225 & ~n20732 ) | ( n12668 & ~n20732 ) ;
  assign n29889 = n15015 ^ n4687 ^ n3937 ;
  assign n29890 = n5740 ^ n508 ^ 1'b0 ;
  assign n29891 = n6903 & n29890 ;
  assign n29892 = n2682 ^ n1315 ^ 1'b0 ;
  assign n29893 = ( n20761 & n29891 ) | ( n20761 & n29892 ) | ( n29891 & n29892 ) ;
  assign n29894 = ( n15892 & n22694 ) | ( n15892 & ~n29893 ) | ( n22694 & ~n29893 ) ;
  assign n29895 = ( n1555 & ~n23320 ) | ( n1555 & n29894 ) | ( ~n23320 & n29894 ) ;
  assign n29900 = n25528 ^ n14322 ^ 1'b0 ;
  assign n29896 = ( ~n9457 & n11630 ) | ( ~n9457 & n20772 ) | ( n11630 & n20772 ) ;
  assign n29897 = n29896 ^ n13717 ^ n9747 ;
  assign n29898 = ( n7486 & ~n8880 ) | ( n7486 & n16886 ) | ( ~n8880 & n16886 ) ;
  assign n29899 = ( n8299 & ~n29897 ) | ( n8299 & n29898 ) | ( ~n29897 & n29898 ) ;
  assign n29901 = n29900 ^ n29899 ^ n5232 ;
  assign n29902 = n9513 ^ n644 ^ 1'b0 ;
  assign n29903 = n4782 | n29902 ;
  assign n29904 = n10990 | n29903 ;
  assign n29905 = ( n3110 & ~n18358 ) | ( n3110 & n29904 ) | ( ~n18358 & n29904 ) ;
  assign n29906 = n24606 | n26543 ;
  assign n29907 = n29906 ^ n7136 ^ 1'b0 ;
  assign n29908 = n17140 ^ n16546 ^ n7576 ;
  assign n29909 = x152 & n3178 ;
  assign n29910 = n29908 & n29909 ;
  assign n29911 = n28078 ^ n8539 ^ 1'b0 ;
  assign n29913 = ~n3138 & n14183 ;
  assign n29912 = ( n5831 & n20100 ) | ( n5831 & n22108 ) | ( n20100 & n22108 ) ;
  assign n29914 = n29913 ^ n29912 ^ n4157 ;
  assign n29915 = ( n9693 & n16652 ) | ( n9693 & ~n29914 ) | ( n16652 & ~n29914 ) ;
  assign n29916 = ~n7198 & n17556 ;
  assign n29917 = ( n20035 & n24556 ) | ( n20035 & n29916 ) | ( n24556 & n29916 ) ;
  assign n29918 = n25494 ^ n17520 ^ n967 ;
  assign n29919 = n24225 ^ n19295 ^ 1'b0 ;
  assign n29920 = n2970 & n29919 ;
  assign n29921 = ( n257 & ~n1197 ) | ( n257 & n29920 ) | ( ~n1197 & n29920 ) ;
  assign n29922 = n29921 ^ n10192 ^ n6750 ;
  assign n29923 = n29922 ^ n26605 ^ 1'b0 ;
  assign n29924 = ~n5514 & n29923 ;
  assign n29925 = ~n16888 & n29924 ;
  assign n29926 = n21432 ^ n13934 ^ 1'b0 ;
  assign n29927 = n5281 & ~n9895 ;
  assign n29928 = n14642 ^ n14380 ^ n10935 ;
  assign n29929 = ~n21341 & n29928 ;
  assign n29930 = n7680 ^ n2991 ^ x117 ;
  assign n29931 = n29930 ^ n29270 ^ n13455 ;
  assign n29932 = ( ~n10778 & n22428 ) | ( ~n10778 & n29931 ) | ( n22428 & n29931 ) ;
  assign n29933 = ( n2664 & n15588 ) | ( n2664 & n29932 ) | ( n15588 & n29932 ) ;
  assign n29934 = n16541 | n21713 ;
  assign n29935 = n5778 | n14185 ;
  assign n29936 = n18709 & n29935 ;
  assign n29937 = ( ~n12884 & n18521 ) | ( ~n12884 & n29936 ) | ( n18521 & n29936 ) ;
  assign n29938 = n26535 ^ n13531 ^ n8676 ;
  assign n29939 = n27081 ^ n5188 ^ n1466 ;
  assign n29940 = n22725 ^ n2476 ^ 1'b0 ;
  assign n29941 = n21824 ^ n6863 ^ 1'b0 ;
  assign n29942 = n11243 | n29941 ;
  assign n29943 = n26812 ^ n1784 ^ 1'b0 ;
  assign n29944 = n25838 & ~n29943 ;
  assign n29945 = ( n27055 & ~n29942 ) | ( n27055 & n29944 ) | ( ~n29942 & n29944 ) ;
  assign n29946 = n9310 ^ n5663 ^ 1'b0 ;
  assign n29947 = n27562 & n28526 ;
  assign n29948 = n4339 & n29947 ;
  assign n29949 = ( n24942 & n29946 ) | ( n24942 & ~n29948 ) | ( n29946 & ~n29948 ) ;
  assign n29950 = ~n12757 & n14492 ;
  assign n29956 = ( n1643 & ~n1708 ) | ( n1643 & n15769 ) | ( ~n1708 & n15769 ) ;
  assign n29955 = n16553 & ~n20039 ;
  assign n29952 = n9469 | n18487 ;
  assign n29953 = n490 & ~n29952 ;
  assign n29951 = n8583 ^ n7544 ^ 1'b0 ;
  assign n29954 = n29953 ^ n29951 ^ n17274 ;
  assign n29957 = n29956 ^ n29955 ^ n29954 ;
  assign n29958 = ~n5119 & n29957 ;
  assign n29959 = n17219 & n29958 ;
  assign n29960 = n8942 ^ n8333 ^ n4208 ;
  assign n29961 = n6662 ^ n2803 ^ 1'b0 ;
  assign n29962 = n29960 | n29961 ;
  assign n29969 = n24520 ^ n2090 ^ 1'b0 ;
  assign n29970 = n10544 & ~n29969 ;
  assign n29965 = n7896 ^ n7040 ^ n5082 ;
  assign n29966 = n29965 ^ n8931 ^ n3810 ;
  assign n29967 = n721 & n29966 ;
  assign n29968 = n29967 ^ n1968 ^ 1'b0 ;
  assign n29963 = n28289 ^ n5757 ^ 1'b0 ;
  assign n29964 = ( n11392 & ~n19095 ) | ( n11392 & n29963 ) | ( ~n19095 & n29963 ) ;
  assign n29971 = n29970 ^ n29968 ^ n29964 ;
  assign n29972 = n27590 ^ n8243 ^ n4077 ;
  assign n29973 = n29972 ^ n15465 ^ 1'b0 ;
  assign n29974 = n1948 ^ n488 ^ 1'b0 ;
  assign n29975 = ( n521 & n4284 ) | ( n521 & ~n29974 ) | ( n4284 & ~n29974 ) ;
  assign n29976 = n26492 ^ n6374 ^ n2343 ;
  assign n29977 = n5587 ^ n1952 ^ 1'b0 ;
  assign n29978 = ~n29976 & n29977 ;
  assign n29979 = n20864 & n28441 ;
  assign n29980 = n14669 ^ n2127 ^ n1076 ;
  assign n29981 = n17795 | n29980 ;
  assign n29982 = n29524 ^ n14906 ^ n4012 ;
  assign n29983 = n7253 ^ n3586 ^ 1'b0 ;
  assign n29984 = ( ~n8627 & n20931 ) | ( ~n8627 & n29983 ) | ( n20931 & n29983 ) ;
  assign n29986 = n4493 & ~n8736 ;
  assign n29987 = n29986 ^ n3728 ^ 1'b0 ;
  assign n29988 = ~n14721 & n29987 ;
  assign n29989 = n15946 & n29988 ;
  assign n29985 = n705 & ~n2651 ;
  assign n29990 = n29989 ^ n29985 ^ 1'b0 ;
  assign n29991 = n5278 & n29990 ;
  assign n29992 = n29991 ^ n7824 ^ 1'b0 ;
  assign n29993 = n1431 & n8561 ;
  assign n29994 = n18737 ^ n5974 ^ n1476 ;
  assign n29995 = ( n5082 & n11966 ) | ( n5082 & n19753 ) | ( n11966 & n19753 ) ;
  assign n29996 = n14300 ^ n5883 ^ n3103 ;
  assign n29997 = n29996 ^ n25359 ^ n9648 ;
  assign n29998 = ( n24397 & ~n29995 ) | ( n24397 & n29997 ) | ( ~n29995 & n29997 ) ;
  assign n29999 = n2866 | n4741 ;
  assign n30000 = n7511 & ~n29999 ;
  assign n30001 = n5863 ^ n1985 ^ n271 ;
  assign n30002 = n30001 ^ n19346 ^ 1'b0 ;
  assign n30003 = n2063 & n8512 ;
  assign n30004 = ( n2014 & n4910 ) | ( n2014 & n27075 ) | ( n4910 & n27075 ) ;
  assign n30005 = n30004 ^ n4753 ^ 1'b0 ;
  assign n30007 = n27224 ^ n21521 ^ n12454 ;
  assign n30006 = n2882 & n8828 ;
  assign n30008 = n30007 ^ n30006 ^ 1'b0 ;
  assign n30009 = ( n30003 & ~n30005 ) | ( n30003 & n30008 ) | ( ~n30005 & n30008 ) ;
  assign n30010 = ( n2851 & n10289 ) | ( n2851 & ~n13867 ) | ( n10289 & ~n13867 ) ;
  assign n30011 = n30010 ^ n4313 ^ 1'b0 ;
  assign n30012 = n7500 & n30011 ;
  assign n30013 = ~n15203 & n22010 ;
  assign n30014 = n14906 ^ n5812 ^ 1'b0 ;
  assign n30015 = ( n8964 & n10153 ) | ( n8964 & ~n30014 ) | ( n10153 & ~n30014 ) ;
  assign n30018 = n13107 ^ n1235 ^ 1'b0 ;
  assign n30019 = n23388 | n30018 ;
  assign n30020 = n12581 | n30019 ;
  assign n30021 = n30020 ^ n17510 ^ 1'b0 ;
  assign n30016 = ~n11555 & n17797 ;
  assign n30017 = n30016 ^ n1905 ^ 1'b0 ;
  assign n30022 = n30021 ^ n30017 ^ n11637 ;
  assign n30023 = ( n16644 & n30015 ) | ( n16644 & n30022 ) | ( n30015 & n30022 ) ;
  assign n30024 = n18566 & ~n25496 ;
  assign n30025 = ~n18280 & n30024 ;
  assign n30026 = n5027 & n30025 ;
  assign n30027 = n30026 ^ n6753 ^ n4451 ;
  assign n30028 = n8743 & n12080 ;
  assign n30029 = n10081 & n30028 ;
  assign n30030 = n358 | n22156 ;
  assign n30031 = n9043 | n30030 ;
  assign n30032 = n6022 | n30031 ;
  assign n30033 = n6443 & n30032 ;
  assign n30034 = ( ~n2506 & n26786 ) | ( ~n2506 & n30033 ) | ( n26786 & n30033 ) ;
  assign n30035 = n30029 | n30034 ;
  assign n30036 = n9505 & ~n28691 ;
  assign n30037 = n12098 | n12874 ;
  assign n30038 = n30036 & ~n30037 ;
  assign n30039 = n5271 ^ n4666 ^ 1'b0 ;
  assign n30040 = ( n8894 & ~n9486 ) | ( n8894 & n30039 ) | ( ~n9486 & n30039 ) ;
  assign n30041 = n10492 | n30040 ;
  assign n30042 = n30041 ^ n14856 ^ 1'b0 ;
  assign n30043 = n4325 ^ n3909 ^ 1'b0 ;
  assign n30044 = n4130 & n30043 ;
  assign n30045 = n2791 & n30044 ;
  assign n30046 = n30045 ^ n10856 ^ n8983 ;
  assign n30047 = n1614 | n6439 ;
  assign n30048 = n25315 & ~n30047 ;
  assign n30049 = n30048 ^ n21562 ^ 1'b0 ;
  assign n30050 = n2440 & ~n12561 ;
  assign n30052 = n5641 & ~n9344 ;
  assign n30053 = n30052 ^ n23072 ^ 1'b0 ;
  assign n30051 = n13152 & ~n29696 ;
  assign n30054 = n30053 ^ n30051 ^ n4373 ;
  assign n30055 = ( ~n4204 & n8772 ) | ( ~n4204 & n11467 ) | ( n8772 & n11467 ) ;
  assign n30056 = ( n7920 & ~n8294 ) | ( n7920 & n30055 ) | ( ~n8294 & n30055 ) ;
  assign n30057 = n10763 ^ n7305 ^ 1'b0 ;
  assign n30058 = n30057 ^ n4786 ^ 1'b0 ;
  assign n30059 = ~n4137 & n30058 ;
  assign n30060 = n24573 ^ n21830 ^ 1'b0 ;
  assign n30061 = n30059 & n30060 ;
  assign n30062 = n17278 & n21943 ;
  assign n30063 = ~n14571 & n30062 ;
  assign n30064 = n10429 & n26843 ;
  assign n30065 = n30064 ^ n8447 ^ 1'b0 ;
  assign n30066 = ( n5543 & ~n7404 ) | ( n5543 & n28103 ) | ( ~n7404 & n28103 ) ;
  assign n30067 = ( x234 & n7478 ) | ( x234 & n20302 ) | ( n7478 & n20302 ) ;
  assign n30068 = n30067 ^ n1851 ^ 1'b0 ;
  assign n30069 = n18126 | n30068 ;
  assign n30070 = n22957 ^ n8835 ^ 1'b0 ;
  assign n30071 = n11362 & ~n30070 ;
  assign n30072 = ( n8577 & ~n18169 ) | ( n8577 & n25331 ) | ( ~n18169 & n25331 ) ;
  assign n30073 = n8943 | n30072 ;
  assign n30074 = ~n5899 & n26254 ;
  assign n30075 = ~n4247 & n30074 ;
  assign n30076 = n8320 ^ n3415 ^ 1'b0 ;
  assign n30077 = ( n2260 & n4981 ) | ( n2260 & ~n30076 ) | ( n4981 & ~n30076 ) ;
  assign n30078 = x203 & n10492 ;
  assign n30079 = n12813 | n30078 ;
  assign n30080 = ( n1526 & n30077 ) | ( n1526 & ~n30079 ) | ( n30077 & ~n30079 ) ;
  assign n30081 = ~n6227 & n19725 ;
  assign n30082 = n8030 ^ n3172 ^ n2962 ;
  assign n30083 = n30082 ^ n19114 ^ n2881 ;
  assign n30084 = n21299 ^ n13147 ^ 1'b0 ;
  assign n30085 = n2280 ^ n678 ^ 1'b0 ;
  assign n30086 = n14544 & ~n30085 ;
  assign n30087 = n4880 | n11685 ;
  assign n30088 = n26645 ^ n17671 ^ n2779 ;
  assign n30089 = n30088 ^ n4591 ^ 1'b0 ;
  assign n30090 = ~n30087 & n30089 ;
  assign n30091 = ( n1359 & n10804 ) | ( n1359 & n17724 ) | ( n10804 & n17724 ) ;
  assign n30092 = n30091 ^ n6544 ^ 1'b0 ;
  assign n30093 = ( ~n11730 & n12778 ) | ( ~n11730 & n30092 ) | ( n12778 & n30092 ) ;
  assign n30094 = n30093 ^ n12509 ^ n11407 ;
  assign n30095 = ( ~n9238 & n16163 ) | ( ~n9238 & n30094 ) | ( n16163 & n30094 ) ;
  assign n30096 = n23678 ^ n16738 ^ n12138 ;
  assign n30097 = ~n2246 & n19409 ;
  assign n30098 = n30096 & n30097 ;
  assign n30099 = n30098 ^ n13581 ^ n3406 ;
  assign n30100 = n14844 & n16724 ;
  assign n30101 = n26131 ^ n15931 ^ n11056 ;
  assign n30102 = n27405 & ~n30101 ;
  assign n30103 = ~n5519 & n30102 ;
  assign n30104 = n30103 ^ n19201 ^ 1'b0 ;
  assign n30105 = ( n4646 & n11288 ) | ( n4646 & n16176 ) | ( n11288 & n16176 ) ;
  assign n30106 = n30105 ^ n7446 ^ 1'b0 ;
  assign n30107 = n30106 ^ n15973 ^ n2485 ;
  assign n30108 = n30107 ^ n28189 ^ x156 ;
  assign n30109 = n10916 ^ n6219 ^ n362 ;
  assign n30110 = n965 | n30109 ;
  assign n30111 = n27733 ^ n18179 ^ n6148 ;
  assign n30112 = ( n6501 & n8546 ) | ( n6501 & ~n30111 ) | ( n8546 & ~n30111 ) ;
  assign n30113 = ( n2970 & n16555 ) | ( n2970 & ~n30112 ) | ( n16555 & ~n30112 ) ;
  assign n30114 = ~n9080 & n14410 ;
  assign n30115 = n1693 & n30114 ;
  assign n30116 = n15545 ^ n14677 ^ n3579 ;
  assign n30117 = n30116 ^ n7266 ^ 1'b0 ;
  assign n30118 = n8548 | n30117 ;
  assign n30119 = n27122 & ~n30118 ;
  assign n30120 = n24283 ^ n22368 ^ 1'b0 ;
  assign n30121 = n30120 ^ n9130 ^ 1'b0 ;
  assign n30122 = ( n11738 & ~n27239 ) | ( n11738 & n30121 ) | ( ~n27239 & n30121 ) ;
  assign n30123 = n4664 & n12938 ;
  assign n30124 = ( ~n7595 & n24378 ) | ( ~n7595 & n30123 ) | ( n24378 & n30123 ) ;
  assign n30125 = ~n20778 & n30124 ;
  assign n30126 = n1184 & ~n27092 ;
  assign n30127 = n30126 ^ n12205 ^ n1941 ;
  assign n30128 = n12066 & ~n12680 ;
  assign n30129 = n11388 ^ n6990 ^ 1'b0 ;
  assign n30130 = n15526 | n30129 ;
  assign n30131 = ( ~n14131 & n30128 ) | ( ~n14131 & n30130 ) | ( n30128 & n30130 ) ;
  assign n30132 = n30131 ^ n28037 ^ 1'b0 ;
  assign n30133 = ( n2176 & ~n9290 ) | ( n2176 & n22360 ) | ( ~n9290 & n22360 ) ;
  assign n30134 = ( n5899 & n19706 ) | ( n5899 & ~n30133 ) | ( n19706 & ~n30133 ) ;
  assign n30135 = ( n10265 & ~n21473 ) | ( n10265 & n30134 ) | ( ~n21473 & n30134 ) ;
  assign n30136 = n14511 ^ n3526 ^ 1'b0 ;
  assign n30137 = n394 & n30136 ;
  assign n30138 = n30137 ^ n29213 ^ n11290 ;
  assign n30139 = n3010 & n3546 ;
  assign n30140 = ( n1463 & n22381 ) | ( n1463 & ~n30139 ) | ( n22381 & ~n30139 ) ;
  assign n30141 = n24413 ^ n9566 ^ 1'b0 ;
  assign n30142 = n2352 & ~n30141 ;
  assign n30143 = n11257 & ~n17110 ;
  assign n30144 = ~n30142 & n30143 ;
  assign n30145 = ~n8270 & n21149 ;
  assign n30146 = ~n8004 & n30145 ;
  assign n30147 = n2904 & ~n23528 ;
  assign n30148 = n258 & n10272 ;
  assign n30149 = n30148 ^ n19238 ^ n4024 ;
  assign n30150 = ~n30147 & n30149 ;
  assign n30151 = n30146 & n30150 ;
  assign n30152 = n18143 ^ n4837 ^ 1'b0 ;
  assign n30153 = n12640 & n30152 ;
  assign n30154 = n753 & ~n903 ;
  assign n30155 = ~n30153 & n30154 ;
  assign n30156 = ( n24507 & n25700 ) | ( n24507 & n30155 ) | ( n25700 & n30155 ) ;
  assign n30157 = n26848 & n30046 ;
  assign n30158 = n18473 ^ n8920 ^ n7743 ;
  assign n30159 = n505 & n30158 ;
  assign n30160 = ~n18504 & n30159 ;
  assign n30161 = n4650 & ~n16567 ;
  assign n30162 = n10384 ^ n2582 ^ 1'b0 ;
  assign n30163 = ( ~n3109 & n8382 ) | ( ~n3109 & n15735 ) | ( n8382 & n15735 ) ;
  assign n30164 = ( ~n4327 & n30162 ) | ( ~n4327 & n30163 ) | ( n30162 & n30163 ) ;
  assign n30165 = ( n3771 & n30161 ) | ( n3771 & ~n30164 ) | ( n30161 & ~n30164 ) ;
  assign n30166 = n17468 ^ n7518 ^ 1'b0 ;
  assign n30167 = ~n17159 & n30166 ;
  assign n30168 = n7116 & n30167 ;
  assign n30169 = n9350 & ~n16007 ;
  assign n30170 = ~n5278 & n30169 ;
  assign n30171 = n30170 ^ n18802 ^ 1'b0 ;
  assign n30172 = n29334 & ~n30171 ;
  assign n30173 = n5451 | n12523 ;
  assign n30174 = ( ~n20643 & n28061 ) | ( ~n20643 & n30173 ) | ( n28061 & n30173 ) ;
  assign n30179 = n8053 ^ n425 ^ n295 ;
  assign n30178 = ( n1953 & n3476 ) | ( n1953 & n19991 ) | ( n3476 & n19991 ) ;
  assign n30180 = n30179 ^ n30178 ^ n10241 ;
  assign n30175 = ( ~n5595 & n17959 ) | ( ~n5595 & n25839 ) | ( n17959 & n25839 ) ;
  assign n30176 = n3021 ^ n1278 ^ 1'b0 ;
  assign n30177 = ~n30175 & n30176 ;
  assign n30181 = n30180 ^ n30177 ^ n20677 ;
  assign n30182 = n15728 ^ n8442 ^ 1'b0 ;
  assign n30183 = n28222 ^ n21676 ^ n9971 ;
  assign n30184 = n21908 & n28148 ;
  assign n30185 = ( ~n30182 & n30183 ) | ( ~n30182 & n30184 ) | ( n30183 & n30184 ) ;
  assign n30186 = n22022 ^ n19809 ^ 1'b0 ;
  assign n30191 = n19139 ^ n3629 ^ 1'b0 ;
  assign n30187 = n5509 & n11996 ;
  assign n30188 = n276 & n30187 ;
  assign n30189 = n18436 ^ n11354 ^ n565 ;
  assign n30190 = ( n3718 & n30188 ) | ( n3718 & ~n30189 ) | ( n30188 & ~n30189 ) ;
  assign n30192 = n30191 ^ n30190 ^ n1699 ;
  assign n30193 = ( n11761 & n17307 ) | ( n11761 & ~n29007 ) | ( n17307 & ~n29007 ) ;
  assign n30194 = ( ~n4017 & n8419 ) | ( ~n4017 & n11527 ) | ( n8419 & n11527 ) ;
  assign n30195 = ~n2712 & n11513 ;
  assign n30196 = n30194 & ~n30195 ;
  assign n30197 = n30196 ^ n1760 ^ 1'b0 ;
  assign n30198 = n4288 ^ n990 ^ n930 ;
  assign n30199 = n6173 | n29071 ;
  assign n30200 = n6510 & ~n30199 ;
  assign n30201 = ~n4201 & n24905 ;
  assign n30202 = ~n16177 & n30201 ;
  assign n30203 = n30202 ^ n3536 ^ 1'b0 ;
  assign n30204 = n30200 | n30203 ;
  assign n30205 = n10534 | n30204 ;
  assign n30206 = ( n21712 & n30198 ) | ( n21712 & ~n30205 ) | ( n30198 & ~n30205 ) ;
  assign n30207 = n2731 | n30206 ;
  assign n30208 = n30207 ^ n13724 ^ 1'b0 ;
  assign n30209 = ~n30197 & n30208 ;
  assign n30210 = n909 & ~n7493 ;
  assign n30214 = n8110 ^ n4475 ^ n4145 ;
  assign n30211 = ( n7845 & n16436 ) | ( n7845 & ~n16936 ) | ( n16436 & ~n16936 ) ;
  assign n30212 = n30211 ^ n25166 ^ n4927 ;
  assign n30213 = ~n17888 & n30212 ;
  assign n30215 = n30214 ^ n30213 ^ n9784 ;
  assign n30216 = ~n3226 & n16501 ;
  assign n30217 = n30216 ^ n15056 ^ 1'b0 ;
  assign n30218 = n23329 ^ n3772 ^ 1'b0 ;
  assign n30219 = ~n18835 & n30218 ;
  assign n30220 = n27812 ^ n18623 ^ n11132 ;
  assign n30221 = n7718 ^ n7249 ^ n3083 ;
  assign n30222 = ( n23026 & ~n24745 ) | ( n23026 & n30221 ) | ( ~n24745 & n30221 ) ;
  assign n30223 = n5018 ^ n3979 ^ 1'b0 ;
  assign n30224 = n30223 ^ n7707 ^ 1'b0 ;
  assign n30225 = n30224 ^ n20593 ^ n9589 ;
  assign n30226 = n1566 & ~n9780 ;
  assign n30227 = ( n3645 & n22134 ) | ( n3645 & n30226 ) | ( n22134 & n30226 ) ;
  assign n30228 = ( n3813 & ~n10328 ) | ( n3813 & n30227 ) | ( ~n10328 & n30227 ) ;
  assign n30229 = n30228 ^ n14021 ^ n8996 ;
  assign n30230 = n18127 ^ n16334 ^ 1'b0 ;
  assign n30231 = n3794 ^ n679 ^ x72 ;
  assign n30232 = ( n3560 & n5684 ) | ( n3560 & ~n30231 ) | ( n5684 & ~n30231 ) ;
  assign n30233 = n30232 ^ n29571 ^ 1'b0 ;
  assign n30235 = n14614 ^ n4124 ^ 1'b0 ;
  assign n30234 = n8906 ^ n6226 ^ n751 ;
  assign n30236 = n30235 ^ n30234 ^ n22061 ;
  assign n30237 = n14021 ^ n9046 ^ 1'b0 ;
  assign n30238 = n936 & n13292 ;
  assign n30239 = n30238 ^ n17058 ^ 1'b0 ;
  assign n30240 = n30239 ^ n20884 ^ n5010 ;
  assign n30241 = ( n5799 & n14789 ) | ( n5799 & n30240 ) | ( n14789 & n30240 ) ;
  assign n30245 = ( n4680 & n7966 ) | ( n4680 & ~n14565 ) | ( n7966 & ~n14565 ) ;
  assign n30242 = ( ~n4328 & n6612 ) | ( ~n4328 & n14249 ) | ( n6612 & n14249 ) ;
  assign n30243 = ~n1682 & n30242 ;
  assign n30244 = n25577 & ~n30243 ;
  assign n30246 = n30245 ^ n30244 ^ 1'b0 ;
  assign n30247 = n12272 ^ n9566 ^ 1'b0 ;
  assign n30248 = ~n21887 & n30247 ;
  assign n30249 = n30248 ^ n29342 ^ n26036 ;
  assign n30250 = ( n8320 & n12979 ) | ( n8320 & ~n14253 ) | ( n12979 & ~n14253 ) ;
  assign n30251 = ( n5558 & ~n10007 ) | ( n5558 & n24003 ) | ( ~n10007 & n24003 ) ;
  assign n30252 = n30251 ^ n672 ^ 1'b0 ;
  assign n30253 = n16410 & ~n24889 ;
  assign n30255 = n15573 ^ n3081 ^ 1'b0 ;
  assign n30254 = ~n2500 & n26728 ;
  assign n30256 = n30255 ^ n30254 ^ 1'b0 ;
  assign n30257 = ~n2924 & n27181 ;
  assign n30258 = ~n20365 & n30257 ;
  assign n30259 = n30256 & n30258 ;
  assign n30260 = ( n4520 & ~n4556 ) | ( n4520 & n8550 ) | ( ~n4556 & n8550 ) ;
  assign n30261 = ( n2121 & n9092 ) | ( n2121 & ~n30260 ) | ( n9092 & ~n30260 ) ;
  assign n30262 = n8472 & n30261 ;
  assign n30263 = n4433 & n30262 ;
  assign n30264 = ~n504 & n11908 ;
  assign n30265 = ( n14121 & ~n24622 ) | ( n14121 & n29022 ) | ( ~n24622 & n29022 ) ;
  assign n30266 = n822 | n2801 ;
  assign n30267 = n30266 ^ n21074 ^ 1'b0 ;
  assign n30270 = n14500 | n23183 ;
  assign n30271 = n5007 | n30270 ;
  assign n30268 = n6463 ^ n4589 ^ n3704 ;
  assign n30269 = n30268 ^ n15336 ^ 1'b0 ;
  assign n30272 = n30271 ^ n30269 ^ n13155 ;
  assign n30273 = n18359 | n30272 ;
  assign n30274 = ~n285 & n5456 ;
  assign n30275 = n10131 ^ n5789 ^ n4951 ;
  assign n30276 = n30275 ^ n7199 ^ 1'b0 ;
  assign n30277 = ( n10989 & ~n30274 ) | ( n10989 & n30276 ) | ( ~n30274 & n30276 ) ;
  assign n30278 = n1560 ^ n950 ^ 1'b0 ;
  assign n30279 = ( n20569 & ~n20939 ) | ( n20569 & n21789 ) | ( ~n20939 & n21789 ) ;
  assign n30280 = ( n638 & n18586 ) | ( n638 & n23118 ) | ( n18586 & n23118 ) ;
  assign n30281 = n7065 ^ n1921 ^ 1'b0 ;
  assign n30282 = n6643 ^ n4985 ^ 1'b0 ;
  assign n30283 = n11003 & n30282 ;
  assign n30284 = ( n21375 & n22910 ) | ( n21375 & n29656 ) | ( n22910 & n29656 ) ;
  assign n30285 = n9936 ^ n3067 ^ n1709 ;
  assign n30286 = n943 | n30285 ;
  assign n30287 = n30286 ^ n1118 ^ 1'b0 ;
  assign n30288 = n30287 ^ n12351 ^ 1'b0 ;
  assign n30289 = n5108 & ~n8375 ;
  assign n30290 = ~n3319 & n30289 ;
  assign n30291 = n2022 | n10013 ;
  assign n30292 = n30290 & ~n30291 ;
  assign n30293 = n30292 ^ n18926 ^ n8682 ;
  assign n30294 = n30293 ^ n20355 ^ n18014 ;
  assign n30295 = ( ~n7531 & n13366 ) | ( ~n7531 & n13878 ) | ( n13366 & n13878 ) ;
  assign n30296 = ( ~n5880 & n20587 ) | ( ~n5880 & n24272 ) | ( n20587 & n24272 ) ;
  assign n30297 = ( ~n12311 & n21025 ) | ( ~n12311 & n30296 ) | ( n21025 & n30296 ) ;
  assign n30300 = n29650 ^ n13094 ^ n4138 ;
  assign n30298 = n7940 ^ x59 ^ 1'b0 ;
  assign n30299 = n26007 & n30298 ;
  assign n30301 = n30300 ^ n30299 ^ n8468 ;
  assign n30302 = ( n30295 & n30297 ) | ( n30295 & ~n30301 ) | ( n30297 & ~n30301 ) ;
  assign n30303 = n10009 ^ n8812 ^ n1313 ;
  assign n30304 = n30303 ^ n14770 ^ n4976 ;
  assign n30305 = n30304 ^ n16244 ^ n6778 ;
  assign n30306 = n16890 & ~n30305 ;
  assign n30307 = n16573 ^ n10041 ^ n1367 ;
  assign n30308 = n30307 ^ n2603 ^ n957 ;
  assign n30309 = n22494 | n30308 ;
  assign n30310 = n30309 ^ n7506 ^ 1'b0 ;
  assign n30314 = n17163 ^ n9269 ^ n1296 ;
  assign n30315 = ( x82 & ~n25306 ) | ( x82 & n30314 ) | ( ~n25306 & n30314 ) ;
  assign n30312 = ( ~n8154 & n17937 ) | ( ~n8154 & n26273 ) | ( n17937 & n26273 ) ;
  assign n30311 = n22619 & ~n23385 ;
  assign n30313 = n30312 ^ n30311 ^ 1'b0 ;
  assign n30316 = n30315 ^ n30313 ^ n29972 ;
  assign n30319 = ~n3554 & n14814 ;
  assign n30320 = ~n5824 & n30319 ;
  assign n30317 = n8889 ^ n2933 ^ n999 ;
  assign n30318 = ( n9437 & n27731 ) | ( n9437 & ~n30317 ) | ( n27731 & ~n30317 ) ;
  assign n30321 = n30320 ^ n30318 ^ n29041 ;
  assign n30322 = ( n10737 & n28321 ) | ( n10737 & n30321 ) | ( n28321 & n30321 ) ;
  assign n30323 = n14422 ^ n9567 ^ n3627 ;
  assign n30324 = ( n12811 & n13633 ) | ( n12811 & ~n30323 ) | ( n13633 & ~n30323 ) ;
  assign n30328 = n18150 ^ n6384 ^ n5894 ;
  assign n30325 = n5924 & ~n22659 ;
  assign n30326 = n30325 ^ n22547 ^ 1'b0 ;
  assign n30327 = n11089 & n30326 ;
  assign n30329 = n30328 ^ n30327 ^ 1'b0 ;
  assign n30330 = ~n13660 & n30329 ;
  assign n30331 = n30330 ^ n29809 ^ n4642 ;
  assign n30332 = ( ~n8371 & n25325 ) | ( ~n8371 & n30331 ) | ( n25325 & n30331 ) ;
  assign n30333 = ( n8243 & ~n9192 ) | ( n8243 & n24828 ) | ( ~n9192 & n24828 ) ;
  assign n30334 = ~n1971 & n30333 ;
  assign n30335 = n7345 & n30334 ;
  assign n30336 = n11039 & n30335 ;
  assign n30337 = n30336 ^ n11881 ^ n858 ;
  assign n30338 = n15971 | n17540 ;
  assign n30339 = n30338 ^ n6359 ^ 1'b0 ;
  assign n30342 = ( n2459 & ~n3303 ) | ( n2459 & n4942 ) | ( ~n3303 & n4942 ) ;
  assign n30341 = n8990 ^ n3485 ^ 1'b0 ;
  assign n30343 = n30342 ^ n30341 ^ n18344 ;
  assign n30340 = n18091 & n18207 ;
  assign n30344 = n30343 ^ n30340 ^ n20154 ;
  assign n30345 = n2511 | n27822 ;
  assign n30346 = ( ~n10980 & n28709 ) | ( ~n10980 & n30345 ) | ( n28709 & n30345 ) ;
  assign n30347 = n15071 ^ n2628 ^ 1'b0 ;
  assign n30348 = n12188 | n30347 ;
  assign n30349 = n1112 | n3835 ;
  assign n30353 = n10380 ^ n2427 ^ 1'b0 ;
  assign n30354 = ~n17924 & n30353 ;
  assign n30352 = n3537 & n9967 ;
  assign n30355 = n30354 ^ n30352 ^ 1'b0 ;
  assign n30350 = ( n561 & n5012 ) | ( n561 & ~n21390 ) | ( n5012 & ~n21390 ) ;
  assign n30351 = n943 | n30350 ;
  assign n30356 = n30355 ^ n30351 ^ 1'b0 ;
  assign n30357 = n17230 ^ n7222 ^ 1'b0 ;
  assign n30358 = n30357 ^ n28857 ^ n3575 ;
  assign n30359 = ( n3579 & n13195 ) | ( n3579 & n30358 ) | ( n13195 & n30358 ) ;
  assign n30360 = n14815 ^ n2605 ^ n2271 ;
  assign n30361 = ( n4142 & n6941 ) | ( n4142 & n24277 ) | ( n6941 & n24277 ) ;
  assign n30362 = n724 & ~n24543 ;
  assign n30363 = n30362 ^ n24622 ^ 1'b0 ;
  assign n30364 = ( n1714 & ~n11494 ) | ( n1714 & n30363 ) | ( ~n11494 & n30363 ) ;
  assign n30365 = n11240 | n30364 ;
  assign n30366 = n30365 ^ n17394 ^ 1'b0 ;
  assign n30368 = ( n11166 & ~n16706 ) | ( n11166 & n17837 ) | ( ~n16706 & n17837 ) ;
  assign n30367 = ~n1671 & n6350 ;
  assign n30369 = n30368 ^ n30367 ^ 1'b0 ;
  assign n30370 = n23535 ^ n3709 ^ n2163 ;
  assign n30371 = n16408 & n30370 ;
  assign n30372 = ~n10788 & n30371 ;
  assign n30373 = n9672 ^ n4176 ^ 1'b0 ;
  assign n30374 = n30373 ^ n4589 ^ 1'b0 ;
  assign n30375 = n16227 & n30374 ;
  assign n30376 = ( ~n29767 & n30372 ) | ( ~n29767 & n30375 ) | ( n30372 & n30375 ) ;
  assign n30377 = ~n1239 & n10491 ;
  assign n30378 = ~n4974 & n21665 ;
  assign n30379 = n20677 | n30378 ;
  assign n30380 = n30379 ^ n24543 ^ n13230 ;
  assign n30381 = n30377 | n30380 ;
  assign n30382 = n30381 ^ n24235 ^ n13906 ;
  assign n30383 = ~n1422 & n19898 ;
  assign n30384 = n27434 ^ n16583 ^ n15540 ;
  assign n30385 = ~n4474 & n11589 ;
  assign n30386 = ~n30384 & n30385 ;
  assign n30387 = n5918 | n7653 ;
  assign n30388 = n30387 ^ n18192 ^ 1'b0 ;
  assign n30389 = n18872 ^ n18601 ^ n5740 ;
  assign n30393 = ~n2060 & n11095 ;
  assign n30394 = n30393 ^ n11339 ^ 1'b0 ;
  assign n30395 = n15616 & n30394 ;
  assign n30396 = n22608 | n30395 ;
  assign n30390 = ( ~x103 & n1646 ) | ( ~x103 & n9216 ) | ( n1646 & n9216 ) ;
  assign n30391 = n13692 & ~n30390 ;
  assign n30392 = n7821 & n30391 ;
  assign n30397 = n30396 ^ n30392 ^ n4612 ;
  assign n30398 = ( n17471 & ~n30389 ) | ( n17471 & n30397 ) | ( ~n30389 & n30397 ) ;
  assign n30399 = ( n14449 & ~n30388 ) | ( n14449 & n30398 ) | ( ~n30388 & n30398 ) ;
  assign n30400 = n1016 & n1927 ;
  assign n30401 = n7169 & n30400 ;
  assign n30402 = n8128 ^ n903 ^ 1'b0 ;
  assign n30403 = n30401 | n30402 ;
  assign n30404 = n30403 ^ n27618 ^ x133 ;
  assign n30405 = n1303 & n16435 ;
  assign n30406 = ~n7486 & n30405 ;
  assign n30407 = n30406 ^ n22748 ^ n14995 ;
  assign n30408 = n19298 ^ n18653 ^ n13192 ;
  assign n30409 = ~n5584 & n5833 ;
  assign n30410 = ~n30408 & n30409 ;
  assign n30411 = n13003 ^ n12844 ^ 1'b0 ;
  assign n30412 = n17910 ^ n16359 ^ n8784 ;
  assign n30413 = n30412 ^ n2613 ^ 1'b0 ;
  assign n30414 = ~n6888 & n30413 ;
  assign n30415 = n6500 | n7070 ;
  assign n30416 = n30415 ^ n3834 ^ n2232 ;
  assign n30417 = n12470 | n30416 ;
  assign n30418 = n22757 & ~n30417 ;
  assign n30419 = n16158 | n30418 ;
  assign n30420 = n3626 | n30419 ;
  assign n30422 = x33 & n5238 ;
  assign n30423 = ~x33 & n30422 ;
  assign n30424 = n10140 | n30423 ;
  assign n30425 = n19187 | n30424 ;
  assign n30426 = n30424 & ~n30425 ;
  assign n30421 = ( n8100 & n19499 ) | ( n8100 & ~n20880 ) | ( n19499 & ~n20880 ) ;
  assign n30427 = n30426 ^ n30421 ^ n397 ;
  assign n30428 = ( n5555 & n13465 ) | ( n5555 & ~n20670 ) | ( n13465 & ~n20670 ) ;
  assign n30429 = n9625 ^ n7033 ^ 1'b0 ;
  assign n30430 = n13893 | n30429 ;
  assign n30431 = n30428 & ~n30430 ;
  assign n30432 = ~n25848 & n30431 ;
  assign n30433 = n7472 ^ n6758 ^ 1'b0 ;
  assign n30434 = x160 & ~n5258 ;
  assign n30435 = ~n30433 & n30434 ;
  assign n30436 = n10855 & n12639 ;
  assign n30437 = n30436 ^ n27132 ^ 1'b0 ;
  assign n30438 = n16983 ^ n11857 ^ n8042 ;
  assign n30439 = n30438 ^ n25437 ^ n15001 ;
  assign n30440 = n5797 ^ n450 ^ 1'b0 ;
  assign n30441 = ( ~n3593 & n5518 ) | ( ~n3593 & n24388 ) | ( n5518 & n24388 ) ;
  assign n30442 = ( n4621 & n15932 ) | ( n4621 & n18853 ) | ( n15932 & n18853 ) ;
  assign n30443 = n18201 ^ n17584 ^ 1'b0 ;
  assign n30444 = n20052 & ~n30443 ;
  assign n30445 = n1310 & n30444 ;
  assign n30446 = n8987 & n30445 ;
  assign n30447 = ( n277 & n1146 ) | ( n277 & n12450 ) | ( n1146 & n12450 ) ;
  assign n30448 = n30447 ^ n12497 ^ 1'b0 ;
  assign n30449 = ~n24509 & n30448 ;
  assign n30450 = ~n13404 & n30449 ;
  assign n30451 = n30450 ^ n15542 ^ 1'b0 ;
  assign n30452 = ( n861 & n7971 ) | ( n861 & ~n19268 ) | ( n7971 & ~n19268 ) ;
  assign n30453 = n20295 | n30452 ;
  assign n30454 = ( ~n2563 & n5830 ) | ( ~n2563 & n8082 ) | ( n5830 & n8082 ) ;
  assign n30455 = n10304 ^ n8245 ^ 1'b0 ;
  assign n30456 = n9219 | n30455 ;
  assign n30457 = ( n3500 & n17862 ) | ( n3500 & ~n30456 ) | ( n17862 & ~n30456 ) ;
  assign n30458 = n30454 & ~n30457 ;
  assign n30459 = n30458 ^ n25640 ^ 1'b0 ;
  assign n30460 = n3661 & ~n23815 ;
  assign n30461 = n5530 & ~n30460 ;
  assign n30462 = n30459 & ~n30461 ;
  assign n30463 = ( n3280 & n3456 ) | ( n3280 & n17057 ) | ( n3456 & n17057 ) ;
  assign n30464 = ( n7791 & n10518 ) | ( n7791 & n11679 ) | ( n10518 & n11679 ) ;
  assign n30465 = n30464 ^ n4214 ^ n1865 ;
  assign n30466 = n30465 ^ x197 ^ 1'b0 ;
  assign n30467 = n30463 | n30466 ;
  assign n30468 = n2404 & n21160 ;
  assign n30469 = ( n13004 & ~n19098 ) | ( n13004 & n30468 ) | ( ~n19098 & n30468 ) ;
  assign n30470 = ~n15307 & n27768 ;
  assign n30471 = n30470 ^ n22049 ^ 1'b0 ;
  assign n30475 = n10611 ^ n9993 ^ n9486 ;
  assign n30476 = n11659 ^ n8946 ^ 1'b0 ;
  assign n30477 = ( n13000 & ~n30475 ) | ( n13000 & n30476 ) | ( ~n30475 & n30476 ) ;
  assign n30478 = ( n270 & ~n10722 ) | ( n270 & n18600 ) | ( ~n10722 & n18600 ) ;
  assign n30479 = ( n27874 & ~n30477 ) | ( n27874 & n30478 ) | ( ~n30477 & n30478 ) ;
  assign n30480 = n30479 ^ n22170 ^ n1275 ;
  assign n30474 = n10218 ^ n5285 ^ n5206 ;
  assign n30481 = n30480 ^ n30474 ^ 1'b0 ;
  assign n30472 = ( n10417 & ~n13614 ) | ( n10417 & n16603 ) | ( ~n13614 & n16603 ) ;
  assign n30473 = n30472 ^ n19063 ^ 1'b0 ;
  assign n30482 = n30481 ^ n30473 ^ n15415 ;
  assign n30483 = ( n13570 & n19235 ) | ( n13570 & n29698 ) | ( n19235 & n29698 ) ;
  assign n30484 = n30483 ^ n16146 ^ n7698 ;
  assign n30485 = ( n2510 & ~n6430 ) | ( n2510 & n20249 ) | ( ~n6430 & n20249 ) ;
  assign n30486 = n30485 ^ n8970 ^ 1'b0 ;
  assign n30487 = n14202 ^ n12008 ^ 1'b0 ;
  assign n30489 = n17539 ^ n3804 ^ 1'b0 ;
  assign n30488 = n16526 | n20593 ;
  assign n30490 = n30489 ^ n30488 ^ 1'b0 ;
  assign n30491 = n18583 ^ n876 ^ 1'b0 ;
  assign n30492 = n2417 & n30491 ;
  assign n30493 = n15217 ^ n6998 ^ n5888 ;
  assign n30494 = n1200 & n19685 ;
  assign n30495 = n30494 ^ n3339 ^ 1'b0 ;
  assign n30496 = ( ~n7382 & n23681 ) | ( ~n7382 & n30495 ) | ( n23681 & n30495 ) ;
  assign n30497 = n24483 ^ n11657 ^ n11521 ;
  assign n30498 = ( n6136 & n23640 ) | ( n6136 & n29421 ) | ( n23640 & n29421 ) ;
  assign n30499 = n16546 | n22502 ;
  assign n30500 = n12675 ^ n10800 ^ n8634 ;
  assign n30501 = ( n11842 & n22134 ) | ( n11842 & n30500 ) | ( n22134 & n30500 ) ;
  assign n30502 = ( n24231 & n24397 ) | ( n24231 & ~n30501 ) | ( n24397 & ~n30501 ) ;
  assign n30503 = n27899 ^ n13822 ^ 1'b0 ;
  assign n30504 = ( n8229 & n15976 ) | ( n8229 & ~n30503 ) | ( n15976 & ~n30503 ) ;
  assign n30505 = n30504 ^ n12119 ^ n7920 ;
  assign n30506 = ( n25059 & n26840 ) | ( n25059 & n30206 ) | ( n26840 & n30206 ) ;
  assign n30507 = n30506 ^ n12578 ^ x38 ;
  assign n30508 = n3865 ^ n1078 ^ 1'b0 ;
  assign n30509 = n3864 & n30508 ;
  assign n30510 = n30509 ^ n16923 ^ n11966 ;
  assign n30511 = n30510 ^ n19013 ^ n11101 ;
  assign n30512 = n6520 & n9248 ;
  assign n30513 = n30512 ^ n29532 ^ n2110 ;
  assign n30514 = ~n3951 & n13450 ;
  assign n30515 = n4373 & n30514 ;
  assign n30516 = n22673 ^ x49 ^ 1'b0 ;
  assign n30517 = n27187 ^ n5999 ^ 1'b0 ;
  assign n30518 = n30516 & ~n30517 ;
  assign n30519 = n24858 ^ n20823 ^ 1'b0 ;
  assign n30520 = n10844 & ~n30519 ;
  assign n30521 = ( n318 & ~n11692 ) | ( n318 & n13195 ) | ( ~n11692 & n13195 ) ;
  assign n30522 = ( n1642 & n26513 ) | ( n1642 & ~n30521 ) | ( n26513 & ~n30521 ) ;
  assign n30523 = n30522 ^ n26599 ^ n3344 ;
  assign n30524 = n12299 & ~n13093 ;
  assign n30528 = ( n2461 & ~n9884 ) | ( n2461 & n10495 ) | ( ~n9884 & n10495 ) ;
  assign n30529 = ( n3761 & n6116 ) | ( n3761 & n30528 ) | ( n6116 & n30528 ) ;
  assign n30530 = n30529 ^ n3840 ^ n2149 ;
  assign n30525 = n6208 ^ n4070 ^ n2653 ;
  assign n30526 = n21653 | n30525 ;
  assign n30527 = n30526 ^ n17379 ^ 1'b0 ;
  assign n30531 = n30530 ^ n30527 ^ n4201 ;
  assign n30532 = n2984 & n25278 ;
  assign n30533 = ~n26724 & n30532 ;
  assign n30534 = n14520 ^ n7873 ^ 1'b0 ;
  assign n30537 = n1894 & ~n3295 ;
  assign n30535 = n18140 ^ n4674 ^ n971 ;
  assign n30536 = n30535 ^ n16101 ^ n2325 ;
  assign n30538 = n30537 ^ n30536 ^ n898 ;
  assign n30539 = n13822 | n28299 ;
  assign n30540 = n30539 ^ n2912 ^ 1'b0 ;
  assign n30541 = n7932 ^ n3958 ^ 1'b0 ;
  assign n30542 = ~n28217 & n30541 ;
  assign n30543 = n30540 & n30542 ;
  assign n30544 = n14355 ^ x73 ^ 1'b0 ;
  assign n30545 = n6025 & n30544 ;
  assign n30546 = n30545 ^ n22476 ^ 1'b0 ;
  assign n30547 = n11393 & ~n30546 ;
  assign n30548 = n10859 & n30547 ;
  assign n30549 = ~n18815 & n30548 ;
  assign n30550 = n30549 ^ n26189 ^ n901 ;
  assign n30551 = n16805 | n30550 ;
  assign n30552 = n22395 | n30551 ;
  assign n30553 = n16738 ^ n1262 ^ 1'b0 ;
  assign n30554 = ( ~n20622 & n30334 ) | ( ~n20622 & n30553 ) | ( n30334 & n30553 ) ;
  assign n30555 = n24220 ^ n8761 ^ 1'b0 ;
  assign n30556 = n4365 & n7060 ;
  assign n30557 = n30556 ^ n13924 ^ 1'b0 ;
  assign n30558 = ( n21002 & n22735 ) | ( n21002 & n29269 ) | ( n22735 & n29269 ) ;
  assign n30559 = n30558 ^ n9071 ^ 1'b0 ;
  assign n30560 = ~n7294 & n19638 ;
  assign n30561 = n30560 ^ n22320 ^ 1'b0 ;
  assign n30562 = ( n11756 & n19283 ) | ( n11756 & n21276 ) | ( n19283 & n21276 ) ;
  assign n30563 = n30562 ^ n17984 ^ 1'b0 ;
  assign n30564 = n18506 ^ n13113 ^ 1'b0 ;
  assign n30565 = n24627 ^ n14622 ^ 1'b0 ;
  assign n30566 = ( n14995 & n17794 ) | ( n14995 & n30565 ) | ( n17794 & n30565 ) ;
  assign n30567 = ( ~n8680 & n30564 ) | ( ~n8680 & n30566 ) | ( n30564 & n30566 ) ;
  assign n30569 = n15494 ^ n5533 ^ 1'b0 ;
  assign n30568 = n12447 & n24283 ;
  assign n30570 = n30569 ^ n30568 ^ 1'b0 ;
  assign n30571 = ( n24586 & n24836 ) | ( n24586 & n30570 ) | ( n24836 & n30570 ) ;
  assign n30572 = n17326 | n24815 ;
  assign n30573 = n19565 & ~n30572 ;
  assign n30574 = n20997 ^ n8218 ^ 1'b0 ;
  assign n30575 = n9752 | n30574 ;
  assign n30576 = ~n3937 & n25030 ;
  assign n30577 = ( n6555 & n14355 ) | ( n6555 & ~n30576 ) | ( n14355 & ~n30576 ) ;
  assign n30578 = n30577 ^ n23410 ^ n6118 ;
  assign n30579 = n25127 ^ n22137 ^ 1'b0 ;
  assign n30580 = n12799 ^ n9381 ^ 1'b0 ;
  assign n30581 = n30580 ^ n14279 ^ n3792 ;
  assign n30582 = n13589 ^ n5211 ^ n4773 ;
  assign n30583 = n18758 & ~n30582 ;
  assign n30584 = n19176 & n30583 ;
  assign n30585 = n30540 ^ n11185 ^ 1'b0 ;
  assign n30586 = n19224 ^ n12698 ^ 1'b0 ;
  assign n30587 = n20739 & n30586 ;
  assign n30588 = n30516 ^ n13096 ^ 1'b0 ;
  assign n30589 = n28976 ^ n23642 ^ n1251 ;
  assign n30590 = n15198 ^ n10524 ^ 1'b0 ;
  assign n30591 = n8435 & ~n30590 ;
  assign n30592 = n29046 ^ n14138 ^ 1'b0 ;
  assign n30593 = ~n12618 & n30592 ;
  assign n30594 = n13292 ^ n2996 ^ n741 ;
  assign n30595 = ~n1739 & n5758 ;
  assign n30596 = n8886 & n30595 ;
  assign n30597 = n5581 | n30596 ;
  assign n30598 = n30597 ^ n2951 ^ 1'b0 ;
  assign n30599 = n30598 ^ n3919 ^ n1469 ;
  assign n30600 = n30594 | n30599 ;
  assign n30601 = n30600 ^ n4337 ^ 1'b0 ;
  assign n30602 = ~n4227 & n28684 ;
  assign n30603 = n19488 ^ n11846 ^ 1'b0 ;
  assign n30604 = n26610 & ~n30603 ;
  assign n30605 = n9216 | n30604 ;
  assign n30606 = n5416 & ~n18013 ;
  assign n30607 = n30606 ^ n5282 ^ 1'b0 ;
  assign n30608 = ~n4507 & n5433 ;
  assign n30609 = ( ~n12243 & n28875 ) | ( ~n12243 & n30608 ) | ( n28875 & n30608 ) ;
  assign n30610 = n26464 & n30609 ;
  assign n30611 = ~n30607 & n30610 ;
  assign n30612 = n24696 ^ n7553 ^ 1'b0 ;
  assign n30613 = n16829 & ~n30612 ;
  assign n30614 = ( ~n9409 & n30121 ) | ( ~n9409 & n30613 ) | ( n30121 & n30613 ) ;
  assign n30615 = ( n8816 & n9117 ) | ( n8816 & ~n11124 ) | ( n9117 & ~n11124 ) ;
  assign n30616 = n28055 ^ n20362 ^ n16530 ;
  assign n30617 = n586 | n30616 ;
  assign n30618 = ( ~n24891 & n30615 ) | ( ~n24891 & n30617 ) | ( n30615 & n30617 ) ;
  assign n30619 = n20126 ^ n3644 ^ 1'b0 ;
  assign n30626 = n16295 ^ n12184 ^ n426 ;
  assign n30620 = ( n3262 & n3956 ) | ( n3262 & ~n5121 ) | ( n3956 & ~n5121 ) ;
  assign n30621 = n30620 ^ n26636 ^ n14288 ;
  assign n30623 = ( n4837 & n14548 ) | ( n4837 & ~n17460 ) | ( n14548 & ~n17460 ) ;
  assign n30622 = n9708 | n10054 ;
  assign n30624 = n30623 ^ n30622 ^ n1712 ;
  assign n30625 = ( n6026 & n30621 ) | ( n6026 & ~n30624 ) | ( n30621 & ~n30624 ) ;
  assign n30627 = n30626 ^ n30625 ^ n12768 ;
  assign n30628 = ( ~n1059 & n6049 ) | ( ~n1059 & n8209 ) | ( n6049 & n8209 ) ;
  assign n30629 = ( n3835 & n9618 ) | ( n3835 & n24539 ) | ( n9618 & n24539 ) ;
  assign n30630 = ~n30628 & n30629 ;
  assign n30631 = ( ~n1476 & n1807 ) | ( ~n1476 & n11467 ) | ( n1807 & n11467 ) ;
  assign n30632 = n12104 ^ n7215 ^ 1'b0 ;
  assign n30633 = n14638 | n30632 ;
  assign n30634 = n30633 ^ n23828 ^ n1648 ;
  assign n30635 = n8011 & n30634 ;
  assign n30636 = n30631 & ~n30635 ;
  assign n30637 = n23540 & n30636 ;
  assign n30638 = n11962 ^ n2502 ^ 1'b0 ;
  assign n30639 = n1883 | n30638 ;
  assign n30640 = n30370 & ~n30639 ;
  assign n30641 = n30640 ^ n29457 ^ 1'b0 ;
  assign n30646 = n3579 & ~n21244 ;
  assign n30647 = n30646 ^ n23492 ^ 1'b0 ;
  assign n30644 = n1669 | n12653 ;
  assign n30645 = n30644 ^ n12923 ^ 1'b0 ;
  assign n30642 = n21460 | n24779 ;
  assign n30643 = n30642 ^ n10046 ^ 1'b0 ;
  assign n30648 = n30647 ^ n30645 ^ n30643 ;
  assign n30649 = n1727 | n13678 ;
  assign n30650 = ~n13780 & n29317 ;
  assign n30651 = ~n30649 & n30650 ;
  assign n30652 = n14004 & ~n30651 ;
  assign n30653 = n30652 ^ n19405 ^ 1'b0 ;
  assign n30654 = ( ~n8015 & n16602 ) | ( ~n8015 & n23839 ) | ( n16602 & n23839 ) ;
  assign n30655 = n13407 & n30654 ;
  assign n30656 = n3965 ^ n519 ^ 1'b0 ;
  assign n30657 = ~n16155 & n24048 ;
  assign n30658 = ( n1759 & n8093 ) | ( n1759 & ~n10364 ) | ( n8093 & ~n10364 ) ;
  assign n30659 = n1164 | n15773 ;
  assign n30660 = n16283 & ~n30659 ;
  assign n30662 = n5696 | n15648 ;
  assign n30663 = n30662 ^ n3630 ^ 1'b0 ;
  assign n30661 = n5347 & ~n19629 ;
  assign n30664 = n30663 ^ n30661 ^ 1'b0 ;
  assign n30665 = n23279 ^ n18461 ^ 1'b0 ;
  assign n30666 = ( n19523 & n23197 ) | ( n19523 & n30665 ) | ( n23197 & n30665 ) ;
  assign n30667 = n2070 ^ x147 ^ 1'b0 ;
  assign n30668 = n8915 & ~n30667 ;
  assign n30669 = n30666 & n30668 ;
  assign n30670 = ( n3092 & n3730 ) | ( n3092 & ~n8995 ) | ( n3730 & ~n8995 ) ;
  assign n30671 = n30670 ^ n16647 ^ n12378 ;
  assign n30672 = n30671 ^ n1152 ^ 1'b0 ;
  assign n30673 = n30669 | n30672 ;
  assign n30674 = n16443 ^ n5126 ^ 1'b0 ;
  assign n30675 = ~n25346 & n30674 ;
  assign n30676 = n7471 & n10369 ;
  assign n30677 = n30676 ^ n16174 ^ 1'b0 ;
  assign n30678 = n30360 ^ n6671 ^ 1'b0 ;
  assign n30679 = n542 & n8057 ;
  assign n30680 = n30679 ^ n21415 ^ n1544 ;
  assign n30681 = ( n1532 & ~n13006 ) | ( n1532 & n23748 ) | ( ~n13006 & n23748 ) ;
  assign n30682 = ( n4755 & n17330 ) | ( n4755 & ~n19510 ) | ( n17330 & ~n19510 ) ;
  assign n30683 = n30682 ^ n26852 ^ 1'b0 ;
  assign n30684 = n8053 & n30683 ;
  assign n30685 = n1598 & n6797 ;
  assign n30686 = n10198 & n30685 ;
  assign n30687 = n29470 & n29565 ;
  assign n30688 = ~n1547 & n30687 ;
  assign n30689 = n26343 ^ n11954 ^ n1694 ;
  assign n30690 = n30689 ^ n13744 ^ 1'b0 ;
  assign n30691 = ~n13290 & n30690 ;
  assign n30695 = n16045 & ~n21020 ;
  assign n30692 = n17963 ^ n10327 ^ 1'b0 ;
  assign n30693 = ( ~n12719 & n21017 ) | ( ~n12719 & n30692 ) | ( n21017 & n30692 ) ;
  assign n30694 = ~n12757 & n30693 ;
  assign n30696 = n30695 ^ n30694 ^ 1'b0 ;
  assign n30697 = n29061 ^ n9991 ^ 1'b0 ;
  assign n30698 = n30697 ^ n24338 ^ n12972 ;
  assign n30699 = n4652 & ~n13534 ;
  assign n30700 = n30699 ^ n3252 ^ 1'b0 ;
  assign n30701 = n30700 ^ n14956 ^ n10675 ;
  assign n30702 = ~n893 & n1197 ;
  assign n30703 = ~n16326 & n30702 ;
  assign n30704 = n30703 ^ n12781 ^ 1'b0 ;
  assign n30705 = ~n22325 & n30704 ;
  assign n30706 = n10976 | n29581 ;
  assign n30707 = n30706 ^ n12207 ^ 1'b0 ;
  assign n30708 = ~n29023 & n30707 ;
  assign n30710 = ~n1833 & n8231 ;
  assign n30709 = n15575 & n21981 ;
  assign n30711 = n30710 ^ n30709 ^ n12177 ;
  assign n30712 = ( n28097 & ~n28582 ) | ( n28097 & n30711 ) | ( ~n28582 & n30711 ) ;
  assign n30714 = n10983 ^ n6831 ^ n926 ;
  assign n30713 = ( n5123 & n7423 ) | ( n5123 & n8219 ) | ( n7423 & n8219 ) ;
  assign n30715 = n30714 ^ n30713 ^ n24360 ;
  assign n30716 = n30715 ^ n20942 ^ n1042 ;
  assign n30717 = n12823 & ~n19476 ;
  assign n30718 = n30717 ^ n14653 ^ 1'b0 ;
  assign n30719 = ( x22 & ~n13590 ) | ( x22 & n28176 ) | ( ~n13590 & n28176 ) ;
  assign n30720 = n30719 ^ n25686 ^ n3195 ;
  assign n30721 = n16743 ^ n5948 ^ 1'b0 ;
  assign n30722 = n30721 ^ n8682 ^ 1'b0 ;
  assign n30723 = ( n793 & ~n22600 ) | ( n793 & n28367 ) | ( ~n22600 & n28367 ) ;
  assign n30724 = ~n2735 & n7890 ;
  assign n30725 = n30724 ^ n2791 ^ 1'b0 ;
  assign n30726 = n8141 & ~n15347 ;
  assign n30727 = ~n901 & n30726 ;
  assign n30728 = n26238 & n30727 ;
  assign n30729 = ~n30725 & n30728 ;
  assign n30730 = n11018 ^ n10139 ^ 1'b0 ;
  assign n30731 = n30730 ^ n13415 ^ 1'b0 ;
  assign n30732 = n30731 ^ n15066 ^ 1'b0 ;
  assign n30733 = n22744 & n25475 ;
  assign n30734 = n30733 ^ n28803 ^ 1'b0 ;
  assign n30735 = n30734 ^ n15989 ^ 1'b0 ;
  assign n30736 = ( ~n1239 & n4420 ) | ( ~n1239 & n29441 ) | ( n4420 & n29441 ) ;
  assign n30737 = ( n15405 & n30667 ) | ( n15405 & n30736 ) | ( n30667 & n30736 ) ;
  assign n30738 = n20729 ^ n4206 ^ 1'b0 ;
  assign n30739 = n15338 ^ n4713 ^ 1'b0 ;
  assign n30740 = n3144 & ~n30739 ;
  assign n30741 = n30740 ^ n8301 ^ 1'b0 ;
  assign n30742 = n17626 & ~n25466 ;
  assign n30744 = n17752 ^ n12073 ^ 1'b0 ;
  assign n30745 = ( n9344 & n21537 ) | ( n9344 & n30744 ) | ( n21537 & n30744 ) ;
  assign n30746 = n30745 ^ n15491 ^ n14523 ;
  assign n30743 = ( n13115 & n20275 ) | ( n13115 & ~n23102 ) | ( n20275 & ~n23102 ) ;
  assign n30747 = n30746 ^ n30743 ^ n30714 ;
  assign n30748 = n12931 ^ n12104 ^ 1'b0 ;
  assign n30749 = n7339 & ~n7965 ;
  assign n30750 = n6509 & n13210 ;
  assign n30751 = ( n18670 & n30749 ) | ( n18670 & n30750 ) | ( n30749 & n30750 ) ;
  assign n30752 = n14183 ^ x65 ^ 1'b0 ;
  assign n30753 = n2955 | n9490 ;
  assign n30754 = ( n6838 & n16739 ) | ( n6838 & ~n30753 ) | ( n16739 & ~n30753 ) ;
  assign n30755 = n27919 & ~n30754 ;
  assign n30756 = n6490 | n17800 ;
  assign n30757 = n13096 | n30756 ;
  assign n30758 = n9248 & n30757 ;
  assign n30759 = n19119 & ~n30758 ;
  assign n30761 = n15612 ^ n14789 ^ 1'b0 ;
  assign n30760 = n19502 ^ n6213 ^ 1'b0 ;
  assign n30762 = n30761 ^ n30760 ^ n1879 ;
  assign n30763 = n18180 ^ n14121 ^ n3060 ;
  assign n30764 = n30763 ^ n17440 ^ 1'b0 ;
  assign n30766 = ( n7539 & n12873 ) | ( n7539 & n19122 ) | ( n12873 & n19122 ) ;
  assign n30765 = n5047 & ~n12070 ;
  assign n30767 = n30766 ^ n30765 ^ 1'b0 ;
  assign n30768 = n30767 ^ n26013 ^ n20413 ;
  assign n30769 = n11622 & ~n27959 ;
  assign n30770 = ~n30768 & n30769 ;
  assign n30771 = n15523 & ~n30770 ;
  assign n30772 = n30764 & n30771 ;
  assign n30773 = n30772 ^ n3031 ^ 1'b0 ;
  assign n30774 = ( n16580 & n23690 ) | ( n16580 & ~n27888 ) | ( n23690 & ~n27888 ) ;
  assign n30775 = ( ~n6289 & n18337 ) | ( ~n6289 & n20293 ) | ( n18337 & n20293 ) ;
  assign n30776 = n3151 ^ n2141 ^ n2020 ;
  assign n30777 = n30776 ^ n21850 ^ 1'b0 ;
  assign n30778 = n25867 & n30777 ;
  assign n30779 = n30778 ^ n10977 ^ 1'b0 ;
  assign n30780 = ( n5278 & n7633 ) | ( n5278 & ~n22337 ) | ( n7633 & ~n22337 ) ;
  assign n30781 = ( n5683 & ~n6115 ) | ( n5683 & n30780 ) | ( ~n6115 & n30780 ) ;
  assign n30782 = n5257 & ~n30781 ;
  assign n30783 = n30782 ^ n11512 ^ 1'b0 ;
  assign n30786 = x189 & n9673 ;
  assign n30787 = n30786 ^ n1572 ^ 1'b0 ;
  assign n30788 = ( n6662 & ~n25107 ) | ( n6662 & n30787 ) | ( ~n25107 & n30787 ) ;
  assign n30784 = n12808 & ~n25797 ;
  assign n30785 = ( n8148 & ~n16392 ) | ( n8148 & n30784 ) | ( ~n16392 & n30784 ) ;
  assign n30789 = n30788 ^ n30785 ^ n3353 ;
  assign n30790 = n22125 | n30789 ;
  assign n30791 = n30783 | n30790 ;
  assign n30792 = ( ~n11823 & n12424 ) | ( ~n11823 & n30791 ) | ( n12424 & n30791 ) ;
  assign n30793 = n30792 ^ n17256 ^ 1'b0 ;
  assign n30794 = n13320 & n20726 ;
  assign n30795 = n29765 & n30794 ;
  assign n30796 = n16021 | n30795 ;
  assign n30801 = n12359 ^ n10915 ^ 1'b0 ;
  assign n30797 = n4632 | n23228 ;
  assign n30798 = n13299 & ~n30797 ;
  assign n30799 = n30798 ^ n26685 ^ 1'b0 ;
  assign n30800 = n6164 & ~n30799 ;
  assign n30802 = n30801 ^ n30800 ^ 1'b0 ;
  assign n30803 = ~n30796 & n30802 ;
  assign n30805 = n4293 | n14919 ;
  assign n30804 = ~n6332 & n9747 ;
  assign n30806 = n30805 ^ n30804 ^ 1'b0 ;
  assign n30807 = ( ~n5320 & n13080 ) | ( ~n5320 & n24768 ) | ( n13080 & n24768 ) ;
  assign n30808 = n30807 ^ n14234 ^ 1'b0 ;
  assign n30809 = ~n11893 & n30808 ;
  assign n30810 = n21592 | n30809 ;
  assign n30811 = ( n16545 & n30806 ) | ( n16545 & ~n30810 ) | ( n30806 & ~n30810 ) ;
  assign n30814 = n25262 ^ n12067 ^ n6613 ;
  assign n30812 = n647 | n14540 ;
  assign n30813 = n30812 ^ n5660 ^ 1'b0 ;
  assign n30815 = n30814 ^ n30813 ^ x206 ;
  assign n30816 = n4850 | n5717 ;
  assign n30817 = n18048 ^ n6883 ^ 1'b0 ;
  assign n30818 = n9061 & ~n30817 ;
  assign n30819 = n11452 ^ n3837 ^ n3117 ;
  assign n30820 = n8226 | n8902 ;
  assign n30821 = n6253 & ~n30820 ;
  assign n30822 = ( n2371 & ~n12017 ) | ( n2371 & n19605 ) | ( ~n12017 & n19605 ) ;
  assign n30823 = ( n11682 & n30821 ) | ( n11682 & ~n30822 ) | ( n30821 & ~n30822 ) ;
  assign n30824 = n26220 ^ n3667 ^ 1'b0 ;
  assign n30825 = n24602 & ~n30824 ;
  assign n30826 = n14382 & n30825 ;
  assign n30827 = n23441 ^ n13262 ^ 1'b0 ;
  assign n30828 = n30827 ^ n16416 ^ 1'b0 ;
  assign n30829 = n7300 & ~n24278 ;
  assign n30832 = n5709 ^ n2080 ^ n1491 ;
  assign n30831 = n17743 ^ n11181 ^ n5962 ;
  assign n30830 = ( n12230 & n12523 ) | ( n12230 & n29524 ) | ( n12523 & n29524 ) ;
  assign n30833 = n30832 ^ n30831 ^ n30830 ;
  assign n30838 = ~n9448 & n12879 ;
  assign n30834 = n15804 ^ n1002 ^ 1'b0 ;
  assign n30835 = ~n14172 & n30834 ;
  assign n30836 = n3065 & n30835 ;
  assign n30837 = n30836 ^ n26074 ^ 1'b0 ;
  assign n30839 = n30838 ^ n30837 ^ n8124 ;
  assign n30840 = n19178 ^ n13481 ^ n2594 ;
  assign n30841 = n30840 ^ n9148 ^ 1'b0 ;
  assign n30842 = n16311 | n30359 ;
  assign n30847 = n21287 ^ n4752 ^ n1645 ;
  assign n30845 = n802 & n14234 ;
  assign n30846 = ~n16762 & n30845 ;
  assign n30843 = ( n10975 & ~n17104 ) | ( n10975 & n27976 ) | ( ~n17104 & n27976 ) ;
  assign n30844 = ( n16961 & n28940 ) | ( n16961 & n30843 ) | ( n28940 & n30843 ) ;
  assign n30848 = n30847 ^ n30846 ^ n30844 ;
  assign n30849 = x17 & n13863 ;
  assign n30850 = n30849 ^ n5785 ^ 1'b0 ;
  assign n30851 = n8939 | n30850 ;
  assign n30852 = n8436 | n21837 ;
  assign n30853 = n30852 ^ n23348 ^ n2623 ;
  assign n30854 = ( n12093 & ~n30851 ) | ( n12093 & n30853 ) | ( ~n30851 & n30853 ) ;
  assign n30855 = n30854 ^ n9799 ^ 1'b0 ;
  assign n30856 = n30848 | n30855 ;
  assign n30857 = n19601 ^ n16351 ^ 1'b0 ;
  assign n30863 = ~n8287 & n15383 ;
  assign n30864 = n30863 ^ n17426 ^ 1'b0 ;
  assign n30858 = ~n4568 & n13781 ;
  assign n30859 = ~n11945 & n30858 ;
  assign n30860 = ( n2424 & n17268 ) | ( n2424 & ~n30859 ) | ( n17268 & ~n30859 ) ;
  assign n30861 = n1701 & ~n30860 ;
  assign n30862 = ( n692 & n28987 ) | ( n692 & n30861 ) | ( n28987 & n30861 ) ;
  assign n30865 = n30864 ^ n30862 ^ n20165 ;
  assign n30867 = n18917 ^ n14113 ^ 1'b0 ;
  assign n30866 = n25165 ^ n16249 ^ 1'b0 ;
  assign n30868 = n30867 ^ n30866 ^ n3624 ;
  assign n30869 = n1892 & ~n26101 ;
  assign n30870 = n30869 ^ n16217 ^ n1474 ;
  assign n30871 = n8168 & ~n25108 ;
  assign n30872 = n30871 ^ n25385 ^ 1'b0 ;
  assign n30873 = n30872 ^ n22968 ^ 1'b0 ;
  assign n30874 = ( ~n6808 & n7776 ) | ( ~n6808 & n18713 ) | ( n7776 & n18713 ) ;
  assign n30875 = ( n15538 & n18087 ) | ( n15538 & ~n20126 ) | ( n18087 & ~n20126 ) ;
  assign n30876 = ( n2099 & n10077 ) | ( n2099 & n30875 ) | ( n10077 & n30875 ) ;
  assign n30877 = ( n18508 & n30874 ) | ( n18508 & n30876 ) | ( n30874 & n30876 ) ;
  assign n30878 = n24285 & ~n30877 ;
  assign n30879 = n30878 ^ n2085 ^ 1'b0 ;
  assign n30882 = n7631 & ~n16071 ;
  assign n30883 = ~n426 & n30882 ;
  assign n30884 = ~n10520 & n22414 ;
  assign n30885 = n30883 & n30884 ;
  assign n30886 = n30885 ^ n15488 ^ n2775 ;
  assign n30880 = n14518 ^ n11204 ^ n2069 ;
  assign n30881 = n30880 ^ n26691 ^ n17433 ;
  assign n30887 = n30886 ^ n30881 ^ 1'b0 ;
  assign n30888 = n12546 ^ n11022 ^ 1'b0 ;
  assign n30889 = n19201 ^ n971 ^ 1'b0 ;
  assign n30890 = n9788 | n12735 ;
  assign n30891 = n11192 & n30890 ;
  assign n30892 = n11637 ^ n7322 ^ 1'b0 ;
  assign n30893 = n27008 & ~n30892 ;
  assign n30894 = n8710 & ~n17562 ;
  assign n30895 = n30894 ^ n28024 ^ 1'b0 ;
  assign n30896 = n30854 ^ n24819 ^ n15884 ;
  assign n30897 = n12493 ^ n735 ^ x152 ;
  assign n30898 = x65 & ~n20367 ;
  assign n30899 = ( n1310 & n2155 ) | ( n1310 & ~n7860 ) | ( n2155 & ~n7860 ) ;
  assign n30900 = n28820 & ~n30899 ;
  assign n30901 = n30900 ^ n3996 ^ 1'b0 ;
  assign n30902 = ~n15966 & n24298 ;
  assign n30903 = n30902 ^ n28254 ^ 1'b0 ;
  assign n30904 = n9217 & n26464 ;
  assign n30905 = ~n15791 & n30904 ;
  assign n30906 = n16702 ^ n15632 ^ n9045 ;
  assign n30907 = n10555 ^ n8842 ^ 1'b0 ;
  assign n30908 = n28983 ^ n2918 ^ 1'b0 ;
  assign n30909 = n5350 & ~n30908 ;
  assign n30911 = n21204 ^ n16266 ^ n1754 ;
  assign n30910 = n5830 & n19785 ;
  assign n30912 = n30911 ^ n30910 ^ 1'b0 ;
  assign n30913 = n28353 ^ n4642 ^ 1'b0 ;
  assign n30914 = ( ~n6862 & n7351 ) | ( ~n6862 & n30913 ) | ( n7351 & n30913 ) ;
  assign n30915 = n15533 ^ n11436 ^ 1'b0 ;
  assign n30917 = n23169 ^ n18998 ^ n9402 ;
  assign n30916 = n30055 ^ n27049 ^ n22651 ;
  assign n30918 = n30917 ^ n30916 ^ n23294 ;
  assign n30919 = n6529 & ~n23207 ;
  assign n30920 = n4373 | n19557 ;
  assign n30921 = n30920 ^ n3339 ^ 1'b0 ;
  assign n30922 = n15725 & n30921 ;
  assign n30923 = n30919 | n30922 ;
  assign n30924 = ( n7531 & n8985 ) | ( n7531 & ~n12891 ) | ( n8985 & ~n12891 ) ;
  assign n30925 = n13935 ^ n13148 ^ 1'b0 ;
  assign n30926 = n14234 & n30925 ;
  assign n30927 = n24929 ^ n13453 ^ 1'b0 ;
  assign n30928 = n30927 ^ n2500 ^ n1977 ;
  assign n30929 = n6472 & n11720 ;
  assign n30930 = ( ~n22121 & n24084 ) | ( ~n22121 & n30929 ) | ( n24084 & n30929 ) ;
  assign n30931 = ( n11060 & n27863 ) | ( n11060 & n29444 ) | ( n27863 & n29444 ) ;
  assign n30932 = n12426 & n21795 ;
  assign n30933 = ~n11653 & n30932 ;
  assign n30934 = n30933 ^ n13183 ^ 1'b0 ;
  assign n30938 = n14501 & n28836 ;
  assign n30939 = ~n7919 & n30938 ;
  assign n30940 = n30939 ^ n29306 ^ 1'b0 ;
  assign n30941 = ~n10856 & n30940 ;
  assign n30935 = ( n7719 & n9292 ) | ( n7719 & ~n11634 ) | ( n9292 & ~n11634 ) ;
  assign n30936 = n20413 ^ n14375 ^ 1'b0 ;
  assign n30937 = ~n30935 & n30936 ;
  assign n30942 = n30941 ^ n30937 ^ 1'b0 ;
  assign n30943 = ~n285 & n15264 ;
  assign n30944 = n30943 ^ n15261 ^ 1'b0 ;
  assign n30945 = ( n5769 & ~n21327 ) | ( n5769 & n27766 ) | ( ~n21327 & n27766 ) ;
  assign n30946 = n324 | n7137 ;
  assign n30947 = n11210 | n30946 ;
  assign n30948 = n23316 & ~n30947 ;
  assign n30949 = ~n4078 & n16573 ;
  assign n30953 = ( n2348 & ~n9007 ) | ( n2348 & n10356 ) | ( ~n9007 & n10356 ) ;
  assign n30950 = n7604 ^ x138 ^ 1'b0 ;
  assign n30951 = n6360 & ~n30950 ;
  assign n30952 = ( ~n10300 & n22242 ) | ( ~n10300 & n30951 ) | ( n22242 & n30951 ) ;
  assign n30954 = n30953 ^ n30952 ^ 1'b0 ;
  assign n30955 = ( n6810 & ~n16486 ) | ( n6810 & n30954 ) | ( ~n16486 & n30954 ) ;
  assign n30956 = n30955 ^ n23333 ^ 1'b0 ;
  assign n30957 = ~n30949 & n30956 ;
  assign n30958 = n18013 ^ n603 ^ 1'b0 ;
  assign n30959 = n25879 ^ n24065 ^ 1'b0 ;
  assign n30960 = n28415 & n30959 ;
  assign n30961 = n30415 ^ n7982 ^ 1'b0 ;
  assign n30962 = n10819 ^ n4998 ^ n2560 ;
  assign n30963 = n14303 ^ n458 ^ 1'b0 ;
  assign n30964 = n30963 ^ n7465 ^ n786 ;
  assign n30965 = ( ~n22438 & n30962 ) | ( ~n22438 & n30964 ) | ( n30962 & n30964 ) ;
  assign n30966 = n8482 & ~n14101 ;
  assign n30967 = n15589 ^ n2780 ^ n405 ;
  assign n30968 = n30967 ^ n13291 ^ n9475 ;
  assign n30969 = n19065 ^ n16292 ^ 1'b0 ;
  assign n30970 = n30968 | n30969 ;
  assign n30971 = ( n1760 & n7047 ) | ( n1760 & ~n17847 ) | ( n7047 & ~n17847 ) ;
  assign n30972 = x249 & ~n12744 ;
  assign n30973 = ~n30971 & n30972 ;
  assign n30974 = n5522 & n16878 ;
  assign n30975 = n27572 ^ n9016 ^ 1'b0 ;
  assign n30976 = n1014 & ~n30975 ;
  assign n30977 = ~n19843 & n30976 ;
  assign n30978 = n19231 ^ n12882 ^ 1'b0 ;
  assign n30979 = ( ~n6132 & n9533 ) | ( ~n6132 & n20076 ) | ( n9533 & n20076 ) ;
  assign n30980 = n13836 ^ n8702 ^ 1'b0 ;
  assign n30981 = ( ~n286 & n16442 ) | ( ~n286 & n18965 ) | ( n16442 & n18965 ) ;
  assign n30982 = ( n16295 & ~n19190 ) | ( n16295 & n23336 ) | ( ~n19190 & n23336 ) ;
  assign n30983 = n30982 ^ n4487 ^ 1'b0 ;
  assign n30984 = n30981 | n30983 ;
  assign n30985 = n22680 & ~n30984 ;
  assign n30994 = n14257 & ~n21600 ;
  assign n30995 = ( n17004 & n25016 ) | ( n17004 & n30994 ) | ( n25016 & n30994 ) ;
  assign n30986 = n14499 & n20913 ;
  assign n30987 = n30986 ^ n13233 ^ n7809 ;
  assign n30988 = n30987 ^ n22042 ^ 1'b0 ;
  assign n30989 = n14192 & ~n30988 ;
  assign n30990 = n28617 ^ n3448 ^ 1'b0 ;
  assign n30991 = n30989 & n30990 ;
  assign n30992 = n28106 & n30991 ;
  assign n30993 = n30992 ^ n12807 ^ 1'b0 ;
  assign n30996 = n30995 ^ n30993 ^ n27291 ;
  assign n30997 = ( n3419 & n6201 ) | ( n3419 & ~n19806 ) | ( n6201 & ~n19806 ) ;
  assign n30998 = n18765 & ~n30997 ;
  assign n30999 = n30998 ^ n3440 ^ n632 ;
  assign n31000 = n4097 & ~n5941 ;
  assign n31001 = n12915 & ~n31000 ;
  assign n31002 = ~n8105 & n31001 ;
  assign n31003 = n19565 ^ n13599 ^ 1'b0 ;
  assign n31004 = ~n4378 & n31003 ;
  assign n31005 = n16894 ^ n5626 ^ 1'b0 ;
  assign n31006 = n31005 ^ n10467 ^ n1333 ;
  assign n31007 = ~n7356 & n14641 ;
  assign n31008 = n31007 ^ n14572 ^ 1'b0 ;
  assign n31009 = ( n18403 & n23908 ) | ( n18403 & n31008 ) | ( n23908 & n31008 ) ;
  assign n31010 = n16351 ^ n7146 ^ 1'b0 ;
  assign n31011 = n16980 | n31010 ;
  assign n31012 = ~n20389 & n31011 ;
  assign n31013 = ( n2764 & n2885 ) | ( n2764 & ~n18237 ) | ( n2885 & ~n18237 ) ;
  assign n31014 = n31013 ^ n20732 ^ 1'b0 ;
  assign n31015 = n31014 ^ n12392 ^ n12368 ;
  assign n31016 = n30887 ^ n6773 ^ n1044 ;
  assign n31017 = ~n5719 & n9881 ;
  assign n31018 = ~n8201 & n31017 ;
  assign n31019 = n10770 ^ n7910 ^ n670 ;
  assign n31020 = n31019 ^ n4256 ^ 1'b0 ;
  assign n31021 = n17077 ^ n13754 ^ 1'b0 ;
  assign n31022 = ( n4789 & n31020 ) | ( n4789 & n31021 ) | ( n31020 & n31021 ) ;
  assign n31023 = n31022 ^ n24618 ^ n4958 ;
  assign n31024 = ( n8484 & n9056 ) | ( n8484 & ~n20343 ) | ( n9056 & ~n20343 ) ;
  assign n31025 = ( n5609 & ~n8798 ) | ( n5609 & n24371 ) | ( ~n8798 & n24371 ) ;
  assign n31026 = n4315 | n13791 ;
  assign n31027 = n21872 & ~n31026 ;
  assign n31028 = ~n21261 & n24170 ;
  assign n31029 = n16670 & n31028 ;
  assign n31030 = n4379 | n11042 ;
  assign n31031 = n31030 ^ n30626 ^ n12670 ;
  assign n31032 = n15898 ^ n11823 ^ n8100 ;
  assign n31033 = n7098 & n14507 ;
  assign n31034 = ~n1570 & n11443 ;
  assign n31035 = n31034 ^ n5316 ^ 1'b0 ;
  assign n31036 = n31035 ^ n21899 ^ 1'b0 ;
  assign n31037 = n31033 | n31036 ;
  assign n31038 = ( n2545 & n23968 ) | ( n2545 & ~n31037 ) | ( n23968 & ~n31037 ) ;
  assign n31039 = ( n11473 & n14419 ) | ( n11473 & ~n16042 ) | ( n14419 & ~n16042 ) ;
  assign n31041 = n25916 ^ n9155 ^ 1'b0 ;
  assign n31040 = n29781 ^ n22854 ^ n735 ;
  assign n31042 = n31041 ^ n31040 ^ n23928 ;
  assign n31043 = n31042 ^ n4592 ^ 1'b0 ;
  assign n31044 = n16588 ^ n12587 ^ 1'b0 ;
  assign n31045 = ~n1779 & n31044 ;
  assign n31047 = n15517 ^ n5535 ^ n4360 ;
  assign n31048 = n31047 ^ n25561 ^ n7108 ;
  assign n31046 = ( n4338 & n16409 ) | ( n4338 & ~n17979 ) | ( n16409 & ~n17979 ) ;
  assign n31049 = n31048 ^ n31046 ^ 1'b0 ;
  assign n31050 = n23214 & ~n31049 ;
  assign n31051 = n14873 ^ n6141 ^ n5456 ;
  assign n31052 = n13490 & ~n31051 ;
  assign n31053 = n31052 ^ x77 ^ 1'b0 ;
  assign n31054 = n21793 ^ n14880 ^ 1'b0 ;
  assign n31055 = n6220 | n31054 ;
  assign n31056 = n31055 ^ n27784 ^ n21034 ;
  assign n31057 = n4817 | n23758 ;
  assign n31058 = n10552 ^ n1163 ^ 1'b0 ;
  assign n31059 = ( n26267 & n31057 ) | ( n26267 & ~n31058 ) | ( n31057 & ~n31058 ) ;
  assign n31061 = ~n3353 & n10891 ;
  assign n31062 = n31061 ^ n7669 ^ 1'b0 ;
  assign n31060 = n14576 ^ n11172 ^ 1'b0 ;
  assign n31063 = n31062 ^ n31060 ^ n25423 ;
  assign n31064 = n9791 | n23324 ;
  assign n31065 = n27493 & n31064 ;
  assign n31066 = ( n3489 & n3636 ) | ( n3489 & n8886 ) | ( n3636 & n8886 ) ;
  assign n31067 = ~n12068 & n31066 ;
  assign n31068 = n1353 & ~n2171 ;
  assign n31069 = n31068 ^ n19009 ^ 1'b0 ;
  assign n31070 = ( n13318 & n29659 ) | ( n13318 & ~n31069 ) | ( n29659 & ~n31069 ) ;
  assign n31078 = x228 & n10299 ;
  assign n31079 = n9872 & n31078 ;
  assign n31076 = n17782 ^ n10415 ^ n10261 ;
  assign n31077 = ( n7791 & ~n21436 ) | ( n7791 & n31076 ) | ( ~n21436 & n31076 ) ;
  assign n31071 = n25867 ^ n6219 ^ n1909 ;
  assign n31072 = n31071 ^ n30649 ^ n11668 ;
  assign n31073 = n31072 ^ n28047 ^ n4063 ;
  assign n31074 = n11416 | n31073 ;
  assign n31075 = n7426 | n31074 ;
  assign n31080 = n31079 ^ n31077 ^ n31075 ;
  assign n31081 = n13096 ^ n9742 ^ n4682 ;
  assign n31082 = n17736 & ~n23955 ;
  assign n31083 = n31082 ^ n25584 ^ 1'b0 ;
  assign n31084 = n25253 ^ n16855 ^ 1'b0 ;
  assign n31085 = n5781 & n31084 ;
  assign n31086 = n24852 ^ n15165 ^ 1'b0 ;
  assign n31087 = n13027 | n16357 ;
  assign n31091 = n5634 & ~n17966 ;
  assign n31092 = ~n4451 & n31091 ;
  assign n31088 = n18161 ^ n601 ^ 1'b0 ;
  assign n31089 = n4416 ^ n562 ^ 1'b0 ;
  assign n31090 = n31088 | n31089 ;
  assign n31093 = n31092 ^ n31090 ^ 1'b0 ;
  assign n31094 = n900 & ~n12495 ;
  assign n31095 = n31094 ^ n10814 ^ 1'b0 ;
  assign n31096 = ~n15585 & n31095 ;
  assign n31097 = n4003 & n31096 ;
  assign n31098 = n9623 ^ n3279 ^ n1886 ;
  assign n31099 = n1468 & n31098 ;
  assign n31100 = n31099 ^ n16431 ^ 1'b0 ;
  assign n31101 = n10635 & ~n13858 ;
  assign n31102 = n31101 ^ n6336 ^ 1'b0 ;
  assign n31103 = ~n14481 & n25228 ;
  assign n31104 = n31103 ^ n18631 ^ 1'b0 ;
  assign n31105 = ( n6805 & n8528 ) | ( n6805 & n31104 ) | ( n8528 & n31104 ) ;
  assign n31106 = ( ~n9694 & n31102 ) | ( ~n9694 & n31105 ) | ( n31102 & n31105 ) ;
  assign n31107 = n15526 ^ n8634 ^ 1'b0 ;
  assign n31108 = n23484 ^ n21866 ^ n19932 ;
  assign n31109 = n31108 ^ n7881 ^ n735 ;
  assign n31110 = n24491 & n31109 ;
  assign n31111 = n26711 ^ n19631 ^ 1'b0 ;
  assign n31112 = n25345 ^ n6592 ^ 1'b0 ;
  assign n31113 = ( n2251 & n15883 ) | ( n2251 & n31112 ) | ( n15883 & n31112 ) ;
  assign n31114 = n31113 ^ n26342 ^ n19368 ;
  assign n31117 = ~n448 & n13328 ;
  assign n31115 = n5814 & ~n13055 ;
  assign n31116 = ( n11954 & n17516 ) | ( n11954 & n31115 ) | ( n17516 & n31115 ) ;
  assign n31118 = n31117 ^ n31116 ^ 1'b0 ;
  assign n31119 = n25912 ^ n4626 ^ 1'b0 ;
  assign n31120 = n7858 & ~n31119 ;
  assign n31121 = n31120 ^ n3497 ^ 1'b0 ;
  assign n31122 = n31118 & n31121 ;
  assign n31125 = n13764 ^ n5944 ^ n5330 ;
  assign n31123 = ~n733 & n6957 ;
  assign n31124 = n20073 | n31123 ;
  assign n31126 = n31125 ^ n31124 ^ n14285 ;
  assign n31127 = n23545 ^ n22096 ^ n4266 ;
  assign n31128 = ( n1625 & n7216 ) | ( n1625 & n11657 ) | ( n7216 & n11657 ) ;
  assign n31129 = n8580 ^ n7387 ^ 1'b0 ;
  assign n31130 = ( n2348 & n25450 ) | ( n2348 & ~n31129 ) | ( n25450 & ~n31129 ) ;
  assign n31131 = ( n14439 & n29071 ) | ( n14439 & n31130 ) | ( n29071 & n31130 ) ;
  assign n31132 = n6285 ^ n740 ^ 1'b0 ;
  assign n31133 = ~n14799 & n31132 ;
  assign n31134 = n31133 ^ n8486 ^ 1'b0 ;
  assign n31135 = ~n14370 & n14677 ;
  assign n31136 = n31135 ^ n20634 ^ 1'b0 ;
  assign n31137 = n9530 ^ n9455 ^ n9270 ;
  assign n31138 = n19298 ^ n10155 ^ n3604 ;
  assign n31139 = n17640 ^ n13780 ^ 1'b0 ;
  assign n31140 = n15466 ^ n5091 ^ 1'b0 ;
  assign n31141 = n4166 & ~n31140 ;
  assign n31143 = n22809 ^ n21526 ^ n15603 ;
  assign n31142 = n13017 | n22355 ;
  assign n31144 = n31143 ^ n31142 ^ 1'b0 ;
  assign n31145 = ~n14462 & n31144 ;
  assign n31146 = ~n4121 & n31145 ;
  assign n31147 = n31146 ^ n11663 ^ 1'b0 ;
  assign n31148 = n31147 ^ n10919 ^ n8228 ;
  assign n31150 = n12048 ^ n1163 ^ 1'b0 ;
  assign n31151 = n1968 & n31150 ;
  assign n31149 = n18310 ^ n5549 ^ n1603 ;
  assign n31152 = n31151 ^ n31149 ^ n23469 ;
  assign n31153 = n7305 & ~n12972 ;
  assign n31154 = n10019 & ~n20326 ;
  assign n31155 = ~n31153 & n31154 ;
  assign n31156 = n27501 ^ n24476 ^ n11819 ;
  assign n31157 = ( n9474 & n9523 ) | ( n9474 & ~n15121 ) | ( n9523 & ~n15121 ) ;
  assign n31158 = ~n1985 & n31157 ;
  assign n31159 = ~n31156 & n31158 ;
  assign n31160 = n22748 ^ n8331 ^ x132 ;
  assign n31161 = ( ~n6326 & n9633 ) | ( ~n6326 & n23758 ) | ( n9633 & n23758 ) ;
  assign n31162 = ~n25464 & n31161 ;
  assign n31163 = ~n31160 & n31162 ;
  assign n31164 = ( n665 & n15842 ) | ( n665 & ~n18620 ) | ( n15842 & ~n18620 ) ;
  assign n31168 = ( n1241 & n10113 ) | ( n1241 & ~n11506 ) | ( n10113 & ~n11506 ) ;
  assign n31165 = n11096 & ~n23166 ;
  assign n31166 = n15546 & ~n31165 ;
  assign n31167 = ~n21609 & n31166 ;
  assign n31169 = n31168 ^ n31167 ^ n27731 ;
  assign n31170 = ( ~n2031 & n5902 ) | ( ~n2031 & n17154 ) | ( n5902 & n17154 ) ;
  assign n31171 = n19133 | n24504 ;
  assign n31172 = n31171 ^ n27759 ^ n7119 ;
  assign n31173 = n31170 | n31172 ;
  assign n31174 = n13500 | n31173 ;
  assign n31175 = n26891 ^ n2432 ^ n2271 ;
  assign n31176 = n13645 & ~n31175 ;
  assign n31177 = n7219 & n9457 ;
  assign n31178 = ( n2511 & n5564 ) | ( n2511 & n31177 ) | ( n5564 & n31177 ) ;
  assign n31179 = n1248 | n19489 ;
  assign n31180 = n14375 ^ n10025 ^ n4880 ;
  assign n31181 = n21888 | n31180 ;
  assign n31182 = n5275 | n25345 ;
  assign n31183 = n31182 ^ n7553 ^ 1'b0 ;
  assign n31184 = ( n3825 & ~n13127 ) | ( n3825 & n31183 ) | ( ~n13127 & n31183 ) ;
  assign n31185 = n3905 ^ n1447 ^ 1'b0 ;
  assign n31186 = ( ~n1714 & n2515 ) | ( ~n1714 & n31185 ) | ( n2515 & n31185 ) ;
  assign n31187 = ~n13478 & n31186 ;
  assign n31188 = ~n18485 & n31187 ;
  assign n31189 = n31188 ^ n26532 ^ n1892 ;
  assign n31190 = n25163 | n31189 ;
  assign n31191 = n4300 | n16603 ;
  assign n31192 = ~n6261 & n8900 ;
  assign n31193 = ~n7736 & n31192 ;
  assign n31194 = n31193 ^ n23084 ^ n551 ;
  assign n31195 = n12999 ^ n1023 ^ 1'b0 ;
  assign n31196 = n2565 | n31195 ;
  assign n31197 = n31196 ^ n24174 ^ n5803 ;
  assign n31198 = ( n4929 & ~n7616 ) | ( n4929 & n30594 ) | ( ~n7616 & n30594 ) ;
  assign n31199 = ~n4575 & n31198 ;
  assign n31200 = n6385 | n10984 ;
  assign n31201 = n31200 ^ n5499 ^ 1'b0 ;
  assign n31202 = ~n24109 & n31201 ;
  assign n31203 = n22688 ^ n16054 ^ 1'b0 ;
  assign n31204 = ~n7035 & n31203 ;
  assign n31205 = n10946 ^ n8810 ^ n5340 ;
  assign n31206 = ( n10155 & n21441 ) | ( n10155 & ~n31205 ) | ( n21441 & ~n31205 ) ;
  assign n31207 = n14382 ^ n12261 ^ n12227 ;
  assign n31208 = n31206 & n31207 ;
  assign n31209 = n8434 & n31208 ;
  assign n31210 = n13408 | n29120 ;
  assign n31211 = n9523 | n31210 ;
  assign n31212 = n17368 ^ n16563 ^ 1'b0 ;
  assign n31213 = n28177 & n31212 ;
  assign n31214 = n10709 ^ n5917 ^ 1'b0 ;
  assign n31215 = ( n8785 & n26247 ) | ( n8785 & ~n31214 ) | ( n26247 & ~n31214 ) ;
  assign n31216 = n3446 & n4010 ;
  assign n31217 = n11816 | n13572 ;
  assign n31218 = n5490 & ~n31217 ;
  assign n31219 = n12551 & ~n31218 ;
  assign n31220 = n31219 ^ n30579 ^ 1'b0 ;
  assign n31221 = n24164 & ~n27871 ;
  assign n31224 = ~n11112 & n19440 ;
  assign n31225 = n31224 ^ n22294 ^ 1'b0 ;
  assign n31222 = n7590 | n25253 ;
  assign n31223 = n31222 ^ n24951 ^ x91 ;
  assign n31226 = n31225 ^ n31223 ^ n25176 ;
  assign n31227 = n7912 | n31117 ;
  assign n31228 = ( n12898 & ~n17926 ) | ( n12898 & n18542 ) | ( ~n17926 & n18542 ) ;
  assign n31229 = n31228 ^ n9086 ^ 1'b0 ;
  assign n31230 = n31227 & n31229 ;
  assign n31231 = n30205 ^ n5184 ^ n3559 ;
  assign n31232 = ~n27108 & n31231 ;
  assign n31233 = ( n7873 & n26259 ) | ( n7873 & n31232 ) | ( n26259 & n31232 ) ;
  assign n31234 = ( n4164 & n6251 ) | ( n4164 & n7614 ) | ( n6251 & n7614 ) ;
  assign n31235 = n31234 ^ n1621 ^ 1'b0 ;
  assign n31236 = n29557 ^ n13593 ^ 1'b0 ;
  assign n31237 = ( ~n6745 & n27169 ) | ( ~n6745 & n31236 ) | ( n27169 & n31236 ) ;
  assign n31238 = n6729 & n26918 ;
  assign n31239 = n6232 & n31238 ;
  assign n31240 = ( ~n14277 & n26979 ) | ( ~n14277 & n31239 ) | ( n26979 & n31239 ) ;
  assign n31241 = n12673 & n31240 ;
  assign n31242 = n25633 & n31241 ;
  assign n31243 = ~n848 & n9702 ;
  assign n31244 = ( ~n7910 & n28639 ) | ( ~n7910 & n31243 ) | ( n28639 & n31243 ) ;
  assign n31245 = ( n467 & n3080 ) | ( n467 & ~n17490 ) | ( n3080 & ~n17490 ) ;
  assign n31246 = n31245 ^ n25412 ^ n20754 ;
  assign n31249 = n1288 | n12948 ;
  assign n31247 = ( n7862 & ~n8189 ) | ( n7862 & n12960 ) | ( ~n8189 & n12960 ) ;
  assign n31248 = ( ~n5719 & n6106 ) | ( ~n5719 & n31247 ) | ( n6106 & n31247 ) ;
  assign n31250 = n31249 ^ n31248 ^ n30707 ;
  assign n31251 = n1604 | n7820 ;
  assign n31252 = n31251 ^ n943 ^ 1'b0 ;
  assign n31253 = n26872 | n27597 ;
  assign n31254 = n31252 & ~n31253 ;
  assign n31255 = ( ~x35 & n6899 ) | ( ~x35 & n17385 ) | ( n6899 & n17385 ) ;
  assign n31256 = n31255 ^ x243 ^ 1'b0 ;
  assign n31257 = ( n3017 & ~n5246 ) | ( n3017 & n31256 ) | ( ~n5246 & n31256 ) ;
  assign n31258 = n8625 & ~n12035 ;
  assign n31259 = ( n23990 & ~n29548 ) | ( n23990 & n31258 ) | ( ~n29548 & n31258 ) ;
  assign n31260 = n16836 & ~n30647 ;
  assign n31261 = n9234 & n31260 ;
  assign n31262 = n3387 & n22799 ;
  assign n31263 = ( ~n4225 & n13740 ) | ( ~n4225 & n13992 ) | ( n13740 & n13992 ) ;
  assign n31264 = ( n4397 & ~n7129 ) | ( n4397 & n9793 ) | ( ~n7129 & n9793 ) ;
  assign n31265 = ( n21810 & n31263 ) | ( n21810 & ~n31264 ) | ( n31263 & ~n31264 ) ;
  assign n31268 = n5192 ^ n4469 ^ n3337 ;
  assign n31266 = ( n467 & n4164 ) | ( n467 & ~n11618 ) | ( n4164 & ~n11618 ) ;
  assign n31267 = n31266 ^ n16927 ^ n6366 ;
  assign n31269 = n31268 ^ n31267 ^ 1'b0 ;
  assign n31270 = n23508 & n31269 ;
  assign n31271 = n15616 | n29049 ;
  assign n31274 = n4038 & n4953 ;
  assign n31275 = n14055 | n31274 ;
  assign n31276 = n31275 ^ n4975 ^ 1'b0 ;
  assign n31272 = ( ~n2939 & n12376 ) | ( ~n2939 & n16440 ) | ( n12376 & n16440 ) ;
  assign n31273 = ( ~n2348 & n6092 ) | ( ~n2348 & n31272 ) | ( n6092 & n31272 ) ;
  assign n31277 = n31276 ^ n31273 ^ n28148 ;
  assign n31278 = n31271 & n31277 ;
  assign n31279 = n14873 ^ n14503 ^ n14471 ;
  assign n31280 = ( n23324 & n28337 ) | ( n23324 & ~n29454 ) | ( n28337 & ~n29454 ) ;
  assign n31281 = ( n15412 & n17639 ) | ( n15412 & ~n18510 ) | ( n17639 & ~n18510 ) ;
  assign n31282 = ( n13088 & n13245 ) | ( n13088 & n16243 ) | ( n13245 & n16243 ) ;
  assign n31283 = ( n15456 & n31281 ) | ( n15456 & ~n31282 ) | ( n31281 & ~n31282 ) ;
  assign n31284 = n10368 ^ n1745 ^ 1'b0 ;
  assign n31285 = n31284 ^ n26618 ^ 1'b0 ;
  assign n31286 = n31285 ^ n23834 ^ n7995 ;
  assign n31287 = n7463 | n9580 ;
  assign n31288 = n31287 ^ n15226 ^ 1'b0 ;
  assign n31289 = ~n31286 & n31288 ;
  assign n31290 = n9157 ^ n1862 ^ 1'b0 ;
  assign n31291 = n6359 & n31290 ;
  assign n31292 = n7620 ^ n3360 ^ 1'b0 ;
  assign n31293 = ~n6059 & n11013 ;
  assign n31294 = n31293 ^ n21991 ^ 1'b0 ;
  assign n31295 = n3948 & n31294 ;
  assign n31296 = ( n22997 & n31292 ) | ( n22997 & ~n31295 ) | ( n31292 & ~n31295 ) ;
  assign n31297 = n16561 ^ n5720 ^ n2229 ;
  assign n31298 = ~n23683 & n26333 ;
  assign n31299 = ~n16730 & n31298 ;
  assign n31300 = ~n6168 & n31299 ;
  assign n31301 = n6080 | n19187 ;
  assign n31302 = n31301 ^ n6476 ^ 1'b0 ;
  assign n31303 = n23871 ^ n847 ^ 1'b0 ;
  assign n31304 = n14257 & ~n31303 ;
  assign n31305 = n14046 ^ n12759 ^ n10173 ;
  assign n31306 = n1582 & n31305 ;
  assign n31307 = ~n5354 & n31306 ;
  assign n31308 = n5509 ^ n1739 ^ 1'b0 ;
  assign n31309 = n31307 | n31308 ;
  assign n31310 = n14369 | n14991 ;
  assign n31311 = ( n5500 & n30350 ) | ( n5500 & ~n31310 ) | ( n30350 & ~n31310 ) ;
  assign n31312 = n678 & n24331 ;
  assign n31313 = n10651 ^ x96 ^ 1'b0 ;
  assign n31314 = n31313 ^ n5472 ^ n2521 ;
  assign n31315 = n31314 ^ n27724 ^ 1'b0 ;
  assign n31317 = ~n2785 & n4298 ;
  assign n31318 = n741 & n31317 ;
  assign n31319 = n31318 ^ n5765 ^ 1'b0 ;
  assign n31316 = n16284 ^ n12756 ^ n4613 ;
  assign n31320 = n31319 ^ n31316 ^ 1'b0 ;
  assign n31321 = ~n4621 & n31320 ;
  assign n31322 = n30875 ^ n13346 ^ n11550 ;
  assign n31323 = n10364 ^ n7502 ^ 1'b0 ;
  assign n31324 = n31323 ^ n17844 ^ n3293 ;
  assign n31325 = n31324 ^ n27528 ^ n13724 ;
  assign n31326 = ( n18567 & ~n24092 ) | ( n18567 & n27701 ) | ( ~n24092 & n27701 ) ;
  assign n31327 = n27845 & ~n30273 ;
  assign n31328 = n1806 & n6301 ;
  assign n31329 = n31328 ^ n12285 ^ 1'b0 ;
  assign n31330 = ~n4129 & n31329 ;
  assign n31331 = ( n1297 & n7674 ) | ( n1297 & n31330 ) | ( n7674 & n31330 ) ;
  assign n31332 = n4807 ^ n4527 ^ n1901 ;
  assign n31333 = ( n5827 & ~n18628 ) | ( n5827 & n31115 ) | ( ~n18628 & n31115 ) ;
  assign n31334 = ~n15379 & n23728 ;
  assign n31335 = n24874 ^ n11824 ^ n5170 ;
  assign n31336 = n14040 ^ n12583 ^ n1635 ;
  assign n31337 = n31335 & ~n31336 ;
  assign n31338 = n2060 | n6999 ;
  assign n31339 = n31338 ^ n5431 ^ 1'b0 ;
  assign n31340 = n570 & n31339 ;
  assign n31341 = n31340 ^ n29107 ^ n27715 ;
  assign n31342 = n14235 ^ n5171 ^ n5072 ;
  assign n31343 = ~n13379 & n31342 ;
  assign n31344 = n22158 & ~n31343 ;
  assign n31345 = n2528 & n11622 ;
  assign n31346 = ~n15666 & n31345 ;
  assign n31347 = n14822 & ~n31346 ;
  assign n31348 = ( n9971 & ~n31344 ) | ( n9971 & n31347 ) | ( ~n31344 & n31347 ) ;
  assign n31349 = n16438 & ~n22853 ;
  assign n31350 = n30957 ^ n11748 ^ 1'b0 ;
  assign n31351 = ~n31349 & n31350 ;
  assign n31352 = ( x238 & ~n4932 ) | ( x238 & n11868 ) | ( ~n4932 & n11868 ) ;
  assign n31353 = n1438 | n31352 ;
  assign n31354 = n31353 ^ n17826 ^ n7139 ;
  assign n31355 = ( ~n3815 & n15272 ) | ( ~n3815 & n31354 ) | ( n15272 & n31354 ) ;
  assign n31356 = n31355 ^ n20823 ^ n4598 ;
  assign n31357 = n21217 ^ n13872 ^ 1'b0 ;
  assign n31358 = ( n26230 & n31356 ) | ( n26230 & ~n31357 ) | ( n31356 & ~n31357 ) ;
  assign n31359 = ( n1684 & n5773 ) | ( n1684 & n31358 ) | ( n5773 & n31358 ) ;
  assign n31360 = ( ~n11366 & n15479 ) | ( ~n11366 & n30228 ) | ( n15479 & n30228 ) ;
  assign n31361 = ( n9845 & n10139 ) | ( n9845 & ~n15336 ) | ( n10139 & ~n15336 ) ;
  assign n31362 = n31361 ^ x140 ^ 1'b0 ;
  assign n31363 = n28576 & ~n31362 ;
  assign n31364 = ( ~n3217 & n31360 ) | ( ~n3217 & n31363 ) | ( n31360 & n31363 ) ;
  assign n31366 = n11040 ^ n2266 ^ 1'b0 ;
  assign n31365 = n5127 | n18839 ;
  assign n31367 = n31366 ^ n31365 ^ 1'b0 ;
  assign n31368 = n1187 | n6844 ;
  assign n31373 = n17393 ^ n9301 ^ n3972 ;
  assign n31372 = ~n9980 & n12573 ;
  assign n31369 = n20221 ^ n746 ^ 1'b0 ;
  assign n31370 = ( n25725 & ~n28179 ) | ( n25725 & n31369 ) | ( ~n28179 & n31369 ) ;
  assign n31371 = ( n3290 & ~n26396 ) | ( n3290 & n31370 ) | ( ~n26396 & n31370 ) ;
  assign n31374 = n31373 ^ n31372 ^ n31371 ;
  assign n31375 = ( ~x5 & n6557 ) | ( ~x5 & n7126 ) | ( n6557 & n7126 ) ;
  assign n31376 = n18344 ^ n6626 ^ n2390 ;
  assign n31377 = n31376 ^ n11066 ^ x38 ;
  assign n31378 = n31377 ^ n15623 ^ 1'b0 ;
  assign n31379 = n31375 & ~n31378 ;
  assign n31380 = n376 | n19375 ;
  assign n31381 = n31380 ^ n26363 ^ 1'b0 ;
  assign n31382 = ( x170 & n16064 ) | ( x170 & n20939 ) | ( n16064 & n20939 ) ;
  assign n31383 = n29397 | n31382 ;
  assign n31384 = n17922 | n31383 ;
  assign n31385 = ( n7516 & n7917 ) | ( n7516 & ~n7922 ) | ( n7917 & ~n7922 ) ;
  assign n31386 = n31385 ^ n6869 ^ n5797 ;
  assign n31387 = ( n540 & ~n8063 ) | ( n540 & n13651 ) | ( ~n8063 & n13651 ) ;
  assign n31388 = n23240 & n31387 ;
  assign n31389 = n7784 & ~n27600 ;
  assign n31390 = n6324 | n12550 ;
  assign n31391 = n31390 ^ n9721 ^ 1'b0 ;
  assign n31392 = ( n9192 & n12456 ) | ( n9192 & ~n12982 ) | ( n12456 & ~n12982 ) ;
  assign n31393 = n31392 ^ n14543 ^ 1'b0 ;
  assign n31394 = n29423 ^ n2254 ^ 1'b0 ;
  assign n31395 = n31394 ^ n21577 ^ 1'b0 ;
  assign n31396 = ~n31393 & n31395 ;
  assign n31397 = n14977 ^ n8678 ^ 1'b0 ;
  assign n31398 = n31397 ^ n12507 ^ 1'b0 ;
  assign n31399 = n7528 & ~n31398 ;
  assign n31400 = n12587 ^ n11737 ^ 1'b0 ;
  assign n31401 = n31400 ^ n6040 ^ 1'b0 ;
  assign n31402 = n18647 ^ n4942 ^ 1'b0 ;
  assign n31403 = n31402 ^ n9732 ^ n4405 ;
  assign n31404 = n11674 ^ n378 ^ 1'b0 ;
  assign n31405 = n23705 | n31404 ;
  assign n31406 = n13865 & n17046 ;
  assign n31407 = n31406 ^ n30164 ^ n8024 ;
  assign n31408 = ~n6564 & n11697 ;
  assign n31409 = n31408 ^ n6031 ^ 1'b0 ;
  assign n31410 = n14010 & ~n24371 ;
  assign n31411 = ~n18658 & n31410 ;
  assign n31412 = ( n21652 & ~n31409 ) | ( n21652 & n31411 ) | ( ~n31409 & n31411 ) ;
  assign n31413 = ( ~n31405 & n31407 ) | ( ~n31405 & n31412 ) | ( n31407 & n31412 ) ;
  assign n31414 = n21999 ^ n8654 ^ 1'b0 ;
  assign n31415 = n12062 ^ n9140 ^ n2669 ;
  assign n31416 = n29207 | n31415 ;
  assign n31417 = n12831 ^ n11754 ^ 1'b0 ;
  assign n31418 = n29078 ^ n26867 ^ 1'b0 ;
  assign n31419 = ~n31417 & n31418 ;
  assign n31420 = n30615 ^ n17469 ^ n7352 ;
  assign n31421 = n31420 ^ n873 ^ 1'b0 ;
  assign n31422 = n22004 ^ n7907 ^ 1'b0 ;
  assign n31423 = ~n31421 & n31422 ;
  assign n31424 = ( ~n16988 & n21355 ) | ( ~n16988 & n26355 ) | ( n21355 & n26355 ) ;
  assign n31425 = n26719 ^ n24064 ^ n12258 ;
  assign n31426 = ( ~n19035 & n31424 ) | ( ~n19035 & n31425 ) | ( n31424 & n31425 ) ;
  assign n31427 = ( ~n10763 & n25345 ) | ( ~n10763 & n26712 ) | ( n25345 & n26712 ) ;
  assign n31428 = n15024 | n19037 ;
  assign n31429 = n31428 ^ n29899 ^ n10587 ;
  assign n31430 = ( n8880 & n14772 ) | ( n8880 & n31429 ) | ( n14772 & n31429 ) ;
  assign n31431 = ( n18409 & ~n23968 ) | ( n18409 & n31430 ) | ( ~n23968 & n31430 ) ;
  assign n31438 = ~n8077 & n18355 ;
  assign n31439 = ~n16760 & n31438 ;
  assign n31436 = n9193 ^ n4848 ^ 1'b0 ;
  assign n31437 = n22191 | n31436 ;
  assign n31440 = n31439 ^ n31437 ^ 1'b0 ;
  assign n31432 = n6877 | n14135 ;
  assign n31433 = n26583 ^ n11514 ^ 1'b0 ;
  assign n31434 = n31433 ^ n16696 ^ 1'b0 ;
  assign n31435 = ~n31432 & n31434 ;
  assign n31441 = n31440 ^ n31435 ^ 1'b0 ;
  assign n31442 = ( n562 & n12065 ) | ( n562 & n17283 ) | ( n12065 & n17283 ) ;
  assign n31443 = n4481 | n31442 ;
  assign n31444 = n31443 ^ n8828 ^ 1'b0 ;
  assign n31445 = n3326 & n31444 ;
  assign n31446 = n20883 & ~n28556 ;
  assign n31447 = n31446 ^ n2537 ^ 1'b0 ;
  assign n31448 = n20883 ^ n16503 ^ 1'b0 ;
  assign n31449 = n18118 & ~n31448 ;
  assign n31450 = n4966 & n9569 ;
  assign n31451 = ~n9569 & n31450 ;
  assign n31452 = n31451 ^ n1814 ^ 1'b0 ;
  assign n31453 = n31449 & ~n31452 ;
  assign n31455 = n1784 | n19620 ;
  assign n31456 = n31455 ^ n3861 ^ 1'b0 ;
  assign n31457 = ( n20317 & n23339 ) | ( n20317 & ~n31456 ) | ( n23339 & ~n31456 ) ;
  assign n31454 = n5325 & ~n16433 ;
  assign n31458 = n31457 ^ n31454 ^ 1'b0 ;
  assign n31461 = n5310 ^ n2118 ^ n2069 ;
  assign n31459 = n7405 ^ x169 ^ 1'b0 ;
  assign n31460 = n1803 | n31459 ;
  assign n31462 = n31461 ^ n31460 ^ n22411 ;
  assign n31463 = ( n10885 & n25369 ) | ( n10885 & n31462 ) | ( n25369 & n31462 ) ;
  assign n31464 = n4798 | n8643 ;
  assign n31465 = n31464 ^ n4315 ^ 1'b0 ;
  assign n31466 = n14073 | n31465 ;
  assign n31467 = ( n4962 & n14594 ) | ( n4962 & n16327 ) | ( n14594 & n16327 ) ;
  assign n31468 = n18935 ^ n5650 ^ 1'b0 ;
  assign n31469 = ( n5752 & ~n9732 ) | ( n5752 & n29714 ) | ( ~n9732 & n29714 ) ;
  assign n31470 = n31469 ^ n7271 ^ 1'b0 ;
  assign n31471 = n8313 & n31470 ;
  assign n31472 = n16329 ^ n16149 ^ n14351 ;
  assign n31473 = ~n6124 & n20403 ;
  assign n31474 = ~n18301 & n31473 ;
  assign n31475 = n31474 ^ x33 ^ 1'b0 ;
  assign n31476 = n31472 & ~n31475 ;
  assign n31477 = n20687 & n26571 ;
  assign n31478 = n10417 & ~n23054 ;
  assign n31479 = n31477 & n31478 ;
  assign n31480 = n3185 & ~n8909 ;
  assign n31481 = n31480 ^ n13723 ^ 1'b0 ;
  assign n31482 = n12805 ^ n8614 ^ 1'b0 ;
  assign n31483 = ( ~n4518 & n4585 ) | ( ~n4518 & n31482 ) | ( n4585 & n31482 ) ;
  assign n31484 = ~n9267 & n31483 ;
  assign n31485 = n31484 ^ n19133 ^ 1'b0 ;
  assign n31486 = n31485 ^ n17139 ^ n11172 ;
  assign n31487 = n5789 & n22437 ;
  assign n31488 = n31487 ^ n16909 ^ 1'b0 ;
  assign n31489 = ~n1510 & n10491 ;
  assign n31490 = ( n4123 & ~n8043 ) | ( n4123 & n22171 ) | ( ~n8043 & n22171 ) ;
  assign n31491 = ( n17369 & n21741 ) | ( n17369 & ~n31490 ) | ( n21741 & ~n31490 ) ;
  assign n31497 = n5075 & n10571 ;
  assign n31495 = n1932 & n8462 ;
  assign n31496 = n31495 ^ n4272 ^ 1'b0 ;
  assign n31492 = n11873 ^ n1277 ^ 1'b0 ;
  assign n31493 = ~n5236 & n31492 ;
  assign n31494 = n1334 & ~n31493 ;
  assign n31498 = n31497 ^ n31496 ^ n31494 ;
  assign n31499 = n9275 & ~n14178 ;
  assign n31500 = n2944 & n31499 ;
  assign n31501 = n22474 | n31500 ;
  assign n31502 = ( ~n8821 & n9836 ) | ( ~n8821 & n13399 ) | ( n9836 & n13399 ) ;
  assign n31503 = n31502 ^ n8582 ^ 1'b0 ;
  assign n31504 = n21686 ^ n3257 ^ 1'b0 ;
  assign n31505 = n5337 & n31504 ;
  assign n31506 = n21737 ^ n4698 ^ 1'b0 ;
  assign n31507 = n2973 | n31506 ;
  assign n31508 = ( n5336 & n15953 ) | ( n5336 & n20186 ) | ( n15953 & n20186 ) ;
  assign n31509 = n31508 ^ n4089 ^ n1637 ;
  assign n31510 = ( n2217 & n13440 ) | ( n2217 & n31509 ) | ( n13440 & n31509 ) ;
  assign n31511 = n12454 | n31510 ;
  assign n31512 = n23963 & ~n31511 ;
  assign n31513 = n31512 ^ n30021 ^ n20581 ;
  assign n31514 = ( n11179 & n18679 ) | ( n11179 & n23424 ) | ( n18679 & n23424 ) ;
  assign n31515 = n14762 ^ n14629 ^ n10976 ;
  assign n31516 = n31515 ^ n19131 ^ n10902 ;
  assign n31517 = n31516 ^ n11068 ^ n5478 ;
  assign n31518 = n31517 ^ n13891 ^ n13767 ;
  assign n31519 = n2152 & ~n26268 ;
  assign n31520 = n31519 ^ n27489 ^ 1'b0 ;
  assign n31521 = n25686 ^ n12143 ^ 1'b0 ;
  assign n31522 = n31521 ^ n20003 ^ n17245 ;
  assign n31523 = ( ~n8205 & n22458 ) | ( ~n8205 & n28605 ) | ( n22458 & n28605 ) ;
  assign n31524 = n20824 ^ n10056 ^ x181 ;
  assign n31525 = ( n3562 & ~n8259 ) | ( n3562 & n10191 ) | ( ~n8259 & n10191 ) ;
  assign n31526 = n1138 | n12083 ;
  assign n31527 = n31525 | n31526 ;
  assign n31528 = n31527 ^ n16654 ^ 1'b0 ;
  assign n31529 = n31528 ^ n15598 ^ n5667 ;
  assign n31530 = n7620 & ~n31529 ;
  assign n31532 = n3522 & n20763 ;
  assign n31533 = n31532 ^ n16572 ^ 1'b0 ;
  assign n31534 = ~n13539 & n31533 ;
  assign n31531 = n10255 | n20791 ;
  assign n31535 = n31534 ^ n31531 ^ 1'b0 ;
  assign n31536 = n15360 | n28824 ;
  assign n31537 = n8509 | n28896 ;
  assign n31538 = n28194 & ~n31537 ;
  assign n31539 = ( ~n6579 & n13432 ) | ( ~n6579 & n15328 ) | ( n13432 & n15328 ) ;
  assign n31540 = n31539 ^ n15626 ^ 1'b0 ;
  assign n31541 = n31540 ^ n10176 ^ 1'b0 ;
  assign n31542 = n27894 ^ n18939 ^ n849 ;
  assign n31543 = n12292 ^ n3999 ^ 1'b0 ;
  assign n31544 = n31543 ^ n1041 ^ 1'b0 ;
  assign n31545 = n11137 ^ n7393 ^ n5660 ;
  assign n31546 = ( ~n11218 & n24749 ) | ( ~n11218 & n31545 ) | ( n24749 & n31545 ) ;
  assign n31547 = n26380 ^ n5180 ^ n4103 ;
  assign n31548 = n21152 ^ n16079 ^ 1'b0 ;
  assign n31549 = n22830 & ~n31548 ;
  assign n31550 = n31549 ^ n29822 ^ 1'b0 ;
  assign n31551 = n15426 ^ n13902 ^ 1'b0 ;
  assign n31552 = ( n1779 & n3363 ) | ( n1779 & n5128 ) | ( n3363 & n5128 ) ;
  assign n31553 = ~n466 & n3638 ;
  assign n31554 = ~n22029 & n31553 ;
  assign n31555 = n31554 ^ n7922 ^ n6536 ;
  assign n31556 = ( n31551 & n31552 ) | ( n31551 & n31555 ) | ( n31552 & n31555 ) ;
  assign n31557 = ( n8724 & n16950 ) | ( n8724 & ~n30153 ) | ( n16950 & ~n30153 ) ;
  assign n31558 = n9130 & n31557 ;
  assign n31559 = n27503 ^ n13846 ^ 1'b0 ;
  assign n31560 = n24667 ^ n17534 ^ n10057 ;
  assign n31561 = n29812 ^ n26927 ^ 1'b0 ;
  assign n31563 = ~n1010 & n14294 ;
  assign n31562 = n7483 & n8437 ;
  assign n31564 = n31563 ^ n31562 ^ 1'b0 ;
  assign n31565 = n31564 ^ n12188 ^ 1'b0 ;
  assign n31566 = n31561 & n31565 ;
  assign n31567 = ( ~n631 & n24526 ) | ( ~n631 & n31566 ) | ( n24526 & n31566 ) ;
  assign n31568 = n14045 | n21379 ;
  assign n31569 = n31568 ^ n7382 ^ 1'b0 ;
  assign n31570 = n17658 ^ n13085 ^ n3725 ;
  assign n31571 = ( n6658 & ~n16136 ) | ( n6658 & n18298 ) | ( ~n16136 & n18298 ) ;
  assign n31572 = n31571 ^ n16898 ^ 1'b0 ;
  assign n31573 = n31572 ^ n9919 ^ n7973 ;
  assign n31574 = n5299 & n11378 ;
  assign n31575 = n2714 & n10597 ;
  assign n31576 = n31575 ^ n22312 ^ 1'b0 ;
  assign n31577 = n31576 ^ n31551 ^ n7506 ;
  assign n31578 = ( ~n6648 & n12618 ) | ( ~n6648 & n28241 ) | ( n12618 & n28241 ) ;
  assign n31579 = n6601 & ~n31578 ;
  assign n31580 = n31579 ^ n3331 ^ 1'b0 ;
  assign n31581 = n31580 ^ n21965 ^ 1'b0 ;
  assign n31582 = n31577 | n31581 ;
  assign n31584 = n5713 ^ n384 ^ 1'b0 ;
  assign n31583 = ~n7812 & n22855 ;
  assign n31585 = n31584 ^ n31583 ^ 1'b0 ;
  assign n31586 = n320 & ~n21310 ;
  assign n31587 = ~n6032 & n31586 ;
  assign n31588 = n1225 & ~n31587 ;
  assign n31589 = ( n6168 & n6181 ) | ( n6168 & n10094 ) | ( n6181 & n10094 ) ;
  assign n31590 = n31589 ^ n29215 ^ n1476 ;
  assign n31591 = ( n1675 & ~n6423 ) | ( n1675 & n11533 ) | ( ~n6423 & n11533 ) ;
  assign n31592 = ( n14928 & n16871 ) | ( n14928 & ~n31591 ) | ( n16871 & ~n31591 ) ;
  assign n31593 = n13651 ^ n5548 ^ 1'b0 ;
  assign n31594 = ~n21132 & n31593 ;
  assign n31595 = ( x84 & n7839 ) | ( x84 & ~n8901 ) | ( n7839 & ~n8901 ) ;
  assign n31596 = ( n6323 & n14236 ) | ( n6323 & ~n31595 ) | ( n14236 & ~n31595 ) ;
  assign n31597 = n31596 ^ n7031 ^ 1'b0 ;
  assign n31598 = ( n17379 & n24943 ) | ( n17379 & ~n31597 ) | ( n24943 & ~n31597 ) ;
  assign n31599 = ( n15410 & n31594 ) | ( n15410 & n31598 ) | ( n31594 & n31598 ) ;
  assign n31600 = n2059 | n31599 ;
  assign n31601 = ( ~n7216 & n10701 ) | ( ~n7216 & n31600 ) | ( n10701 & n31600 ) ;
  assign n31602 = n1760 & n3989 ;
  assign n31603 = ~n12740 & n31602 ;
  assign n31604 = n31603 ^ n20655 ^ n11627 ;
  assign n31605 = ( n6265 & n7218 ) | ( n6265 & n31604 ) | ( n7218 & n31604 ) ;
  assign n31606 = ( ~n18909 & n20579 ) | ( ~n18909 & n31605 ) | ( n20579 & n31605 ) ;
  assign n31607 = n8059 ^ n7062 ^ 1'b0 ;
  assign n31608 = ~n6956 & n12237 ;
  assign n31609 = n31608 ^ n16435 ^ 1'b0 ;
  assign n31610 = n20733 ^ n10742 ^ 1'b0 ;
  assign n31611 = n2003 & ~n31610 ;
  assign n31612 = ( n15434 & ~n16053 ) | ( n15434 & n16198 ) | ( ~n16053 & n16198 ) ;
  assign n31613 = ( n3515 & ~n10577 ) | ( n3515 & n11529 ) | ( ~n10577 & n11529 ) ;
  assign n31614 = n8309 & ~n31613 ;
  assign n31615 = n17973 ^ n5909 ^ n2671 ;
  assign n31616 = ( n7258 & n31614 ) | ( n7258 & n31615 ) | ( n31614 & n31615 ) ;
  assign n31617 = n13374 ^ n5121 ^ 1'b0 ;
  assign n31618 = n3569 | n4638 ;
  assign n31619 = n16232 ^ n12798 ^ n6787 ;
  assign n31620 = ( n5513 & n12163 ) | ( n5513 & n31619 ) | ( n12163 & n31619 ) ;
  assign n31621 = ( n11494 & n31618 ) | ( n11494 & ~n31620 ) | ( n31618 & ~n31620 ) ;
  assign n31622 = n18151 ^ n10072 ^ 1'b0 ;
  assign n31623 = n19944 | n31622 ;
  assign n31624 = n13937 ^ n13002 ^ n10551 ;
  assign n31625 = n31624 ^ n6520 ^ n4078 ;
  assign n31626 = n8067 | n31625 ;
  assign n31627 = ( n3810 & n31623 ) | ( n3810 & n31626 ) | ( n31623 & n31626 ) ;
  assign n31628 = ~n7859 & n18672 ;
  assign n31629 = n8442 & ~n11335 ;
  assign n31630 = n26231 | n31629 ;
  assign n31631 = n21048 | n31630 ;
  assign n31632 = n26472 ^ n6599 ^ 1'b0 ;
  assign n31633 = n4598 & ~n31632 ;
  assign n31634 = n2879 & n4991 ;
  assign n31635 = ~n27193 & n31634 ;
  assign n31636 = n11448 & n31635 ;
  assign n31638 = ~n2764 & n6479 ;
  assign n31637 = n28499 ^ n27140 ^ n23140 ;
  assign n31639 = n31638 ^ n31637 ^ n31624 ;
  assign n31640 = x162 & ~n14821 ;
  assign n31641 = n17800 & n31640 ;
  assign n31642 = n27784 ^ n4358 ^ n3827 ;
  assign n31643 = n4390 | n13746 ;
  assign n31644 = n31642 | n31643 ;
  assign n31645 = x220 & n23583 ;
  assign n31646 = ~n31644 & n31645 ;
  assign n31647 = n2624 & n8616 ;
  assign n31648 = ( n22244 & n31340 ) | ( n22244 & n31647 ) | ( n31340 & n31647 ) ;
  assign n31649 = n13801 & n20882 ;
  assign n31650 = n5643 & n16785 ;
  assign n31651 = ~n31649 & n31650 ;
  assign n31652 = ( n17211 & n31576 ) | ( n17211 & ~n31651 ) | ( n31576 & ~n31651 ) ;
  assign n31653 = n23843 ^ n14973 ^ n1822 ;
  assign n31655 = n18549 ^ n10795 ^ 1'b0 ;
  assign n31656 = ( ~n1829 & n14112 ) | ( ~n1829 & n31655 ) | ( n14112 & n31655 ) ;
  assign n31654 = n29966 ^ n15589 ^ 1'b0 ;
  assign n31657 = n31656 ^ n31654 ^ n4649 ;
  assign n31658 = ( n2662 & n15020 ) | ( n2662 & ~n31657 ) | ( n15020 & ~n31657 ) ;
  assign n31659 = n31658 ^ n5195 ^ 1'b0 ;
  assign n31660 = n27700 ^ n26558 ^ n670 ;
  assign n31662 = n2943 ^ n1644 ^ 1'b0 ;
  assign n31663 = ~n4313 & n31662 ;
  assign n31661 = n13960 ^ n2288 ^ n1669 ;
  assign n31664 = n31663 ^ n31661 ^ n23244 ;
  assign n31665 = n5474 & ~n25779 ;
  assign n31666 = n23152 & n31665 ;
  assign n31667 = n3997 & n7091 ;
  assign n31668 = n31667 ^ n5090 ^ 1'b0 ;
  assign n31669 = n394 | n9167 ;
  assign n31670 = n623 & n31669 ;
  assign n31671 = ~n31668 & n31670 ;
  assign n31672 = n21298 | n26780 ;
  assign n31673 = n5944 & n31267 ;
  assign n31674 = n22680 ^ n13523 ^ n2930 ;
  assign n31675 = n31674 ^ n17466 ^ 1'b0 ;
  assign n31676 = ( n6695 & n22439 ) | ( n6695 & ~n31675 ) | ( n22439 & ~n31675 ) ;
  assign n31677 = n26826 ^ n21810 ^ n2850 ;
  assign n31678 = ( n3568 & ~n12455 ) | ( n3568 & n19167 ) | ( ~n12455 & n19167 ) ;
  assign n31680 = n21950 ^ n14088 ^ n9832 ;
  assign n31679 = x234 & n28397 ;
  assign n31681 = n31680 ^ n31679 ^ 1'b0 ;
  assign n31682 = n9817 & ~n27938 ;
  assign n31683 = ~n475 & n31682 ;
  assign n31684 = n11397 & n31683 ;
  assign n31685 = n26950 & n31684 ;
  assign n31686 = n25672 ^ n20516 ^ n5411 ;
  assign n31687 = n12046 & ~n14941 ;
  assign n31688 = n31687 ^ n4275 ^ 1'b0 ;
  assign n31689 = ( n19674 & n21851 ) | ( n19674 & n31688 ) | ( n21851 & n31688 ) ;
  assign n31690 = ( n6714 & ~n11035 ) | ( n6714 & n26621 ) | ( ~n11035 & n26621 ) ;
  assign n31691 = n11255 ^ n5759 ^ 1'b0 ;
  assign n31692 = ( n2638 & ~n31690 ) | ( n2638 & n31691 ) | ( ~n31690 & n31691 ) ;
  assign n31693 = n17553 ^ n16862 ^ n5593 ;
  assign n31694 = n31693 ^ n25247 ^ n16341 ;
  assign n31695 = n25870 ^ n15055 ^ n3956 ;
  assign n31696 = n31695 ^ n26074 ^ n8539 ;
  assign n31699 = ~n1549 & n16691 ;
  assign n31700 = n31699 ^ n15472 ^ 1'b0 ;
  assign n31701 = n8254 & n31700 ;
  assign n31697 = n23485 ^ n2426 ^ 1'b0 ;
  assign n31698 = n25626 & n31697 ;
  assign n31702 = n31701 ^ n31698 ^ n14161 ;
  assign n31703 = n16844 ^ n12017 ^ n6671 ;
  assign n31704 = n22708 ^ n17879 ^ 1'b0 ;
  assign n31705 = n17635 & ~n31704 ;
  assign n31706 = ( n10993 & n31703 ) | ( n10993 & ~n31705 ) | ( n31703 & ~n31705 ) ;
  assign n31707 = n8956 ^ n891 ^ 1'b0 ;
  assign n31708 = n22825 & n31707 ;
  assign n31709 = n4070 & ~n17465 ;
  assign n31710 = n4741 & n31709 ;
  assign n31711 = n17400 | n31710 ;
  assign n31712 = x196 & n16883 ;
  assign n31713 = n31712 ^ n22522 ^ 1'b0 ;
  assign n31714 = n20478 ^ n12275 ^ 1'b0 ;
  assign n31715 = n7999 | n31714 ;
  assign n31716 = n1428 | n4763 ;
  assign n31717 = n31716 ^ n545 ^ 1'b0 ;
  assign n31718 = n22061 ^ n17396 ^ n2785 ;
  assign n31719 = n31718 ^ n7693 ^ 1'b0 ;
  assign n31720 = n10786 | n17466 ;
  assign n31721 = ( n10177 & n26702 ) | ( n10177 & ~n28443 ) | ( n26702 & ~n28443 ) ;
  assign n31722 = n17706 ^ n2882 ^ 1'b0 ;
  assign n31723 = n7335 & ~n26939 ;
  assign n31724 = n12219 ^ n11209 ^ n2920 ;
  assign n31725 = ( n7386 & n19425 ) | ( n7386 & n31724 ) | ( n19425 & n31724 ) ;
  assign n31726 = ( ~n7325 & n15576 ) | ( ~n7325 & n31725 ) | ( n15576 & n31725 ) ;
  assign n31727 = n31726 ^ n27977 ^ n4001 ;
  assign n31728 = ~n4834 & n23675 ;
  assign n31729 = n31728 ^ n25348 ^ 1'b0 ;
  assign n31730 = n15723 | n31729 ;
  assign n31731 = n5910 & ~n31730 ;
  assign n31732 = n31731 ^ n25349 ^ 1'b0 ;
  assign n31733 = n5351 | n12083 ;
  assign n31734 = n8657 & ~n31733 ;
  assign n31735 = n8656 ^ n5456 ^ 1'b0 ;
  assign n31736 = n31734 | n31735 ;
  assign n31737 = ( n991 & n13483 ) | ( n991 & n19754 ) | ( n13483 & n19754 ) ;
  assign n31738 = n31737 ^ n29003 ^ 1'b0 ;
  assign n31739 = ( n3648 & ~n12587 ) | ( n3648 & n25589 ) | ( ~n12587 & n25589 ) ;
  assign n31740 = n31739 ^ n13199 ^ n500 ;
  assign n31741 = ( ~n2794 & n10989 ) | ( ~n2794 & n31740 ) | ( n10989 & n31740 ) ;
  assign n31742 = n31741 ^ n6863 ^ 1'b0 ;
  assign n31743 = n28185 & ~n31742 ;
  assign n31744 = n9512 & ~n15323 ;
  assign n31745 = n27888 ^ n19183 ^ n8221 ;
  assign n31746 = n23469 ^ n8247 ^ n7247 ;
  assign n31747 = ~n2910 & n7714 ;
  assign n31748 = n31747 ^ n2208 ^ 1'b0 ;
  assign n31749 = n30785 ^ n19880 ^ 1'b0 ;
  assign n31750 = n31748 & ~n31749 ;
  assign n31751 = n19478 ^ n326 ^ 1'b0 ;
  assign n31752 = n31750 & ~n31751 ;
  assign n31753 = n29891 ^ n21005 ^ n13379 ;
  assign n31754 = n31753 ^ n17427 ^ 1'b0 ;
  assign n31756 = n585 | n9280 ;
  assign n31757 = n6430 ^ n5441 ^ 1'b0 ;
  assign n31758 = n31756 & n31757 ;
  assign n31755 = n22323 ^ n20964 ^ n10418 ;
  assign n31759 = n31758 ^ n31755 ^ n21063 ;
  assign n31760 = n9921 ^ n1104 ^ 1'b0 ;
  assign n31761 = n7652 | n31760 ;
  assign n31762 = n31761 ^ n12148 ^ 1'b0 ;
  assign n31763 = n8985 | n16642 ;
  assign n31764 = ( n2560 & ~n3632 ) | ( n2560 & n12185 ) | ( ~n3632 & n12185 ) ;
  assign n31765 = n7485 | n10021 ;
  assign n31766 = n28610 & ~n31765 ;
  assign n31767 = ( n22050 & n31764 ) | ( n22050 & n31766 ) | ( n31764 & n31766 ) ;
  assign n31768 = n9475 | n31767 ;
  assign n31769 = n29711 | n31768 ;
  assign n31770 = n31769 ^ n27259 ^ n8435 ;
  assign n31771 = n30380 ^ n27862 ^ 1'b0 ;
  assign n31772 = n12525 ^ n3247 ^ 1'b0 ;
  assign n31773 = n22437 & ~n31772 ;
  assign n31774 = n11326 ^ n10642 ^ 1'b0 ;
  assign n31775 = ~n8637 & n31774 ;
  assign n31776 = n11172 ^ n9623 ^ 1'b0 ;
  assign n31777 = ~n7113 & n31776 ;
  assign n31778 = ( n7152 & n9319 ) | ( n7152 & n31777 ) | ( n9319 & n31777 ) ;
  assign n31779 = n1271 & ~n16329 ;
  assign n31780 = n31779 ^ n10784 ^ 1'b0 ;
  assign n31781 = n1465 & ~n31780 ;
  assign n31782 = n31781 ^ n18798 ^ 1'b0 ;
  assign n31783 = n31778 & n31782 ;
  assign n31785 = n25610 ^ n4611 ^ n558 ;
  assign n31784 = n2040 & ~n6645 ;
  assign n31786 = n31785 ^ n31784 ^ n6783 ;
  assign n31787 = ~n3080 & n24375 ;
  assign n31788 = n31787 ^ n14065 ^ 1'b0 ;
  assign n31789 = n31786 | n31788 ;
  assign n31790 = n30649 ^ n23894 ^ 1'b0 ;
  assign n31791 = n31790 ^ n24650 ^ n6269 ;
  assign n31792 = n15276 & ~n24075 ;
  assign n31793 = n5760 & n31792 ;
  assign n31794 = ( ~n3933 & n11266 ) | ( ~n3933 & n31793 ) | ( n11266 & n31793 ) ;
  assign n31795 = n5378 ^ n2498 ^ 1'b0 ;
  assign n31796 = ~n18421 & n24797 ;
  assign n31797 = n31796 ^ n3003 ^ 1'b0 ;
  assign n31798 = n18883 ^ n17817 ^ n12832 ;
  assign n31799 = n30203 ^ n22325 ^ n4682 ;
  assign n31800 = ( n8179 & ~n19163 ) | ( n8179 & n22381 ) | ( ~n19163 & n22381 ) ;
  assign n31801 = n18278 ^ n13988 ^ 1'b0 ;
  assign n31802 = n6711 & ~n31801 ;
  assign n31803 = n31800 & n31802 ;
  assign n31804 = n31799 & n31803 ;
  assign n31805 = n28005 ^ n23649 ^ n10215 ;
  assign n31806 = ~n3563 & n5549 ;
  assign n31807 = n31806 ^ n8562 ^ 1'b0 ;
  assign n31808 = n31807 ^ n29632 ^ n5489 ;
  assign n31809 = ( n9405 & ~n14951 ) | ( n9405 & n25769 ) | ( ~n14951 & n25769 ) ;
  assign n31810 = ( n3301 & n16097 ) | ( n3301 & n17147 ) | ( n16097 & n17147 ) ;
  assign n31811 = n31810 ^ n16567 ^ n4192 ;
  assign n31812 = ( n3430 & ~n4494 ) | ( n3430 & n16652 ) | ( ~n4494 & n16652 ) ;
  assign n31813 = n5567 | n31812 ;
  assign n31814 = n31811 & ~n31813 ;
  assign n31815 = n12677 ^ n10111 ^ 1'b0 ;
  assign n31816 = n31815 ^ n30814 ^ n12861 ;
  assign n31817 = n5468 & ~n31816 ;
  assign n31818 = n2991 | n17261 ;
  assign n31819 = n31818 ^ n1884 ^ 1'b0 ;
  assign n31820 = n4030 & ~n5271 ;
  assign n31821 = n31820 ^ n15089 ^ 1'b0 ;
  assign n31822 = n7800 & ~n31821 ;
  assign n31823 = ~n14721 & n31822 ;
  assign n31824 = n31823 ^ n15144 ^ 1'b0 ;
  assign n31825 = n8857 & n31824 ;
  assign n31826 = n9161 ^ n650 ^ 1'b0 ;
  assign n31827 = n31826 ^ n28078 ^ n25119 ;
  assign n31828 = n6219 & ~n11910 ;
  assign n31829 = n31827 & n31828 ;
  assign n31831 = n17914 & n25448 ;
  assign n31832 = n31831 ^ n10597 ^ 1'b0 ;
  assign n31830 = n9781 & n20052 ;
  assign n31833 = n31832 ^ n31830 ^ 1'b0 ;
  assign n31834 = ~n5033 & n6471 ;
  assign n31835 = n31834 ^ n9180 ^ n3678 ;
  assign n31836 = n31835 ^ n15442 ^ 1'b0 ;
  assign n31837 = ( n11185 & ~n12385 ) | ( n11185 & n21986 ) | ( ~n12385 & n21986 ) ;
  assign n31838 = n31252 ^ n10765 ^ n3879 ;
  assign n31839 = n26471 ^ n9246 ^ 1'b0 ;
  assign n31840 = n21814 | n31839 ;
  assign n31841 = n24771 ^ n4899 ^ 1'b0 ;
  assign n31842 = n23364 & ~n31841 ;
  assign n31849 = n12757 ^ n12750 ^ n11789 ;
  assign n31843 = n15087 ^ n5317 ^ n652 ;
  assign n31844 = ( n3358 & n10055 ) | ( n3358 & n31843 ) | ( n10055 & n31843 ) ;
  assign n31845 = n16724 & ~n31844 ;
  assign n31846 = n31845 ^ n15167 ^ 1'b0 ;
  assign n31847 = n9626 | n17759 ;
  assign n31848 = ( n14611 & ~n31846 ) | ( n14611 & n31847 ) | ( ~n31846 & n31847 ) ;
  assign n31850 = n31849 ^ n31848 ^ n7746 ;
  assign n31851 = ( n3335 & n10885 ) | ( n3335 & n29383 ) | ( n10885 & n29383 ) ;
  assign n31852 = n7712 & ~n20892 ;
  assign n31853 = ~n18844 & n31852 ;
  assign n31854 = n31853 ^ n14540 ^ n7809 ;
  assign n31855 = n23851 ^ n15544 ^ 1'b0 ;
  assign n31856 = n7541 & n31855 ;
  assign n31857 = n23430 ^ n18428 ^ n17757 ;
  assign n31858 = n31857 ^ n15078 ^ 1'b0 ;
  assign n31859 = n21531 & n31858 ;
  assign n31861 = n29155 ^ n6299 ^ 1'b0 ;
  assign n31860 = ( ~n405 & n3670 ) | ( ~n405 & n8053 ) | ( n3670 & n8053 ) ;
  assign n31862 = n31861 ^ n31860 ^ n13066 ;
  assign n31863 = n3377 & n8199 ;
  assign n31864 = n31863 ^ n27281 ^ 1'b0 ;
  assign n31865 = n6589 & n29378 ;
  assign n31866 = n31865 ^ n11427 ^ 1'b0 ;
  assign n31867 = n29320 & n31866 ;
  assign n31868 = ~n31864 & n31867 ;
  assign n31869 = n5385 | n5482 ;
  assign n31870 = n7924 ^ n3285 ^ 1'b0 ;
  assign n31871 = n13608 | n29285 ;
  assign n31872 = n31870 | n31871 ;
  assign n31873 = n17606 ^ n3997 ^ 1'b0 ;
  assign n31874 = n31872 & ~n31873 ;
  assign n31875 = ( n1351 & ~n31869 ) | ( n1351 & n31874 ) | ( ~n31869 & n31874 ) ;
  assign n31876 = ( n5662 & n5682 ) | ( n5662 & ~n13731 ) | ( n5682 & ~n13731 ) ;
  assign n31877 = n995 & ~n31876 ;
  assign n31878 = n27727 ^ n17905 ^ n15200 ;
  assign n31879 = n4541 & ~n12797 ;
  assign n31880 = ( ~n7127 & n10821 ) | ( ~n7127 & n31879 ) | ( n10821 & n31879 ) ;
  assign n31881 = ( ~n490 & n31878 ) | ( ~n490 & n31880 ) | ( n31878 & n31880 ) ;
  assign n31882 = n16961 & ~n26000 ;
  assign n31883 = n9418 ^ n499 ^ 1'b0 ;
  assign n31884 = n31883 ^ n9206 ^ x95 ;
  assign n31885 = x77 & n10497 ;
  assign n31886 = n31884 & n31885 ;
  assign n31887 = n5690 ^ n2528 ^ n1545 ;
  assign n31890 = n1091 | n19823 ;
  assign n31888 = ( n2145 & ~n3217 ) | ( n2145 & n9128 ) | ( ~n3217 & n9128 ) ;
  assign n31889 = ( n25799 & n26007 ) | ( n25799 & n31888 ) | ( n26007 & n31888 ) ;
  assign n31891 = n31890 ^ n31889 ^ 1'b0 ;
  assign n31892 = ( ~n4682 & n31887 ) | ( ~n4682 & n31891 ) | ( n31887 & n31891 ) ;
  assign n31893 = n31892 ^ n19564 ^ n6196 ;
  assign n31894 = n31633 ^ n11438 ^ n9380 ;
  assign n31895 = ( n3659 & ~n6483 ) | ( n3659 & n7824 ) | ( ~n6483 & n7824 ) ;
  assign n31896 = ( n3984 & n21366 ) | ( n3984 & ~n31895 ) | ( n21366 & ~n31895 ) ;
  assign n31897 = n21546 | n31896 ;
  assign n31899 = n28174 ^ n14854 ^ n13211 ;
  assign n31898 = n9804 & n19527 ;
  assign n31900 = n31899 ^ n31898 ^ 1'b0 ;
  assign n31901 = n31900 ^ n2506 ^ 1'b0 ;
  assign n31902 = n23267 ^ n17613 ^ n14153 ;
  assign n31903 = n2333 & n31902 ;
  assign n31904 = n31903 ^ n1014 ^ 1'b0 ;
  assign n31905 = n12538 & ~n31904 ;
  assign n31906 = n21694 ^ n7483 ^ 1'b0 ;
  assign n31907 = n1478 & n31906 ;
  assign n31908 = ~n1133 & n31907 ;
  assign n31909 = n12899 & n31908 ;
  assign n31910 = n4671 & n18697 ;
  assign n31911 = n11395 ^ n8947 ^ 1'b0 ;
  assign n31913 = ( n3015 & n7091 ) | ( n3015 & n10596 ) | ( n7091 & n10596 ) ;
  assign n31912 = ~n3117 & n29842 ;
  assign n31914 = n31913 ^ n31912 ^ n586 ;
  assign n31915 = ~n22675 & n22710 ;
  assign n31917 = n7565 | n13059 ;
  assign n31918 = n11048 | n31917 ;
  assign n31916 = n18241 & n26784 ;
  assign n31919 = n31918 ^ n31916 ^ 1'b0 ;
  assign n31920 = n31919 ^ n26760 ^ n5638 ;
  assign n31921 = n14813 & n17067 ;
  assign n31922 = n31921 ^ n6861 ^ 1'b0 ;
  assign n31923 = ( n4523 & ~n10381 ) | ( n4523 & n31922 ) | ( ~n10381 & n31922 ) ;
  assign n31924 = ( n3490 & ~n10497 ) | ( n3490 & n15560 ) | ( ~n10497 & n15560 ) ;
  assign n31925 = ( n24928 & n31923 ) | ( n24928 & n31924 ) | ( n31923 & n31924 ) ;
  assign n31926 = n26887 ^ n16334 ^ 1'b0 ;
  assign n31927 = n9009 & ~n19879 ;
  assign n31928 = n15479 & n31927 ;
  assign n31929 = ( ~n4421 & n16469 ) | ( ~n4421 & n31928 ) | ( n16469 & n31928 ) ;
  assign n31930 = n28211 & ~n30795 ;
  assign n31931 = n31929 & n31930 ;
  assign n31932 = n3529 & ~n10669 ;
  assign n31933 = n31932 ^ n24067 ^ n20285 ;
  assign n31934 = ( n933 & n7092 ) | ( n933 & n29168 ) | ( n7092 & n29168 ) ;
  assign n31935 = ( n3322 & n19895 ) | ( n3322 & n31934 ) | ( n19895 & n31934 ) ;
  assign n31937 = n21270 ^ n15567 ^ n14073 ;
  assign n31936 = n18840 | n29600 ;
  assign n31938 = n31937 ^ n31936 ^ 1'b0 ;
  assign n31939 = ( n14942 & n31935 ) | ( n14942 & ~n31938 ) | ( n31935 & ~n31938 ) ;
  assign n31940 = n31248 ^ n20964 ^ x147 ;
  assign n31941 = ( n933 & n6367 ) | ( n933 & n11655 ) | ( n6367 & n11655 ) ;
  assign n31942 = n31941 ^ n22188 ^ n634 ;
  assign n31943 = n31942 ^ n9188 ^ 1'b0 ;
  assign n31944 = n28964 ^ n20113 ^ 1'b0 ;
  assign n31945 = ~n13084 & n31944 ;
  assign n31946 = n31945 ^ n26372 ^ n19157 ;
  assign n31947 = n11351 ^ n636 ^ 1'b0 ;
  assign n31948 = ~n31946 & n31947 ;
  assign n31949 = n16422 ^ n12108 ^ n10820 ;
  assign n31950 = n4139 ^ n3813 ^ n2097 ;
  assign n31951 = n28592 ^ n19741 ^ 1'b0 ;
  assign n31952 = n31950 & n31951 ;
  assign n31953 = ( n3233 & n8147 ) | ( n3233 & ~n31952 ) | ( n8147 & ~n31952 ) ;
  assign n31954 = n31064 ^ n13274 ^ n4520 ;
  assign n31955 = ~n463 & n4471 ;
  assign n31963 = n18564 ^ n16160 ^ n15316 ;
  assign n31956 = n30406 ^ n9420 ^ 1'b0 ;
  assign n31957 = ( n8964 & n21650 ) | ( n8964 & n31956 ) | ( n21650 & n31956 ) ;
  assign n31958 = ~n5771 & n9684 ;
  assign n31959 = ~n31957 & n31958 ;
  assign n31960 = n31959 ^ n11270 ^ 1'b0 ;
  assign n31961 = n22483 & ~n31960 ;
  assign n31962 = n31961 ^ n1189 ^ 1'b0 ;
  assign n31964 = n31963 ^ n31962 ^ n22822 ;
  assign n31965 = n13848 & ~n15402 ;
  assign n31966 = ( n7778 & ~n27288 ) | ( n7778 & n31965 ) | ( ~n27288 & n31965 ) ;
  assign n31967 = n19509 ^ n4778 ^ 1'b0 ;
  assign n31968 = n31966 & ~n31967 ;
  assign n31969 = n14577 & n23724 ;
  assign n31970 = n17680 ^ n10800 ^ n5102 ;
  assign n31971 = ( n4404 & n30183 ) | ( n4404 & n31970 ) | ( n30183 & n31970 ) ;
  assign n31972 = n9819 ^ n8601 ^ n4200 ;
  assign n31973 = ( n8804 & n26046 ) | ( n8804 & ~n31972 ) | ( n26046 & ~n31972 ) ;
  assign n31974 = ~n2482 & n5427 ;
  assign n31975 = n12329 & n31974 ;
  assign n31976 = n3310 ^ n1528 ^ 1'b0 ;
  assign n31977 = n31976 ^ n15659 ^ n12723 ;
  assign n31978 = n31975 & ~n31977 ;
  assign n31979 = n31978 ^ n19084 ^ n1713 ;
  assign n31980 = n2250 & n20146 ;
  assign n31981 = n31980 ^ n19738 ^ n9185 ;
  assign n31982 = ( ~n2427 & n4412 ) | ( ~n2427 & n24008 ) | ( n4412 & n24008 ) ;
  assign n31983 = n31982 ^ n12514 ^ n10787 ;
  assign n31984 = n3991 & ~n31983 ;
  assign n31985 = ( ~n2017 & n25068 ) | ( ~n2017 & n31984 ) | ( n25068 & n31984 ) ;
  assign n31986 = ~n8775 & n31985 ;
  assign n31987 = n7379 & n25260 ;
  assign n31988 = n31987 ^ n29038 ^ 1'b0 ;
  assign n31989 = n24578 ^ n14537 ^ 1'b0 ;
  assign n31990 = n6169 | n21033 ;
  assign n31991 = n31990 ^ n11801 ^ 1'b0 ;
  assign n31992 = n6771 | n14053 ;
  assign n31993 = ( n11595 & n20399 ) | ( n11595 & ~n31992 ) | ( n20399 & ~n31992 ) ;
  assign n31994 = ~n9046 & n31993 ;
  assign n31995 = n31994 ^ n1198 ^ 1'b0 ;
  assign n31996 = ( n9048 & n31991 ) | ( n9048 & ~n31995 ) | ( n31991 & ~n31995 ) ;
  assign n31997 = ( n11461 & n15225 ) | ( n11461 & n31996 ) | ( n15225 & n31996 ) ;
  assign n31998 = n12993 | n24268 ;
  assign n31999 = ( n596 & n20900 ) | ( n596 & ~n31998 ) | ( n20900 & ~n31998 ) ;
  assign n32000 = n19119 & ~n31999 ;
  assign n32001 = n1184 & ~n15024 ;
  assign n32002 = n32001 ^ n15464 ^ 1'b0 ;
  assign n32003 = ( n8781 & n19667 ) | ( n8781 & ~n32002 ) | ( n19667 & ~n32002 ) ;
  assign n32006 = n15318 ^ n3495 ^ 1'b0 ;
  assign n32007 = n1505 & n32006 ;
  assign n32008 = n32007 ^ n2993 ^ 1'b0 ;
  assign n32004 = ( n12060 & ~n13950 ) | ( n12060 & n19801 ) | ( ~n13950 & n19801 ) ;
  assign n32005 = n12078 & n32004 ;
  assign n32009 = n32008 ^ n32005 ^ 1'b0 ;
  assign n32010 = n16726 & ~n30665 ;
  assign n32019 = n6517 | n29169 ;
  assign n32020 = n32019 ^ n3475 ^ 1'b0 ;
  assign n32017 = n20227 ^ n16567 ^ n8466 ;
  assign n32018 = n32017 ^ n18011 ^ n17440 ;
  assign n32015 = ( ~n5517 & n13529 ) | ( ~n5517 & n24863 ) | ( n13529 & n24863 ) ;
  assign n32011 = n692 ^ n304 ^ 1'b0 ;
  assign n32012 = n21365 ^ n10773 ^ 1'b0 ;
  assign n32013 = n32012 ^ n18208 ^ 1'b0 ;
  assign n32014 = ~n32011 & n32013 ;
  assign n32016 = n32015 ^ n32014 ^ 1'b0 ;
  assign n32021 = n32020 ^ n32018 ^ n32016 ;
  assign n32022 = n2114 | n10045 ;
  assign n32023 = n32022 ^ n18578 ^ n1361 ;
  assign n32024 = n1713 ^ n1396 ^ n818 ;
  assign n32025 = n31798 ^ n15366 ^ 1'b0 ;
  assign n32026 = n32024 & n32025 ;
  assign n32027 = ( n13980 & n20454 ) | ( n13980 & ~n30937 ) | ( n20454 & ~n30937 ) ;
  assign n32028 = n13300 ^ n12291 ^ n2570 ;
  assign n32029 = ( n6562 & n30120 ) | ( n6562 & n32028 ) | ( n30120 & n32028 ) ;
  assign n32030 = n32029 ^ n28043 ^ 1'b0 ;
  assign n32031 = ~n32027 & n32030 ;
  assign n32032 = n15678 ^ n5708 ^ 1'b0 ;
  assign n32033 = ( n1046 & n21521 ) | ( n1046 & n32032 ) | ( n21521 & n32032 ) ;
  assign n32034 = ( ~n5522 & n20687 ) | ( ~n5522 & n26208 ) | ( n20687 & n26208 ) ;
  assign n32035 = n26488 ^ n12896 ^ 1'b0 ;
  assign n32036 = n28467 ^ n27159 ^ 1'b0 ;
  assign n32037 = n32035 & ~n32036 ;
  assign n32038 = n21287 & n32037 ;
  assign n32039 = n14129 & n32038 ;
  assign n32040 = n9357 & ~n27353 ;
  assign n32041 = n32040 ^ n13646 ^ n1622 ;
  assign n32043 = n18878 ^ n8904 ^ 1'b0 ;
  assign n32044 = ~n25131 & n32043 ;
  assign n32042 = n7471 ^ n799 ^ 1'b0 ;
  assign n32045 = n32044 ^ n32042 ^ n20926 ;
  assign n32046 = n11513 & n31907 ;
  assign n32047 = ~n4586 & n32046 ;
  assign n32048 = n26945 ^ n8205 ^ 1'b0 ;
  assign n32049 = n32048 ^ n8702 ^ 1'b0 ;
  assign n32050 = n32047 | n32049 ;
  assign n32051 = n15429 ^ n14928 ^ 1'b0 ;
  assign n32052 = ~n17191 & n32051 ;
  assign n32053 = n28993 & n32052 ;
  assign n32054 = n32053 ^ n12512 ^ 1'b0 ;
  assign n32055 = n7280 | n32054 ;
  assign n32056 = n32055 ^ n21355 ^ 1'b0 ;
  assign n32057 = ( n3823 & n26041 ) | ( n3823 & ~n27900 ) | ( n26041 & ~n27900 ) ;
  assign n32058 = n32057 ^ n17638 ^ n15770 ;
  assign n32059 = ( n10727 & ~n16530 ) | ( n10727 & n32058 ) | ( ~n16530 & n32058 ) ;
  assign n32060 = n4884 | n15433 ;
  assign n32061 = n32060 ^ n13859 ^ 1'b0 ;
  assign n32062 = ( ~n15850 & n32059 ) | ( ~n15850 & n32061 ) | ( n32059 & n32061 ) ;
  assign n32063 = ( n9564 & ~n10179 ) | ( n9564 & n15542 ) | ( ~n10179 & n15542 ) ;
  assign n32064 = n24965 ^ n18631 ^ 1'b0 ;
  assign n32065 = ~n22656 & n30623 ;
  assign n32066 = n32065 ^ n6902 ^ 1'b0 ;
  assign n32067 = n25524 | n32066 ;
  assign n32068 = ~x88 & n32067 ;
  assign n32069 = n26154 ^ n5156 ^ n1709 ;
  assign n32070 = x39 & ~n15423 ;
  assign n32071 = n32069 | n32070 ;
  assign n32072 = n32071 ^ n20807 ^ 1'b0 ;
  assign n32073 = n32072 ^ n5899 ^ 1'b0 ;
  assign n32074 = ~n11153 & n32073 ;
  assign n32075 = n31373 ^ n21683 ^ n18268 ;
  assign n32076 = ( n9390 & n11378 ) | ( n9390 & ~n28801 ) | ( n11378 & ~n28801 ) ;
  assign n32077 = n17523 & n23339 ;
  assign n32079 = ( n4255 & n10914 ) | ( n4255 & n16621 ) | ( n10914 & n16621 ) ;
  assign n32078 = ~n3459 & n22694 ;
  assign n32080 = n32079 ^ n32078 ^ n15332 ;
  assign n32081 = ( ~n4922 & n18157 ) | ( ~n4922 & n27074 ) | ( n18157 & n27074 ) ;
  assign n32082 = ~n13665 & n15053 ;
  assign n32083 = ~n32081 & n32082 ;
  assign n32084 = n8684 | n13980 ;
  assign n32085 = n15482 | n32084 ;
  assign n32087 = n7868 ^ n3235 ^ 1'b0 ;
  assign n32088 = n12432 & ~n32087 ;
  assign n32086 = n14192 & n15632 ;
  assign n32089 = n32088 ^ n32086 ^ 1'b0 ;
  assign n32092 = ~n962 & n8992 ;
  assign n32093 = n32092 ^ n7912 ^ 1'b0 ;
  assign n32090 = n8484 ^ n1089 ^ 1'b0 ;
  assign n32091 = n14548 | n32090 ;
  assign n32094 = n32093 ^ n32091 ^ 1'b0 ;
  assign n32095 = n32094 ^ n29641 ^ 1'b0 ;
  assign n32096 = ~n32089 & n32095 ;
  assign n32097 = n30667 ^ n8509 ^ 1'b0 ;
  assign n32098 = ~n7670 & n29956 ;
  assign n32099 = n14881 & ~n32098 ;
  assign n32100 = n32099 ^ n23633 ^ n13538 ;
  assign n32101 = ( n2667 & ~n3476 ) | ( n2667 & n24514 ) | ( ~n3476 & n24514 ) ;
  assign n32102 = n18506 | n32101 ;
  assign n32103 = ( n14900 & n15129 ) | ( n14900 & n28076 ) | ( n15129 & n28076 ) ;
  assign n32104 = n19801 ^ n7550 ^ n3081 ;
  assign n32105 = n32104 ^ n25496 ^ 1'b0 ;
  assign n32106 = ( n14728 & n32103 ) | ( n14728 & ~n32105 ) | ( n32103 & ~n32105 ) ;
  assign n32110 = n3252 | n15035 ;
  assign n32111 = n2885 | n32110 ;
  assign n32107 = n12513 & ~n15502 ;
  assign n32108 = ~n6731 & n32107 ;
  assign n32109 = n16470 & ~n32108 ;
  assign n32112 = n32111 ^ n32109 ^ n14985 ;
  assign n32113 = n15614 ^ n4990 ^ 1'b0 ;
  assign n32114 = n7220 & ~n14097 ;
  assign n32115 = n8803 & n32114 ;
  assign n32116 = n28246 ^ n21514 ^ n3142 ;
  assign n32117 = ( n358 & n9142 ) | ( n358 & n28427 ) | ( n9142 & n28427 ) ;
  assign n32118 = ( n2350 & n22133 ) | ( n2350 & ~n22412 ) | ( n22133 & ~n22412 ) ;
  assign n32119 = n29446 ^ n27381 ^ n15426 ;
  assign n32120 = ( x23 & n18487 ) | ( x23 & ~n25520 ) | ( n18487 & ~n25520 ) ;
  assign n32121 = n10093 & n15024 ;
  assign n32122 = n10374 | n32121 ;
  assign n32123 = n3184 | n32122 ;
  assign n32124 = n31822 ^ n8389 ^ 1'b0 ;
  assign n32125 = ~n25009 & n32124 ;
  assign n32126 = n19643 ^ n5057 ^ 1'b0 ;
  assign n32127 = n28507 | n32126 ;
  assign n32130 = n19568 ^ n9531 ^ n2162 ;
  assign n32128 = n18323 ^ n17413 ^ n11567 ;
  assign n32129 = n32128 ^ n23579 ^ n4208 ;
  assign n32131 = n32130 ^ n32129 ^ n11158 ;
  assign n32132 = n20709 ^ n6279 ^ 1'b0 ;
  assign n32133 = n4028 ^ n3234 ^ n286 ;
  assign n32134 = ( n7736 & n17853 ) | ( n7736 & ~n32133 ) | ( n17853 & ~n32133 ) ;
  assign n32135 = n16399 ^ n14142 ^ 1'b0 ;
  assign n32136 = ~n7534 & n32135 ;
  assign n32137 = ( ~n20433 & n21422 ) | ( ~n20433 & n22180 ) | ( n21422 & n22180 ) ;
  assign n32138 = ( n19639 & n32136 ) | ( n19639 & ~n32137 ) | ( n32136 & ~n32137 ) ;
  assign n32139 = n10076 & ~n32138 ;
  assign n32140 = n32134 & n32139 ;
  assign n32146 = n681 | n9461 ;
  assign n32147 = n32146 ^ n25691 ^ 1'b0 ;
  assign n32148 = n32147 ^ x100 ^ 1'b0 ;
  assign n32149 = n427 | n32148 ;
  assign n32144 = n22615 ^ n8127 ^ x230 ;
  assign n32142 = n7805 ^ n6563 ^ n473 ;
  assign n32143 = ( n5435 & n22773 ) | ( n5435 & n32142 ) | ( n22773 & n32142 ) ;
  assign n32145 = n32144 ^ n32143 ^ n4393 ;
  assign n32141 = n12515 ^ n11527 ^ n2878 ;
  assign n32150 = n32149 ^ n32145 ^ n32141 ;
  assign n32151 = n29850 ^ n22659 ^ n21766 ;
  assign n32152 = n30670 ^ n19077 ^ n10743 ;
  assign n32153 = ( n24213 & n28669 ) | ( n24213 & n32152 ) | ( n28669 & n32152 ) ;
  assign n32154 = ( n21217 & n26228 ) | ( n21217 & n32153 ) | ( n26228 & n32153 ) ;
  assign n32155 = n7980 ^ n5875 ^ n3007 ;
  assign n32156 = n32155 ^ n7036 ^ 1'b0 ;
  assign n32157 = ( ~n4490 & n5913 ) | ( ~n4490 & n32156 ) | ( n5913 & n32156 ) ;
  assign n32158 = n25803 ^ n19275 ^ 1'b0 ;
  assign n32159 = n21264 ^ n3548 ^ 1'b0 ;
  assign n32160 = n25594 ^ n15402 ^ 1'b0 ;
  assign n32161 = ( n2326 & n25599 ) | ( n2326 & ~n32160 ) | ( n25599 & ~n32160 ) ;
  assign n32162 = n287 & ~n922 ;
  assign n32163 = ~x204 & n32162 ;
  assign n32164 = ( n20001 & ~n25088 ) | ( n20001 & n32163 ) | ( ~n25088 & n32163 ) ;
  assign n32165 = n9064 | n18937 ;
  assign n32166 = n32165 ^ n25933 ^ 1'b0 ;
  assign n32167 = n505 & ~n7641 ;
  assign n32168 = n8452 ^ n3329 ^ 1'b0 ;
  assign n32169 = n32168 ^ n25214 ^ n10516 ;
  assign n32170 = n18002 | n32169 ;
  assign n32171 = n32170 ^ n16494 ^ 1'b0 ;
  assign n32172 = n32167 & n32171 ;
  assign n32173 = n32172 ^ n8145 ^ 1'b0 ;
  assign n32174 = ( n9946 & ~n22951 ) | ( n9946 & n26493 ) | ( ~n22951 & n26493 ) ;
  assign n32175 = ( n12429 & n17403 ) | ( n12429 & ~n18687 ) | ( n17403 & ~n18687 ) ;
  assign n32176 = n8278 & n20235 ;
  assign n32177 = ~x96 & n32176 ;
  assign n32178 = n32177 ^ n21731 ^ n9980 ;
  assign n32179 = n12024 ^ n6763 ^ n256 ;
  assign n32180 = n32179 ^ n14349 ^ 1'b0 ;
  assign n32181 = ( n3559 & n5341 ) | ( n3559 & n7789 ) | ( n5341 & n7789 ) ;
  assign n32182 = n17912 ^ n701 ^ 1'b0 ;
  assign n32183 = n22083 ^ x254 ^ 1'b0 ;
  assign n32184 = n32182 & ~n32183 ;
  assign n32185 = n32181 & n32184 ;
  assign n32186 = n32180 & n32185 ;
  assign n32187 = n7759 & ~n15824 ;
  assign n32188 = ~n26121 & n29334 ;
  assign n32189 = n805 | n25548 ;
  assign n32190 = n28097 & ~n32189 ;
  assign n32191 = n23373 ^ n15008 ^ 1'b0 ;
  assign n32194 = n6945 ^ n4564 ^ n2111 ;
  assign n32192 = n15427 ^ n10403 ^ 1'b0 ;
  assign n32193 = n3807 & ~n32192 ;
  assign n32195 = n32194 ^ n32193 ^ 1'b0 ;
  assign n32196 = n8684 & n29201 ;
  assign n32197 = n786 & ~n28900 ;
  assign n32198 = ~n1629 & n32197 ;
  assign n32199 = n2022 | n14506 ;
  assign n32200 = n21363 & ~n32199 ;
  assign n32201 = n7270 & ~n10569 ;
  assign n32202 = n32201 ^ n4951 ^ 1'b0 ;
  assign n32203 = n32200 | n32202 ;
  assign n32204 = n28081 ^ n27832 ^ n8510 ;
  assign n32205 = ( n1122 & ~n8633 ) | ( n1122 & n29663 ) | ( ~n8633 & n29663 ) ;
  assign n32206 = n32205 ^ n19982 ^ n14619 ;
  assign n32207 = n29104 ^ n16676 ^ n8294 ;
  assign n32208 = n32207 ^ n14370 ^ n10854 ;
  assign n32210 = n18442 ^ n13292 ^ 1'b0 ;
  assign n32211 = ~n12178 & n32210 ;
  assign n32209 = ~n6472 & n12064 ;
  assign n32212 = n32211 ^ n32209 ^ 1'b0 ;
  assign n32213 = n13578 & n30370 ;
  assign n32214 = n32213 ^ n22955 ^ 1'b0 ;
  assign n32215 = n14413 | n24436 ;
  assign n32216 = ( ~n740 & n960 ) | ( ~n740 & n6195 ) | ( n960 & n6195 ) ;
  assign n32217 = n21271 ^ n19742 ^ n10411 ;
  assign n32218 = n1302 | n27416 ;
  assign n32219 = ( n11065 & n32217 ) | ( n11065 & ~n32218 ) | ( n32217 & ~n32218 ) ;
  assign n32223 = n8331 ^ n702 ^ 1'b0 ;
  assign n32224 = ( ~n10073 & n13864 ) | ( ~n10073 & n32223 ) | ( n13864 & n32223 ) ;
  assign n32220 = n23896 ^ n14805 ^ n4381 ;
  assign n32221 = ( n4582 & ~n6005 ) | ( n4582 & n32220 ) | ( ~n6005 & n32220 ) ;
  assign n32222 = n32221 ^ n23116 ^ n5971 ;
  assign n32225 = n32224 ^ n32222 ^ n3829 ;
  assign n32231 = n25581 ^ n20636 ^ n11858 ;
  assign n32232 = n4716 & ~n32231 ;
  assign n32226 = n7144 & ~n8827 ;
  assign n32227 = n6532 ^ n4562 ^ n4440 ;
  assign n32228 = n11709 ^ n7221 ^ n2609 ;
  assign n32229 = ( n10801 & ~n32227 ) | ( n10801 & n32228 ) | ( ~n32227 & n32228 ) ;
  assign n32230 = n32226 & n32229 ;
  assign n32233 = n32232 ^ n32230 ^ 1'b0 ;
  assign n32234 = n28589 ^ n2808 ^ 1'b0 ;
  assign n32235 = n4905 & ~n16595 ;
  assign n32236 = n26284 | n28238 ;
  assign n32237 = n20395 ^ n6219 ^ 1'b0 ;
  assign n32238 = ~n6392 & n32237 ;
  assign n32239 = n32238 ^ n16275 ^ n10576 ;
  assign n32240 = ~n1803 & n1985 ;
  assign n32241 = n32240 ^ n7851 ^ n5904 ;
  assign n32244 = n10653 ^ n7638 ^ 1'b0 ;
  assign n32242 = n26595 ^ n14302 ^ 1'b0 ;
  assign n32243 = n21874 | n32242 ;
  assign n32245 = n32244 ^ n32243 ^ 1'b0 ;
  assign n32246 = n19892 ^ n12070 ^ 1'b0 ;
  assign n32247 = n15787 ^ n9581 ^ 1'b0 ;
  assign n32248 = n32247 ^ n18592 ^ n13813 ;
  assign n32249 = n15960 ^ n6055 ^ n2962 ;
  assign n32250 = ~n3004 & n5934 ;
  assign n32251 = ~n4533 & n32250 ;
  assign n32252 = n32251 ^ n13024 ^ n8552 ;
  assign n32253 = n9775 ^ n2198 ^ 1'b0 ;
  assign n32254 = n32253 ^ n11769 ^ 1'b0 ;
  assign n32255 = n20446 & ~n32254 ;
  assign n32256 = ( n3793 & n10124 ) | ( n3793 & ~n13914 ) | ( n10124 & ~n13914 ) ;
  assign n32257 = n16640 ^ n4899 ^ 1'b0 ;
  assign n32258 = n32256 & n32257 ;
  assign n32259 = ~n6068 & n32258 ;
  assign n32260 = n3586 | n15615 ;
  assign n32261 = n29515 ^ n22731 ^ n11123 ;
  assign n32262 = n21359 ^ n15360 ^ n7133 ;
  assign n32263 = ( n9959 & n25459 ) | ( n9959 & ~n32262 ) | ( n25459 & ~n32262 ) ;
  assign n32264 = n27510 ^ n25898 ^ 1'b0 ;
  assign n32265 = ~n32263 & n32264 ;
  assign n32266 = n32265 ^ n11428 ^ 1'b0 ;
  assign n32268 = ( n16078 & n16729 ) | ( n16078 & ~n20247 ) | ( n16729 & ~n20247 ) ;
  assign n32267 = n28512 ^ n8007 ^ 1'b0 ;
  assign n32269 = n32268 ^ n32267 ^ n14909 ;
  assign n32270 = ( n8890 & n12075 ) | ( n8890 & n30944 ) | ( n12075 & n30944 ) ;
  assign n32273 = n6677 & ~n30147 ;
  assign n32271 = ( n10112 & n13950 ) | ( n10112 & ~n15802 ) | ( n13950 & ~n15802 ) ;
  assign n32272 = n19528 | n32271 ;
  assign n32274 = n32273 ^ n32272 ^ 1'b0 ;
  assign n32275 = n29898 ^ n18430 ^ 1'b0 ;
  assign n32276 = n14767 | n32275 ;
  assign n32277 = ~n5038 & n32276 ;
  assign n32278 = n32277 ^ n8018 ^ 1'b0 ;
  assign n32280 = n6308 | n20711 ;
  assign n32281 = n32280 ^ n16703 ^ 1'b0 ;
  assign n32282 = n22325 ^ n10035 ^ 1'b0 ;
  assign n32283 = n533 | n32282 ;
  assign n32284 = n32283 ^ n17807 ^ 1'b0 ;
  assign n32285 = ~n32281 & n32284 ;
  assign n32279 = n3568 & n11411 ;
  assign n32286 = n32285 ^ n32279 ^ 1'b0 ;
  assign n32287 = n5717 | n5814 ;
  assign n32288 = n32287 ^ n2637 ^ 1'b0 ;
  assign n32289 = n32288 ^ n15453 ^ n735 ;
  assign n32290 = n5335 & n31330 ;
  assign n32291 = ( ~n1248 & n19315 ) | ( ~n1248 & n32290 ) | ( n19315 & n32290 ) ;
  assign n32292 = n2243 | n5645 ;
  assign n32293 = n2411 & ~n22247 ;
  assign n32294 = n32293 ^ n2163 ^ 1'b0 ;
  assign n32295 = ( ~n10090 & n17492 ) | ( ~n10090 & n32294 ) | ( n17492 & n32294 ) ;
  assign n32296 = n4724 | n21919 ;
  assign n32297 = n14149 & n32296 ;
  assign n32298 = n32295 & n32297 ;
  assign n32299 = n24979 ^ n23401 ^ n19905 ;
  assign n32300 = n32299 ^ n30852 ^ n8627 ;
  assign n32301 = n27148 ^ n17687 ^ n2565 ;
  assign n32302 = n23587 ^ n6095 ^ n343 ;
  assign n32303 = n693 & ~n14108 ;
  assign n32304 = n32303 ^ n5390 ^ 1'b0 ;
  assign n32305 = ( ~n18011 & n25772 ) | ( ~n18011 & n30608 ) | ( n25772 & n30608 ) ;
  assign n32306 = ( ~n32302 & n32304 ) | ( ~n32302 & n32305 ) | ( n32304 & n32305 ) ;
  assign n32307 = n21483 ^ n18961 ^ 1'b0 ;
  assign n32309 = n7912 ^ n7241 ^ 1'b0 ;
  assign n32308 = ~n4196 & n13473 ;
  assign n32310 = n32309 ^ n32308 ^ 1'b0 ;
  assign n32311 = n5469 | n13581 ;
  assign n32312 = n15984 | n32311 ;
  assign n32313 = n32312 ^ n25833 ^ 1'b0 ;
  assign n32314 = n16844 & ~n32313 ;
  assign n32315 = n15533 & n28398 ;
  assign n32316 = ~n32314 & n32315 ;
  assign n32317 = ( ~n3509 & n16295 ) | ( ~n3509 & n16825 ) | ( n16295 & n16825 ) ;
  assign n32318 = n14280 ^ n546 ^ n317 ;
  assign n32319 = x157 ^ x125 ^ 1'b0 ;
  assign n32320 = n32318 & n32319 ;
  assign n32321 = n32320 ^ n24436 ^ n19187 ;
  assign n32322 = n5978 ^ n1688 ^ 1'b0 ;
  assign n32323 = n32322 ^ n27049 ^ n8596 ;
  assign n32324 = n21885 ^ n13723 ^ 1'b0 ;
  assign n32325 = x229 & ~n1299 ;
  assign n32326 = ~n668 & n32325 ;
  assign n32327 = n3894 | n32326 ;
  assign n32328 = n20925 & ~n32327 ;
  assign n32329 = n27670 ^ n15244 ^ n8024 ;
  assign n32330 = ( n8893 & ~n9832 ) | ( n8893 & n32329 ) | ( ~n9832 & n32329 ) ;
  assign n32331 = n32330 ^ n1100 ^ 1'b0 ;
  assign n32332 = ~n10499 & n10916 ;
  assign n32333 = ~n18037 & n32332 ;
  assign n32334 = n9089 | n32333 ;
  assign n32335 = n32334 ^ n14749 ^ 1'b0 ;
  assign n32336 = ( ~n5686 & n17363 ) | ( ~n5686 & n32335 ) | ( n17363 & n32335 ) ;
  assign n32337 = n2602 & n7044 ;
  assign n32338 = n3992 & n32337 ;
  assign n32339 = n20557 & ~n32338 ;
  assign n32340 = ~n7513 & n32339 ;
  assign n32341 = ( n4489 & n10631 ) | ( n4489 & ~n16874 ) | ( n10631 & ~n16874 ) ;
  assign n32342 = n32341 ^ n32103 ^ n18892 ;
  assign n32345 = n22152 & ~n28812 ;
  assign n32343 = n13029 ^ n6982 ^ 1'b0 ;
  assign n32344 = n32083 | n32343 ;
  assign n32346 = n32345 ^ n32344 ^ 1'b0 ;
  assign n32348 = n14096 ^ n11357 ^ n2775 ;
  assign n32347 = n5368 | n24268 ;
  assign n32349 = n32348 ^ n32347 ^ 1'b0 ;
  assign n32350 = n14815 & ~n15263 ;
  assign n32351 = n13862 ^ n3799 ^ 1'b0 ;
  assign n32352 = n8137 & n32351 ;
  assign n32353 = n32352 ^ n23077 ^ 1'b0 ;
  assign n32354 = n32353 ^ n30886 ^ n15300 ;
  assign n32355 = ( n10749 & n32350 ) | ( n10749 & ~n32354 ) | ( n32350 & ~n32354 ) ;
  assign n32356 = ( n7474 & ~n11031 ) | ( n7474 & n21025 ) | ( ~n11031 & n21025 ) ;
  assign n32357 = n17900 & ~n20229 ;
  assign n32358 = n5500 & n18602 ;
  assign n32359 = n32358 ^ n15926 ^ 1'b0 ;
  assign n32360 = n6884 & ~n30719 ;
  assign n32361 = n32360 ^ n2651 ^ 1'b0 ;
  assign n32362 = n17393 ^ n16416 ^ n14033 ;
  assign n32363 = n32362 ^ n15270 ^ n6418 ;
  assign n32364 = n24318 ^ n22066 ^ 1'b0 ;
  assign n32365 = n9147 | n32364 ;
  assign n32366 = n6682 & ~n32365 ;
  assign n32367 = n21442 & ~n29424 ;
  assign n32368 = n27227 ^ n3229 ^ 1'b0 ;
  assign n32369 = ( ~n10702 & n25264 ) | ( ~n10702 & n31526 ) | ( n25264 & n31526 ) ;
  assign n32376 = n26681 ^ n25881 ^ n14728 ;
  assign n32370 = n18982 ^ n3503 ^ 1'b0 ;
  assign n32371 = x57 & n32370 ;
  assign n32372 = n32371 ^ n12812 ^ n6858 ;
  assign n32373 = n9747 & ~n32372 ;
  assign n32374 = n32373 ^ n6158 ^ 1'b0 ;
  assign n32375 = ( n11991 & n23995 ) | ( n11991 & n32374 ) | ( n23995 & n32374 ) ;
  assign n32377 = n32376 ^ n32375 ^ n15623 ;
  assign n32378 = ( n15877 & n16953 ) | ( n15877 & n30010 ) | ( n16953 & n30010 ) ;
  assign n32379 = n21503 ^ n15876 ^ 1'b0 ;
  assign n32380 = n17935 ^ n14399 ^ 1'b0 ;
  assign n32381 = n32380 ^ n5818 ^ n5098 ;
  assign n32382 = n6049 ^ n852 ^ 1'b0 ;
  assign n32383 = n6860 & ~n16238 ;
  assign n32384 = ~n32382 & n32383 ;
  assign n32385 = n26389 ^ n7923 ^ n4738 ;
  assign n32386 = n2512 & ~n32385 ;
  assign n32387 = ( x148 & n3673 ) | ( x148 & n15632 ) | ( n3673 & n15632 ) ;
  assign n32388 = n3004 ^ x64 ^ 1'b0 ;
  assign n32389 = n30438 | n32388 ;
  assign n32390 = n32389 ^ n14503 ^ n11757 ;
  assign n32391 = n4425 & n17134 ;
  assign n32392 = ( ~n5520 & n10432 ) | ( ~n5520 & n13672 ) | ( n10432 & n13672 ) ;
  assign n32393 = n32392 ^ n22631 ^ n13730 ;
  assign n32394 = n14757 ^ n7836 ^ 1'b0 ;
  assign n32395 = ~n32393 & n32394 ;
  assign n32396 = n32391 & n32395 ;
  assign n32397 = ( n3873 & ~n5081 ) | ( n3873 & n30662 ) | ( ~n5081 & n30662 ) ;
  assign n32398 = n7520 & ~n16939 ;
  assign n32399 = ~n1268 & n32398 ;
  assign n32400 = n21076 ^ n19499 ^ n12764 ;
  assign n32401 = n32400 ^ n21034 ^ 1'b0 ;
  assign n32402 = n16709 & ~n32401 ;
  assign n32403 = n2003 & n15549 ;
  assign n32404 = n32403 ^ n10823 ^ 1'b0 ;
  assign n32405 = n13385 ^ n12122 ^ n920 ;
  assign n32406 = n18150 ^ n3736 ^ 1'b0 ;
  assign n32407 = n32405 | n32406 ;
  assign n32408 = n2602 & ~n7588 ;
  assign n32409 = ~n7163 & n32408 ;
  assign n32410 = ( ~n28609 & n32407 ) | ( ~n28609 & n32409 ) | ( n32407 & n32409 ) ;
  assign n32411 = n1376 & ~n32410 ;
  assign n32412 = n32411 ^ n10300 ^ 1'b0 ;
  assign n32413 = n24593 ^ n5944 ^ n5764 ;
  assign n32414 = ( n10359 & ~n21497 ) | ( n10359 & n32413 ) | ( ~n21497 & n32413 ) ;
  assign n32415 = ( n12050 & n26283 ) | ( n12050 & n31997 ) | ( n26283 & n31997 ) ;
  assign n32416 = n2945 ^ n2799 ^ 1'b0 ;
  assign n32417 = n1122 | n19931 ;
  assign n32418 = n32417 ^ n10206 ^ n4007 ;
  assign n32419 = ~n851 & n9655 ;
  assign n32420 = n27721 ^ n22878 ^ 1'b0 ;
  assign n32421 = ( n2739 & n3047 ) | ( n2739 & ~n10681 ) | ( n3047 & ~n10681 ) ;
  assign n32422 = ( n14946 & n29487 ) | ( n14946 & n32421 ) | ( n29487 & n32421 ) ;
  assign n32423 = n4464 & n11935 ;
  assign n32424 = n32423 ^ n20918 ^ n18604 ;
  assign n32425 = ~n1825 & n8032 ;
  assign n32426 = ( ~n4150 & n19064 ) | ( ~n4150 & n32425 ) | ( n19064 & n32425 ) ;
  assign n32427 = n32426 ^ n22324 ^ n2110 ;
  assign n32428 = n20456 & ~n32427 ;
  assign n32431 = n19111 ^ n10685 ^ n5999 ;
  assign n32429 = n15866 | n21578 ;
  assign n32430 = n32429 ^ n12190 ^ 1'b0 ;
  assign n32432 = n32431 ^ n32430 ^ n17783 ;
  assign n32433 = n3069 & ~n4006 ;
  assign n32434 = n32432 & n32433 ;
  assign n32435 = n17599 ^ n4271 ^ n2914 ;
  assign n32436 = n24941 ^ n2426 ^ 1'b0 ;
  assign n32437 = ~n31760 & n32436 ;
  assign n32438 = ~n32435 & n32437 ;
  assign n32439 = n29689 ^ n16957 ^ 1'b0 ;
  assign n32440 = n8366 | n32439 ;
  assign n32441 = n23767 ^ n11414 ^ 1'b0 ;
  assign n32442 = ( n14125 & ~n23908 ) | ( n14125 & n29605 ) | ( ~n23908 & n29605 ) ;
  assign n32443 = n1765 & ~n7384 ;
  assign n32444 = n32443 ^ n4801 ^ 1'b0 ;
  assign n32445 = n15613 | n32444 ;
  assign n32446 = n20569 | n26935 ;
  assign n32447 = n4980 & n21750 ;
  assign n32448 = n32447 ^ n10272 ^ 1'b0 ;
  assign n32449 = n32448 ^ n25891 ^ n18902 ;
  assign n32450 = ( n32445 & n32446 ) | ( n32445 & n32449 ) | ( n32446 & n32449 ) ;
  assign n32451 = n7812 & ~n12630 ;
  assign n32452 = n9418 | n23009 ;
  assign n32453 = n32452 ^ x138 ^ 1'b0 ;
  assign n32454 = ( n3947 & n32451 ) | ( n3947 & n32453 ) | ( n32451 & n32453 ) ;
  assign n32458 = n12129 ^ n8655 ^ n6393 ;
  assign n32459 = n32458 ^ n18367 ^ n6420 ;
  assign n32455 = x42 & ~n2108 ;
  assign n32456 = n32455 ^ n2695 ^ 1'b0 ;
  assign n32457 = n31457 & n32456 ;
  assign n32460 = n32459 ^ n32457 ^ 1'b0 ;
  assign n32461 = ~n26479 & n32460 ;
  assign n32462 = n5556 & n32461 ;
  assign n32463 = n32249 ^ n16323 ^ 1'b0 ;
  assign n32464 = n3217 & ~n32463 ;
  assign n32465 = ~n17050 & n20845 ;
  assign n32466 = n32465 ^ x122 ^ 1'b0 ;
  assign n32467 = ~n10589 & n32466 ;
  assign n32468 = n13347 ^ n6274 ^ n3084 ;
  assign n32469 = n9576 & n21078 ;
  assign n32470 = ( n7946 & n9324 ) | ( n7946 & ~n32469 ) | ( n9324 & ~n32469 ) ;
  assign n32472 = n30671 ^ n27196 ^ n9096 ;
  assign n32471 = ~n19566 & n26987 ;
  assign n32473 = n32472 ^ n32471 ^ 1'b0 ;
  assign n32474 = n1823 & ~n2575 ;
  assign n32475 = n32474 ^ n10728 ^ 1'b0 ;
  assign n32476 = ~n3715 & n32475 ;
  assign n32477 = n18156 ^ n10929 ^ n8260 ;
  assign n32478 = n7632 ^ n6849 ^ 1'b0 ;
  assign n32479 = ~n17412 & n32478 ;
  assign n32480 = ( n14707 & n32477 ) | ( n14707 & n32479 ) | ( n32477 & n32479 ) ;
  assign n32481 = ( n11082 & n32476 ) | ( n11082 & ~n32480 ) | ( n32476 & ~n32480 ) ;
  assign n32482 = n2017 | n13168 ;
  assign n32483 = ~n20564 & n25650 ;
  assign n32484 = ( n14740 & n32482 ) | ( n14740 & ~n32483 ) | ( n32482 & ~n32483 ) ;
  assign n32485 = n21009 ^ n4917 ^ 1'b0 ;
  assign n32486 = ( n13381 & ~n24436 ) | ( n13381 & n31811 ) | ( ~n24436 & n31811 ) ;
  assign n32487 = n32486 ^ n14921 ^ 1'b0 ;
  assign n32488 = n10260 & n22129 ;
  assign n32489 = ~n26691 & n32488 ;
  assign n32490 = n29629 ^ n12508 ^ 1'b0 ;
  assign n32491 = ( n1465 & ~n19937 ) | ( n1465 & n32490 ) | ( ~n19937 & n32490 ) ;
  assign n32492 = n25296 ^ n16944 ^ n2798 ;
  assign n32493 = ~n9162 & n32492 ;
  assign n32494 = n32493 ^ n7163 ^ 1'b0 ;
  assign n32495 = n5723 | n13850 ;
  assign n32496 = n2374 & ~n32495 ;
  assign n32497 = n27158 ^ n11139 ^ 1'b0 ;
  assign n32498 = n25897 | n32497 ;
  assign n32499 = ( n22649 & n32496 ) | ( n22649 & n32498 ) | ( n32496 & n32498 ) ;
  assign n32500 = n32499 ^ n29407 ^ n1783 ;
  assign n32501 = ( n14590 & n16332 ) | ( n14590 & n18308 ) | ( n16332 & n18308 ) ;
  assign n32502 = n6993 & ~n8677 ;
  assign n32503 = n32502 ^ n1378 ^ 1'b0 ;
  assign n32504 = n32503 ^ n31361 ^ n27784 ;
  assign n32505 = n7739 | n21502 ;
  assign n32506 = n5884 & n32505 ;
  assign n32507 = ~n32504 & n32506 ;
  assign n32508 = n26276 ^ n4828 ^ 1'b0 ;
  assign n32511 = n13204 ^ n3172 ^ 1'b0 ;
  assign n32512 = n17051 | n32511 ;
  assign n32509 = n10930 & ~n20314 ;
  assign n32510 = n32509 ^ n5854 ^ 1'b0 ;
  assign n32513 = n32512 ^ n32510 ^ 1'b0 ;
  assign n32514 = ( ~n9210 & n16360 ) | ( ~n9210 & n32513 ) | ( n16360 & n32513 ) ;
  assign n32515 = n20875 | n32514 ;
  assign n32516 = n32515 ^ n7968 ^ 1'b0 ;
  assign n32517 = n32516 ^ n25884 ^ n9490 ;
  assign n32518 = n32517 ^ n7597 ^ n6391 ;
  assign n32519 = ~n4633 & n17870 ;
  assign n32520 = ( n3655 & n6673 ) | ( n3655 & ~n31618 ) | ( n6673 & ~n31618 ) ;
  assign n32521 = n32520 ^ n30080 ^ 1'b0 ;
  assign n32522 = n6277 & n32521 ;
  assign n32523 = n31945 ^ n11287 ^ 1'b0 ;
  assign n32524 = ~n1884 & n32523 ;
  assign n32525 = n31729 ^ n20272 ^ 1'b0 ;
  assign n32526 = ~n27465 & n32525 ;
  assign n32527 = n32526 ^ n23257 ^ 1'b0 ;
  assign n32528 = n32524 & n32527 ;
  assign n32529 = n32528 ^ n31945 ^ n15887 ;
  assign n32530 = ~n6584 & n7587 ;
  assign n32531 = n10696 ^ n8994 ^ 1'b0 ;
  assign n32532 = n32530 & n32531 ;
  assign n32533 = n32532 ^ n6334 ^ 1'b0 ;
  assign n32534 = n2046 & n32533 ;
  assign n32535 = n32534 ^ n24803 ^ n8139 ;
  assign n32536 = n32535 ^ n28541 ^ n14422 ;
  assign n32537 = n20354 ^ n19251 ^ n15504 ;
  assign n32538 = n22037 ^ n8593 ^ 1'b0 ;
  assign n32539 = n25774 | n32538 ;
  assign n32540 = n32539 ^ n5420 ^ 1'b0 ;
  assign n32541 = ~n5246 & n32540 ;
  assign n32542 = n24480 & n32541 ;
  assign n32543 = ~n6760 & n8053 ;
  assign n32544 = n32543 ^ n21824 ^ 1'b0 ;
  assign n32547 = n5098 ^ n3314 ^ n1943 ;
  assign n32545 = n16026 ^ n5945 ^ 1'b0 ;
  assign n32546 = n2034 | n32545 ;
  assign n32548 = n32547 ^ n32546 ^ 1'b0 ;
  assign n32549 = ~n5783 & n32548 ;
  assign n32550 = n19133 ^ n12624 ^ n9301 ;
  assign n32551 = n32550 ^ n25898 ^ n14067 ;
  assign n32552 = n26874 ^ n18504 ^ n2793 ;
  assign n32553 = n20425 & n28943 ;
  assign n32554 = n32553 ^ x5 ^ 1'b0 ;
  assign n32559 = n10540 | n29530 ;
  assign n32560 = n11400 & ~n32559 ;
  assign n32561 = n16739 ^ n9911 ^ 1'b0 ;
  assign n32562 = ~n32560 & n32561 ;
  assign n32563 = n32562 ^ n9698 ^ n4334 ;
  assign n32555 = n11179 ^ n7496 ^ 1'b0 ;
  assign n32556 = x123 & ~n32555 ;
  assign n32557 = n32556 ^ n22436 ^ 1'b0 ;
  assign n32558 = n6643 | n32557 ;
  assign n32564 = n32563 ^ n32558 ^ 1'b0 ;
  assign n32565 = ( n538 & n3159 ) | ( n538 & ~n8638 ) | ( n3159 & ~n8638 ) ;
  assign n32566 = n32565 ^ n25233 ^ 1'b0 ;
  assign n32567 = n17929 & ~n30326 ;
  assign n32568 = n32567 ^ n15137 ^ 1'b0 ;
  assign n32569 = ~n3789 & n6602 ;
  assign n32570 = n16484 & n32569 ;
  assign n32571 = n7134 & ~n13275 ;
  assign n32572 = n32571 ^ n25849 ^ 1'b0 ;
  assign n32573 = n19314 & ~n32572 ;
  assign n32574 = n32573 ^ n17985 ^ n12576 ;
  assign n32575 = n9581 & n32574 ;
  assign n32576 = n7391 & n32575 ;
  assign n32577 = n32570 & n32576 ;
  assign n32578 = n11782 ^ n6214 ^ n2438 ;
  assign n32579 = ( ~n12786 & n22620 ) | ( ~n12786 & n32578 ) | ( n22620 & n32578 ) ;
  assign n32581 = n15153 ^ n1042 ^ 1'b0 ;
  assign n32580 = n11895 & n19214 ;
  assign n32582 = n32581 ^ n32580 ^ 1'b0 ;
  assign n32585 = n8707 & ~n14851 ;
  assign n32586 = n14309 & n32585 ;
  assign n32583 = n11250 & n32159 ;
  assign n32584 = n32583 ^ n26648 ^ 1'b0 ;
  assign n32587 = n32586 ^ n32584 ^ n17556 ;
  assign n32588 = n23732 ^ n13173 ^ 1'b0 ;
  assign n32589 = n1135 & n32588 ;
  assign n32590 = n7157 & n32589 ;
  assign n32591 = n9750 ^ n2711 ^ 1'b0 ;
  assign n32592 = ~n702 & n32591 ;
  assign n32593 = n32592 ^ n22939 ^ n9823 ;
  assign n32595 = ( n771 & n1125 ) | ( n771 & ~n24351 ) | ( n1125 & ~n24351 ) ;
  assign n32594 = n9203 & ~n30789 ;
  assign n32596 = n32595 ^ n32594 ^ 1'b0 ;
  assign n32597 = n23293 ^ n10710 ^ n10449 ;
  assign n32599 = ( ~n3793 & n8419 ) | ( ~n3793 & n10755 ) | ( n8419 & n10755 ) ;
  assign n32600 = ( ~n1806 & n31035 ) | ( ~n1806 & n32599 ) | ( n31035 & n32599 ) ;
  assign n32598 = n573 & n7428 ;
  assign n32601 = n32600 ^ n32598 ^ n25605 ;
  assign n32602 = ~n9344 & n25070 ;
  assign n32603 = n32602 ^ n30234 ^ 1'b0 ;
  assign n32604 = n5069 & n32603 ;
  assign n32605 = n6338 | n11686 ;
  assign n32606 = n20682 & ~n32605 ;
  assign n32607 = ~n10385 & n14415 ;
  assign n32608 = n32607 ^ n18689 ^ 1'b0 ;
  assign n32609 = x217 & n426 ;
  assign n32610 = ( n4197 & n10406 ) | ( n4197 & n32609 ) | ( n10406 & n32609 ) ;
  assign n32611 = n3725 ^ n3658 ^ 1'b0 ;
  assign n32612 = n32611 ^ n19651 ^ 1'b0 ;
  assign n32613 = n32610 & n32612 ;
  assign n32614 = n32608 & n32613 ;
  assign n32615 = ~n13863 & n32614 ;
  assign n32616 = n29865 ^ n18601 ^ 1'b0 ;
  assign n32617 = ( n17462 & ~n22055 ) | ( n17462 & n24505 ) | ( ~n22055 & n24505 ) ;
  assign n32618 = ( n2311 & ~n5592 ) | ( n2311 & n21356 ) | ( ~n5592 & n21356 ) ;
  assign n32619 = n30474 | n32618 ;
  assign n32620 = ( n1702 & n5112 ) | ( n1702 & n12013 ) | ( n5112 & n12013 ) ;
  assign n32621 = ~n18228 & n32620 ;
  assign n32622 = ~n32619 & n32621 ;
  assign n32623 = n32622 ^ n29364 ^ 1'b0 ;
  assign n32624 = n28569 ^ n20516 ^ 1'b0 ;
  assign n32625 = ~n1592 & n32624 ;
  assign n32626 = n3958 | n8173 ;
  assign n32627 = ( n20066 & ~n32625 ) | ( n20066 & n32626 ) | ( ~n32625 & n32626 ) ;
  assign n32628 = n25452 ^ n15890 ^ n15164 ;
  assign n32629 = ~n21161 & n32628 ;
  assign n32630 = ( ~n1004 & n13924 ) | ( ~n1004 & n16679 ) | ( n13924 & n16679 ) ;
  assign n32631 = n32630 ^ n31807 ^ 1'b0 ;
  assign n32632 = n27940 ^ n6189 ^ 1'b0 ;
  assign n32633 = n32632 ^ n14842 ^ n14683 ;
  assign n32634 = n28498 ^ n25890 ^ n2577 ;
  assign n32635 = ( ~n7737 & n8858 ) | ( ~n7737 & n23390 ) | ( n8858 & n23390 ) ;
  assign n32636 = n1068 & ~n32635 ;
  assign n32637 = n8575 | n19722 ;
  assign n32638 = n7446 & ~n13833 ;
  assign n32639 = n32638 ^ n14233 ^ n1671 ;
  assign n32640 = ~n17210 & n32639 ;
  assign n32642 = n13502 ^ x204 ^ 1'b0 ;
  assign n32643 = n21913 & ~n32642 ;
  assign n32641 = n11387 | n24006 ;
  assign n32644 = n32643 ^ n32641 ^ 1'b0 ;
  assign n32645 = n6058 & ~n29378 ;
  assign n32646 = n7487 & n32645 ;
  assign n32647 = ~n4728 & n25303 ;
  assign n32648 = ( ~n2020 & n32646 ) | ( ~n2020 & n32647 ) | ( n32646 & n32647 ) ;
  assign n32649 = n2515 | n12794 ;
  assign n32650 = n5264 | n32649 ;
  assign n32651 = ( n23609 & n32648 ) | ( n23609 & ~n32650 ) | ( n32648 & ~n32650 ) ;
  assign n32652 = n18248 ^ n15569 ^ 1'b0 ;
  assign n32653 = n7669 & ~n32652 ;
  assign n32654 = ( ~n10523 & n13554 ) | ( ~n10523 & n32653 ) | ( n13554 & n32653 ) ;
  assign n32655 = n17272 & ~n27237 ;
  assign n32656 = n22840 | n25148 ;
  assign n32657 = n18682 & ~n32656 ;
  assign n32658 = ~n15444 & n26352 ;
  assign n32659 = n12896 & n30076 ;
  assign n32660 = ( ~n9136 & n13348 ) | ( ~n9136 & n32659 ) | ( n13348 & n32659 ) ;
  assign n32664 = ( n3699 & n3789 ) | ( n3699 & ~n28292 ) | ( n3789 & ~n28292 ) ;
  assign n32665 = n32664 ^ n21994 ^ n12214 ;
  assign n32666 = ~n14469 & n32665 ;
  assign n32662 = ~n1783 & n25882 ;
  assign n32661 = ( ~n18345 & n22045 ) | ( ~n18345 & n24001 ) | ( n22045 & n24001 ) ;
  assign n32663 = n32662 ^ n32661 ^ 1'b0 ;
  assign n32667 = n32666 ^ n32663 ^ n25231 ;
  assign n32668 = n16217 ^ n14004 ^ n10717 ;
  assign n32669 = n12169 & ~n32668 ;
  assign n32670 = n6742 & n13608 ;
  assign n32671 = n5369 & ~n20186 ;
  assign n32672 = n17629 ^ n8296 ^ 1'b0 ;
  assign n32673 = n10497 & n32672 ;
  assign n32674 = n32671 & n32673 ;
  assign n32675 = n30761 ^ n15626 ^ 1'b0 ;
  assign n32676 = ~n7199 & n12887 ;
  assign n32677 = n20310 & ~n21606 ;
  assign n32678 = ~n4290 & n32677 ;
  assign n32679 = n32678 ^ n22736 ^ 1'b0 ;
  assign n32680 = ( n5504 & n20761 ) | ( n5504 & n32679 ) | ( n20761 & n32679 ) ;
  assign n32681 = ( n5904 & n15504 ) | ( n5904 & n32680 ) | ( n15504 & n32680 ) ;
  assign n32682 = n18752 ^ n8305 ^ n4754 ;
  assign n32683 = n32682 ^ n22635 ^ 1'b0 ;
  assign n32684 = ( ~n3199 & n10996 ) | ( ~n3199 & n15677 ) | ( n10996 & n15677 ) ;
  assign n32685 = n32684 ^ n6478 ^ 1'b0 ;
  assign n32686 = ( ~n2775 & n6647 ) | ( ~n2775 & n32685 ) | ( n6647 & n32685 ) ;
  assign n32687 = ( n5741 & n12224 ) | ( n5741 & ~n22485 ) | ( n12224 & ~n22485 ) ;
  assign n32688 = ~n2376 & n32687 ;
  assign n32689 = n5314 & n13799 ;
  assign n32690 = n32689 ^ n8579 ^ 1'b0 ;
  assign n32691 = n29671 ^ n12467 ^ 1'b0 ;
  assign n32692 = n21864 & ~n32691 ;
  assign n32693 = n32692 ^ n10409 ^ 1'b0 ;
  assign n32694 = ~n8646 & n9667 ;
  assign n32695 = n1628 & n32694 ;
  assign n32696 = n32695 ^ n16743 ^ n14859 ;
  assign n32697 = ~n1387 & n26339 ;
  assign n32698 = ~n29524 & n32697 ;
  assign n32699 = ( ~n6323 & n32696 ) | ( ~n6323 & n32698 ) | ( n32696 & n32698 ) ;
  assign n32700 = n24154 ^ n5190 ^ 1'b0 ;
  assign n32701 = ~n10585 & n28837 ;
  assign n32703 = ( x51 & n5886 ) | ( x51 & ~n6431 ) | ( n5886 & ~n6431 ) ;
  assign n32704 = n17910 & n32703 ;
  assign n32702 = n3155 & ~n23892 ;
  assign n32705 = n32704 ^ n32702 ^ 1'b0 ;
  assign n32706 = n32705 ^ n29953 ^ 1'b0 ;
  assign n32707 = n3858 & ~n26887 ;
  assign n32708 = ~n19646 & n32707 ;
  assign n32709 = n11964 | n13258 ;
  assign n32710 = ~n23114 & n24354 ;
  assign n32711 = ~n32709 & n32710 ;
  assign n32712 = n1600 & n31850 ;
  assign n32713 = ( n11638 & n17727 ) | ( n11638 & ~n23900 ) | ( n17727 & ~n23900 ) ;
  assign n32714 = n9204 ^ n1183 ^ n310 ;
  assign n32715 = n17926 ^ n4476 ^ 1'b0 ;
  assign n32716 = n32714 & ~n32715 ;
  assign n32717 = n21375 ^ n13002 ^ n991 ;
  assign n32720 = n16105 ^ n1416 ^ 1'b0 ;
  assign n32721 = n8772 | n32720 ;
  assign n32718 = ~n9824 & n15167 ;
  assign n32719 = n28787 & n32718 ;
  assign n32722 = n32721 ^ n32719 ^ n10104 ;
  assign n32723 = n19910 ^ n15706 ^ n11455 ;
  assign n32725 = ~n13965 & n15577 ;
  assign n32726 = n13353 & n32725 ;
  assign n32724 = ~n3562 & n17317 ;
  assign n32727 = n32726 ^ n32724 ^ 1'b0 ;
  assign n32728 = n23692 ^ n6776 ^ n1015 ;
  assign n32729 = ( n15300 & n31509 ) | ( n15300 & ~n32728 ) | ( n31509 & ~n32728 ) ;
  assign n32730 = n32729 ^ n15845 ^ n12516 ;
  assign n32732 = n6607 & ~n26686 ;
  assign n32733 = n32732 ^ n1569 ^ 1'b0 ;
  assign n32731 = ~n12630 & n16078 ;
  assign n32734 = n32733 ^ n32731 ^ 1'b0 ;
  assign n32735 = ~n8530 & n29042 ;
  assign n32736 = n32734 & n32735 ;
  assign n32737 = n32736 ^ n17381 ^ n6398 ;
  assign n32738 = n19530 ^ n18952 ^ 1'b0 ;
  assign n32739 = n7885 & n32738 ;
  assign n32740 = n32739 ^ n22651 ^ n7679 ;
  assign n32741 = ( n20553 & ~n32737 ) | ( n20553 & n32740 ) | ( ~n32737 & n32740 ) ;
  assign n32742 = ~n17047 & n27248 ;
  assign n32743 = ~n2940 & n32742 ;
  assign n32744 = ( ~n22869 & n31790 ) | ( ~n22869 & n32743 ) | ( n31790 & n32743 ) ;
  assign n32745 = n14518 ^ n7213 ^ 1'b0 ;
  assign n32746 = n7246 | n32745 ;
  assign n32747 = ( ~n25046 & n28321 ) | ( ~n25046 & n32746 ) | ( n28321 & n32746 ) ;
  assign n32748 = n20225 | n27780 ;
  assign n32749 = ~n8344 & n32748 ;
  assign n32750 = n17043 ^ n5524 ^ 1'b0 ;
  assign n32751 = n9793 ^ n3325 ^ n1158 ;
  assign n32752 = n32750 & n32751 ;
  assign n32753 = n8484 & ~n32752 ;
  assign n32754 = n32753 ^ n25565 ^ n13629 ;
  assign n32755 = n18654 & ~n32754 ;
  assign n32756 = n32571 & n32755 ;
  assign n32757 = n2962 & ~n25391 ;
  assign n32758 = ~n3484 & n32757 ;
  assign n32759 = n32758 ^ n11188 ^ 1'b0 ;
  assign n32760 = ~n32756 & n32759 ;
  assign n32761 = ( ~n7092 & n32749 ) | ( ~n7092 & n32760 ) | ( n32749 & n32760 ) ;
  assign n32762 = ( n4848 & n8639 ) | ( n4848 & n11446 ) | ( n8639 & n11446 ) ;
  assign n32763 = n32762 ^ n11324 ^ n7891 ;
  assign n32764 = ~n1054 & n32763 ;
  assign n32765 = n14555 ^ n13754 ^ n13129 ;
  assign n32766 = n32765 ^ n11077 ^ n2837 ;
  assign n32767 = ( ~n394 & n3991 ) | ( ~n394 & n13922 ) | ( n3991 & n13922 ) ;
  assign n32768 = ( ~n15579 & n21526 ) | ( ~n15579 & n32767 ) | ( n21526 & n32767 ) ;
  assign n32769 = ~n14595 & n32768 ;
  assign n32770 = n32766 & n32769 ;
  assign n32771 = n3598 & ~n4662 ;
  assign n32772 = n32771 ^ n5999 ^ 1'b0 ;
  assign n32773 = ~n11752 & n32772 ;
  assign n32774 = n32773 ^ n9260 ^ 1'b0 ;
  assign n32775 = n32774 ^ n2528 ^ 1'b0 ;
  assign n32776 = n16451 ^ n15783 ^ n8221 ;
  assign n32777 = n32776 ^ n10889 ^ 1'b0 ;
  assign n32778 = ~n32775 & n32777 ;
  assign n32779 = x210 & ~n6929 ;
  assign n32780 = ~n30255 & n32779 ;
  assign n32781 = n30195 | n32780 ;
  assign n32782 = n2866 | n29035 ;
  assign n32783 = ( n19895 & ~n22710 ) | ( n19895 & n32782 ) | ( ~n22710 & n32782 ) ;
  assign n32784 = ( n32052 & n32781 ) | ( n32052 & ~n32783 ) | ( n32781 & ~n32783 ) ;
  assign n32785 = n25300 ^ n15188 ^ n8516 ;
  assign n32786 = ~n8635 & n22140 ;
  assign n32787 = ( ~n6421 & n25621 ) | ( ~n6421 & n32136 ) | ( n25621 & n32136 ) ;
  assign n32788 = ( n12798 & ~n29417 ) | ( n12798 & n32787 ) | ( ~n29417 & n32787 ) ;
  assign n32789 = n2748 | n11492 ;
  assign n32790 = n12717 ^ n4951 ^ n1604 ;
  assign n32791 = ( n15700 & n24174 ) | ( n15700 & ~n32790 ) | ( n24174 & ~n32790 ) ;
  assign n32792 = n19820 ^ n14821 ^ n10572 ;
  assign n32793 = ( ~n14874 & n20190 ) | ( ~n14874 & n29844 ) | ( n20190 & n29844 ) ;
  assign n32794 = ( n16999 & n21789 ) | ( n16999 & ~n32793 ) | ( n21789 & ~n32793 ) ;
  assign n32798 = ~n1434 & n14281 ;
  assign n32795 = ( n9437 & n13523 ) | ( n9437 & n15886 ) | ( n13523 & n15886 ) ;
  assign n32796 = n32795 ^ n27442 ^ n23587 ;
  assign n32797 = n32500 | n32796 ;
  assign n32799 = n32798 ^ n32797 ^ 1'b0 ;
  assign n32801 = n29844 ^ n19780 ^ 1'b0 ;
  assign n32802 = n16622 & n32801 ;
  assign n32803 = n32802 ^ n27957 ^ n11441 ;
  assign n32804 = n25984 ^ n5580 ^ n2674 ;
  assign n32805 = ~n5385 & n32804 ;
  assign n32806 = ~n2106 & n32805 ;
  assign n32807 = n32803 & n32806 ;
  assign n32800 = n4263 & ~n10151 ;
  assign n32808 = n32807 ^ n32800 ^ 1'b0 ;
  assign n32809 = n511 & n4773 ;
  assign n32810 = n29227 & n32809 ;
  assign n32811 = ~n29752 & n32810 ;
  assign n32812 = n32811 ^ n8329 ^ 1'b0 ;
  assign n32813 = ~n3290 & n4065 ;
  assign n32814 = n32813 ^ n29816 ^ 1'b0 ;
  assign n32815 = n5327 & n11515 ;
  assign n32826 = n826 ^ x74 ^ 1'b0 ;
  assign n32825 = ~n15039 & n15413 ;
  assign n32816 = n9571 ^ n9295 ^ 1'b0 ;
  assign n32817 = n10153 | n32816 ;
  assign n32818 = n8282 & ~n32817 ;
  assign n32819 = ( n7824 & ~n7944 ) | ( n7824 & n12040 ) | ( ~n7944 & n12040 ) ;
  assign n32820 = n13475 ^ n4463 ^ 1'b0 ;
  assign n32821 = ~n7120 & n32820 ;
  assign n32822 = n32821 ^ n4720 ^ 1'b0 ;
  assign n32823 = n32819 | n32822 ;
  assign n32824 = ( n11646 & n32818 ) | ( n11646 & ~n32823 ) | ( n32818 & ~n32823 ) ;
  assign n32827 = n32826 ^ n32825 ^ n32824 ;
  assign n32828 = n32815 & ~n32827 ;
  assign n32829 = n5397 ^ n4688 ^ 1'b0 ;
  assign n32830 = ( n6071 & n20816 ) | ( n6071 & n32829 ) | ( n20816 & n32829 ) ;
  assign n32834 = n19178 ^ n16060 ^ n15942 ;
  assign n32831 = n20425 & n27247 ;
  assign n32832 = n32831 ^ n12874 ^ 1'b0 ;
  assign n32833 = ( n7675 & n11440 ) | ( n7675 & n32832 ) | ( n11440 & n32832 ) ;
  assign n32835 = n32834 ^ n32833 ^ n23861 ;
  assign n32836 = n32741 ^ n7337 ^ 1'b0 ;
  assign n32837 = ( n5303 & n17107 ) | ( n5303 & n18516 ) | ( n17107 & n18516 ) ;
  assign n32838 = n29598 ^ n12072 ^ 1'b0 ;
  assign n32839 = n29893 ^ n25913 ^ n18560 ;
  assign n32840 = n17844 ^ n10318 ^ 1'b0 ;
  assign n32841 = n27288 | n32840 ;
  assign n32842 = n32841 ^ n8646 ^ 1'b0 ;
  assign n32843 = ( n18288 & ~n23732 ) | ( n18288 & n32842 ) | ( ~n23732 & n32842 ) ;
  assign n32844 = n27706 ^ n16946 ^ 1'b0 ;
  assign n32845 = n14984 & n24841 ;
  assign n32846 = n7749 ^ n7411 ^ 1'b0 ;
  assign n32847 = ( n14747 & ~n22930 ) | ( n14747 & n32846 ) | ( ~n22930 & n32846 ) ;
  assign n32848 = ( n20447 & ~n21453 ) | ( n20447 & n32847 ) | ( ~n21453 & n32847 ) ;
  assign n32849 = ~n7910 & n25030 ;
  assign n32850 = n32849 ^ n18121 ^ n11680 ;
  assign n32851 = n9819 ^ n6633 ^ 1'b0 ;
  assign n32852 = n7846 & ~n32851 ;
  assign n32853 = n26833 ^ n6018 ^ 1'b0 ;
  assign n32854 = n32853 ^ n28044 ^ 1'b0 ;
  assign n32855 = x37 & n2269 ;
  assign n32856 = n32855 ^ n3416 ^ 1'b0 ;
  assign n32857 = n32856 ^ n29814 ^ n12509 ;
  assign n32858 = ( n32852 & n32854 ) | ( n32852 & n32857 ) | ( n32854 & n32857 ) ;
  assign n32859 = ( n1395 & n10488 ) | ( n1395 & ~n20953 ) | ( n10488 & ~n20953 ) ;
  assign n32860 = ( n6143 & ~n20450 ) | ( n6143 & n32859 ) | ( ~n20450 & n32859 ) ;
  assign n32861 = n15735 | n28443 ;
  assign n32862 = n25209 ^ n5885 ^ 1'b0 ;
  assign n32863 = n12683 ^ n2056 ^ 1'b0 ;
  assign n32864 = n15889 & n32863 ;
  assign n32865 = ( n11674 & n22280 ) | ( n11674 & ~n32864 ) | ( n22280 & ~n32864 ) ;
  assign n32866 = ~n549 & n30223 ;
  assign n32867 = n31976 ^ n22495 ^ 1'b0 ;
  assign n32868 = ( n12344 & n32866 ) | ( n12344 & ~n32867 ) | ( n32866 & ~n32867 ) ;
  assign n32869 = n30198 & n32868 ;
  assign n32870 = n2595 & ~n9003 ;
  assign n32872 = n7260 ^ n2575 ^ 1'b0 ;
  assign n32873 = n7133 | n32872 ;
  assign n32871 = ~n1294 & n26164 ;
  assign n32874 = n32873 ^ n32871 ^ 1'b0 ;
  assign n32875 = ( ~n10294 & n17195 ) | ( ~n10294 & n31563 ) | ( n17195 & n31563 ) ;
  assign n32876 = ( n8561 & n11489 ) | ( n8561 & ~n19101 ) | ( n11489 & ~n19101 ) ;
  assign n32877 = n2123 & n18093 ;
  assign n32878 = ~n32876 & n32877 ;
  assign n32879 = n9552 | n32878 ;
  assign n32880 = n32879 ^ n23043 ^ 1'b0 ;
  assign n32881 = n32880 ^ n6612 ^ 1'b0 ;
  assign n32882 = n16255 & n32881 ;
  assign n32883 = n23650 ^ n1028 ^ 1'b0 ;
  assign n32884 = n5403 ^ n1031 ^ 1'b0 ;
  assign n32885 = n32883 | n32884 ;
  assign n32886 = n18077 ^ n1198 ^ 1'b0 ;
  assign n32887 = n1221 | n32886 ;
  assign n32888 = n24026 ^ n7232 ^ n6815 ;
  assign n32889 = ( n12129 & n32887 ) | ( n12129 & n32888 ) | ( n32887 & n32888 ) ;
  assign n32890 = n5189 | n12362 ;
  assign n32891 = n32890 ^ n4245 ^ 1'b0 ;
  assign n32892 = n32891 ^ n18176 ^ n3684 ;
  assign n32893 = n3791 & ~n32892 ;
  assign n32894 = n30328 ^ n7030 ^ 1'b0 ;
  assign n32895 = n7846 & ~n32894 ;
  assign n32896 = ( n2296 & ~n12048 ) | ( n2296 & n20033 ) | ( ~n12048 & n20033 ) ;
  assign n32897 = ~n4931 & n32896 ;
  assign n32898 = n32897 ^ n5830 ^ 1'b0 ;
  assign n32899 = ( n6096 & n13733 ) | ( n6096 & n32898 ) | ( n13733 & n32898 ) ;
  assign n32900 = ( ~n1900 & n22039 ) | ( ~n1900 & n32899 ) | ( n22039 & n32899 ) ;
  assign n32901 = n32895 & ~n32900 ;
  assign n32902 = ~n22382 & n32901 ;
  assign n32903 = n32902 ^ n19713 ^ n5572 ;
  assign n32904 = n17941 & n32903 ;
  assign n32905 = n27673 ^ n20235 ^ 1'b0 ;
  assign n32906 = ~n29095 & n32905 ;
  assign n32907 = n32906 ^ n11989 ^ n2247 ;
  assign n32908 = n10560 ^ n2759 ^ n1012 ;
  assign n32909 = ( n6238 & n6308 ) | ( n6238 & ~n32908 ) | ( n6308 & ~n32908 ) ;
  assign n32910 = n32909 ^ n18173 ^ n13347 ;
  assign n32911 = n23145 ^ n19840 ^ n15409 ;
  assign n32912 = ( n10417 & ~n16046 ) | ( n10417 & n19111 ) | ( ~n16046 & n19111 ) ;
  assign n32913 = n32912 ^ n7674 ^ 1'b0 ;
  assign n32914 = n32911 & n32913 ;
  assign n32915 = n13482 | n32914 ;
  assign n32916 = n11618 ^ n3354 ^ 1'b0 ;
  assign n32917 = ~n1760 & n2043 ;
  assign n32918 = ~n29932 & n32917 ;
  assign n32919 = n20883 ^ n18644 ^ 1'b0 ;
  assign n32920 = ~n7654 & n9193 ;
  assign n32921 = ~n32919 & n32920 ;
  assign n32922 = n6045 & ~n28813 ;
  assign n32923 = n25916 ^ n16999 ^ 1'b0 ;
  assign n32924 = n4022 & ~n32923 ;
  assign n32925 = n7398 & n32924 ;
  assign n32926 = n32922 & n32925 ;
  assign n32927 = n3996 & n9844 ;
  assign n32933 = n27193 ^ n14674 ^ 1'b0 ;
  assign n32929 = ( n4943 & n5638 ) | ( n4943 & n6185 ) | ( n5638 & n6185 ) ;
  assign n32930 = n8955 ^ n7609 ^ 1'b0 ;
  assign n32931 = n342 | n32930 ;
  assign n32932 = ( n937 & n32929 ) | ( n937 & ~n32931 ) | ( n32929 & ~n32931 ) ;
  assign n32934 = n32933 ^ n32932 ^ n7182 ;
  assign n32928 = n12984 | n22591 ;
  assign n32935 = n32934 ^ n32928 ^ 1'b0 ;
  assign n32936 = x192 & n16141 ;
  assign n32937 = n32935 & n32936 ;
  assign n32938 = ~n13665 & n28307 ;
  assign n32939 = n28916 ^ n11395 ^ n5901 ;
  assign n32940 = n32939 ^ n5361 ^ 1'b0 ;
  assign n32941 = n31995 ^ n12614 ^ n9135 ;
  assign n32942 = n4963 & ~n15409 ;
  assign n32943 = ( ~n8444 & n11038 ) | ( ~n8444 & n11112 ) | ( n11038 & n11112 ) ;
  assign n32944 = ~n13363 & n32943 ;
  assign n32945 = ( n4058 & n32942 ) | ( n4058 & n32944 ) | ( n32942 & n32944 ) ;
  assign n32946 = ( n2892 & ~n4316 ) | ( n2892 & n30623 ) | ( ~n4316 & n30623 ) ;
  assign n32947 = ~n27892 & n32946 ;
  assign n32948 = n17594 ^ n3092 ^ 1'b0 ;
  assign n32949 = n26287 & n32948 ;
  assign n32950 = n11057 & n32949 ;
  assign n32951 = n7376 & n32950 ;
  assign n32952 = n13899 | n22331 ;
  assign n32953 = n32952 ^ n16055 ^ 1'b0 ;
  assign n32954 = n18868 ^ n13007 ^ 1'b0 ;
  assign n32955 = n21088 | n32954 ;
  assign n32956 = n27498 ^ n8138 ^ 1'b0 ;
  assign n32957 = ( n13688 & n26128 ) | ( n13688 & n32956 ) | ( n26128 & n32956 ) ;
  assign n32958 = n32957 ^ n31229 ^ n3340 ;
  assign n32959 = ~n14433 & n20987 ;
  assign n32960 = n24935 ^ n16011 ^ n3534 ;
  assign n32961 = n17482 ^ n15366 ^ n6569 ;
  assign n32962 = ~n19382 & n32961 ;
  assign n32963 = n16877 ^ n301 ^ 1'b0 ;
  assign n32964 = n15780 | n32963 ;
  assign n32965 = n4723 | n32964 ;
  assign n32966 = ( n425 & n542 ) | ( n425 & ~n6986 ) | ( n542 & ~n6986 ) ;
  assign n32967 = n22410 ^ n16883 ^ 1'b0 ;
  assign n32968 = n32966 & ~n32967 ;
  assign n32969 = ~n21319 & n24981 ;
  assign n32970 = n6298 | n11994 ;
  assign n32971 = n2475 & ~n32970 ;
  assign n32972 = n16983 ^ n15608 ^ x229 ;
  assign n32973 = ( n11509 & n18335 ) | ( n11509 & n32972 ) | ( n18335 & n32972 ) ;
  assign n32974 = n11206 | n32973 ;
  assign n32975 = n4441 & ~n32974 ;
  assign n32976 = ( n5587 & ~n32971 ) | ( n5587 & n32975 ) | ( ~n32971 & n32975 ) ;
  assign n32977 = ~n23449 & n27642 ;
  assign n32978 = ( ~n1606 & n7057 ) | ( ~n1606 & n7644 ) | ( n7057 & n7644 ) ;
  assign n32979 = ~n2066 & n11705 ;
  assign n32980 = n32979 ^ n20304 ^ 1'b0 ;
  assign n32981 = ( n3099 & ~n24894 ) | ( n3099 & n32980 ) | ( ~n24894 & n32980 ) ;
  assign n32984 = n28499 ^ n11374 ^ n1573 ;
  assign n32982 = n9575 | n24521 ;
  assign n32983 = n9844 & ~n32982 ;
  assign n32985 = n32984 ^ n32983 ^ 1'b0 ;
  assign n32986 = n32067 & n32985 ;
  assign n32987 = ~n32981 & n32986 ;
  assign n32988 = ( ~n1145 & n4198 ) | ( ~n1145 & n6554 ) | ( n4198 & n6554 ) ;
  assign n32989 = n32988 ^ n16602 ^ n1651 ;
  assign n32990 = n32989 ^ n10979 ^ 1'b0 ;
  assign n32991 = n10545 | n32990 ;
  assign n32992 = n14123 ^ n5218 ^ 1'b0 ;
  assign n32993 = n12386 ^ n11661 ^ 1'b0 ;
  assign n32994 = n31822 ^ n4166 ^ n2796 ;
  assign n32995 = ( n18575 & n32993 ) | ( n18575 & n32994 ) | ( n32993 & n32994 ) ;
  assign n32996 = n14036 & n23517 ;
  assign n32997 = n32996 ^ n10193 ^ 1'b0 ;
  assign n32998 = n17202 ^ n15321 ^ n12219 ;
  assign n32999 = ( n32458 & n32997 ) | ( n32458 & n32998 ) | ( n32997 & n32998 ) ;
  assign n33000 = n2014 | n32999 ;
  assign n33001 = ( n19361 & ~n22421 ) | ( n19361 & n33000 ) | ( ~n22421 & n33000 ) ;
  assign n33002 = n6455 & ~n22502 ;
  assign n33003 = n33002 ^ n11161 ^ 1'b0 ;
  assign n33004 = n21487 ^ n4972 ^ 1'b0 ;
  assign n33005 = ~n33003 & n33004 ;
  assign n33006 = n33005 ^ n20273 ^ n6109 ;
  assign n33007 = ( ~n3707 & n31087 ) | ( ~n3707 & n33006 ) | ( n31087 & n33006 ) ;
  assign n33009 = ~n601 & n11023 ;
  assign n33010 = ~n10065 & n33009 ;
  assign n33011 = n33010 ^ n16153 ^ 1'b0 ;
  assign n33008 = n3881 & ~n13552 ;
  assign n33012 = n33011 ^ n33008 ^ 1'b0 ;
  assign n33013 = n10994 ^ n8487 ^ 1'b0 ;
  assign n33014 = ~x130 & n7369 ;
  assign n33015 = n33014 ^ n26178 ^ n18779 ;
  assign n33016 = ~n11950 & n33015 ;
  assign n33017 = ~n33013 & n33016 ;
  assign n33018 = n32142 ^ n4326 ^ n954 ;
  assign n33019 = n33018 ^ n28956 ^ n27058 ;
  assign n33020 = n2015 ^ n1813 ^ 1'b0 ;
  assign n33021 = n1570 | n33020 ;
  assign n33022 = ( ~n17757 & n33019 ) | ( ~n17757 & n33021 ) | ( n33019 & n33021 ) ;
  assign n33023 = ~n10794 & n21789 ;
  assign n33024 = n33023 ^ n9688 ^ 1'b0 ;
  assign n33025 = ( ~n1294 & n4422 ) | ( ~n1294 & n9220 ) | ( n4422 & n9220 ) ;
  assign n33026 = n5924 | n33025 ;
  assign n33027 = ( ~n13396 & n33024 ) | ( ~n13396 & n33026 ) | ( n33024 & n33026 ) ;
  assign n33028 = ( ~n2546 & n8689 ) | ( ~n2546 & n15772 ) | ( n8689 & n15772 ) ;
  assign n33029 = ~n3899 & n7531 ;
  assign n33030 = n33029 ^ n5729 ^ 1'b0 ;
  assign n33031 = n33030 ^ n12947 ^ 1'b0 ;
  assign n33032 = n13594 ^ n4589 ^ 1'b0 ;
  assign n33033 = ( n19168 & n25081 ) | ( n19168 & n33032 ) | ( n25081 & n33032 ) ;
  assign n33034 = n33033 ^ n3366 ^ 1'b0 ;
  assign n33035 = n15851 & ~n33034 ;
  assign n33036 = n3186 & ~n8874 ;
  assign n33037 = ~n4710 & n33036 ;
  assign n33038 = ~n32600 & n33037 ;
  assign n33039 = n33038 ^ n7278 ^ 1'b0 ;
  assign n33040 = n16530 & n33039 ;
  assign n33041 = n24626 ^ n17413 ^ 1'b0 ;
  assign n33042 = n29840 & n33041 ;
  assign n33043 = n12310 & n28302 ;
  assign n33044 = n33043 ^ n26342 ^ n20224 ;
  assign n33045 = n15880 ^ n14844 ^ n12995 ;
  assign n33046 = n33045 ^ n9491 ^ n2575 ;
  assign n33047 = n33046 ^ n24033 ^ n14681 ;
  assign n33048 = n33044 | n33047 ;
  assign n33049 = n14309 ^ n11220 ^ 1'b0 ;
  assign n33050 = n33049 ^ n32909 ^ n11715 ;
  assign n33051 = n16114 ^ n7082 ^ 1'b0 ;
  assign n33053 = n15601 & n19835 ;
  assign n33052 = x117 & n1678 ;
  assign n33054 = n33053 ^ n33052 ^ 1'b0 ;
  assign n33055 = n9195 & n11335 ;
  assign n33056 = n339 & n17571 ;
  assign n33057 = n33055 & n33056 ;
  assign n33058 = n4706 | n33057 ;
  assign n33059 = n33054 & ~n33058 ;
  assign n33060 = ~n4546 & n14789 ;
  assign n33061 = n12703 & ~n14666 ;
  assign n33062 = n33061 ^ n17115 ^ n15851 ;
  assign n33063 = n33062 ^ n14749 ^ 1'b0 ;
  assign n33064 = ~n33060 & n33063 ;
  assign n33065 = ( n8215 & n10235 ) | ( n8215 & ~n19624 ) | ( n10235 & ~n19624 ) ;
  assign n33066 = n15063 ^ n9810 ^ 1'b0 ;
  assign n33067 = n6297 & ~n33066 ;
  assign n33068 = n33067 ^ n18981 ^ n7700 ;
  assign n33069 = n22891 ^ n17836 ^ 1'b0 ;
  assign n33070 = ~n26044 & n30949 ;
  assign n33071 = n10208 & n14831 ;
  assign n33072 = ~n33070 & n33071 ;
  assign n33073 = n10780 | n11059 ;
  assign n33074 = n28078 ^ n25061 ^ n15781 ;
  assign n33075 = ( n21414 & n24661 ) | ( n21414 & ~n33074 ) | ( n24661 & ~n33074 ) ;
  assign n33076 = ( n9566 & n33073 ) | ( n9566 & ~n33075 ) | ( n33073 & ~n33075 ) ;
  assign n33077 = ( ~n6326 & n9092 ) | ( ~n6326 & n13320 ) | ( n9092 & n13320 ) ;
  assign n33078 = ~n1305 & n32318 ;
  assign n33079 = ~n19530 & n33078 ;
  assign n33080 = n33079 ^ n28272 ^ n16630 ;
  assign n33081 = n11090 & ~n14360 ;
  assign n33082 = ( n3061 & n4315 ) | ( n3061 & ~n4996 ) | ( n4315 & ~n4996 ) ;
  assign n33083 = n33082 ^ n21490 ^ n325 ;
  assign n33084 = ~n22795 & n33083 ;
  assign n33085 = n12812 & n33084 ;
  assign n33086 = ~x144 & n5729 ;
  assign n33087 = ~n8780 & n33086 ;
  assign n33088 = n6546 ^ n3730 ^ 1'b0 ;
  assign n33089 = n1642 | n33088 ;
  assign n33090 = ( n15917 & ~n21713 ) | ( n15917 & n33089 ) | ( ~n21713 & n33089 ) ;
  assign n33091 = n2684 & n4437 ;
  assign n33095 = n1623 & n6534 ;
  assign n33094 = n3188 & n10063 ;
  assign n33096 = n33095 ^ n33094 ^ 1'b0 ;
  assign n33097 = n4671 & ~n7083 ;
  assign n33098 = n33097 ^ n11511 ^ 1'b0 ;
  assign n33099 = n33098 ^ n21717 ^ 1'b0 ;
  assign n33100 = n33096 & ~n33099 ;
  assign n33092 = n25107 ^ n9736 ^ 1'b0 ;
  assign n33093 = ( n20804 & ~n30200 ) | ( n20804 & n33092 ) | ( ~n30200 & n33092 ) ;
  assign n33101 = n33100 ^ n33093 ^ n11589 ;
  assign n33102 = n24248 | n31940 ;
  assign n33103 = n19371 ^ n12847 ^ n5190 ;
  assign n33104 = ~n3910 & n33103 ;
  assign n33105 = n19697 & n33104 ;
  assign n33106 = ( n3049 & ~n23467 ) | ( n3049 & n27670 ) | ( ~n23467 & n27670 ) ;
  assign n33107 = ~n23499 & n33106 ;
  assign n33108 = n30667 ^ n26858 ^ 1'b0 ;
  assign n33109 = n12544 ^ n11470 ^ n7466 ;
  assign n33110 = ( n13322 & n16886 ) | ( n13322 & ~n33109 ) | ( n16886 & ~n33109 ) ;
  assign n33111 = ~n364 & n6828 ;
  assign n33112 = ~n15814 & n33111 ;
  assign n33113 = n17555 | n33112 ;
  assign n33114 = n10507 & ~n33113 ;
  assign n33115 = n22499 | n33114 ;
  assign n33116 = n33110 | n33115 ;
  assign n33117 = n15964 & n33116 ;
  assign n33118 = ( n30577 & n31962 ) | ( n30577 & n33117 ) | ( n31962 & n33117 ) ;
  assign n33119 = n1962 | n32647 ;
  assign n33120 = n33119 ^ n14085 ^ n1555 ;
  assign n33121 = n6608 | n10075 ;
  assign n33122 = n33121 ^ n4585 ^ 1'b0 ;
  assign n33123 = ( ~n6094 & n16894 ) | ( ~n6094 & n33122 ) | ( n16894 & n33122 ) ;
  assign n33124 = n959 & n25890 ;
  assign n33125 = n33124 ^ n1771 ^ 1'b0 ;
  assign n33126 = ( n3174 & ~n33123 ) | ( n3174 & n33125 ) | ( ~n33123 & n33125 ) ;
  assign n33127 = n17225 ^ n17206 ^ n5947 ;
  assign n33128 = n24470 ^ n18374 ^ n6963 ;
  assign n33129 = n8224 & ~n10397 ;
  assign n33130 = n33129 ^ n1669 ^ 1'b0 ;
  assign n33131 = ( ~n33127 & n33128 ) | ( ~n33127 & n33130 ) | ( n33128 & n33130 ) ;
  assign n33132 = ~n8551 & n17360 ;
  assign n33133 = n28357 & n33132 ;
  assign n33134 = n3626 & n5693 ;
  assign n33135 = n12887 ^ n2562 ^ 1'b0 ;
  assign n33136 = n14394 & ~n33135 ;
  assign n33137 = n3269 & ~n18827 ;
  assign n33138 = n33137 ^ n26430 ^ 1'b0 ;
  assign n33139 = n1264 & n19535 ;
  assign n33140 = n33139 ^ x108 ^ 1'b0 ;
  assign n33141 = n5492 | n33140 ;
  assign n33142 = n33138 | n33141 ;
  assign n33143 = ~n11671 & n24957 ;
  assign n33144 = x34 & n33143 ;
  assign n33145 = ~x34 & n33144 ;
  assign n33146 = n9896 ^ n6373 ^ n1545 ;
  assign n33147 = ( ~n5803 & n27874 ) | ( ~n5803 & n33146 ) | ( n27874 & n33146 ) ;
  assign n33148 = n4483 | n33147 ;
  assign n33149 = n5616 | n13338 ;
  assign n33150 = n33149 ^ n5098 ^ 1'b0 ;
  assign n33151 = n23808 & n27422 ;
  assign n33154 = n30091 ^ n12457 ^ 1'b0 ;
  assign n33155 = n2673 & ~n33154 ;
  assign n33152 = ( n416 & n1884 ) | ( n416 & ~n3145 ) | ( n1884 & ~n3145 ) ;
  assign n33153 = n29528 & n33152 ;
  assign n33156 = n33155 ^ n33153 ^ 1'b0 ;
  assign n33157 = ( n1415 & ~n16570 ) | ( n1415 & n32746 ) | ( ~n16570 & n32746 ) ;
  assign n33158 = ( n6446 & n15053 ) | ( n6446 & ~n33157 ) | ( n15053 & ~n33157 ) ;
  assign n33159 = ( n3340 & ~n19271 ) | ( n3340 & n19803 ) | ( ~n19271 & n19803 ) ;
  assign n33160 = n27917 ^ n5775 ^ n1677 ;
  assign n33161 = ( ~n5596 & n10643 ) | ( ~n5596 & n13175 ) | ( n10643 & n13175 ) ;
  assign n33162 = n14917 & ~n16760 ;
  assign n33163 = ( ~n1666 & n33161 ) | ( ~n1666 & n33162 ) | ( n33161 & n33162 ) ;
  assign n33164 = n1597 | n29931 ;
  assign n33165 = n29488 | n33164 ;
  assign n33166 = n22058 ^ n7351 ^ 1'b0 ;
  assign n33167 = ~n4775 & n33166 ;
  assign n33168 = n6471 & n16182 ;
  assign n33169 = ~n33167 & n33168 ;
  assign n33170 = ( n472 & ~n12959 ) | ( n472 & n17251 ) | ( ~n12959 & n17251 ) ;
  assign n33171 = ~n18054 & n33170 ;
  assign n33172 = ~n14708 & n33171 ;
  assign n33173 = ~n1783 & n3351 ;
  assign n33174 = n33173 ^ n12960 ^ 1'b0 ;
  assign n33175 = ( n14394 & ~n23719 ) | ( n14394 & n33174 ) | ( ~n23719 & n33174 ) ;
  assign n33176 = n21481 ^ n11827 ^ n3078 ;
  assign n33177 = n33176 ^ n26283 ^ 1'b0 ;
  assign n33178 = ~n31033 & n33177 ;
  assign n33179 = n5244 ^ n696 ^ n256 ;
  assign n33180 = n33179 ^ n15835 ^ n9441 ;
  assign n33181 = n14029 & n25315 ;
  assign n33182 = n775 | n22748 ;
  assign n33183 = n20978 ^ n14772 ^ n8119 ;
  assign n33184 = n1086 & ~n11527 ;
  assign n33185 = ~n257 & n33184 ;
  assign n33186 = n33183 & n33185 ;
  assign n33187 = n10057 ^ n7296 ^ 1'b0 ;
  assign n33188 = n10103 | n33187 ;
  assign n33189 = n4651 & ~n33188 ;
  assign n33190 = n33189 ^ n12636 ^ 1'b0 ;
  assign n33191 = n27198 ^ n5900 ^ 1'b0 ;
  assign n33192 = n30514 ^ n9520 ^ n8784 ;
  assign n33193 = n13658 ^ n9610 ^ 1'b0 ;
  assign n33195 = n14590 ^ n13278 ^ 1'b0 ;
  assign n33196 = ( n9754 & n20875 ) | ( n9754 & ~n33195 ) | ( n20875 & ~n33195 ) ;
  assign n33194 = ~n3141 & n30516 ;
  assign n33197 = n33196 ^ n33194 ^ 1'b0 ;
  assign n33198 = n10415 ^ x225 ^ 1'b0 ;
  assign n33199 = n20073 | n33198 ;
  assign n33200 = n2808 | n33199 ;
  assign n33201 = n13183 | n16252 ;
  assign n33202 = n19732 & ~n33201 ;
  assign n33203 = ( n965 & n3097 ) | ( n965 & ~n11585 ) | ( n3097 & ~n11585 ) ;
  assign n33204 = n10221 & ~n25888 ;
  assign n33205 = n6215 | n28864 ;
  assign n33206 = n9208 & ~n33205 ;
  assign n33207 = ( n11838 & n14228 ) | ( n11838 & n16659 ) | ( n14228 & n16659 ) ;
  assign n33208 = ( n18046 & n33206 ) | ( n18046 & ~n33207 ) | ( n33206 & ~n33207 ) ;
  assign n33209 = ( n7563 & n27638 ) | ( n7563 & n33208 ) | ( n27638 & n33208 ) ;
  assign n33210 = ( n6704 & n6934 ) | ( n6704 & ~n11028 ) | ( n6934 & ~n11028 ) ;
  assign n33212 = ~n10673 & n17699 ;
  assign n33211 = ( n1113 & n14901 ) | ( n1113 & n18910 ) | ( n14901 & n18910 ) ;
  assign n33213 = n33212 ^ n33211 ^ n7179 ;
  assign n33214 = n3686 & n33213 ;
  assign n33215 = ~n33210 & n33214 ;
  assign n33216 = n33215 ^ n7851 ^ 1'b0 ;
  assign n33217 = n13400 ^ n2606 ^ n499 ;
  assign n33218 = ( n2213 & ~n2325 ) | ( n2213 & n33217 ) | ( ~n2325 & n33217 ) ;
  assign n33219 = n33218 ^ n3320 ^ 1'b0 ;
  assign n33220 = n5264 & ~n33219 ;
  assign n33221 = ( n18173 & ~n25127 ) | ( n18173 & n25988 ) | ( ~n25127 & n25988 ) ;
  assign n33222 = n13033 & ~n33221 ;
  assign n33223 = n33222 ^ n21748 ^ 1'b0 ;
  assign n33224 = n17523 | n33223 ;
  assign n33225 = n12640 ^ n10746 ^ n3044 ;
  assign n33226 = ( n4510 & n29874 ) | ( n4510 & n31800 ) | ( n29874 & n31800 ) ;
  assign n33227 = ( n5933 & n9413 ) | ( n5933 & ~n33226 ) | ( n9413 & ~n33226 ) ;
  assign n33228 = ( ~n14834 & n25391 ) | ( ~n14834 & n26422 ) | ( n25391 & n26422 ) ;
  assign n33229 = n33228 ^ n1039 ^ 1'b0 ;
  assign n33230 = ( n12205 & n21309 ) | ( n12205 & ~n33229 ) | ( n21309 & ~n33229 ) ;
  assign n33231 = n1793 | n17712 ;
  assign n33232 = n33231 ^ n5901 ^ 1'b0 ;
  assign n33233 = n33232 ^ n20343 ^ n6683 ;
  assign n33234 = n33233 ^ n24580 ^ n19670 ;
  assign n33235 = n18518 ^ n3307 ^ n1445 ;
  assign n33236 = n22770 & n28371 ;
  assign n33237 = ( n6266 & ~n33235 ) | ( n6266 & n33236 ) | ( ~n33235 & n33236 ) ;
  assign n33238 = n14046 ^ n8266 ^ 1'b0 ;
  assign n33239 = n33237 | n33238 ;
  assign n33240 = n3646 | n14139 ;
  assign n33241 = n33239 & ~n33240 ;
  assign n33242 = n32218 ^ n7923 ^ 1'b0 ;
  assign n33243 = n6460 & n33242 ;
  assign n33244 = ~n4157 & n11944 ;
  assign n33245 = ( ~n6339 & n30268 ) | ( ~n6339 & n33244 ) | ( n30268 & n33244 ) ;
  assign n33246 = n27504 ^ n1538 ^ 1'b0 ;
  assign n33247 = ( n19008 & n29243 ) | ( n19008 & n33246 ) | ( n29243 & n33246 ) ;
  assign n33248 = n28179 ^ n22484 ^ n11310 ;
  assign n33249 = ( n2489 & n8813 ) | ( n2489 & ~n12995 ) | ( n8813 & ~n12995 ) ;
  assign n33250 = n33249 ^ n31654 ^ n26206 ;
  assign n33251 = ( n8021 & ~n14063 ) | ( n8021 & n27579 ) | ( ~n14063 & n27579 ) ;
  assign n33252 = n8139 & ~n27575 ;
  assign n33253 = ~n33251 & n33252 ;
  assign n33255 = n6277 & n13545 ;
  assign n33256 = n12697 & n33255 ;
  assign n33254 = n17246 & n31317 ;
  assign n33257 = n33256 ^ n33254 ^ n7942 ;
  assign n33258 = n15831 ^ n12568 ^ n8316 ;
  assign n33259 = n25494 ^ n23906 ^ n20091 ;
  assign n33260 = n33259 ^ n24110 ^ n22710 ;
  assign n33262 = ( n2199 & n9898 ) | ( n2199 & ~n19703 ) | ( n9898 & ~n19703 ) ;
  assign n33261 = ( n1555 & n15698 ) | ( n1555 & n29143 ) | ( n15698 & n29143 ) ;
  assign n33263 = n33262 ^ n33261 ^ n13899 ;
  assign n33264 = n11012 ^ n4024 ^ 1'b0 ;
  assign n33265 = ~n3419 & n16893 ;
  assign n33266 = n33265 ^ n17937 ^ 1'b0 ;
  assign n33267 = n32039 ^ n2206 ^ 1'b0 ;
  assign n33272 = ( n3514 & ~n4226 ) | ( n3514 & n5295 ) | ( ~n4226 & n5295 ) ;
  assign n33268 = n2960 ^ n1955 ^ 1'b0 ;
  assign n33269 = n20395 | n33268 ;
  assign n33270 = n33269 ^ n18545 ^ n14189 ;
  assign n33271 = ~n14645 & n33270 ;
  assign n33273 = n33272 ^ n33271 ^ n759 ;
  assign n33275 = ~n14975 & n20720 ;
  assign n33276 = ( ~n15976 & n18502 ) | ( ~n15976 & n33275 ) | ( n18502 & n33275 ) ;
  assign n33274 = n23372 | n29819 ;
  assign n33277 = n33276 ^ n33274 ^ n19937 ;
  assign n33278 = n33277 ^ n33162 ^ n21399 ;
  assign n33279 = ( n11848 & n12777 ) | ( n11848 & n22253 ) | ( n12777 & n22253 ) ;
  assign n33280 = ~n12917 & n33279 ;
  assign n33281 = n9815 & n22110 ;
  assign n33282 = n33281 ^ n24366 ^ 1'b0 ;
  assign n33283 = n9802 & n15482 ;
  assign n33284 = n33283 ^ n2600 ^ 1'b0 ;
  assign n33286 = n24005 | n27324 ;
  assign n33287 = n3806 | n33286 ;
  assign n33285 = n4266 & n18578 ;
  assign n33288 = n33287 ^ n33285 ^ 1'b0 ;
  assign n33289 = ( n2397 & ~n33284 ) | ( n2397 & n33288 ) | ( ~n33284 & n33288 ) ;
  assign n33290 = n13573 | n16271 ;
  assign n33291 = n8672 | n33290 ;
  assign n33292 = n33291 ^ n6270 ^ n2442 ;
  assign n33293 = n33292 ^ n27453 ^ 1'b0 ;
  assign n33295 = ( n458 & ~n495 ) | ( n458 & n7541 ) | ( ~n495 & n7541 ) ;
  assign n33294 = n12624 ^ n8032 ^ n312 ;
  assign n33296 = n33295 ^ n33294 ^ n26162 ;
  assign n33297 = ( n14934 & n15660 ) | ( n14934 & n33296 ) | ( n15660 & n33296 ) ;
  assign n33298 = n11692 ^ n721 ^ 1'b0 ;
  assign n33299 = n15683 | n26736 ;
  assign n33300 = n30226 ^ n8501 ^ 1'b0 ;
  assign n33301 = n5953 | n33300 ;
  assign n33302 = ( ~n15552 & n15701 ) | ( ~n15552 & n33301 ) | ( n15701 & n33301 ) ;
  assign n33303 = n662 & n7697 ;
  assign n33304 = n33303 ^ n4816 ^ 1'b0 ;
  assign n33305 = n1073 & ~n33304 ;
  assign n33306 = n33302 & n33305 ;
  assign n33307 = ( ~n14968 & n26748 ) | ( ~n14968 & n32768 ) | ( n26748 & n32768 ) ;
  assign n33308 = n12196 ^ n2975 ^ n1087 ;
  assign n33309 = ( n14220 & n18982 ) | ( n14220 & ~n33308 ) | ( n18982 & ~n33308 ) ;
  assign n33310 = n16195 ^ n8045 ^ n2533 ;
  assign n33311 = n21348 ^ n5844 ^ n5568 ;
  assign n33314 = ~n4052 & n11271 ;
  assign n33315 = n33314 ^ n24199 ^ n3909 ;
  assign n33316 = ~n11381 & n33315 ;
  assign n33317 = n6899 & n33316 ;
  assign n33312 = n21230 ^ n12133 ^ n6150 ;
  assign n33313 = n8787 | n33312 ;
  assign n33318 = n33317 ^ n33313 ^ 1'b0 ;
  assign n33319 = n16950 ^ n13238 ^ 1'b0 ;
  assign n33320 = ( n9192 & n14349 ) | ( n9192 & n33319 ) | ( n14349 & n33319 ) ;
  assign n33321 = n32931 ^ n397 ^ 1'b0 ;
  assign n33322 = n5764 & n6293 ;
  assign n33323 = n660 & n33322 ;
  assign n33324 = n33323 ^ n19515 ^ n5465 ;
  assign n33325 = n27246 | n33324 ;
  assign n33326 = n31793 ^ n16463 ^ n8114 ;
  assign n33327 = n33326 ^ n26140 ^ n610 ;
  assign n33328 = n33060 ^ n5662 ^ 1'b0 ;
  assign n33329 = n23420 | n33328 ;
  assign n33330 = n25584 ^ n16744 ^ 1'b0 ;
  assign n33331 = ( ~n9889 & n29159 ) | ( ~n9889 & n33330 ) | ( n29159 & n33330 ) ;
  assign n33332 = n13906 ^ n9171 ^ 1'b0 ;
  assign n33333 = ~n5783 & n19670 ;
  assign n33334 = n33333 ^ n8895 ^ 1'b0 ;
  assign n33335 = n33334 ^ n15912 ^ n8354 ;
  assign n33336 = n23552 & ~n33335 ;
  assign n33338 = n10700 ^ n6269 ^ 1'b0 ;
  assign n33339 = n3994 & ~n33338 ;
  assign n33340 = n10247 & ~n33339 ;
  assign n33341 = n33340 ^ n17847 ^ n6903 ;
  assign n33337 = ~n11221 & n30500 ;
  assign n33342 = n33341 ^ n33337 ^ 1'b0 ;
  assign n33343 = n31344 ^ n27877 ^ 1'b0 ;
  assign n33344 = n4659 ^ n3679 ^ 1'b0 ;
  assign n33345 = ~n15452 & n33344 ;
  assign n33346 = ~n7327 & n33345 ;
  assign n33347 = n33346 ^ n10744 ^ n1507 ;
  assign n33348 = n20339 & n28373 ;
  assign n33353 = n3914 | n8013 ;
  assign n33354 = n26202 & ~n33353 ;
  assign n33350 = n26154 ^ n7412 ^ 1'b0 ;
  assign n33351 = ~n25050 & n33350 ;
  assign n33352 = n22280 & n33351 ;
  assign n33349 = n6219 ^ n1184 ^ n789 ;
  assign n33355 = n33354 ^ n33352 ^ n33349 ;
  assign n33357 = n2118 ^ x169 ^ 1'b0 ;
  assign n33358 = n14550 | n33357 ;
  assign n33356 = ( ~x142 & n529 ) | ( ~x142 & n19233 ) | ( n529 & n19233 ) ;
  assign n33359 = n33358 ^ n33356 ^ 1'b0 ;
  assign n33360 = n30296 ^ n14565 ^ 1'b0 ;
  assign n33361 = ( n2188 & ~n21356 ) | ( n2188 & n33360 ) | ( ~n21356 & n33360 ) ;
  assign n33362 = n7600 & ~n24290 ;
  assign n33363 = n25231 & n33362 ;
  assign n33364 = n33363 ^ n20067 ^ 1'b0 ;
  assign n33365 = n33364 ^ n9266 ^ 1'b0 ;
  assign n33366 = n33361 & ~n33365 ;
  assign n33367 = n9669 & ~n25196 ;
  assign n33368 = ~n14206 & n21833 ;
  assign n33369 = n33367 & n33368 ;
  assign n33370 = n6928 & ~n9627 ;
  assign n33371 = n33370 ^ n5831 ^ 1'b0 ;
  assign n33372 = n33371 ^ n19644 ^ 1'b0 ;
  assign n33373 = n27935 | n33372 ;
  assign n33374 = n33373 ^ n7493 ^ 1'b0 ;
  assign n33375 = n12198 ^ n10055 ^ n1303 ;
  assign n33376 = ( n13806 & n24915 ) | ( n13806 & n30240 ) | ( n24915 & n30240 ) ;
  assign n33377 = n14120 ^ n10176 ^ n6973 ;
  assign n33378 = n33377 ^ n6342 ^ n2736 ;
  assign n33379 = n313 & ~n19200 ;
  assign n33380 = ~n32703 & n33379 ;
  assign n33381 = n33380 ^ n14432 ^ n2497 ;
  assign n33382 = n33381 ^ n7668 ^ 1'b0 ;
  assign n33383 = n6657 ^ n770 ^ 1'b0 ;
  assign n33384 = n7345 & ~n33383 ;
  assign n33385 = n33384 ^ n7432 ^ 1'b0 ;
  assign n33386 = n33385 ^ n12045 ^ 1'b0 ;
  assign n33387 = n5660 & n33386 ;
  assign n33388 = ( n7498 & n9918 ) | ( n7498 & n33387 ) | ( n9918 & n33387 ) ;
  assign n33389 = n6390 & n9285 ;
  assign n33390 = n33389 ^ n5781 ^ 1'b0 ;
  assign n33391 = ( ~n33382 & n33388 ) | ( ~n33382 & n33390 ) | ( n33388 & n33390 ) ;
  assign n33392 = n13105 | n33391 ;
  assign n33393 = n33392 ^ n30599 ^ 1'b0 ;
  assign n33394 = n3958 ^ n1198 ^ 1'b0 ;
  assign n33395 = n2417 & ~n33394 ;
  assign n33396 = n20091 ^ n13250 ^ 1'b0 ;
  assign n33397 = n33395 & n33396 ;
  assign n33398 = ( n2071 & n10382 ) | ( n2071 & ~n32318 ) | ( n10382 & ~n32318 ) ;
  assign n33399 = n21359 & n33398 ;
  assign n33400 = n18514 ^ n1699 ^ 1'b0 ;
  assign n33401 = n33400 ^ n7681 ^ n4307 ;
  assign n33402 = ( n18296 & n19585 ) | ( n18296 & n33401 ) | ( n19585 & n33401 ) ;
  assign n33403 = n2595 & ~n32163 ;
  assign n33404 = ( n268 & n1084 ) | ( n268 & ~n33403 ) | ( n1084 & ~n33403 ) ;
  assign n33405 = n33404 ^ n32291 ^ n30001 ;
  assign n33406 = n32318 ^ n18755 ^ n15057 ;
  assign n33417 = n17091 | n23331 ;
  assign n33413 = n1330 | n3138 ;
  assign n33414 = n6322 | n23840 ;
  assign n33415 = n33413 | n33414 ;
  assign n33407 = ( n6850 & n7436 ) | ( n6850 & ~n16857 ) | ( n7436 & ~n16857 ) ;
  assign n33408 = n4080 ^ n604 ^ 1'b0 ;
  assign n33409 = n3889 & ~n33408 ;
  assign n33410 = n14297 & n33409 ;
  assign n33411 = ~n13814 & n33410 ;
  assign n33412 = ( n7935 & ~n33407 ) | ( n7935 & n33411 ) | ( ~n33407 & n33411 ) ;
  assign n33416 = n33415 ^ n33412 ^ 1'b0 ;
  assign n33418 = n33417 ^ n33416 ^ n19231 ;
  assign n33419 = x234 & ~n5927 ;
  assign n33421 = ~n26567 & n27093 ;
  assign n33420 = n5791 & ~n12147 ;
  assign n33422 = n33421 ^ n33420 ^ 1'b0 ;
  assign n33428 = n32876 ^ n16923 ^ n6670 ;
  assign n33423 = n10802 ^ n7325 ^ 1'b0 ;
  assign n33424 = n8854 | n33423 ;
  assign n33425 = n3794 ^ n2349 ^ 1'b0 ;
  assign n33426 = n33425 ^ n22194 ^ 1'b0 ;
  assign n33427 = n33424 | n33426 ;
  assign n33429 = n33428 ^ n33427 ^ n14410 ;
  assign n33430 = n14603 | n25375 ;
  assign n33431 = ( ~n1721 & n3898 ) | ( ~n1721 & n6488 ) | ( n3898 & n6488 ) ;
  assign n33432 = n1356 & n26026 ;
  assign n33433 = n29213 & n33432 ;
  assign n33434 = n6762 & ~n33433 ;
  assign n33435 = ( n12272 & ~n33431 ) | ( n12272 & n33434 ) | ( ~n33431 & n33434 ) ;
  assign n33436 = n6666 ^ n926 ^ 1'b0 ;
  assign n33437 = n20255 & n33436 ;
  assign n33438 = n11033 & ~n33437 ;
  assign n33439 = n19441 | n33438 ;
  assign n33440 = n4078 & ~n33439 ;
  assign n33441 = n2174 & ~n14900 ;
  assign n33442 = n33441 ^ n16195 ^ 1'b0 ;
  assign n33443 = n33442 ^ n23204 ^ n492 ;
  assign n33444 = ( ~n2142 & n30109 ) | ( ~n2142 & n30949 ) | ( n30109 & n30949 ) ;
  assign n33445 = n26464 & ~n30707 ;
  assign n33446 = n5856 ^ n3317 ^ 1'b0 ;
  assign n33447 = n20795 ^ n2067 ^ 1'b0 ;
  assign n33448 = n9604 & n11954 ;
  assign n33449 = ~n13937 & n33448 ;
  assign n33450 = n28635 | n33449 ;
  assign n33451 = n33450 ^ n20051 ^ 1'b0 ;
  assign n33452 = n849 & n7919 ;
  assign n33453 = n33451 & n33452 ;
  assign n33454 = n15413 ^ n12249 ^ n9461 ;
  assign n33455 = ~n16101 & n33454 ;
  assign n33456 = n28336 ^ n6589 ^ 1'b0 ;
  assign n33457 = n1846 & n33456 ;
  assign n33458 = ( ~n5996 & n6549 ) | ( ~n5996 & n29036 ) | ( n6549 & n29036 ) ;
  assign n33459 = n33457 & ~n33458 ;
  assign n33460 = n15016 & n33459 ;
  assign n33461 = n31361 ^ n6323 ^ 1'b0 ;
  assign n33462 = ( n8311 & n27670 ) | ( n8311 & n32281 ) | ( n27670 & n32281 ) ;
  assign n33463 = ( n8669 & n9823 ) | ( n8669 & ~n33462 ) | ( n9823 & ~n33462 ) ;
  assign n33464 = n30564 & ~n33463 ;
  assign n33465 = n33464 ^ n5778 ^ 1'b0 ;
  assign n33466 = n32023 ^ n30454 ^ 1'b0 ;
  assign n33467 = n19523 ^ n13917 ^ n7386 ;
  assign n33468 = ( n6102 & ~n6825 ) | ( n6102 & n27440 ) | ( ~n6825 & n27440 ) ;
  assign n33469 = n1028 & ~n5097 ;
  assign n33470 = n26505 & n33469 ;
  assign n33471 = n33470 ^ n22394 ^ 1'b0 ;
  assign n33473 = n2280 & ~n22136 ;
  assign n33474 = n25438 ^ n2782 ^ 1'b0 ;
  assign n33475 = n33473 | n33474 ;
  assign n33472 = n9085 ^ n701 ^ 1'b0 ;
  assign n33476 = n33475 ^ n33472 ^ n545 ;
  assign n33477 = ~n3040 & n23866 ;
  assign n33478 = ( n2144 & n12797 ) | ( n2144 & n16348 ) | ( n12797 & n16348 ) ;
  assign n33479 = n4814 ^ n1182 ^ 1'b0 ;
  assign n33480 = n19275 ^ n6881 ^ n3500 ;
  assign n33481 = n33480 ^ n9744 ^ n6569 ;
  assign n33482 = n33481 ^ n25699 ^ n10902 ;
  assign n33483 = ( n16622 & n33479 ) | ( n16622 & ~n33482 ) | ( n33479 & ~n33482 ) ;
  assign n33484 = n33483 ^ n21743 ^ 1'b0 ;
  assign n33488 = ~n8280 & n11477 ;
  assign n33489 = n21393 & n33488 ;
  assign n33485 = n4847 | n8017 ;
  assign n33486 = n33485 ^ n20160 ^ 1'b0 ;
  assign n33487 = n16137 & ~n33486 ;
  assign n33490 = n33489 ^ n33487 ^ n27965 ;
  assign n33491 = n21847 & ~n33490 ;
  assign n33492 = n21773 ^ n10654 ^ 1'b0 ;
  assign n33493 = n33491 & n33492 ;
  assign n33494 = n7625 & ~n22677 ;
  assign n33495 = n25018 ^ n20849 ^ 1'b0 ;
  assign n33496 = n18077 ^ n12860 ^ 1'b0 ;
  assign n33497 = ~n10520 & n33496 ;
  assign n33498 = ~n12220 & n33497 ;
  assign n33499 = n33498 ^ n6028 ^ 1'b0 ;
  assign n33500 = n4004 | n13906 ;
  assign n33501 = n33500 ^ n19692 ^ 1'b0 ;
  assign n33502 = n26446 ^ n23640 ^ n5529 ;
  assign n33503 = n26257 ^ n11642 ^ 1'b0 ;
  assign n33504 = n19461 & ~n33503 ;
  assign n33505 = n4656 | n15122 ;
  assign n33506 = n33505 ^ n19588 ^ 1'b0 ;
  assign n33507 = ( n5346 & n26429 ) | ( n5346 & ~n33506 ) | ( n26429 & ~n33506 ) ;
  assign n33508 = n33507 ^ n33312 ^ n21892 ;
  assign n33509 = n308 | n31057 ;
  assign n33510 = ( n7903 & n13587 ) | ( n7903 & ~n33509 ) | ( n13587 & ~n33509 ) ;
  assign n33511 = n33508 & n33510 ;
  assign n33512 = n33511 ^ n425 ^ 1'b0 ;
  assign n33513 = n3371 ^ n710 ^ 1'b0 ;
  assign n33514 = n22570 | n33513 ;
  assign n33515 = n33514 ^ n13720 ^ n7125 ;
  assign n33516 = n33515 ^ n19385 ^ x152 ;
  assign n33517 = ~n24409 & n27621 ;
  assign n33518 = n20932 | n22210 ;
  assign n33519 = ( ~n6360 & n16521 ) | ( ~n6360 & n20523 ) | ( n16521 & n20523 ) ;
  assign n33520 = ( n8607 & ~n18179 ) | ( n8607 & n28050 ) | ( ~n18179 & n28050 ) ;
  assign n33521 = ( ~n8288 & n33519 ) | ( ~n8288 & n33520 ) | ( n33519 & n33520 ) ;
  assign n33522 = n4245 | n12964 ;
  assign n33523 = n24320 & ~n33522 ;
  assign n33524 = n15203 ^ n10060 ^ 1'b0 ;
  assign n33525 = ~n32367 & n33524 ;
  assign n33526 = n33525 ^ n30005 ^ 1'b0 ;
  assign n33527 = n17806 & ~n28684 ;
  assign n33528 = ~n20565 & n33527 ;
  assign n33529 = n2050 | n2632 ;
  assign n33530 = n17783 | n33529 ;
  assign n33531 = n28163 ^ n21577 ^ n19949 ;
  assign n33532 = n4371 | n18046 ;
  assign n33533 = n33532 ^ n2272 ^ 1'b0 ;
  assign n33534 = n24928 & ~n33533 ;
  assign n33535 = n14643 | n33534 ;
  assign n33536 = ( ~n852 & n8778 ) | ( ~n852 & n33535 ) | ( n8778 & n33535 ) ;
  assign n33537 = n4418 ^ n994 ^ 1'b0 ;
  assign n33538 = n33537 ^ n24573 ^ n19566 ;
  assign n33539 = n16938 ^ n10691 ^ 1'b0 ;
  assign n33540 = n1761 | n33539 ;
  assign n33541 = n13932 & ~n33540 ;
  assign n33542 = n33541 ^ n9767 ^ 1'b0 ;
  assign n33543 = n30412 ^ n16970 ^ n12512 ;
  assign n33544 = ( n9595 & ~n21222 ) | ( n9595 & n30007 ) | ( ~n21222 & n30007 ) ;
  assign n33545 = n33543 & n33544 ;
  assign n33547 = n7120 ^ n6811 ^ n513 ;
  assign n33546 = ~n665 & n12416 ;
  assign n33548 = n33547 ^ n33546 ^ 1'b0 ;
  assign n33549 = n20501 ^ n11185 ^ n3210 ;
  assign n33550 = ~n1050 & n23882 ;
  assign n33551 = n6009 | n19829 ;
  assign n33552 = n33551 ^ n4228 ^ 1'b0 ;
  assign n33553 = ( ~n14739 & n33550 ) | ( ~n14739 & n33552 ) | ( n33550 & n33552 ) ;
  assign n33554 = n33553 ^ n9357 ^ n1183 ;
  assign n33555 = n18543 ^ n10571 ^ n8272 ;
  assign n33556 = ( ~n1219 & n23001 ) | ( ~n1219 & n33555 ) | ( n23001 & n33555 ) ;
  assign n33557 = ( ~n3832 & n9580 ) | ( ~n3832 & n18275 ) | ( n9580 & n18275 ) ;
  assign n33558 = n24643 | n28291 ;
  assign n33559 = n33558 ^ n4757 ^ 1'b0 ;
  assign n33560 = n20226 ^ n17251 ^ 1'b0 ;
  assign n33561 = n3193 & ~n33560 ;
  assign n33562 = n33561 ^ n30479 ^ 1'b0 ;
  assign n33563 = n26948 ^ n8608 ^ n2495 ;
  assign n33564 = ( n1538 & n2569 ) | ( n1538 & n3253 ) | ( n2569 & n3253 ) ;
  assign n33565 = ( n1249 & ~n22248 ) | ( n1249 & n33564 ) | ( ~n22248 & n33564 ) ;
  assign n33566 = ( ~n2688 & n10943 ) | ( ~n2688 & n26988 ) | ( n10943 & n26988 ) ;
  assign n33567 = n1398 | n33566 ;
  assign n33568 = n33567 ^ x96 ^ 1'b0 ;
  assign n33569 = ( n5282 & n6960 ) | ( n5282 & ~n12681 ) | ( n6960 & ~n12681 ) ;
  assign n33570 = ~n2087 & n33569 ;
  assign n33571 = n15622 & n33570 ;
  assign n33572 = n13336 ^ n11025 ^ n2406 ;
  assign n33573 = n33572 ^ n30375 ^ n26392 ;
  assign n33574 = n33573 ^ n10432 ^ n386 ;
  assign n33575 = ( ~n4685 & n9176 ) | ( ~n4685 & n9425 ) | ( n9176 & n9425 ) ;
  assign n33576 = n33575 ^ n28784 ^ n8842 ;
  assign n33577 = ( n13756 & n29643 ) | ( n13756 & ~n33576 ) | ( n29643 & ~n33576 ) ;
  assign n33578 = n8309 & ~n19601 ;
  assign n33579 = n28070 & n33578 ;
  assign n33581 = ( n613 & n3832 ) | ( n613 & ~n33082 ) | ( n3832 & ~n33082 ) ;
  assign n33580 = n15725 ^ n14840 ^ n1923 ;
  assign n33582 = n33581 ^ n33580 ^ 1'b0 ;
  assign n33583 = n13135 | n33582 ;
  assign n33584 = ~n6020 & n11493 ;
  assign n33585 = ( n17718 & ~n28185 ) | ( n17718 & n33584 ) | ( ~n28185 & n33584 ) ;
  assign n33586 = ( n14235 & n29855 ) | ( n14235 & n33585 ) | ( n29855 & n33585 ) ;
  assign n33588 = n21005 ^ n4446 ^ 1'b0 ;
  assign n33589 = n10677 & n33588 ;
  assign n33590 = n33589 ^ n13399 ^ 1'b0 ;
  assign n33587 = ( x170 & ~n9688 ) | ( x170 & n21039 ) | ( ~n9688 & n21039 ) ;
  assign n33591 = n33590 ^ n33587 ^ n31658 ;
  assign n33592 = n33591 ^ n14194 ^ n14144 ;
  assign n33593 = n2207 | n10970 ;
  assign n33594 = n24674 | n33593 ;
  assign n33595 = x148 & n4507 ;
  assign n33596 = n33595 ^ x175 ^ 1'b0 ;
  assign n33597 = n20366 ^ n4061 ^ n2858 ;
  assign n33598 = n33597 ^ n12362 ^ 1'b0 ;
  assign n33599 = n33598 ^ n6410 ^ n5298 ;
  assign n33600 = n19617 ^ n9220 ^ n3864 ;
  assign n33601 = ( n9661 & ~n11702 ) | ( n9661 & n33600 ) | ( ~n11702 & n33600 ) ;
  assign n33602 = n20738 ^ n5976 ^ n3211 ;
  assign n33603 = ( n559 & n5935 ) | ( n559 & n30776 ) | ( n5935 & n30776 ) ;
  assign n33604 = ( n1176 & ~n11919 ) | ( n1176 & n18127 ) | ( ~n11919 & n18127 ) ;
  assign n33605 = ( n7511 & n23945 ) | ( n7511 & n33604 ) | ( n23945 & n33604 ) ;
  assign n33606 = n1803 & n8224 ;
  assign n33607 = ( n20403 & ~n30398 ) | ( n20403 & n33606 ) | ( ~n30398 & n33606 ) ;
  assign n33608 = ( ~n9571 & n13346 ) | ( ~n9571 & n18992 ) | ( n13346 & n18992 ) ;
  assign n33609 = n10856 & ~n33608 ;
  assign n33610 = n33609 ^ n15620 ^ 1'b0 ;
  assign n33611 = n16697 & n33610 ;
  assign n33612 = n33611 ^ n3696 ^ 1'b0 ;
  assign n33613 = n2031 | n15023 ;
  assign n33614 = n33210 & ~n33613 ;
  assign n33615 = n16034 & ~n33614 ;
  assign n33616 = n10549 & n33615 ;
  assign n33617 = n347 & n32812 ;
  assign n33618 = n13664 ^ n12680 ^ 1'b0 ;
  assign n33619 = n26851 ^ n26173 ^ n16240 ;
  assign n33620 = n5707 & ~n14593 ;
  assign n33621 = n33620 ^ n4007 ^ 1'b0 ;
  assign n33622 = ( n509 & n33619 ) | ( n509 & n33621 ) | ( n33619 & n33621 ) ;
  assign n33625 = ~n3518 & n5273 ;
  assign n33623 = n3440 | n31983 ;
  assign n33624 = n28010 & ~n33623 ;
  assign n33626 = n33625 ^ n33624 ^ n24945 ;
  assign n33627 = ~n3362 & n7332 ;
  assign n33628 = ~n21620 & n33627 ;
  assign n33629 = n29853 ^ n27886 ^ n6871 ;
  assign n33630 = n33629 ^ n22331 ^ x207 ;
  assign n33631 = n29486 ^ n11619 ^ 1'b0 ;
  assign n33632 = ~n7102 & n8051 ;
  assign n33633 = n18755 ^ n17059 ^ n15938 ;
  assign n33636 = n13736 & ~n32022 ;
  assign n33637 = ( n18286 & n18748 ) | ( n18286 & n33636 ) | ( n18748 & n33636 ) ;
  assign n33638 = n33637 ^ n23580 ^ n3569 ;
  assign n33634 = n27620 ^ n10304 ^ n9864 ;
  assign n33635 = n6865 & n33634 ;
  assign n33639 = n33638 ^ n33635 ^ 1'b0 ;
  assign n33640 = n32685 ^ n23711 ^ 1'b0 ;
  assign n33641 = n5455 & ~n33640 ;
  assign n33642 = n8062 & n13636 ;
  assign n33643 = ( n2750 & n5583 ) | ( n2750 & n31274 ) | ( n5583 & n31274 ) ;
  assign n33644 = n33643 ^ n9754 ^ 1'b0 ;
  assign n33645 = n24033 & ~n33644 ;
  assign n33646 = n33645 ^ n10532 ^ n5020 ;
  assign n33647 = n33642 | n33646 ;
  assign n33648 = n11514 | n33647 ;
  assign n33649 = n7280 & n24182 ;
  assign n33650 = n1016 & n6673 ;
  assign n33651 = n3047 & ~n33650 ;
  assign n33652 = n33651 ^ n25630 ^ 1'b0 ;
  assign n33653 = n10659 & n29042 ;
  assign n33654 = n33653 ^ n9344 ^ 1'b0 ;
  assign n33655 = ( ~x94 & n3248 ) | ( ~x94 & n6413 ) | ( n3248 & n6413 ) ;
  assign n33656 = n33655 ^ n18605 ^ n8111 ;
  assign n33657 = n26948 & n32972 ;
  assign n33658 = n33657 ^ n22818 ^ 1'b0 ;
  assign n33659 = n33656 & ~n33658 ;
  assign n33660 = ~n2735 & n6323 ;
  assign n33661 = n29033 & n33660 ;
  assign n33662 = n14199 ^ n6550 ^ n3999 ;
  assign n33663 = n3392 | n7311 ;
  assign n33664 = n5467 & ~n33663 ;
  assign n33665 = n33664 ^ n27691 ^ 1'b0 ;
  assign n33666 = n22261 & n33665 ;
  assign n33667 = n29775 ^ n24732 ^ 1'b0 ;
  assign n33669 = n16247 ^ n13849 ^ 1'b0 ;
  assign n33670 = n2799 | n33669 ;
  assign n33668 = ( n1351 & n25073 ) | ( n1351 & n28418 ) | ( n25073 & n28418 ) ;
  assign n33671 = n33670 ^ n33668 ^ n4522 ;
  assign n33672 = ( n7885 & n18423 ) | ( n7885 & n33671 ) | ( n18423 & n33671 ) ;
  assign n33673 = n4111 | n13025 ;
  assign n33674 = n33673 ^ n10665 ^ 1'b0 ;
  assign n33675 = n12108 | n33674 ;
  assign n33676 = n33675 ^ n18604 ^ n6840 ;
  assign n33677 = ~n2651 & n14885 ;
  assign n33678 = n33677 ^ n5515 ^ 1'b0 ;
  assign n33679 = ( n25416 & n31748 ) | ( n25416 & ~n33678 ) | ( n31748 & ~n33678 ) ;
  assign n33680 = n19043 ^ n13190 ^ 1'b0 ;
  assign n33681 = n10108 & ~n33680 ;
  assign n33682 = n15963 ^ n12157 ^ 1'b0 ;
  assign n33683 = n33681 & ~n33682 ;
  assign n33684 = n33683 ^ n2198 ^ 1'b0 ;
  assign n33688 = n12642 ^ n6035 ^ n1251 ;
  assign n33689 = ( ~n4214 & n7172 ) | ( ~n4214 & n33688 ) | ( n7172 & n33688 ) ;
  assign n33685 = n30217 ^ n10897 ^ 1'b0 ;
  assign n33686 = n1648 & ~n33685 ;
  assign n33687 = n2681 & n33686 ;
  assign n33690 = n33689 ^ n33687 ^ n25331 ;
  assign n33692 = ( ~n10415 & n18892 ) | ( ~n10415 & n26296 ) | ( n18892 & n26296 ) ;
  assign n33691 = ~n3625 & n5268 ;
  assign n33693 = n33692 ^ n33691 ^ 1'b0 ;
  assign n33696 = n14112 & n19290 ;
  assign n33697 = n33696 ^ n7213 ^ 1'b0 ;
  assign n33698 = n33697 ^ n32510 ^ 1'b0 ;
  assign n33694 = ~n4237 & n7590 ;
  assign n33695 = ~n20443 & n33694 ;
  assign n33699 = n33698 ^ n33695 ^ 1'b0 ;
  assign n33700 = n16491 & ~n28745 ;
  assign n33701 = n3588 & n33700 ;
  assign n33702 = n18569 ^ n4855 ^ 1'b0 ;
  assign n33703 = n9212 & ~n33702 ;
  assign n33704 = n25765 & n33703 ;
  assign n33705 = n23624 & ~n33704 ;
  assign n33706 = ( n14497 & n16434 ) | ( n14497 & ~n17665 ) | ( n16434 & ~n17665 ) ;
  assign n33707 = n835 ^ n454 ^ 1'b0 ;
  assign n33708 = n33707 ^ n29469 ^ 1'b0 ;
  assign n33709 = n29900 ^ n7212 ^ 1'b0 ;
  assign n33710 = n9155 & n9947 ;
  assign n33711 = n33710 ^ n27347 ^ 1'b0 ;
  assign n33712 = ~n4812 & n33711 ;
  assign n33713 = n29003 ^ n24606 ^ n16601 ;
  assign n33714 = n8700 | n13917 ;
  assign n33715 = n10363 ^ x174 ^ 1'b0 ;
  assign n33716 = n3426 & n20105 ;
  assign n33717 = ~n33715 & n33716 ;
  assign n33718 = n13203 & n29381 ;
  assign n33719 = n13593 & n14391 ;
  assign n33720 = n31993 ^ n15607 ^ n11642 ;
  assign n33721 = n11560 ^ n730 ^ x15 ;
  assign n33722 = n33721 ^ n9623 ^ n3717 ;
  assign n33723 = ( n7693 & n28679 ) | ( n7693 & n33722 ) | ( n28679 & n33722 ) ;
  assign n33724 = n22213 ^ n16020 ^ n10106 ;
  assign n33725 = n15214 ^ n3364 ^ 1'b0 ;
  assign n33726 = n3537 & n32687 ;
  assign n33727 = n33726 ^ n9925 ^ 1'b0 ;
  assign n33728 = n2898 & n10490 ;
  assign n33729 = n27915 ^ n23050 ^ 1'b0 ;
  assign n33730 = ~n33728 & n33729 ;
  assign n33731 = ( n3249 & n10380 ) | ( n3249 & ~n33730 ) | ( n10380 & ~n33730 ) ;
  assign n33732 = ~n9087 & n21795 ;
  assign n33733 = n16873 | n26806 ;
  assign n33734 = ( ~n25421 & n30355 ) | ( ~n25421 & n33733 ) | ( n30355 & n33733 ) ;
  assign n33735 = n12374 & ~n29834 ;
  assign n33736 = n33735 ^ n11805 ^ 1'b0 ;
  assign n33737 = n33736 ^ n29916 ^ n6471 ;
  assign n33738 = n33737 ^ n33044 ^ n4082 ;
  assign n33739 = n25940 & ~n33738 ;
  assign n33740 = n11132 ^ n1887 ^ 1'b0 ;
  assign n33741 = n10008 & ~n33740 ;
  assign n33742 = n7759 & ~n33741 ;
  assign n33743 = n21600 ^ n13705 ^ 1'b0 ;
  assign n33744 = n29852 | n33743 ;
  assign n33745 = n9266 & ~n33744 ;
  assign n33746 = n19896 ^ n4241 ^ 1'b0 ;
  assign n33749 = ( n3278 & n6950 ) | ( n3278 & n15573 ) | ( n6950 & n15573 ) ;
  assign n33747 = ( ~n995 & n1241 ) | ( ~n995 & n15059 ) | ( n1241 & n15059 ) ;
  assign n33748 = n33747 ^ n26365 ^ n5081 ;
  assign n33750 = n33749 ^ n33748 ^ 1'b0 ;
  assign n33751 = n33746 & n33750 ;
  assign n33752 = n14877 & ~n33751 ;
  assign n33753 = n23292 ^ n9895 ^ 1'b0 ;
  assign n33754 = n9016 | n33753 ;
  assign n33755 = n33754 ^ n5295 ^ 1'b0 ;
  assign n33756 = n18841 & n33755 ;
  assign n33758 = n24620 ^ n24070 ^ n4160 ;
  assign n33757 = n3217 & n4874 ;
  assign n33759 = n33758 ^ n33757 ^ 1'b0 ;
  assign n33760 = n9593 & ~n10259 ;
  assign n33761 = n24606 & n33760 ;
  assign n33762 = n33761 ^ n13115 ^ n5685 ;
  assign n33763 = ( n1574 & n11313 ) | ( n1574 & n24319 ) | ( n11313 & n24319 ) ;
  assign n33764 = ( ~n8606 & n16528 ) | ( ~n8606 & n33763 ) | ( n16528 & n33763 ) ;
  assign n33766 = n27125 ^ n23923 ^ 1'b0 ;
  assign n33767 = ~n17843 & n33766 ;
  assign n33765 = n29659 ^ n18498 ^ 1'b0 ;
  assign n33768 = n33767 ^ n33765 ^ n25698 ;
  assign n33769 = ~n660 & n4040 ;
  assign n33770 = ( n19101 & n29839 ) | ( n19101 & n33769 ) | ( n29839 & n33769 ) ;
  assign n33771 = n4948 ^ n2889 ^ n1232 ;
  assign n33772 = n33771 ^ n6673 ^ n1023 ;
  assign n33773 = n2416 & n33772 ;
  assign n33774 = n33773 ^ n17865 ^ 1'b0 ;
  assign n33775 = ( n16885 & n20357 ) | ( n16885 & ~n22839 ) | ( n20357 & ~n22839 ) ;
  assign n33776 = n7478 & ~n33775 ;
  assign n33777 = n24435 ^ n15966 ^ n2308 ;
  assign n33778 = ( n23804 & n29156 ) | ( n23804 & n33777 ) | ( n29156 & n33777 ) ;
  assign n33779 = ( ~n10357 & n19052 ) | ( ~n10357 & n22138 ) | ( n19052 & n22138 ) ;
  assign n33780 = n24144 ^ n16663 ^ n15751 ;
  assign n33781 = n32699 ^ n32665 ^ n9436 ;
  assign n33782 = n5208 & ~n18929 ;
  assign n33783 = n12535 & n14132 ;
  assign n33784 = ~n33782 & n33783 ;
  assign n33786 = ~n6712 & n29259 ;
  assign n33787 = ~n11023 & n33786 ;
  assign n33788 = ( n3943 & ~n24026 ) | ( n3943 & n33787 ) | ( ~n24026 & n33787 ) ;
  assign n33785 = n9371 & ~n24718 ;
  assign n33789 = n33788 ^ n33785 ^ 1'b0 ;
  assign n33793 = n15086 ^ n12889 ^ 1'b0 ;
  assign n33794 = n33793 ^ n23576 ^ 1'b0 ;
  assign n33795 = n6539 & ~n33794 ;
  assign n33790 = n3659 & n13594 ;
  assign n33791 = n8113 ^ n7063 ^ n834 ;
  assign n33792 = n33790 | n33791 ;
  assign n33796 = n33795 ^ n33792 ^ 1'b0 ;
  assign n33797 = n10180 ^ n807 ^ 1'b0 ;
  assign n33798 = n33797 ^ n10457 ^ n1122 ;
  assign n33799 = n24075 | n24937 ;
  assign n33800 = ~n12984 & n27904 ;
  assign n33801 = n10559 & ~n33800 ;
  assign n33802 = n33801 ^ n16444 ^ 1'b0 ;
  assign n33803 = n27187 & n33802 ;
  assign n33804 = n3897 & n6256 ;
  assign n33805 = n33804 ^ n25741 ^ 1'b0 ;
  assign n33806 = n19904 ^ n13565 ^ n12415 ;
  assign n33807 = ( ~n22820 & n33304 ) | ( ~n22820 & n33806 ) | ( n33304 & n33806 ) ;
  assign n33808 = n26378 ^ n3408 ^ 1'b0 ;
  assign n33809 = ~n10733 & n21340 ;
  assign n33810 = n33809 ^ n31019 ^ 1'b0 ;
  assign n33811 = n24447 & ~n33810 ;
  assign n33812 = n33811 ^ n428 ^ 1'b0 ;
  assign n33813 = ~n33010 & n33812 ;
  assign n33814 = ( n26263 & n29380 ) | ( n26263 & ~n33813 ) | ( n29380 & ~n33813 ) ;
  assign n33815 = n13773 ^ n8452 ^ n6305 ;
  assign n33816 = ( n24718 & ~n26851 ) | ( n24718 & n33815 ) | ( ~n26851 & n33815 ) ;
  assign n33817 = ~n32027 & n33816 ;
  assign n33820 = n5044 | n7381 ;
  assign n33818 = n13587 ^ n10162 ^ n2260 ;
  assign n33819 = n33818 ^ n11618 ^ n6489 ;
  assign n33821 = n33820 ^ n33819 ^ 1'b0 ;
  assign n33822 = ~n12559 & n26571 ;
  assign n33823 = n33822 ^ n14744 ^ 1'b0 ;
  assign n33824 = n8771 & n33823 ;
  assign n33825 = ~n8037 & n33824 ;
  assign n33826 = n18543 ^ n11108 ^ 1'b0 ;
  assign n33827 = ~n33825 & n33826 ;
  assign n33828 = n16360 ^ n2589 ^ 1'b0 ;
  assign n33829 = ~n15955 & n33828 ;
  assign n33830 = n14309 & n20938 ;
  assign n33831 = n11461 ^ n626 ^ 1'b0 ;
  assign n33832 = ( n7618 & ~n27324 ) | ( n7618 & n33831 ) | ( ~n27324 & n33831 ) ;
  assign n33833 = n9593 | n18444 ;
  assign n33834 = ~n352 & n32453 ;
  assign n33838 = ( n6981 & n11884 ) | ( n6981 & ~n25988 ) | ( n11884 & ~n25988 ) ;
  assign n33835 = ( ~n2718 & n13183 ) | ( ~n2718 & n13430 ) | ( n13183 & n13430 ) ;
  assign n33836 = n3187 & n30825 ;
  assign n33837 = n33835 | n33836 ;
  assign n33839 = n33838 ^ n33837 ^ 1'b0 ;
  assign n33840 = n6056 | n14258 ;
  assign n33841 = n33840 ^ n4263 ^ 1'b0 ;
  assign n33842 = n20709 ^ n10941 ^ n9010 ;
  assign n33843 = ( n3729 & n19101 ) | ( n3729 & n33842 ) | ( n19101 & n33842 ) ;
  assign n33844 = n32479 ^ n21602 ^ 1'b0 ;
  assign n33845 = ~n33843 & n33844 ;
  assign n33854 = ~n9877 & n20449 ;
  assign n33848 = n8092 ^ n2614 ^ 1'b0 ;
  assign n33849 = n10457 & ~n33848 ;
  assign n33850 = n5025 ^ n3606 ^ 1'b0 ;
  assign n33851 = n6052 | n33850 ;
  assign n33852 = ( ~n6497 & n12898 ) | ( ~n6497 & n33851 ) | ( n12898 & n33851 ) ;
  assign n33853 = ( ~n17774 & n33849 ) | ( ~n17774 & n33852 ) | ( n33849 & n33852 ) ;
  assign n33846 = n6146 | n8612 ;
  assign n33847 = n30040 & ~n33846 ;
  assign n33855 = n33854 ^ n33853 ^ n33847 ;
  assign n33856 = ( n9928 & ~n20686 ) | ( n9928 & n21271 ) | ( ~n20686 & n21271 ) ;
  assign n33858 = n15561 | n19854 ;
  assign n33857 = n5596 & n25674 ;
  assign n33859 = n33858 ^ n33857 ^ n17120 ;
  assign n33860 = ( n13781 & ~n33856 ) | ( n13781 & n33859 ) | ( ~n33856 & n33859 ) ;
  assign n33861 = ( n12188 & n17012 ) | ( n12188 & n24792 ) | ( n17012 & n24792 ) ;
  assign n33862 = ( n707 & ~n4132 ) | ( n707 & n8703 ) | ( ~n4132 & n8703 ) ;
  assign n33863 = n31976 | n33862 ;
  assign n33864 = n33863 ^ n3977 ^ 1'b0 ;
  assign n33865 = n1199 & ~n12017 ;
  assign n33866 = n33865 ^ n26143 ^ 1'b0 ;
  assign n33867 = n16855 & ~n33866 ;
  assign n33868 = ~n25489 & n33867 ;
  assign n33869 = n2924 & n33868 ;
  assign n33870 = ( n8937 & n25322 ) | ( n8937 & n31965 ) | ( n25322 & n31965 ) ;
  assign n33871 = n33870 ^ n8013 ^ 1'b0 ;
  assign n33872 = n27334 | n33871 ;
  assign n33873 = n2362 ^ n315 ^ 1'b0 ;
  assign n33874 = n26202 | n33873 ;
  assign n33875 = n19265 | n33874 ;
  assign n33876 = n1364 | n4863 ;
  assign n33877 = n15059 ^ n9010 ^ n6014 ;
  assign n33878 = n11328 & n33877 ;
  assign n33879 = ~n32171 & n33878 ;
  assign n33881 = n17604 & ~n29062 ;
  assign n33880 = n1791 & ~n31242 ;
  assign n33882 = n33881 ^ n33880 ^ 1'b0 ;
  assign n33883 = n25294 ^ n313 ^ 1'b0 ;
  assign n33884 = n33883 ^ n20330 ^ n7311 ;
  assign n33885 = n33884 ^ n7378 ^ 1'b0 ;
  assign n33886 = n2571 & n32672 ;
  assign n33887 = n33886 ^ n18730 ^ 1'b0 ;
  assign n33888 = n16807 | n33887 ;
  assign n33889 = n2553 | n33888 ;
  assign n33890 = n33885 | n33889 ;
  assign n33891 = ( ~n6481 & n9058 ) | ( ~n6481 & n22877 ) | ( n9058 & n22877 ) ;
  assign n33892 = n5513 ^ n5188 ^ n586 ;
  assign n33893 = n33892 ^ n24428 ^ n16530 ;
  assign n33894 = n32513 ^ n31108 ^ n1617 ;
  assign n33895 = n12512 & ~n21861 ;
  assign n33896 = ~x205 & n33895 ;
  assign n33897 = ( ~n16472 & n29231 ) | ( ~n16472 & n33896 ) | ( n29231 & n33896 ) ;
  assign n33898 = n13021 ^ n3807 ^ n705 ;
  assign n33899 = n3618 & ~n33898 ;
  assign n33900 = ( n28573 & ~n32448 ) | ( n28573 & n33899 ) | ( ~n32448 & n33899 ) ;
  assign n33901 = ( ~x89 & n3511 ) | ( ~x89 & n9969 ) | ( n3511 & n9969 ) ;
  assign n33902 = n33900 & n33901 ;
  assign n33903 = n28348 ^ n19955 ^ n407 ;
  assign n33904 = n33903 ^ n18858 ^ 1'b0 ;
  assign n33905 = n27063 ^ n15579 ^ n2095 ;
  assign n33906 = ( n358 & n1050 ) | ( n358 & ~n24136 ) | ( n1050 & ~n24136 ) ;
  assign n33907 = n6776 & ~n6929 ;
  assign n33908 = ~n3806 & n33907 ;
  assign n33909 = n33908 ^ n6495 ^ 1'b0 ;
  assign n33910 = n17220 & ~n28801 ;
  assign n33911 = n15979 & ~n22339 ;
  assign n33912 = n33911 ^ x83 ^ 1'b0 ;
  assign n33913 = n33741 ^ n27689 ^ n5703 ;
  assign n33914 = n13306 ^ n10537 ^ 1'b0 ;
  assign n33915 = n895 & n33914 ;
  assign n33916 = n33913 & n33915 ;
  assign n33917 = ~n11123 & n33916 ;
  assign n33918 = n16343 ^ n10790 ^ n10706 ;
  assign n33920 = n2607 ^ x71 ^ 1'b0 ;
  assign n33919 = n2377 | n17172 ;
  assign n33921 = n33920 ^ n33919 ^ 1'b0 ;
  assign n33922 = n28409 & ~n33921 ;
  assign n33923 = n1636 & n15250 ;
  assign n33924 = n29288 ^ n23386 ^ 1'b0 ;
  assign n33925 = n29564 & ~n33924 ;
  assign n33926 = ( n754 & ~n31993 ) | ( n754 & n33117 ) | ( ~n31993 & n33117 ) ;
  assign n33927 = n33926 ^ n33581 ^ n10060 ;
  assign n33928 = n26847 ^ n2265 ^ 1'b0 ;
  assign n33929 = n20599 & ~n29055 ;
  assign n33930 = n33929 ^ n30553 ^ 1'b0 ;
  assign n33931 = ( n24482 & n33928 ) | ( n24482 & ~n33930 ) | ( n33928 & ~n33930 ) ;
  assign n33932 = ~n1614 & n5119 ;
  assign n33933 = n33932 ^ n29007 ^ n7901 ;
  assign n33934 = ( n5312 & n29317 ) | ( n5312 & n33933 ) | ( n29317 & n33933 ) ;
  assign n33935 = n5092 ^ n3532 ^ 1'b0 ;
  assign n33936 = ( n15364 & n19957 ) | ( n15364 & ~n32512 ) | ( n19957 & ~n32512 ) ;
  assign n33937 = n29320 & ~n33936 ;
  assign n33938 = n33937 ^ n5281 ^ 1'b0 ;
  assign n33939 = n2117 | n2827 ;
  assign n33940 = n25630 ^ n20613 ^ 1'b0 ;
  assign n33941 = ~n33939 & n33940 ;
  assign n33942 = ~n33938 & n33941 ;
  assign n33943 = ~n3439 & n33942 ;
  assign n33944 = ~n7051 & n19703 ;
  assign n33945 = n11827 ^ n3283 ^ n3202 ;
  assign n33946 = n10638 & n28175 ;
  assign n33947 = ( x90 & n33945 ) | ( x90 & ~n33946 ) | ( n33945 & ~n33946 ) ;
  assign n33948 = n22498 ^ n6001 ^ 1'b0 ;
  assign n33949 = n2637 & ~n19220 ;
  assign n33950 = n33949 ^ n8802 ^ 1'b0 ;
  assign n33951 = n33950 ^ n25913 ^ n17043 ;
  assign n33955 = ( n6594 & n12891 ) | ( n6594 & n22278 ) | ( n12891 & n22278 ) ;
  assign n33953 = n26273 ^ n12289 ^ 1'b0 ;
  assign n33952 = n16918 ^ n16338 ^ 1'b0 ;
  assign n33954 = n33953 ^ n33952 ^ n16330 ;
  assign n33956 = n33955 ^ n33954 ^ 1'b0 ;
  assign n33960 = ( ~n10015 & n10786 ) | ( ~n10015 & n10861 ) | ( n10786 & n10861 ) ;
  assign n33957 = n4333 ^ n1620 ^ n1205 ;
  assign n33958 = ( n7233 & ~n15057 ) | ( n7233 & n33957 ) | ( ~n15057 & n33957 ) ;
  assign n33959 = n20182 | n33958 ;
  assign n33961 = n33960 ^ n33959 ^ 1'b0 ;
  assign n33962 = n31833 ^ n10633 ^ 1'b0 ;
  assign n33963 = n16821 ^ n12483 ^ 1'b0 ;
  assign n33964 = n6318 | n33963 ;
  assign n33965 = n17327 & n20490 ;
  assign n33966 = ~n5638 & n33965 ;
  assign n33967 = n33966 ^ n10538 ^ 1'b0 ;
  assign n33968 = n9872 | n33967 ;
  assign n33969 = n28085 ^ n2648 ^ 1'b0 ;
  assign n33970 = n3887 & n21949 ;
  assign n33971 = n33970 ^ n14543 ^ 1'b0 ;
  assign n33972 = ( n26208 & n33969 ) | ( n26208 & n33971 ) | ( n33969 & n33971 ) ;
  assign n33973 = x224 & ~n5309 ;
  assign n33974 = n33973 ^ n14148 ^ 1'b0 ;
  assign n33975 = n21063 | n33974 ;
  assign n33976 = n33975 ^ n8357 ^ 1'b0 ;
  assign n33977 = n17352 ^ n550 ^ 1'b0 ;
  assign n33978 = ( ~n1600 & n8396 ) | ( ~n1600 & n16745 ) | ( n8396 & n16745 ) ;
  assign n33979 = ~n33977 & n33978 ;
  assign n33980 = n3210 ^ n1833 ^ 1'b0 ;
  assign n33981 = ~n18266 & n33980 ;
  assign n33982 = n33981 ^ n13581 ^ n8306 ;
  assign n33983 = n25396 ^ n14260 ^ n9601 ;
  assign n33984 = n6932 ^ n5817 ^ 1'b0 ;
  assign n33985 = ~n4403 & n33984 ;
  assign n33986 = n11364 & n33985 ;
  assign n33987 = n33986 ^ n865 ^ 1'b0 ;
  assign n33988 = n33987 ^ n18929 ^ 1'b0 ;
  assign n33989 = ( ~n18374 & n33983 ) | ( ~n18374 & n33988 ) | ( n33983 & n33988 ) ;
  assign n33990 = ( n4611 & n16314 ) | ( n4611 & ~n25746 ) | ( n16314 & ~n25746 ) ;
  assign n33991 = n16705 & ~n33990 ;
  assign n33993 = n8985 ^ n2036 ^ n705 ;
  assign n33994 = n33636 ^ n4572 ^ 1'b0 ;
  assign n33995 = n33993 & n33994 ;
  assign n33992 = n19511 ^ n11737 ^ n5500 ;
  assign n33996 = n33995 ^ n33992 ^ n3561 ;
  assign n33997 = n33996 ^ n31417 ^ n15976 ;
  assign n33998 = n28237 ^ n15211 ^ 1'b0 ;
  assign n33999 = ~n2775 & n9765 ;
  assign n34000 = n27162 ^ n15088 ^ 1'b0 ;
  assign n34001 = ~n33999 & n34000 ;
  assign n34002 = n7047 & n9246 ;
  assign n34003 = n34002 ^ n9167 ^ 1'b0 ;
  assign n34004 = n10069 & n27255 ;
  assign n34005 = n10138 & n34004 ;
  assign n34008 = n9669 ^ n6562 ^ 1'b0 ;
  assign n34009 = n15883 & ~n34008 ;
  assign n34006 = n25515 ^ n8646 ^ 1'b0 ;
  assign n34007 = n6839 & n34006 ;
  assign n34010 = n34009 ^ n34007 ^ n7410 ;
  assign n34011 = ( n12346 & ~n23545 ) | ( n12346 & n34010 ) | ( ~n23545 & n34010 ) ;
  assign n34012 = n17940 ^ n17819 ^ n12197 ;
  assign n34013 = n28675 ^ n6095 ^ 1'b0 ;
  assign n34014 = n32586 | n34013 ;
  assign n34015 = ( n34011 & n34012 ) | ( n34011 & n34014 ) | ( n34012 & n34014 ) ;
  assign n34016 = n34015 ^ n28837 ^ n14725 ;
  assign n34017 = ( n9526 & ~n12206 ) | ( n9526 & n27617 ) | ( ~n12206 & n27617 ) ;
  assign n34018 = ~n3394 & n34017 ;
  assign n34019 = ( ~n1585 & n16078 ) | ( ~n1585 & n34018 ) | ( n16078 & n34018 ) ;
  assign n34020 = n17368 ^ n13715 ^ n1378 ;
  assign n34021 = ( n2727 & n5071 ) | ( n2727 & n5258 ) | ( n5071 & n5258 ) ;
  assign n34022 = n17514 & ~n25624 ;
  assign n34023 = n1400 & n10382 ;
  assign n34024 = n3650 & n34023 ;
  assign n34028 = n5604 & n23104 ;
  assign n34029 = n16620 & n34028 ;
  assign n34030 = n34029 ^ n14744 ^ n7579 ;
  assign n34025 = n5498 & ~n29636 ;
  assign n34026 = n34025 ^ n29289 ^ 1'b0 ;
  assign n34027 = n18182 | n34026 ;
  assign n34031 = n34030 ^ n34027 ^ 1'b0 ;
  assign n34034 = x254 & ~n21532 ;
  assign n34035 = n7891 & n34034 ;
  assign n34032 = ~n15521 & n17024 ;
  assign n34033 = n34032 ^ n15137 ^ 1'b0 ;
  assign n34036 = n34035 ^ n34033 ^ 1'b0 ;
  assign n34037 = n12313 & n18156 ;
  assign n34038 = n34037 ^ n16836 ^ 1'b0 ;
  assign n34039 = ( n893 & n6653 ) | ( n893 & ~n34038 ) | ( n6653 & ~n34038 ) ;
  assign n34040 = n15126 ^ n10149 ^ 1'b0 ;
  assign n34041 = n22294 ^ n8311 ^ 1'b0 ;
  assign n34042 = x23 & ~n34041 ;
  assign n34043 = n7703 | n12493 ;
  assign n34044 = n14001 & ~n34043 ;
  assign n34045 = n34044 ^ n23770 ^ 1'b0 ;
  assign n34046 = ~n8577 & n34045 ;
  assign n34047 = ( n3182 & ~n34042 ) | ( n3182 & n34046 ) | ( ~n34042 & n34046 ) ;
  assign n34048 = n33383 ^ n8406 ^ n1721 ;
  assign n34049 = n29280 & n34048 ;
  assign n34050 = n22390 ^ n21262 ^ 1'b0 ;
  assign n34051 = n34050 ^ n11489 ^ 1'b0 ;
  assign n34052 = n6512 | n23310 ;
  assign n34053 = n19017 ^ n18112 ^ n6621 ;
  assign n34054 = n34053 ^ n13867 ^ n11426 ;
  assign n34055 = ~n6220 & n11328 ;
  assign n34056 = n34055 ^ n19875 ^ 1'b0 ;
  assign n34057 = n34056 ^ n12701 ^ 1'b0 ;
  assign n34058 = n1673 | n9473 ;
  assign n34059 = n7372 | n34058 ;
  assign n34060 = n15338 & ~n34043 ;
  assign n34061 = n23852 & n34060 ;
  assign n34062 = x69 & ~n14793 ;
  assign n34063 = n20881 & n34062 ;
  assign n34064 = n9160 & n11271 ;
  assign n34065 = n34064 ^ n28816 ^ n24798 ;
  assign n34067 = x208 & ~n3070 ;
  assign n34068 = n34067 ^ n12358 ^ 1'b0 ;
  assign n34066 = n15663 | n27084 ;
  assign n34069 = n34068 ^ n34066 ^ 1'b0 ;
  assign n34070 = n34069 ^ n25079 ^ n8669 ;
  assign n34071 = n8849 ^ n3848 ^ 1'b0 ;
  assign n34072 = n34071 ^ n19961 ^ 1'b0 ;
  assign n34073 = n8436 & ~n34072 ;
  assign n34074 = n20540 ^ n15089 ^ 1'b0 ;
  assign n34075 = n13196 & n25990 ;
  assign n34076 = ~n34074 & n34075 ;
  assign n34077 = n3996 ^ n3071 ^ 1'b0 ;
  assign n34078 = n20240 ^ n10924 ^ 1'b0 ;
  assign n34079 = n1886 & n34078 ;
  assign n34080 = n34077 & n34079 ;
  assign n34081 = ( n20962 & n29632 ) | ( n20962 & n34080 ) | ( n29632 & n34080 ) ;
  assign n34082 = n34081 ^ n15105 ^ n4078 ;
  assign n34083 = ( n1985 & n3886 ) | ( n1985 & n22178 ) | ( n3886 & n22178 ) ;
  assign n34084 = ( n10223 & ~n11689 ) | ( n10223 & n17463 ) | ( ~n11689 & n17463 ) ;
  assign n34085 = n2195 ^ n2049 ^ 1'b0 ;
  assign n34086 = ( n865 & n8193 ) | ( n865 & ~n34085 ) | ( n8193 & ~n34085 ) ;
  assign n34087 = n28462 ^ n18752 ^ n285 ;
  assign n34088 = ( ~n16660 & n34086 ) | ( ~n16660 & n34087 ) | ( n34086 & n34087 ) ;
  assign n34089 = ~n21965 & n34088 ;
  assign n34090 = n1918 | n34089 ;
  assign n34091 = n21263 & ~n28750 ;
  assign n34092 = ~n3489 & n34091 ;
  assign n34093 = n34092 ^ n9418 ^ 1'b0 ;
  assign n34094 = n30893 & n34093 ;
  assign n34095 = n8013 ^ n5947 ^ 1'b0 ;
  assign n34096 = n12146 ^ n536 ^ 1'b0 ;
  assign n34098 = ( n2398 & n16645 ) | ( n2398 & n20610 ) | ( n16645 & n20610 ) ;
  assign n34097 = ( n1157 & n1516 ) | ( n1157 & n21174 ) | ( n1516 & n21174 ) ;
  assign n34099 = n34098 ^ n34097 ^ 1'b0 ;
  assign n34100 = n34096 | n34099 ;
  assign n34101 = n20511 ^ n1585 ^ 1'b0 ;
  assign n34102 = n6092 & ~n34101 ;
  assign n34103 = ~n4121 & n16893 ;
  assign n34104 = ~n23528 & n34103 ;
  assign n34105 = n34104 ^ n30626 ^ n516 ;
  assign n34106 = n13581 ^ n5111 ^ 1'b0 ;
  assign n34107 = n5042 & n34106 ;
  assign n34108 = n34107 ^ n29914 ^ 1'b0 ;
  assign n34109 = n30955 & ~n33999 ;
  assign n34110 = n11944 ^ n2444 ^ 1'b0 ;
  assign n34111 = ~n922 & n34110 ;
  assign n34112 = n16330 ^ n6521 ^ n4984 ;
  assign n34113 = n34111 & ~n34112 ;
  assign n34116 = ( n2098 & ~n18239 ) | ( n2098 & n26343 ) | ( ~n18239 & n26343 ) ;
  assign n34114 = ~n492 & n33946 ;
  assign n34115 = n34114 ^ n7369 ^ 1'b0 ;
  assign n34117 = n34116 ^ n34115 ^ 1'b0 ;
  assign n34118 = n25340 ^ n24401 ^ 1'b0 ;
  assign n34119 = n31878 ^ n12032 ^ 1'b0 ;
  assign n34121 = ( n3988 & n6553 ) | ( n3988 & n22111 ) | ( n6553 & n22111 ) ;
  assign n34120 = n5118 | n24509 ;
  assign n34122 = n34121 ^ n34120 ^ 1'b0 ;
  assign n34123 = n7989 ^ n6463 ^ x175 ;
  assign n34124 = n8791 | n34123 ;
  assign n34125 = n34124 ^ n2154 ^ 1'b0 ;
  assign n34126 = n23213 & ~n34125 ;
  assign n34127 = n34122 & n34126 ;
  assign n34128 = n25749 | n30899 ;
  assign n34129 = n3037 & ~n34128 ;
  assign n34130 = ( n1756 & ~n1830 ) | ( n1756 & n25565 ) | ( ~n1830 & n25565 ) ;
  assign n34131 = n11327 & ~n34130 ;
  assign n34132 = n34129 & n34131 ;
  assign n34133 = n25438 ^ n10977 ^ n7504 ;
  assign n34134 = n18784 ^ n13741 ^ 1'b0 ;
  assign n34135 = n34133 | n34134 ;
  assign n34136 = ( n3798 & n21235 ) | ( n3798 & n34135 ) | ( n21235 & n34135 ) ;
  assign n34137 = ( n14339 & n28642 ) | ( n14339 & n34136 ) | ( n28642 & n34136 ) ;
  assign n34138 = n16883 ^ n10138 ^ 1'b0 ;
  assign n34139 = ( n3247 & ~n26847 ) | ( n3247 & n30580 ) | ( ~n26847 & n30580 ) ;
  assign n34140 = n13899 | n32309 ;
  assign n34141 = n14116 | n33629 ;
  assign n34142 = n34141 ^ n20027 ^ 1'b0 ;
  assign n34144 = ~n13382 & n21594 ;
  assign n34145 = ~n4033 & n34144 ;
  assign n34146 = ( n10188 & n31688 ) | ( n10188 & n34145 ) | ( n31688 & n34145 ) ;
  assign n34143 = ~n8130 & n14909 ;
  assign n34147 = n34146 ^ n34143 ^ 1'b0 ;
  assign n34148 = n16626 & ~n20759 ;
  assign n34150 = ( n3399 & n8821 ) | ( n3399 & n8940 ) | ( n8821 & n8940 ) ;
  assign n34149 = n11865 | n21994 ;
  assign n34151 = n34150 ^ n34149 ^ 1'b0 ;
  assign n34152 = ( n3472 & n34148 ) | ( n3472 & n34151 ) | ( n34148 & n34151 ) ;
  assign n34153 = ( x5 & n6768 ) | ( x5 & ~n34152 ) | ( n6768 & ~n34152 ) ;
  assign n34154 = n27426 ^ n7636 ^ 1'b0 ;
  assign n34155 = n34154 ^ n19131 ^ n1424 ;
  assign n34156 = n26324 ^ n7435 ^ n6416 ;
  assign n34157 = n34156 ^ n15554 ^ 1'b0 ;
  assign n34158 = n23633 & n33019 ;
  assign n34159 = n32449 & n34158 ;
  assign n34160 = ~n34157 & n34159 ;
  assign n34161 = ( n3824 & ~n5722 ) | ( n3824 & n15347 ) | ( ~n5722 & n15347 ) ;
  assign n34162 = n34161 ^ n16186 ^ n6736 ;
  assign n34168 = ~n5132 & n8320 ;
  assign n34166 = ~n10054 & n25186 ;
  assign n34167 = n34166 ^ n18612 ^ 1'b0 ;
  assign n34163 = n882 & n15243 ;
  assign n34164 = ~n8854 & n34163 ;
  assign n34165 = n34164 ^ n9766 ^ 1'b0 ;
  assign n34169 = n34168 ^ n34167 ^ n34165 ;
  assign n34170 = n32729 ^ n9613 ^ 1'b0 ;
  assign n34171 = n31552 ^ n12612 ^ 1'b0 ;
  assign n34172 = ( x39 & n6385 ) | ( x39 & n27417 ) | ( n6385 & n27417 ) ;
  assign n34173 = ~n3125 & n34172 ;
  assign n34174 = n34173 ^ n28337 ^ n15683 ;
  assign n34176 = ( n4300 & n5744 ) | ( n4300 & n9895 ) | ( n5744 & n9895 ) ;
  assign n34177 = n34176 ^ n5949 ^ 1'b0 ;
  assign n34178 = ( ~n3399 & n5712 ) | ( ~n3399 & n6903 ) | ( n5712 & n6903 ) ;
  assign n34179 = n3339 & ~n15194 ;
  assign n34180 = ~n34178 & n34179 ;
  assign n34181 = ( n9268 & ~n34177 ) | ( n9268 & n34180 ) | ( ~n34177 & n34180 ) ;
  assign n34175 = n14527 | n24511 ;
  assign n34182 = n34181 ^ n34175 ^ 1'b0 ;
  assign n34183 = n34182 ^ n21087 ^ 1'b0 ;
  assign n34184 = ~n8880 & n22788 ;
  assign n34185 = n34184 ^ n10381 ^ n6121 ;
  assign n34188 = n29725 ^ n15118 ^ 1'b0 ;
  assign n34189 = n12975 | n34188 ;
  assign n34186 = n12300 ^ n9652 ^ 1'b0 ;
  assign n34187 = n3709 & n34186 ;
  assign n34190 = n34189 ^ n34187 ^ n2724 ;
  assign n34191 = n16527 & n31503 ;
  assign n34195 = ~n5166 & n29819 ;
  assign n34192 = ( n2430 & ~n2733 ) | ( n2430 & n7664 ) | ( ~n2733 & n7664 ) ;
  assign n34193 = n34192 ^ n9925 ^ 1'b0 ;
  assign n34194 = n7800 & ~n34193 ;
  assign n34196 = n34195 ^ n34194 ^ 1'b0 ;
  assign n34197 = n32595 ^ n18173 ^ n7899 ;
  assign n34198 = n34197 ^ n7439 ^ 1'b0 ;
  assign n34199 = n10345 | n23205 ;
  assign n34200 = n34199 ^ n2806 ^ 1'b0 ;
  assign n34201 = n34200 ^ n24492 ^ n17333 ;
  assign n34202 = n8665 & n33304 ;
  assign n34203 = n8704 ^ n2393 ^ 1'b0 ;
  assign n34204 = ~n3132 & n34203 ;
  assign n34205 = n6756 ^ n3351 ^ 1'b0 ;
  assign n34206 = n14320 & ~n34205 ;
  assign n34208 = n16741 ^ n10749 ^ 1'b0 ;
  assign n34209 = n13235 | n34208 ;
  assign n34207 = n27698 ^ n24828 ^ n2054 ;
  assign n34210 = n34209 ^ n34207 ^ n8132 ;
  assign n34211 = n22479 ^ n9964 ^ 1'b0 ;
  assign n34212 = n11381 ^ n8957 ^ 1'b0 ;
  assign n34213 = n9132 & ~n11386 ;
  assign n34214 = n3354 ^ x203 ^ 1'b0 ;
  assign n34217 = n11760 ^ n5189 ^ 1'b0 ;
  assign n34218 = n34217 ^ n22324 ^ n18421 ;
  assign n34215 = n18926 ^ n15855 ^ 1'b0 ;
  assign n34216 = n34215 ^ n1777 ^ 1'b0 ;
  assign n34219 = n34218 ^ n34216 ^ n33903 ;
  assign n34220 = n2551 & n20453 ;
  assign n34221 = n13788 & n34220 ;
  assign n34222 = n21999 | n34221 ;
  assign n34223 = n30017 ^ n4635 ^ 1'b0 ;
  assign n34224 = ~n3042 & n9622 ;
  assign n34225 = ~n12274 & n27117 ;
  assign n34226 = ( n1789 & ~n11043 ) | ( n1789 & n12457 ) | ( ~n11043 & n12457 ) ;
  assign n34227 = ~n22593 & n34226 ;
  assign n34228 = ~x222 & n34227 ;
  assign n34239 = n17963 ^ n14914 ^ n7551 ;
  assign n34229 = ( n634 & ~n4611 ) | ( n634 & n11666 ) | ( ~n4611 & n11666 ) ;
  assign n34230 = n13068 | n21366 ;
  assign n34231 = n34230 ^ n9147 ^ 1'b0 ;
  assign n34232 = ( n2567 & ~n13272 ) | ( n2567 & n34231 ) | ( ~n13272 & n34231 ) ;
  assign n34233 = n34232 ^ n17819 ^ n15359 ;
  assign n34234 = ( ~n11675 & n27653 ) | ( ~n11675 & n34233 ) | ( n27653 & n34233 ) ;
  assign n34235 = n22130 ^ n10261 ^ n9126 ;
  assign n34236 = n34235 ^ n8942 ^ n4217 ;
  assign n34237 = n34236 ^ n33361 ^ n20612 ;
  assign n34238 = ( n34229 & n34234 ) | ( n34229 & n34237 ) | ( n34234 & n34237 ) ;
  assign n34240 = n34239 ^ n34238 ^ n23694 ;
  assign n34241 = n14149 ^ n560 ^ 1'b0 ;
  assign n34242 = n32609 ^ x2 ^ 1'b0 ;
  assign n34243 = n34242 ^ n6913 ^ n460 ;
  assign n34244 = ( n10297 & n10661 ) | ( n10297 & n12564 ) | ( n10661 & n12564 ) ;
  assign n34245 = n34244 ^ n29650 ^ 1'b0 ;
  assign n34246 = n34243 & ~n34245 ;
  assign n34247 = n31440 ^ n12590 ^ n4807 ;
  assign n34248 = ( n34241 & n34246 ) | ( n34241 & ~n34247 ) | ( n34246 & ~n34247 ) ;
  assign n34249 = n27771 ^ n19053 ^ n3721 ;
  assign n34250 = ( ~n9611 & n11766 ) | ( ~n9611 & n33284 ) | ( n11766 & n33284 ) ;
  assign n34251 = n34250 ^ n15499 ^ 1'b0 ;
  assign n34252 = n9951 & n21037 ;
  assign n34253 = n16868 ^ n9270 ^ 1'b0 ;
  assign n34254 = ~n13045 & n33854 ;
  assign n34255 = n29519 ^ n28387 ^ 1'b0 ;
  assign n34256 = n1966 & n34255 ;
  assign n34257 = n34256 ^ n20263 ^ 1'b0 ;
  assign n34258 = ( n422 & n4546 ) | ( n422 & n34257 ) | ( n4546 & n34257 ) ;
  assign n34259 = n34258 ^ n14073 ^ 1'b0 ;
  assign n34260 = n9946 & n20485 ;
  assign n34261 = n34260 ^ n19898 ^ n7814 ;
  assign n34263 = n3828 ^ n3821 ^ 1'b0 ;
  assign n34262 = n8008 | n11132 ;
  assign n34264 = n34263 ^ n34262 ^ 1'b0 ;
  assign n34266 = n22522 ^ n18721 ^ n15762 ;
  assign n34267 = n9397 & ~n14704 ;
  assign n34268 = ~n34266 & n34267 ;
  assign n34265 = n31389 ^ n12162 ^ n5592 ;
  assign n34269 = n34268 ^ n34265 ^ n21001 ;
  assign n34271 = n5273 ^ n3517 ^ 1'b0 ;
  assign n34272 = n3005 & n34271 ;
  assign n34270 = n20249 ^ n5764 ^ 1'b0 ;
  assign n34273 = n34272 ^ n34270 ^ n15594 ;
  assign n34274 = n25310 ^ n23516 ^ 1'b0 ;
  assign n34275 = n5838 & ~n19149 ;
  assign n34276 = n29584 | n34275 ;
  assign n34277 = n34274 & ~n34276 ;
  assign n34279 = ( ~n3061 & n6428 ) | ( ~n3061 & n9604 ) | ( n6428 & n9604 ) ;
  assign n34278 = n8565 & n19765 ;
  assign n34280 = n34279 ^ n34278 ^ 1'b0 ;
  assign n34281 = n1026 & ~n28936 ;
  assign n34282 = ~n3044 & n34281 ;
  assign n34283 = n4078 & n17549 ;
  assign n34284 = ( n1034 & n28562 ) | ( n1034 & n34283 ) | ( n28562 & n34283 ) ;
  assign n34285 = n20471 | n30497 ;
  assign n34286 = n34197 & n34285 ;
  assign n34287 = n30158 ^ n16333 ^ n1720 ;
  assign n34288 = n34287 ^ n21294 ^ 1'b0 ;
  assign n34290 = ( n7627 & n8337 ) | ( n7627 & ~n16049 ) | ( n8337 & ~n16049 ) ;
  assign n34289 = n16047 ^ n15288 ^ n8575 ;
  assign n34291 = n34290 ^ n34289 ^ n7618 ;
  assign n34292 = n30045 ^ n17369 ^ n12365 ;
  assign n34293 = n6717 ^ n4156 ^ 1'b0 ;
  assign n34294 = n13677 & n34293 ;
  assign n34295 = n20269 & ~n28702 ;
  assign n34296 = ~n16078 & n34295 ;
  assign n34297 = n27249 & ~n34296 ;
  assign n34298 = n26674 & n34297 ;
  assign n34299 = n12840 & ~n34298 ;
  assign n34300 = ( n1122 & n7642 ) | ( n1122 & ~n15926 ) | ( n7642 & ~n15926 ) ;
  assign n34301 = n34300 ^ n31888 ^ n30009 ;
  assign n34302 = ( n5192 & n7220 ) | ( n5192 & ~n10859 ) | ( n7220 & ~n10859 ) ;
  assign n34303 = n25519 ^ n1924 ^ 1'b0 ;
  assign n34304 = n34303 ^ n12692 ^ n5172 ;
  assign n34305 = ( ~n34255 & n34302 ) | ( ~n34255 & n34304 ) | ( n34302 & n34304 ) ;
  assign n34306 = n30740 ^ n22991 ^ n17358 ;
  assign n34307 = ( n277 & n25149 ) | ( n277 & ~n34306 ) | ( n25149 & ~n34306 ) ;
  assign n34308 = n20273 & ~n21911 ;
  assign n34309 = n840 & ~n5077 ;
  assign n34310 = n34309 ^ n14431 ^ 1'b0 ;
  assign n34311 = n23763 ^ n18281 ^ 1'b0 ;
  assign n34312 = n34310 | n34311 ;
  assign n34313 = n34312 ^ n948 ^ 1'b0 ;
  assign n34314 = n34308 & ~n34313 ;
  assign n34315 = ( n2930 & ~n10524 ) | ( n2930 & n16888 ) | ( ~n10524 & n16888 ) ;
  assign n34316 = n34315 ^ n15472 ^ n6039 ;
  assign n34317 = n13687 ^ n2560 ^ 1'b0 ;
  assign n34318 = n33246 & ~n34317 ;
  assign n34319 = ( n29392 & n31282 ) | ( n29392 & n34318 ) | ( n31282 & n34318 ) ;
  assign n34320 = n16163 | n16214 ;
  assign n34321 = n5049 | n12220 ;
  assign n34322 = ( n7114 & n23022 ) | ( n7114 & n30191 ) | ( n23022 & n30191 ) ;
  assign n34323 = x189 & n34322 ;
  assign n34324 = ~n34321 & n34323 ;
  assign n34325 = n6333 | n30040 ;
  assign n34326 = n3295 | n34325 ;
  assign n34327 = n34326 ^ n25751 ^ 1'b0 ;
  assign n34328 = n18712 ^ n792 ^ 1'b0 ;
  assign n34329 = n9108 & n11644 ;
  assign n34330 = ~n5784 & n34329 ;
  assign n34331 = n34330 ^ n20643 ^ n389 ;
  assign n34332 = n2422 & n7036 ;
  assign n34333 = n34332 ^ n12510 ^ 1'b0 ;
  assign n34334 = n8007 ^ n5242 ^ x204 ;
  assign n34335 = ( ~n33188 & n34333 ) | ( ~n33188 & n34334 ) | ( n34333 & n34334 ) ;
  assign n34336 = n17882 ^ n10526 ^ n3226 ;
  assign n34337 = ( n32993 & ~n34335 ) | ( n32993 & n34336 ) | ( ~n34335 & n34336 ) ;
  assign n34338 = ( n3918 & ~n4450 ) | ( n3918 & n19881 ) | ( ~n4450 & n19881 ) ;
  assign n34339 = n34338 ^ n23680 ^ n20707 ;
  assign n34340 = n1678 & n4676 ;
  assign n34341 = ( ~n13371 & n27175 ) | ( ~n13371 & n34340 ) | ( n27175 & n34340 ) ;
  assign n34342 = n2896 ^ n1822 ^ x101 ;
  assign n34343 = ~n2049 & n12959 ;
  assign n34344 = ( n1230 & n17164 ) | ( n1230 & ~n34343 ) | ( n17164 & ~n34343 ) ;
  assign n34345 = n4729 ^ n1166 ^ 1'b0 ;
  assign n34346 = ( n13305 & n23038 ) | ( n13305 & n34345 ) | ( n23038 & n34345 ) ;
  assign n34347 = n34346 ^ n23968 ^ n11205 ;
  assign n34348 = ( n13596 & n28512 ) | ( n13596 & n28829 ) | ( n28512 & n28829 ) ;
  assign n34349 = ~n5654 & n7958 ;
  assign n34350 = n34349 ^ n963 ^ 1'b0 ;
  assign n34351 = n2757 & n18999 ;
  assign n34352 = ~n30015 & n34351 ;
  assign n34356 = n1824 & ~n5234 ;
  assign n34357 = ( n20685 & ~n25528 ) | ( n20685 & n34356 ) | ( ~n25528 & n34356 ) ;
  assign n34353 = n14078 ^ n12863 ^ n2053 ;
  assign n34354 = n34353 ^ n12996 ^ 1'b0 ;
  assign n34355 = n1534 | n34354 ;
  assign n34358 = n34357 ^ n34355 ^ n5509 ;
  assign n34359 = n7820 | n10969 ;
  assign n34360 = n6901 ^ n748 ^ 1'b0 ;
  assign n34361 = n34360 ^ n19361 ^ n14919 ;
  assign n34362 = ( n6774 & n14980 ) | ( n6774 & ~n28423 ) | ( n14980 & ~n28423 ) ;
  assign n34363 = n30510 ^ n15476 ^ 1'b0 ;
  assign n34364 = n14269 ^ n9833 ^ 1'b0 ;
  assign n34365 = ~n25419 & n34364 ;
  assign n34366 = n29581 ^ n23935 ^ n17653 ;
  assign n34367 = n2864 & n19283 ;
  assign n34368 = ~n19744 & n34367 ;
  assign n34369 = ( n11397 & n16606 ) | ( n11397 & ~n34368 ) | ( n16606 & ~n34368 ) ;
  assign n34370 = ( n2809 & n7979 ) | ( n2809 & n9744 ) | ( n7979 & n9744 ) ;
  assign n34371 = n34370 ^ n15568 ^ n3965 ;
  assign n34372 = n25581 & n30768 ;
  assign n34373 = n8124 & n34372 ;
  assign n34374 = ( n11488 & n15183 ) | ( n11488 & n30777 ) | ( n15183 & n30777 ) ;
  assign n34375 = n8895 & n34374 ;
  assign n34376 = n3920 ^ n2707 ^ n2425 ;
  assign n34377 = n34376 ^ n31161 ^ n16347 ;
  assign n34378 = n34377 ^ n4064 ^ 1'b0 ;
  assign n34379 = ~n24676 & n34378 ;
  assign n34380 = n24283 ^ n4960 ^ n2057 ;
  assign n34383 = n5279 ^ n3394 ^ x158 ;
  assign n34384 = n34383 ^ n32703 ^ n15862 ;
  assign n34381 = n11617 ^ n9039 ^ n1131 ;
  assign n34382 = n34381 ^ n9879 ^ 1'b0 ;
  assign n34385 = n34384 ^ n34382 ^ n24801 ;
  assign n34386 = n11306 & ~n15048 ;
  assign n34387 = n34386 ^ n25440 ^ 1'b0 ;
  assign n34388 = ( n928 & n15347 ) | ( n928 & ~n34387 ) | ( n15347 & ~n34387 ) ;
  assign n34389 = n4638 | n18473 ;
  assign n34390 = ( n15866 & n24394 ) | ( n15866 & n34389 ) | ( n24394 & n34389 ) ;
  assign n34391 = n5562 ^ n2002 ^ 1'b0 ;
  assign n34392 = n16551 & n34391 ;
  assign n34393 = ( n3313 & n8150 ) | ( n3313 & ~n13635 ) | ( n8150 & ~n13635 ) ;
  assign n34394 = n34393 ^ n2048 ^ 1'b0 ;
  assign n34395 = n34392 & n34394 ;
  assign n34396 = n34395 ^ n6815 ^ n826 ;
  assign n34397 = ~n5944 & n18280 ;
  assign n34398 = n3457 & ~n20924 ;
  assign n34399 = ~n28354 & n34398 ;
  assign n34400 = n18306 ^ n16414 ^ n10481 ;
  assign n34401 = n2590 & n34400 ;
  assign n34402 = ( n22260 & n25422 ) | ( n22260 & n26744 ) | ( n25422 & n26744 ) ;
  assign n34403 = ( n9765 & ~n23888 ) | ( n9765 & n34402 ) | ( ~n23888 & n34402 ) ;
  assign n34404 = n10701 ^ n8037 ^ 1'b0 ;
  assign n34405 = n31526 | n34404 ;
  assign n34406 = x100 | n34405 ;
  assign n34407 = n14903 ^ n3586 ^ n2035 ;
  assign n34410 = ( n4720 & n8834 ) | ( n4720 & ~n12495 ) | ( n8834 & ~n12495 ) ;
  assign n34411 = ( n12267 & n17327 ) | ( n12267 & ~n34410 ) | ( n17327 & ~n34410 ) ;
  assign n34412 = n34411 ^ n7820 ^ 1'b0 ;
  assign n34408 = ~n32223 & n34263 ;
  assign n34409 = ( n4220 & ~n24347 ) | ( n4220 & n34408 ) | ( ~n24347 & n34408 ) ;
  assign n34413 = n34412 ^ n34409 ^ n8463 ;
  assign n34414 = ~n633 & n9645 ;
  assign n34415 = n34414 ^ n1381 ^ 1'b0 ;
  assign n34416 = n21606 ^ n19976 ^ n14249 ;
  assign n34417 = n8158 ^ n2327 ^ 1'b0 ;
  assign n34418 = n18795 ^ n14783 ^ 1'b0 ;
  assign n34419 = n5272 & ~n34418 ;
  assign n34420 = n34419 ^ n18508 ^ 1'b0 ;
  assign n34421 = n34417 | n34420 ;
  assign n34422 = n34421 ^ n23280 ^ 1'b0 ;
  assign n34423 = ( n2384 & n3823 ) | ( n2384 & n34422 ) | ( n3823 & n34422 ) ;
  assign n34424 = n26220 ^ n16766 ^ n2971 ;
  assign n34425 = ( n34416 & n34423 ) | ( n34416 & ~n34424 ) | ( n34423 & ~n34424 ) ;
  assign n34426 = n34425 ^ n28724 ^ 1'b0 ;
  assign n34427 = ( n27869 & n28663 ) | ( n27869 & n33856 ) | ( n28663 & n33856 ) ;
  assign n34428 = ( n6416 & n24299 ) | ( n6416 & ~n34427 ) | ( n24299 & ~n34427 ) ;
  assign n34429 = n18070 ^ n6526 ^ x124 ;
  assign n34430 = ~n30789 & n34429 ;
  assign n34431 = n8946 & ~n13272 ;
  assign n34432 = n34431 ^ n18266 ^ 1'b0 ;
  assign n34433 = n34432 ^ n13042 ^ 1'b0 ;
  assign n34434 = ( x6 & ~n18119 ) | ( x6 & n34433 ) | ( ~n18119 & n34433 ) ;
  assign n34435 = ~n9527 & n9857 ;
  assign n34437 = ( ~n2539 & n7157 ) | ( ~n2539 & n13608 ) | ( n7157 & n13608 ) ;
  assign n34436 = n22371 ^ n16935 ^ 1'b0 ;
  assign n34438 = n34437 ^ n34436 ^ n5595 ;
  assign n34439 = n24776 & ~n34438 ;
  assign n34440 = n9353 & n34439 ;
  assign n34441 = n12037 ^ n395 ^ 1'b0 ;
  assign n34442 = ~n27806 & n34441 ;
  assign n34443 = ( n6737 & ~n8119 ) | ( n6737 & n34442 ) | ( ~n8119 & n34442 ) ;
  assign n34444 = n34443 ^ n31827 ^ n13823 ;
  assign n34445 = ( ~n9291 & n11683 ) | ( ~n9291 & n13167 ) | ( n11683 & n13167 ) ;
  assign n34446 = ~n7795 & n34445 ;
  assign n34447 = ~n2330 & n9675 ;
  assign n34448 = n16107 & n34447 ;
  assign n34449 = ( ~n5005 & n9349 ) | ( ~n5005 & n34448 ) | ( n9349 & n34448 ) ;
  assign n34450 = n8276 ^ n4858 ^ 1'b0 ;
  assign n34451 = n14197 & n34450 ;
  assign n34452 = n7897 ^ n5392 ^ 1'b0 ;
  assign n34453 = n34451 & ~n34452 ;
  assign n34454 = ~n5040 & n34453 ;
  assign n34455 = n34454 ^ n3394 ^ 1'b0 ;
  assign n34456 = ( ~n293 & n3900 ) | ( ~n293 & n20237 ) | ( n3900 & n20237 ) ;
  assign n34457 = n34456 ^ n5443 ^ 1'b0 ;
  assign n34458 = n12626 & ~n34457 ;
  assign n34459 = n6182 & ~n14727 ;
  assign n34460 = ~n4574 & n34459 ;
  assign n34461 = ~n34458 & n34460 ;
  assign n34462 = n12372 ^ n536 ^ 1'b0 ;
  assign n34463 = n34462 ^ n27722 ^ n12365 ;
  assign n34464 = n13017 & n18505 ;
  assign n34467 = n1518 ^ n1034 ^ 1'b0 ;
  assign n34468 = ~n5608 & n34467 ;
  assign n34469 = n34468 ^ n1884 ^ 1'b0 ;
  assign n34470 = n19470 & ~n34469 ;
  assign n34465 = ~n2364 & n21720 ;
  assign n34466 = n34465 ^ n2475 ^ 1'b0 ;
  assign n34471 = n34470 ^ n34466 ^ 1'b0 ;
  assign n34472 = ~n761 & n25404 ;
  assign n34473 = ( n12783 & n14951 ) | ( n12783 & n34472 ) | ( n14951 & n34472 ) ;
  assign n34474 = ( n30899 & n34471 ) | ( n30899 & n34473 ) | ( n34471 & n34473 ) ;
  assign n34475 = ( ~n4934 & n5064 ) | ( ~n4934 & n21578 ) | ( n5064 & n21578 ) ;
  assign n34476 = ( n7469 & n9524 ) | ( n7469 & ~n34475 ) | ( n9524 & ~n34475 ) ;
  assign n34477 = n5921 ^ n3956 ^ 1'b0 ;
  assign n34478 = n11071 | n34477 ;
  assign n34479 = ~n12179 & n34478 ;
  assign n34480 = n25199 | n27410 ;
  assign n34481 = n34480 ^ n11642 ^ 1'b0 ;
  assign n34482 = ~n10128 & n34481 ;
  assign n34483 = n34479 & n34482 ;
  assign n34484 = n31546 ^ n26014 ^ 1'b0 ;
  assign n34485 = ~n10549 & n34484 ;
  assign n34486 = ( n9560 & n10104 ) | ( n9560 & ~n19284 ) | ( n10104 & ~n19284 ) ;
  assign n34487 = ( n10936 & n33364 ) | ( n10936 & ~n34486 ) | ( n33364 & ~n34486 ) ;
  assign n34488 = n34487 ^ n4437 ^ 1'b0 ;
  assign n34489 = n2793 & ~n3004 ;
  assign n34490 = n20446 | n34489 ;
  assign n34491 = ~n4846 & n6935 ;
  assign n34492 = n34491 ^ n11157 ^ 1'b0 ;
  assign n34493 = n9564 ^ n2748 ^ 1'b0 ;
  assign n34494 = ~n34492 & n34493 ;
  assign n34495 = n30475 ^ n6182 ^ 1'b0 ;
  assign n34496 = n27834 & ~n34495 ;
  assign n34497 = n34496 ^ n18340 ^ 1'b0 ;
  assign n34498 = n29066 | n34497 ;
  assign n34499 = n27430 ^ n24869 ^ n9148 ;
  assign n34500 = n22729 ^ n13990 ^ n10430 ;
  assign n34501 = ( n9850 & n15579 ) | ( n9850 & ~n34500 ) | ( n15579 & ~n34500 ) ;
  assign n34502 = ( ~n2591 & n10858 ) | ( ~n2591 & n34501 ) | ( n10858 & n34501 ) ;
  assign n34514 = n5200 | n15486 ;
  assign n34515 = n34514 ^ n17812 ^ 1'b0 ;
  assign n34508 = n871 | n15118 ;
  assign n34509 = n10831 & ~n33449 ;
  assign n34510 = n34509 ^ n698 ^ 1'b0 ;
  assign n34511 = ( n17279 & ~n27438 ) | ( n17279 & n34510 ) | ( ~n27438 & n34510 ) ;
  assign n34512 = n34508 | n34511 ;
  assign n34513 = n9075 | n34512 ;
  assign n34503 = ~n11744 & n29380 ;
  assign n34504 = ~n5494 & n34503 ;
  assign n34505 = n29855 | n34504 ;
  assign n34506 = n24382 ^ n8586 ^ n2017 ;
  assign n34507 = ( ~n6230 & n34505 ) | ( ~n6230 & n34506 ) | ( n34505 & n34506 ) ;
  assign n34516 = n34515 ^ n34513 ^ n34507 ;
  assign n34517 = ( n1023 & n1567 ) | ( n1023 & n27697 ) | ( n1567 & n27697 ) ;
  assign n34518 = ( ~n14047 & n18445 ) | ( ~n14047 & n34517 ) | ( n18445 & n34517 ) ;
  assign n34519 = n13181 ^ n6863 ^ 1'b0 ;
  assign n34520 = n5032 & n9464 ;
  assign n34521 = ( n34518 & n34519 ) | ( n34518 & n34520 ) | ( n34519 & n34520 ) ;
  assign n34522 = n8254 ^ n1722 ^ 1'b0 ;
  assign n34523 = ( n12354 & n19368 ) | ( n12354 & ~n21157 ) | ( n19368 & ~n21157 ) ;
  assign n34524 = ( n6366 & n34522 ) | ( n6366 & n34523 ) | ( n34522 & n34523 ) ;
  assign n34525 = ~n12296 & n34524 ;
  assign n34526 = n34525 ^ n28867 ^ 1'b0 ;
  assign n34527 = ~n8774 & n12576 ;
  assign n34528 = n34527 ^ n2567 ^ 1'b0 ;
  assign n34529 = n16676 ^ n12891 ^ n3173 ;
  assign n34530 = n34528 & n34529 ;
  assign n34531 = n4512 & n34530 ;
  assign n34532 = n27921 ^ n12244 ^ 1'b0 ;
  assign n34533 = ( n4356 & n9174 ) | ( n4356 & ~n12991 ) | ( n9174 & ~n12991 ) ;
  assign n34534 = n34533 ^ n10490 ^ n4284 ;
  assign n34535 = ( n701 & n2001 ) | ( n701 & n22480 ) | ( n2001 & n22480 ) ;
  assign n34536 = n6171 ^ x37 ^ 1'b0 ;
  assign n34537 = n4239 & ~n34536 ;
  assign n34538 = n34537 ^ n2198 ^ 1'b0 ;
  assign n34539 = n34535 & ~n34538 ;
  assign n34540 = n9997 & ~n17658 ;
  assign n34541 = n34540 ^ n10285 ^ 1'b0 ;
  assign n34542 = ~n4220 & n34541 ;
  assign n34543 = n4950 & n34542 ;
  assign n34544 = ( n34534 & n34539 ) | ( n34534 & ~n34543 ) | ( n34539 & ~n34543 ) ;
  assign n34545 = n2746 & n2871 ;
  assign n34546 = n4078 & n34545 ;
  assign n34547 = ( n8507 & n15008 ) | ( n8507 & ~n34546 ) | ( n15008 & ~n34546 ) ;
  assign n34548 = n3400 | n11114 ;
  assign n34549 = n18868 | n34548 ;
  assign n34550 = n11599 | n15568 ;
  assign n34551 = n34550 ^ n14859 ^ 1'b0 ;
  assign n34552 = n27913 ^ n19882 ^ 1'b0 ;
  assign n34553 = ~n7222 & n7360 ;
  assign n34554 = n34553 ^ n24181 ^ n13950 ;
  assign n34555 = n22063 ^ n12066 ^ n4518 ;
  assign n34556 = n5818 & n13489 ;
  assign n34557 = ( n1236 & n12714 ) | ( n1236 & n20546 ) | ( n12714 & n20546 ) ;
  assign n34560 = n2637 | n12507 ;
  assign n34558 = ( ~n6776 & n11269 ) | ( ~n6776 & n26412 ) | ( n11269 & n26412 ) ;
  assign n34559 = n34558 ^ n19953 ^ n3111 ;
  assign n34561 = n34560 ^ n34559 ^ n28134 ;
  assign n34562 = ( n11991 & n21269 ) | ( n11991 & n27827 ) | ( n21269 & n27827 ) ;
  assign n34563 = n34562 ^ n19763 ^ n13160 ;
  assign n34564 = n25248 ^ n14921 ^ n9835 ;
  assign n34565 = n16195 | n34564 ;
  assign n34566 = n20330 & ~n34565 ;
  assign n34568 = n19698 ^ n13543 ^ n11250 ;
  assign n34567 = ( ~n15494 & n17190 ) | ( ~n15494 & n18639 ) | ( n17190 & n18639 ) ;
  assign n34569 = n34568 ^ n34567 ^ 1'b0 ;
  assign n34570 = ~n4569 & n27622 ;
  assign n34571 = ~n2820 & n10188 ;
  assign n34572 = n34571 ^ n18744 ^ 1'b0 ;
  assign n34573 = n8805 | n34572 ;
  assign n34574 = n34573 ^ n5948 ^ 1'b0 ;
  assign n34575 = ~n34570 & n34574 ;
  assign n34576 = ( n349 & n1266 ) | ( n349 & ~n10608 ) | ( n1266 & ~n10608 ) ;
  assign n34577 = ( ~n3487 & n9577 ) | ( ~n3487 & n34576 ) | ( n9577 & n34576 ) ;
  assign n34578 = n21380 ^ n11883 ^ n1309 ;
  assign n34579 = n28866 ^ n18578 ^ n11829 ;
  assign n34580 = n11185 & ~n31647 ;
  assign n34581 = n34580 ^ n16289 ^ 1'b0 ;
  assign n34582 = n34579 | n34581 ;
  assign n34583 = n4030 | n11062 ;
  assign n34584 = n34583 ^ n10926 ^ 1'b0 ;
  assign n34585 = ( n6563 & n23978 ) | ( n6563 & n31149 ) | ( n23978 & n31149 ) ;
  assign n34586 = n24514 ^ n20051 ^ n17811 ;
  assign n34587 = ( n2106 & n19730 ) | ( n2106 & ~n34586 ) | ( n19730 & ~n34586 ) ;
  assign n34588 = ( n4204 & n17082 ) | ( n4204 & n18769 ) | ( n17082 & n18769 ) ;
  assign n34589 = n26645 ^ n695 ^ 1'b0 ;
  assign n34590 = ( n5930 & n19621 ) | ( n5930 & ~n33319 ) | ( n19621 & ~n33319 ) ;
  assign n34591 = n34590 ^ n13722 ^ 1'b0 ;
  assign n34592 = n34589 | n34591 ;
  assign n34593 = n34592 ^ n26363 ^ n18863 ;
  assign n34594 = n24656 ^ n3330 ^ 1'b0 ;
  assign n34595 = n8802 & n34594 ;
  assign n34596 = n34595 ^ n4481 ^ 1'b0 ;
  assign n34597 = ~n9993 & n26212 ;
  assign n34598 = n24672 ^ x158 ^ 1'b0 ;
  assign n34599 = n19370 & ~n26714 ;
  assign n34600 = n34599 ^ n10827 ^ 1'b0 ;
  assign n34601 = n662 & n34600 ;
  assign n34602 = ~n34598 & n34601 ;
  assign n34603 = ( ~n744 & n33424 ) | ( ~n744 & n34602 ) | ( n33424 & n34602 ) ;
  assign n34604 = n2290 & ~n6400 ;
  assign n34605 = n34604 ^ n1108 ^ 1'b0 ;
  assign n34606 = n26111 & ~n34605 ;
  assign n34607 = n34606 ^ n558 ^ 1'b0 ;
  assign n34608 = n34607 ^ n30211 ^ n14784 ;
  assign n34609 = n16487 ^ n7721 ^ n2525 ;
  assign n34610 = n15657 ^ n7308 ^ 1'b0 ;
  assign n34611 = n24919 & n34610 ;
  assign n34612 = n5302 & n10799 ;
  assign n34613 = n34612 ^ n11415 ^ 1'b0 ;
  assign n34614 = ( n6188 & ~n13147 ) | ( n6188 & n34613 ) | ( ~n13147 & n34613 ) ;
  assign n34615 = n24562 ^ n16803 ^ 1'b0 ;
  assign n34616 = n7009 & n34615 ;
  assign n34617 = n34616 ^ n27406 ^ 1'b0 ;
  assign n34618 = n34614 & ~n34617 ;
  assign n34619 = n22194 ^ n21240 ^ n18421 ;
  assign n34620 = n33689 & n34619 ;
  assign n34621 = n23240 & n34620 ;
  assign n34622 = n16787 ^ n12919 ^ 1'b0 ;
  assign n34623 = n19193 & n34622 ;
  assign n34626 = n1340 | n4366 ;
  assign n34627 = n34626 ^ n4576 ^ 1'b0 ;
  assign n34624 = n21742 ^ n10062 ^ 1'b0 ;
  assign n34625 = n5554 | n34624 ;
  assign n34628 = n34627 ^ n34625 ^ n7370 ;
  assign n34629 = ( n10218 & ~n16513 ) | ( n10218 & n26854 ) | ( ~n16513 & n26854 ) ;
  assign n34630 = n33985 ^ n1776 ^ x24 ;
  assign n34631 = ( n3036 & n5816 ) | ( n3036 & n34630 ) | ( n5816 & n34630 ) ;
  assign n34632 = n14906 ^ n8745 ^ 1'b0 ;
  assign n34633 = x227 & n22595 ;
  assign n34634 = n34633 ^ n25581 ^ 1'b0 ;
  assign n34635 = n7761 | n15671 ;
  assign n34640 = n4730 ^ n4633 ^ 1'b0 ;
  assign n34636 = n766 & ~n17966 ;
  assign n34637 = n34636 ^ n1621 ^ 1'b0 ;
  assign n34638 = n6558 | n34637 ;
  assign n34639 = n34638 ^ n3476 ^ 1'b0 ;
  assign n34641 = n34640 ^ n34639 ^ x41 ;
  assign n34642 = n13884 ^ n13559 ^ n11402 ;
  assign n34643 = n34642 ^ n9306 ^ n4858 ;
  assign n34644 = n14885 ^ n9984 ^ n6464 ;
  assign n34645 = ( n8678 & n8928 ) | ( n8678 & ~n34644 ) | ( n8928 & ~n34644 ) ;
  assign n34646 = ~n17935 & n34645 ;
  assign n34647 = n9772 & n34646 ;
  assign n34648 = ( ~n1041 & n2250 ) | ( ~n1041 & n2796 ) | ( n2250 & n2796 ) ;
  assign n34649 = n2329 & n7491 ;
  assign n34650 = ( n34647 & n34648 ) | ( n34647 & n34649 ) | ( n34648 & n34649 ) ;
  assign n34651 = n24188 ^ n3755 ^ 1'b0 ;
  assign n34652 = ( n6515 & n19984 ) | ( n6515 & n20113 ) | ( n19984 & n20113 ) ;
  assign n34653 = n6393 ^ n1952 ^ 1'b0 ;
  assign n34654 = n17379 & n34653 ;
  assign n34655 = n33896 & n34654 ;
  assign n34656 = n34655 ^ n12626 ^ 1'b0 ;
  assign n34657 = n34652 & ~n34656 ;
  assign n34659 = n4492 & n25766 ;
  assign n34658 = n5837 | n18238 ;
  assign n34660 = n34659 ^ n34658 ^ 1'b0 ;
  assign n34661 = n20669 ^ n19409 ^ n1059 ;
  assign n34662 = n15345 ^ n14078 ^ n11817 ;
  assign n34663 = n34662 ^ n13411 ^ n4418 ;
  assign n34664 = n34663 ^ n26660 ^ n4376 ;
  assign n34665 = n29354 ^ n27567 ^ n13478 ;
  assign n34666 = n34665 ^ n7628 ^ 1'b0 ;
  assign n34667 = ( ~n3460 & n4313 ) | ( ~n3460 & n6211 ) | ( n4313 & n6211 ) ;
  assign n34668 = ( ~n1192 & n9126 ) | ( ~n1192 & n15740 ) | ( n9126 & n15740 ) ;
  assign n34669 = n16190 ^ n11885 ^ n4937 ;
  assign n34670 = n2873 | n34669 ;
  assign n34671 = n34668 & ~n34670 ;
  assign n34672 = n8318 ^ n1969 ^ 1'b0 ;
  assign n34673 = n909 & n34672 ;
  assign n34674 = ~n10232 & n34673 ;
  assign n34675 = n34674 ^ n1364 ^ 1'b0 ;
  assign n34676 = n632 & ~n12501 ;
  assign n34677 = ~n34675 & n34676 ;
  assign n34678 = ( ~n4004 & n4362 ) | ( ~n4004 & n34677 ) | ( n4362 & n34677 ) ;
  assign n34679 = n19628 ^ n11956 ^ n5713 ;
  assign n34681 = n5084 ^ n4674 ^ n335 ;
  assign n34682 = n32859 | n34681 ;
  assign n34680 = n17050 | n25384 ;
  assign n34683 = n34682 ^ n34680 ^ 1'b0 ;
  assign n34684 = ( ~n3550 & n32405 ) | ( ~n3550 & n34683 ) | ( n32405 & n34683 ) ;
  assign n34685 = n12891 ^ n12803 ^ 1'b0 ;
  assign n34686 = n34685 ^ n23908 ^ n13249 ;
  assign n34687 = n32599 ^ n20696 ^ 1'b0 ;
  assign n34688 = n26429 & ~n34687 ;
  assign n34689 = ~n3920 & n5302 ;
  assign n34690 = n34689 ^ n28609 ^ 1'b0 ;
  assign n34691 = n27950 ^ n14669 ^ n3489 ;
  assign n34692 = n34691 ^ n16200 ^ n2539 ;
  assign n34693 = n33629 ^ n18893 ^ 1'b0 ;
  assign n34694 = ( n928 & n7611 ) | ( n928 & n7791 ) | ( n7611 & n7791 ) ;
  assign n34695 = ( n18151 & ~n30911 ) | ( n18151 & n34694 ) | ( ~n30911 & n34694 ) ;
  assign n34696 = n34695 ^ n27277 ^ n26178 ;
  assign n34697 = n6045 & ~n7152 ;
  assign n34698 = ~n33548 & n34697 ;
  assign n34699 = n34698 ^ n28089 ^ n5899 ;
  assign n34700 = n3985 & ~n23874 ;
  assign n34701 = ( ~n10990 & n28827 ) | ( ~n10990 & n34700 ) | ( n28827 & n34700 ) ;
  assign n34702 = n21693 ^ n9066 ^ 1'b0 ;
  assign n34703 = n28774 | n30288 ;
  assign n34704 = n34702 | n34703 ;
  assign n34705 = n22543 ^ n18272 ^ 1'b0 ;
  assign n34709 = n2864 & ~n6711 ;
  assign n34706 = n20466 ^ n7694 ^ 1'b0 ;
  assign n34707 = n34706 ^ n15321 ^ n1444 ;
  assign n34708 = ~n15015 & n34707 ;
  assign n34710 = n34709 ^ n34708 ^ n17279 ;
  assign n34711 = n13312 & n14657 ;
  assign n34712 = ~n2664 & n34711 ;
  assign n34713 = n5732 & n18889 ;
  assign n34714 = n34713 ^ n25338 ^ n14603 ;
  assign n34715 = n18469 ^ n2208 ^ 1'b0 ;
  assign n34716 = n28942 & ~n34715 ;
  assign n34717 = ( n12634 & ~n20694 ) | ( n12634 & n34716 ) | ( ~n20694 & n34716 ) ;
  assign n34718 = ~n13723 & n18481 ;
  assign n34719 = ( ~n8220 & n17439 ) | ( ~n8220 & n21924 ) | ( n17439 & n21924 ) ;
  assign n34720 = ( ~n1429 & n4123 ) | ( ~n1429 & n8840 ) | ( n4123 & n8840 ) ;
  assign n34721 = n17570 & ~n34720 ;
  assign n34722 = n29893 ^ n25805 ^ n4636 ;
  assign n34723 = n28576 ^ n8987 ^ n2940 ;
  assign n34724 = n10676 | n31999 ;
  assign n34725 = n2092 & n34724 ;
  assign n34726 = n19106 ^ n5352 ^ n2601 ;
  assign n34727 = n4041 | n34726 ;
  assign n34728 = n5430 & n21093 ;
  assign n34729 = ~n1524 & n24592 ;
  assign n34730 = n34729 ^ n7443 ^ 1'b0 ;
  assign n34731 = ( n8150 & n17526 ) | ( n8150 & ~n24529 ) | ( n17526 & ~n24529 ) ;
  assign n34732 = ( n13872 & n15889 ) | ( n13872 & n34731 ) | ( n15889 & n34731 ) ;
  assign n34733 = n1129 | n5211 ;
  assign n34734 = x118 | n34733 ;
  assign n34735 = n34734 ^ n14772 ^ 1'b0 ;
  assign n34736 = n28617 ^ n2620 ^ 1'b0 ;
  assign n34737 = n27158 ^ n21347 ^ 1'b0 ;
  assign n34738 = n34737 ^ n29771 ^ n7193 ;
  assign n34739 = ( n2319 & n18783 ) | ( n2319 & n24822 ) | ( n18783 & n24822 ) ;
  assign n34740 = n22339 ^ n10251 ^ n8509 ;
  assign n34741 = n34740 ^ n19409 ^ n9991 ;
  assign n34742 = n26858 ^ n3705 ^ 1'b0 ;
  assign n34743 = n12570 ^ n1730 ^ 1'b0 ;
  assign n34744 = n34279 & n34743 ;
  assign n34745 = n10368 ^ n8640 ^ n6268 ;
  assign n34746 = n34744 & n34745 ;
  assign n34747 = n34746 ^ n6720 ^ 1'b0 ;
  assign n34749 = ( n4474 & ~n11277 ) | ( n4474 & n17585 ) | ( ~n11277 & n17585 ) ;
  assign n34750 = n7392 | n34749 ;
  assign n34751 = n3520 | n34750 ;
  assign n34748 = n879 & ~n916 ;
  assign n34752 = n34751 ^ n34748 ^ 1'b0 ;
  assign n34753 = n34752 ^ n27056 ^ n7662 ;
  assign n34754 = n29765 ^ n18539 ^ n18352 ;
  assign n34755 = ~n34753 & n34754 ;
  assign n34756 = n27885 ^ n14985 ^ n6422 ;
  assign n34757 = ( n10206 & n29827 ) | ( n10206 & ~n34756 ) | ( n29827 & ~n34756 ) ;
  assign n34758 = ( x9 & ~n8181 ) | ( x9 & n17377 ) | ( ~n8181 & n17377 ) ;
  assign n34759 = n34758 ^ n16079 ^ n11485 ;
  assign n34760 = n14222 ^ n5707 ^ 1'b0 ;
  assign n34761 = n28007 & ~n34760 ;
  assign n34762 = n29357 ^ n5966 ^ 1'b0 ;
  assign n34763 = n17430 ^ n6334 ^ n4858 ;
  assign n34765 = n824 & n16849 ;
  assign n34766 = n34765 ^ n7527 ^ 1'b0 ;
  assign n34764 = n4926 & n25332 ;
  assign n34767 = n34766 ^ n34764 ^ 1'b0 ;
  assign n34768 = n3653 & n8459 ;
  assign n34769 = n34768 ^ n27808 ^ 1'b0 ;
  assign n34770 = ( n13406 & ~n18926 ) | ( n13406 & n23551 ) | ( ~n18926 & n23551 ) ;
  assign n34771 = ( n15479 & n24471 ) | ( n15479 & ~n31105 ) | ( n24471 & ~n31105 ) ;
  assign n34772 = ~n5152 & n18294 ;
  assign n34773 = n34772 ^ n17320 ^ 1'b0 ;
  assign n34774 = ( n29961 & n34771 ) | ( n29961 & n34773 ) | ( n34771 & n34773 ) ;
  assign n34775 = ( ~n9684 & n12921 ) | ( ~n9684 & n23773 ) | ( n12921 & n23773 ) ;
  assign n34776 = ( n4464 & n4864 ) | ( n4464 & n31529 ) | ( n4864 & n31529 ) ;
  assign n34777 = n16746 ^ n7448 ^ 1'b0 ;
  assign n34778 = ~n14857 & n34777 ;
  assign n34779 = n29616 ^ n3220 ^ 1'b0 ;
  assign n34780 = n10743 | n34779 ;
  assign n34781 = n34778 & ~n34780 ;
  assign n34782 = n34781 ^ n21065 ^ 1'b0 ;
  assign n34783 = ( n13111 & n22084 ) | ( n13111 & n22758 ) | ( n22084 & n22758 ) ;
  assign n34784 = ( x102 & n25406 ) | ( x102 & ~n34783 ) | ( n25406 & ~n34783 ) ;
  assign n34786 = ( n16063 & n17436 ) | ( n16063 & ~n26020 ) | ( n17436 & ~n26020 ) ;
  assign n34785 = n1011 & n17783 ;
  assign n34787 = n34786 ^ n34785 ^ 1'b0 ;
  assign n34788 = n1508 & n34787 ;
  assign n34789 = ~n34784 & n34788 ;
  assign n34790 = n3753 | n25153 ;
  assign n34791 = n34790 ^ n25751 ^ n6720 ;
  assign n34792 = ~n24509 & n34791 ;
  assign n34793 = n16330 ^ n12213 ^ n3601 ;
  assign n34794 = n10590 | n34793 ;
  assign n34795 = ( n4409 & ~n10981 ) | ( n4409 & n16431 ) | ( ~n10981 & n16431 ) ;
  assign n34796 = n10366 | n29068 ;
  assign n34797 = n34796 ^ n22391 ^ 1'b0 ;
  assign n34798 = n34797 ^ n9159 ^ 1'b0 ;
  assign n34799 = ( n32271 & n32466 ) | ( n32271 & ~n34798 ) | ( n32466 & ~n34798 ) ;
  assign n34800 = n31549 ^ n11795 ^ 1'b0 ;
  assign n34801 = n21662 ^ n9795 ^ 1'b0 ;
  assign n34802 = n2803 & n34801 ;
  assign n34803 = ~n320 & n34802 ;
  assign n34804 = n31284 ^ n13046 ^ n6222 ;
  assign n34805 = ~n7502 & n18130 ;
  assign n34806 = ( n492 & n7044 ) | ( n492 & n12305 ) | ( n7044 & n12305 ) ;
  assign n34807 = n4795 & n34806 ;
  assign n34808 = ~n34805 & n34807 ;
  assign n34809 = ( ~n8856 & n34804 ) | ( ~n8856 & n34808 ) | ( n34804 & n34808 ) ;
  assign n34810 = n22368 ^ n1713 ^ 1'b0 ;
  assign n34811 = n13595 & n34810 ;
  assign n34812 = x124 & n34811 ;
  assign n34813 = ~n4661 & n34812 ;
  assign n34814 = ( n14562 & n31799 ) | ( n14562 & n34813 ) | ( n31799 & n34813 ) ;
  assign n34815 = ( n18141 & ~n26390 ) | ( n18141 & n34814 ) | ( ~n26390 & n34814 ) ;
  assign n34816 = ( n3117 & n6981 ) | ( n3117 & n25286 ) | ( n6981 & n25286 ) ;
  assign n34817 = n638 & n10664 ;
  assign n34818 = n17216 & ~n34817 ;
  assign n34819 = ( ~n8090 & n20564 ) | ( ~n8090 & n34818 ) | ( n20564 & n34818 ) ;
  assign n34820 = n20069 ^ n8619 ^ n7250 ;
  assign n34821 = n34820 ^ n28934 ^ 1'b0 ;
  assign n34822 = n2688 & n16306 ;
  assign n34823 = n34822 ^ n903 ^ 1'b0 ;
  assign n34824 = n20014 ^ n3516 ^ 1'b0 ;
  assign n34825 = n23526 ^ n15134 ^ 1'b0 ;
  assign n34826 = n24332 | n34825 ;
  assign n34827 = n20232 & n30869 ;
  assign n34828 = n6762 ^ n2601 ^ 1'b0 ;
  assign n34829 = n16219 | n34828 ;
  assign n34830 = n26857 & ~n34829 ;
  assign n34831 = n34830 ^ n29954 ^ n13495 ;
  assign n34832 = n8579 ^ n3263 ^ 1'b0 ;
  assign n34833 = n1553 & n28011 ;
  assign n34834 = n34832 & n34833 ;
  assign n34835 = ( n24188 & ~n32002 ) | ( n24188 & n34834 ) | ( ~n32002 & n34834 ) ;
  assign n34836 = n1551 | n34835 ;
  assign n34837 = n14043 ^ n10274 ^ 1'b0 ;
  assign n34838 = n25549 | n34837 ;
  assign n34839 = n34838 ^ n29430 ^ n19542 ;
  assign n34840 = n19932 ^ n8696 ^ 1'b0 ;
  assign n34847 = n12435 & ~n18552 ;
  assign n34848 = n34847 ^ n4279 ^ 1'b0 ;
  assign n34843 = ( n8657 & n16423 ) | ( n8657 & n20898 ) | ( n16423 & n20898 ) ;
  assign n34841 = n10606 | n18169 ;
  assign n34842 = n14832 & ~n34841 ;
  assign n34844 = n34843 ^ n34842 ^ n12063 ;
  assign n34845 = n12642 & n34844 ;
  assign n34846 = ~n28836 & n34845 ;
  assign n34849 = n34848 ^ n34846 ^ n15020 ;
  assign n34853 = n8886 ^ n4942 ^ n2930 ;
  assign n34850 = ~n1407 & n4171 ;
  assign n34851 = n34850 ^ n17237 ^ n453 ;
  assign n34852 = n955 & n34851 ;
  assign n34854 = n34853 ^ n34852 ^ 1'b0 ;
  assign n34855 = n28695 ^ n15284 ^ 1'b0 ;
  assign n34856 = n15368 & ~n34855 ;
  assign n34857 = n34856 ^ n29332 ^ 1'b0 ;
  assign n34858 = ( ~n3547 & n6618 ) | ( ~n3547 & n23948 ) | ( n6618 & n23948 ) ;
  assign n34859 = n30594 ^ n13557 ^ n5046 ;
  assign n34860 = ( n14015 & n19461 ) | ( n14015 & ~n34859 ) | ( n19461 & ~n34859 ) ;
  assign n34861 = ~n25981 & n34860 ;
  assign n34862 = ~n7928 & n34861 ;
  assign n34863 = n34862 ^ n28359 ^ n26638 ;
  assign n34864 = n31193 ^ n16962 ^ x65 ;
  assign n34865 = n18289 | n22096 ;
  assign n34866 = n5049 | n34865 ;
  assign n34867 = n1755 | n34602 ;
  assign n34868 = n16606 | n34867 ;
  assign n34869 = n5278 & n11430 ;
  assign n34870 = n34869 ^ n16756 ^ 1'b0 ;
  assign n34871 = ( n5965 & n21422 ) | ( n5965 & n31124 ) | ( n21422 & n31124 ) ;
  assign n34872 = n23059 | n31705 ;
  assign n34873 = n19638 | n34872 ;
  assign n34874 = n24828 ^ n19371 ^ n3323 ;
  assign n34875 = n29444 ^ n27055 ^ 1'b0 ;
  assign n34876 = ( n30727 & ~n34874 ) | ( n30727 & n34875 ) | ( ~n34874 & n34875 ) ;
  assign n34877 = n34876 ^ n27565 ^ 1'b0 ;
  assign n34878 = n32984 ^ n14593 ^ 1'b0 ;
  assign n34879 = ( ~n4900 & n17407 ) | ( ~n4900 & n28157 ) | ( n17407 & n28157 ) ;
  assign n34880 = n4027 & n18679 ;
  assign n34881 = ~x192 & n34880 ;
  assign n34882 = ~n15289 & n34881 ;
  assign n34883 = n34882 ^ n10165 ^ n9643 ;
  assign n34884 = ~n13081 & n26151 ;
  assign n34885 = n34883 & n34884 ;
  assign n34886 = n34879 | n34885 ;
  assign n34887 = ( n6181 & n6542 ) | ( n6181 & ~n34886 ) | ( n6542 & ~n34886 ) ;
  assign n34888 = ~n22997 & n34887 ;
  assign n34889 = ( ~n6070 & n13075 ) | ( ~n6070 & n21785 ) | ( n13075 & n21785 ) ;
  assign n34890 = n17783 ^ n1421 ^ 1'b0 ;
  assign n34891 = ~n27218 & n34890 ;
  assign n34892 = n34891 ^ n32906 ^ n4286 ;
  assign n34893 = ( n21842 & ~n27619 ) | ( n21842 & n34892 ) | ( ~n27619 & n34892 ) ;
  assign n34895 = ~n10570 & n22382 ;
  assign n34894 = ( n6313 & n23373 ) | ( n6313 & n27744 ) | ( n23373 & n27744 ) ;
  assign n34896 = n34895 ^ n34894 ^ 1'b0 ;
  assign n34897 = n19348 & ~n22191 ;
  assign n34898 = n15048 & n34897 ;
  assign n34899 = n13907 ^ n7497 ^ 1'b0 ;
  assign n34900 = n1201 & n34899 ;
  assign n34901 = n27497 & ~n34900 ;
  assign n34902 = n34901 ^ n3465 ^ 1'b0 ;
  assign n34903 = ~n10235 & n31869 ;
  assign n34904 = n34903 ^ n18284 ^ 1'b0 ;
  assign n34905 = n27426 ^ n22222 ^ n4913 ;
  assign n34906 = n29536 ^ n28563 ^ n24948 ;
  assign n34907 = n19661 ^ n14800 ^ n7014 ;
  assign n34908 = ( ~n674 & n12630 ) | ( ~n674 & n22638 ) | ( n12630 & n22638 ) ;
  assign n34909 = n17814 & ~n34908 ;
  assign n34910 = n34909 ^ n31517 ^ 1'b0 ;
  assign n34911 = n20273 & ~n27032 ;
  assign n34912 = n34911 ^ n17627 ^ 1'b0 ;
  assign n34913 = ~n18682 & n20488 ;
  assign n34914 = n27977 ^ n2791 ^ 1'b0 ;
  assign n34915 = n14788 & n34914 ;
  assign n34916 = n356 & ~n3919 ;
  assign n34917 = ( n5690 & n7080 ) | ( n5690 & n34916 ) | ( n7080 & n34916 ) ;
  assign n34918 = n5548 | n34917 ;
  assign n34919 = n8781 ^ n440 ^ 1'b0 ;
  assign n34920 = n30379 ^ n9684 ^ n8920 ;
  assign n34921 = n34919 | n34920 ;
  assign n34922 = n6129 | n14799 ;
  assign n34923 = ~n6328 & n20100 ;
  assign n34924 = ~n34922 & n34923 ;
  assign n34925 = n28564 ^ n9980 ^ 1'b0 ;
  assign n34926 = n705 & n34925 ;
  assign n34927 = n9077 ^ n7994 ^ n1563 ;
  assign n34928 = n29839 & ~n34927 ;
  assign n34929 = ~n30623 & n34928 ;
  assign n34935 = n7255 ^ n3841 ^ 1'b0 ;
  assign n34936 = n9542 ^ n4161 ^ n1937 ;
  assign n34937 = n34936 ^ n27504 ^ 1'b0 ;
  assign n34938 = n34935 & ~n34937 ;
  assign n34930 = n22660 ^ n6930 ^ 1'b0 ;
  assign n34931 = n692 | n3431 ;
  assign n34932 = n11583 & ~n34931 ;
  assign n34933 = n34930 | n34932 ;
  assign n34934 = n18159 & ~n34933 ;
  assign n34939 = n34938 ^ n34934 ^ n2398 ;
  assign n34940 = ( n3677 & n7244 ) | ( n3677 & ~n27900 ) | ( n7244 & ~n27900 ) ;
  assign n34941 = n9715 & ~n26138 ;
  assign n34942 = n12504 & ~n34941 ;
  assign n34943 = ~n34940 & n34942 ;
  assign n34944 = ( ~n2604 & n5159 ) | ( ~n2604 & n34943 ) | ( n5159 & n34943 ) ;
  assign n34945 = n34944 ^ n29038 ^ n9258 ;
  assign n34946 = n15828 ^ n5224 ^ 1'b0 ;
  assign n34947 = ( n10809 & n10967 ) | ( n10809 & n15543 ) | ( n10967 & n15543 ) ;
  assign n34948 = n7771 & n34947 ;
  assign n34949 = n1570 | n5707 ;
  assign n34950 = n31105 | n34949 ;
  assign n34951 = n33000 ^ x75 ^ 1'b0 ;
  assign n34952 = ( n13740 & ~n15190 ) | ( n13740 & n31704 ) | ( ~n15190 & n31704 ) ;
  assign n34953 = n21843 & ~n34952 ;
  assign n34954 = n15667 & ~n23988 ;
  assign n34955 = n24765 ^ n13279 ^ 1'b0 ;
  assign n34956 = n34954 | n34955 ;
  assign n34957 = ( n10534 & n15677 ) | ( n10534 & n34353 ) | ( n15677 & n34353 ) ;
  assign n34958 = ~n3122 & n13407 ;
  assign n34959 = ~n2702 & n34958 ;
  assign n34960 = n7266 | n34959 ;
  assign n34961 = n10139 | n34960 ;
  assign n34962 = ( n4761 & n18890 ) | ( n4761 & ~n34961 ) | ( n18890 & ~n34961 ) ;
  assign n34963 = n25203 | n34962 ;
  assign n34964 = n5905 | n34963 ;
  assign n34965 = ( n12221 & ~n17795 ) | ( n12221 & n23816 ) | ( ~n17795 & n23816 ) ;
  assign n34966 = n13856 & ~n13905 ;
  assign n34967 = n34965 & n34966 ;
  assign n34968 = ( n862 & ~n12063 ) | ( n862 & n15066 ) | ( ~n12063 & n15066 ) ;
  assign n34969 = ( ~n5862 & n11406 ) | ( ~n5862 & n32971 ) | ( n11406 & n32971 ) ;
  assign n34970 = n5437 & ~n7578 ;
  assign n34971 = ( n26500 & n34969 ) | ( n26500 & ~n34970 ) | ( n34969 & ~n34970 ) ;
  assign n34972 = ~n8579 & n10260 ;
  assign n34973 = ~n2936 & n34972 ;
  assign n34974 = n34973 ^ n20473 ^ 1'b0 ;
  assign n34975 = ~n27805 & n34974 ;
  assign n34976 = x30 & ~n34975 ;
  assign n34977 = n7895 ^ n698 ^ 1'b0 ;
  assign n34978 = n7686 ^ n5248 ^ 1'b0 ;
  assign n34979 = n34977 & ~n34978 ;
  assign n34980 = n16481 ^ n14657 ^ 1'b0 ;
  assign n34983 = n17592 ^ n8683 ^ n3977 ;
  assign n34982 = n10945 ^ n8270 ^ n4349 ;
  assign n34984 = n34983 ^ n34982 ^ 1'b0 ;
  assign n34985 = n14043 | n34984 ;
  assign n34981 = n5142 | n17764 ;
  assign n34986 = n34985 ^ n34981 ^ 1'b0 ;
  assign n34987 = n13342 & ~n19317 ;
  assign n34988 = n17445 & n34987 ;
  assign n34989 = ( n20698 & ~n28728 ) | ( n20698 & n34988 ) | ( ~n28728 & n34988 ) ;
  assign n34990 = n16296 & n34989 ;
  assign n34991 = n10809 ^ n5824 ^ n1128 ;
  assign n34992 = ( ~n19303 & n30307 ) | ( ~n19303 & n34991 ) | ( n30307 & n34991 ) ;
  assign n34993 = n34992 ^ n11786 ^ 1'b0 ;
  assign n34994 = ( n3010 & ~n3720 ) | ( n3010 & n34993 ) | ( ~n3720 & n34993 ) ;
  assign n34995 = n34994 ^ n22883 ^ n21732 ;
  assign n34996 = ~n544 & n11697 ;
  assign n34997 = n34996 ^ n15609 ^ 1'b0 ;
  assign n34998 = ( ~n15700 & n16095 ) | ( ~n15700 & n19602 ) | ( n16095 & n19602 ) ;
  assign n35000 = ( n2768 & n19873 ) | ( n2768 & n21412 ) | ( n19873 & n21412 ) ;
  assign n34999 = n17710 | n21787 ;
  assign n35001 = n35000 ^ n34999 ^ 1'b0 ;
  assign n35002 = n6440 & n8344 ;
  assign n35003 = n35002 ^ n22875 ^ 1'b0 ;
  assign n35004 = n14193 & n21204 ;
  assign n35005 = ( n13843 & n35003 ) | ( n13843 & n35004 ) | ( n35003 & n35004 ) ;
  assign n35006 = ~n6955 & n18924 ;
  assign n35007 = n35006 ^ n24258 ^ 1'b0 ;
  assign n35008 = n35005 & n35007 ;
  assign n35009 = n7389 ^ n2561 ^ 1'b0 ;
  assign n35010 = n35009 ^ n1200 ^ 1'b0 ;
  assign n35011 = n16234 & n35010 ;
  assign n35012 = ~n12891 & n35011 ;
  assign n35013 = n2590 & n8251 ;
  assign n35014 = ( n29454 & n32187 ) | ( n29454 & n35013 ) | ( n32187 & n35013 ) ;
  assign n35015 = ~n11785 & n27004 ;
  assign n35016 = ( n2426 & ~n9394 ) | ( n2426 & n35015 ) | ( ~n9394 & n35015 ) ;
  assign n35017 = ( ~n7230 & n27487 ) | ( ~n7230 & n35016 ) | ( n27487 & n35016 ) ;
  assign n35018 = n5214 ^ n4368 ^ 1'b0 ;
  assign n35019 = n7091 & ~n35018 ;
  assign n35020 = n25952 | n27311 ;
  assign n35021 = n35019 | n35020 ;
  assign n35024 = n33851 ^ n5033 ^ 1'b0 ;
  assign n35025 = n15521 | n35024 ;
  assign n35022 = n7410 & ~n10790 ;
  assign n35023 = n35022 ^ n22668 ^ 1'b0 ;
  assign n35026 = n35025 ^ n35023 ^ n34159 ;
  assign n35028 = n16051 | n31778 ;
  assign n35027 = ( ~n20687 & n24872 ) | ( ~n20687 & n25042 ) | ( n24872 & n25042 ) ;
  assign n35029 = n35028 ^ n35027 ^ 1'b0 ;
  assign n35030 = ( ~n1548 & n3352 ) | ( ~n1548 & n7172 ) | ( n3352 & n7172 ) ;
  assign n35031 = n35030 ^ n12857 ^ 1'b0 ;
  assign n35032 = n2582 & n24169 ;
  assign n35033 = n7993 & n35032 ;
  assign n35034 = n35033 ^ n11970 ^ 1'b0 ;
  assign n35035 = n16244 & n24044 ;
  assign n35036 = ( n14579 & ~n14630 ) | ( n14579 & n35035 ) | ( ~n14630 & n35035 ) ;
  assign n35037 = n32158 | n35036 ;
  assign n35038 = n9019 & ~n35037 ;
  assign n35041 = n25913 ^ n16678 ^ 1'b0 ;
  assign n35042 = n22809 & ~n35041 ;
  assign n35043 = n35042 ^ n31660 ^ 1'b0 ;
  assign n35039 = n28558 ^ n3673 ^ 1'b0 ;
  assign n35040 = ~n11742 & n35039 ;
  assign n35044 = n35043 ^ n35040 ^ 1'b0 ;
  assign n35045 = ~n7040 & n21342 ;
  assign n35046 = ( ~n12769 & n15914 ) | ( ~n12769 & n23959 ) | ( n15914 & n23959 ) ;
  assign n35047 = n35046 ^ n22458 ^ n12301 ;
  assign n35048 = n35047 ^ n25374 ^ 1'b0 ;
  assign n35049 = n35048 ^ n14412 ^ n3892 ;
  assign n35050 = n35049 ^ n10657 ^ 1'b0 ;
  assign n35051 = n35045 & n35050 ;
  assign n35052 = n17079 ^ n11738 ^ n9846 ;
  assign n35053 = n35052 ^ n5351 ^ n625 ;
  assign n35054 = ~n8567 & n35053 ;
  assign n35055 = n15492 & ~n23064 ;
  assign n35056 = ( n8988 & n11686 ) | ( n8988 & n35055 ) | ( n11686 & n35055 ) ;
  assign n35057 = n33859 ^ n22875 ^ n1916 ;
  assign n35058 = ( n2354 & n13680 ) | ( n2354 & ~n29846 ) | ( n13680 & ~n29846 ) ;
  assign n35059 = n35058 ^ n20826 ^ n17795 ;
  assign n35060 = n29628 ^ n13455 ^ 1'b0 ;
  assign n35061 = ( ~n2620 & n11818 ) | ( ~n2620 & n16274 ) | ( n11818 & n16274 ) ;
  assign n35062 = n35061 ^ n27659 ^ n17952 ;
  assign n35063 = ( n1829 & n2515 ) | ( n1829 & n6842 ) | ( n2515 & n6842 ) ;
  assign n35064 = n35062 | n35063 ;
  assign n35065 = n26973 ^ n24938 ^ n2739 ;
  assign n35067 = n20082 & n20457 ;
  assign n35066 = n12739 | n24005 ;
  assign n35068 = n35067 ^ n35066 ^ n24707 ;
  assign n35069 = n6564 & n6848 ;
  assign n35070 = n35069 ^ n4523 ^ 1'b0 ;
  assign n35071 = n35070 ^ n10384 ^ n1751 ;
  assign n35072 = n35071 ^ n35016 ^ n6236 ;
  assign n35073 = n6114 & n29831 ;
  assign n35074 = ~n26014 & n35073 ;
  assign n35075 = n21512 ^ n8262 ^ 1'b0 ;
  assign n35076 = ~n6570 & n35075 ;
  assign n35077 = n35076 ^ n16267 ^ 1'b0 ;
  assign n35078 = n33624 ^ n29524 ^ n5672 ;
  assign n35079 = n35078 ^ n32705 ^ 1'b0 ;
  assign n35080 = n20308 & ~n22483 ;
  assign n35081 = ( n6196 & ~n8426 ) | ( n6196 & n12715 ) | ( ~n8426 & n12715 ) ;
  assign n35082 = n35081 ^ n28922 ^ n10620 ;
  assign n35083 = ( n11065 & ~n13105 ) | ( n11065 & n26967 ) | ( ~n13105 & n26967 ) ;
  assign n35084 = ~n349 & n4348 ;
  assign n35085 = n35084 ^ n3237 ^ 1'b0 ;
  assign n35087 = n3892 | n14224 ;
  assign n35088 = n35087 ^ n258 ^ 1'b0 ;
  assign n35086 = n10314 | n23223 ;
  assign n35089 = n35088 ^ n35086 ^ n15589 ;
  assign n35090 = ( n25196 & ~n35085 ) | ( n25196 & n35089 ) | ( ~n35085 & n35089 ) ;
  assign n35095 = n32864 ^ n16023 ^ n13552 ;
  assign n35091 = ( ~n688 & n6279 ) | ( ~n688 & n13733 ) | ( n6279 & n13733 ) ;
  assign n35092 = n9117 & n35091 ;
  assign n35093 = n35092 ^ n14611 ^ 1'b0 ;
  assign n35094 = n12909 & n35093 ;
  assign n35096 = n35095 ^ n35094 ^ 1'b0 ;
  assign n35097 = n27008 ^ n11059 ^ n6577 ;
  assign n35098 = n5827 & n35097 ;
  assign n35099 = ~n35096 & n35098 ;
  assign n35100 = n14234 ^ x94 ^ 1'b0 ;
  assign n35101 = ~n8754 & n35100 ;
  assign n35102 = n35101 ^ n10332 ^ 1'b0 ;
  assign n35103 = n35099 | n35102 ;
  assign n35104 = ~n16538 & n29911 ;
  assign n35105 = n3443 & n35104 ;
  assign n35108 = n14867 ^ n9538 ^ 1'b0 ;
  assign n35109 = ~n1901 & n35108 ;
  assign n35106 = n15580 ^ n7809 ^ n397 ;
  assign n35107 = n1534 | n35106 ;
  assign n35110 = n35109 ^ n35107 ^ 1'b0 ;
  assign n35111 = ( n6868 & ~n11301 ) | ( n6868 & n12277 ) | ( ~n11301 & n12277 ) ;
  assign n35112 = ~n11668 & n20793 ;
  assign n35113 = ( n12293 & n32238 ) | ( n12293 & n35112 ) | ( n32238 & n35112 ) ;
  assign n35114 = n14415 & ~n35113 ;
  assign n35115 = n25699 & n35114 ;
  assign n35116 = n35111 | n35115 ;
  assign n35117 = n10858 ^ n6728 ^ 1'b0 ;
  assign n35118 = n35117 ^ n33075 ^ 1'b0 ;
  assign n35119 = n2873 | n25731 ;
  assign n35121 = n7557 ^ n2207 ^ n2086 ;
  assign n35122 = n35121 ^ n20847 ^ x24 ;
  assign n35120 = n14737 ^ n5633 ^ n4753 ;
  assign n35123 = n35122 ^ n35120 ^ 1'b0 ;
  assign n35124 = ( n9924 & n14139 ) | ( n9924 & n30378 ) | ( n14139 & n30378 ) ;
  assign n35125 = n35124 ^ n17600 ^ n2279 ;
  assign n35126 = ~n6847 & n21743 ;
  assign n35127 = ~n25325 & n35126 ;
  assign n35128 = n35127 ^ n22840 ^ n21986 ;
  assign n35129 = ~n7791 & n32688 ;
  assign n35130 = n35129 ^ n16513 ^ 1'b0 ;
  assign n35131 = n13294 & ~n14253 ;
  assign n35132 = n35131 ^ n18586 ^ 1'b0 ;
  assign n35133 = n18508 | n32547 ;
  assign n35134 = n15375 & ~n35133 ;
  assign n35135 = ( ~n3772 & n15523 ) | ( ~n3772 & n29306 ) | ( n15523 & n29306 ) ;
  assign n35136 = ( n13716 & n35134 ) | ( n13716 & n35135 ) | ( n35134 & n35135 ) ;
  assign n35137 = n25610 ^ n23174 ^ 1'b0 ;
  assign n35138 = n35137 ^ n22166 ^ n5392 ;
  assign n35139 = n24026 ^ n9120 ^ n6326 ;
  assign n35140 = ~n6158 & n33457 ;
  assign n35141 = n26832 & n35140 ;
  assign n35142 = n5816 | n6325 ;
  assign n35143 = n12243 & n35142 ;
  assign n35144 = n31618 & n35143 ;
  assign n35145 = ( n9073 & n35141 ) | ( n9073 & ~n35144 ) | ( n35141 & ~n35144 ) ;
  assign n35146 = n23659 ^ x0 ^ 1'b0 ;
  assign n35147 = ~n6548 & n35146 ;
  assign n35148 = n5232 & ~n14885 ;
  assign n35149 = n11635 ^ n8696 ^ n2556 ;
  assign n35150 = n35149 ^ n589 ^ 1'b0 ;
  assign n35151 = ~n35148 & n35150 ;
  assign n35152 = n20088 ^ n14697 ^ 1'b0 ;
  assign n35153 = n23726 ^ n18767 ^ 1'b0 ;
  assign n35154 = ( n791 & n14978 ) | ( n791 & ~n20318 ) | ( n14978 & ~n20318 ) ;
  assign n35155 = n7568 | n11466 ;
  assign n35156 = n18627 | n35155 ;
  assign n35157 = n351 | n28345 ;
  assign n35158 = n35157 ^ n23087 ^ 1'b0 ;
  assign n35159 = ( n35154 & ~n35156 ) | ( n35154 & n35158 ) | ( ~n35156 & n35158 ) ;
  assign n35160 = ( ~n18650 & n22811 ) | ( ~n18650 & n35159 ) | ( n22811 & n35159 ) ;
  assign n35161 = n4362 ^ x89 ^ 1'b0 ;
  assign n35162 = ~n17508 & n35161 ;
  assign n35163 = n35162 ^ n20956 ^ 1'b0 ;
  assign n35164 = n35163 ^ n24609 ^ n19815 ;
  assign n35165 = n33685 ^ n31118 ^ 1'b0 ;
  assign n35166 = n22168 & n23818 ;
  assign n35167 = n5450 & n35166 ;
  assign n35168 = n35167 ^ n20625 ^ n13715 ;
  assign n35169 = n10270 ^ n8669 ^ n5222 ;
  assign n35170 = ( x238 & ~n6100 ) | ( x238 & n35169 ) | ( ~n6100 & n35169 ) ;
  assign n35171 = ( n8123 & n10373 ) | ( n8123 & ~n35170 ) | ( n10373 & ~n35170 ) ;
  assign n35172 = n11990 & ~n30557 ;
  assign n35173 = ~n6045 & n35172 ;
  assign n35174 = n30195 ^ n27137 ^ n5309 ;
  assign n35176 = ( n12553 & n15703 ) | ( n12553 & n32609 ) | ( n15703 & n32609 ) ;
  assign n35175 = n17363 ^ n1295 ^ 1'b0 ;
  assign n35177 = n35176 ^ n35175 ^ n27413 ;
  assign n35178 = ( n8514 & ~n23202 ) | ( n8514 & n29502 ) | ( ~n23202 & n29502 ) ;
  assign n35179 = ( n15491 & ~n23269 ) | ( n15491 & n29874 ) | ( ~n23269 & n29874 ) ;
  assign n35180 = n20882 ^ n10280 ^ 1'b0 ;
  assign n35181 = ~n32426 & n35180 ;
  assign n35182 = ( ~n6826 & n7044 ) | ( ~n6826 & n19128 ) | ( n7044 & n19128 ) ;
  assign n35183 = n32827 ^ n30850 ^ n9702 ;
  assign n35184 = n21442 ^ n14852 ^ n5513 ;
  assign n35185 = ( n13802 & n29234 ) | ( n13802 & n29362 ) | ( n29234 & n29362 ) ;
  assign n35186 = ~n5522 & n13735 ;
  assign n35187 = n11164 & n35186 ;
  assign n35188 = ( n4195 & ~n8332 ) | ( n4195 & n35187 ) | ( ~n8332 & n35187 ) ;
  assign n35189 = n19222 ^ n4262 ^ n2808 ;
  assign n35190 = n2096 | n35189 ;
  assign n35191 = n35188 | n35190 ;
  assign n35192 = n9720 & ~n10283 ;
  assign n35193 = n35192 ^ n31411 ^ 1'b0 ;
  assign n35194 = n23386 ^ n2329 ^ 1'b0 ;
  assign n35195 = ( n7753 & n29671 ) | ( n7753 & n35194 ) | ( n29671 & n35194 ) ;
  assign n35196 = n7175 ^ n6035 ^ 1'b0 ;
  assign n35197 = n19588 & n35196 ;
  assign n35198 = n14158 & n15795 ;
  assign n35199 = n35198 ^ n25334 ^ 1'b0 ;
  assign n35200 = n35199 ^ n18454 ^ n10984 ;
  assign n35201 = n35200 ^ n31822 ^ n30330 ;
  assign n35202 = n9879 ^ n8290 ^ 1'b0 ;
  assign n35203 = ( n4052 & ~n6226 ) | ( n4052 & n7199 ) | ( ~n6226 & n7199 ) ;
  assign n35204 = n21244 | n35203 ;
  assign n35205 = n29288 | n35204 ;
  assign n35206 = ( ~n20845 & n35202 ) | ( ~n20845 & n35205 ) | ( n35202 & n35205 ) ;
  assign n35207 = n1583 & n11178 ;
  assign n35208 = n19753 | n20003 ;
  assign n35209 = n9956 | n25924 ;
  assign n35210 = n15696 ^ n2924 ^ 1'b0 ;
  assign n35211 = n10958 & ~n35210 ;
  assign n35213 = ~n7344 & n12723 ;
  assign n35214 = n35213 ^ n8529 ^ 1'b0 ;
  assign n35212 = n22192 ^ n14898 ^ 1'b0 ;
  assign n35215 = n35214 ^ n35212 ^ n2283 ;
  assign n35216 = n9507 ^ n1592 ^ 1'b0 ;
  assign n35217 = ( n8538 & ~n35215 ) | ( n8538 & n35216 ) | ( ~n35215 & n35216 ) ;
  assign n35218 = n35217 ^ n33650 ^ n15762 ;
  assign n35219 = ( n2900 & n18861 ) | ( n2900 & n18974 ) | ( n18861 & n18974 ) ;
  assign n35221 = n25670 & n29557 ;
  assign n35220 = ( n3154 & n3633 ) | ( n3154 & n8489 ) | ( n3633 & n8489 ) ;
  assign n35222 = n35221 ^ n35220 ^ n399 ;
  assign n35223 = n8460 & ~n35222 ;
  assign n35224 = ~n8086 & n35223 ;
  assign n35225 = n27099 ^ n5216 ^ 1'b0 ;
  assign n35226 = n29317 & ~n35225 ;
  assign n35227 = n19275 ^ n7428 ^ n6726 ;
  assign n35228 = ( n9385 & n34010 ) | ( n9385 & ~n35227 ) | ( n34010 & ~n35227 ) ;
  assign n35229 = n35228 ^ n27632 ^ n9993 ;
  assign n35230 = n10546 ^ n4385 ^ 1'b0 ;
  assign n35231 = n7549 & ~n16438 ;
  assign n35232 = n30019 ^ n16281 ^ 1'b0 ;
  assign n35233 = n35231 | n35232 ;
  assign n35234 = n7797 ^ n5616 ^ n3003 ;
  assign n35235 = n19849 ^ n5212 ^ 1'b0 ;
  assign n35236 = n35234 | n35235 ;
  assign n35237 = n32221 ^ n28719 ^ n1494 ;
  assign n35238 = n33236 & n35237 ;
  assign n35239 = n35238 ^ n665 ^ 1'b0 ;
  assign n35240 = ~n19892 & n35239 ;
  assign n35241 = n3874 & ~n31440 ;
  assign n35242 = n35241 ^ n9535 ^ 1'b0 ;
  assign n35243 = n35242 ^ n23978 ^ n19952 ;
  assign n35244 = n19176 ^ n12682 ^ n10401 ;
  assign n35245 = ( ~n1217 & n16078 ) | ( ~n1217 & n18677 ) | ( n16078 & n18677 ) ;
  assign n35246 = n10374 | n30550 ;
  assign n35247 = ( n14418 & ~n24514 ) | ( n14418 & n35246 ) | ( ~n24514 & n35246 ) ;
  assign n35248 = ~n3103 & n6046 ;
  assign n35249 = ( n12944 & n14679 ) | ( n12944 & ~n35248 ) | ( n14679 & ~n35248 ) ;
  assign n35250 = n776 & n12113 ;
  assign n35252 = ~n5560 & n7141 ;
  assign n35251 = n5504 ^ n4012 ^ 1'b0 ;
  assign n35253 = n35252 ^ n35251 ^ n30079 ;
  assign n35254 = n35250 | n35253 ;
  assign n35255 = n15829 ^ n13107 ^ n4630 ;
  assign n35256 = n12885 & n35255 ;
  assign n35257 = ~n24441 & n35256 ;
  assign n35258 = ( n4760 & ~n12775 ) | ( n4760 & n34050 ) | ( ~n12775 & n34050 ) ;
  assign n35259 = n35258 ^ n13384 ^ 1'b0 ;
  assign n35260 = n26380 & ~n35259 ;
  assign n35261 = n4625 & ~n10349 ;
  assign n35262 = ~n14873 & n35261 ;
  assign n35263 = n16552 ^ n11477 ^ 1'b0 ;
  assign n35264 = ( n13573 & ~n14299 ) | ( n13573 & n17585 ) | ( ~n14299 & n17585 ) ;
  assign n35265 = n3339 & ~n7938 ;
  assign n35266 = n17864 & ~n31732 ;
  assign n35267 = n35266 ^ n11035 ^ 1'b0 ;
  assign n35269 = n14896 ^ n4083 ^ n2733 ;
  assign n35270 = n35269 ^ n8766 ^ n6132 ;
  assign n35268 = n10658 | n12980 ;
  assign n35271 = n35270 ^ n35268 ^ 1'b0 ;
  assign n35272 = n31596 ^ n11186 ^ n1154 ;
  assign n35273 = n35272 ^ n22583 ^ n2946 ;
  assign n35274 = n19190 ^ n4649 ^ 1'b0 ;
  assign n35275 = n21703 ^ n6948 ^ 1'b0 ;
  assign n35276 = n19270 & n25207 ;
  assign n35277 = n35276 ^ n31331 ^ 1'b0 ;
  assign n35278 = n35275 & n35277 ;
  assign n35279 = n35278 ^ n6620 ^ n6230 ;
  assign n35280 = n17284 ^ n7771 ^ n2458 ;
  assign n35281 = n11083 | n35280 ;
  assign n35282 = n35281 ^ n34524 ^ n8782 ;
  assign n35285 = n8321 & ~n10713 ;
  assign n35286 = n5377 & n35285 ;
  assign n35287 = n35286 ^ n6190 ^ 1'b0 ;
  assign n35288 = n19035 & ~n35287 ;
  assign n35283 = n2930 & n18390 ;
  assign n35284 = n35283 ^ n19427 ^ 1'b0 ;
  assign n35289 = n35288 ^ n35284 ^ 1'b0 ;
  assign n35290 = ( ~n5561 & n11510 ) | ( ~n5561 & n18542 ) | ( n11510 & n18542 ) ;
  assign n35294 = n22957 ^ n5246 ^ 1'b0 ;
  assign n35291 = n20283 ^ n7241 ^ 1'b0 ;
  assign n35292 = n35291 ^ n32273 ^ n25196 ;
  assign n35293 = n6185 & n35292 ;
  assign n35295 = n35294 ^ n35293 ^ 1'b0 ;
  assign n35296 = n2944 & n17098 ;
  assign n35297 = ( ~n3853 & n6015 ) | ( ~n3853 & n34272 ) | ( n6015 & n34272 ) ;
  assign n35298 = n35297 ^ n10263 ^ n768 ;
  assign n35299 = n35298 ^ n31788 ^ 1'b0 ;
  assign n35300 = ~n6237 & n35299 ;
  assign n35301 = ~n7117 & n23347 ;
  assign n35302 = n35301 ^ n13738 ^ 1'b0 ;
  assign n35303 = n32054 ^ n29068 ^ n932 ;
  assign n35304 = ( ~n4018 & n19353 ) | ( ~n4018 & n30251 ) | ( n19353 & n30251 ) ;
  assign n35305 = n12936 | n28793 ;
  assign n35306 = n35305 ^ n10505 ^ 1'b0 ;
  assign n35307 = n35306 ^ n21415 ^ n3608 ;
  assign n35308 = n1096 & n9231 ;
  assign n35309 = ~n20346 & n35308 ;
  assign n35310 = ( n9438 & n23382 ) | ( n9438 & n35309 ) | ( n23382 & n35309 ) ;
  assign n35311 = n19972 ^ n12620 ^ 1'b0 ;
  assign n35312 = n6027 & ~n35311 ;
  assign n35313 = ~n15204 & n35312 ;
  assign n35314 = ~n25827 & n35313 ;
  assign n35315 = n2057 & ~n35314 ;
  assign n35317 = n12473 ^ n4822 ^ 1'b0 ;
  assign n35316 = ~n18121 & n31800 ;
  assign n35318 = n35317 ^ n35316 ^ n25940 ;
  assign n35319 = n35318 ^ n16284 ^ n8637 ;
  assign n35320 = n8455 ^ n4735 ^ n4367 ;
  assign n35321 = ( ~n5855 & n17815 ) | ( ~n5855 & n35320 ) | ( n17815 & n35320 ) ;
  assign n35322 = n35321 ^ n5275 ^ 1'b0 ;
  assign n35327 = n11335 ^ n5583 ^ n2168 ;
  assign n35325 = n6219 | n25789 ;
  assign n35326 = n4591 & ~n35325 ;
  assign n35323 = n3327 & ~n24579 ;
  assign n35324 = n24826 & n35323 ;
  assign n35328 = n35327 ^ n35326 ^ n35324 ;
  assign n35330 = ( n2541 & ~n2627 ) | ( n2541 & n18549 ) | ( ~n2627 & n18549 ) ;
  assign n35331 = n22323 ^ n7223 ^ n1205 ;
  assign n35332 = ( n21831 & ~n35330 ) | ( n21831 & n35331 ) | ( ~n35330 & n35331 ) ;
  assign n35329 = ~n10088 & n20431 ;
  assign n35333 = n35332 ^ n35329 ^ 1'b0 ;
  assign n35334 = ( n35322 & n35328 ) | ( n35322 & ~n35333 ) | ( n35328 & ~n35333 ) ;
  assign n35335 = ~n2118 & n30966 ;
  assign n35336 = n23032 ^ n3958 ^ 1'b0 ;
  assign n35337 = ( ~n2655 & n9661 ) | ( ~n2655 & n28875 ) | ( n9661 & n28875 ) ;
  assign n35338 = ~n10935 & n35337 ;
  assign n35339 = n35336 | n35338 ;
  assign n35340 = n21415 ^ n7988 ^ 1'b0 ;
  assign n35341 = n35340 ^ n20242 ^ 1'b0 ;
  assign n35342 = n17626 & n35341 ;
  assign n35343 = n5513 | n22411 ;
  assign n35344 = n35343 ^ n26260 ^ 1'b0 ;
  assign n35345 = ( n1727 & n24679 ) | ( n1727 & ~n35344 ) | ( n24679 & ~n35344 ) ;
  assign n35346 = ( n8635 & n17566 ) | ( n8635 & n21567 ) | ( n17566 & n21567 ) ;
  assign n35347 = n8835 ^ n5729 ^ 1'b0 ;
  assign n35348 = n13332 | n22673 ;
  assign n35349 = ( ~n35346 & n35347 ) | ( ~n35346 & n35348 ) | ( n35347 & n35348 ) ;
  assign n35350 = ( ~x203 & n12299 ) | ( ~x203 & n25912 ) | ( n12299 & n25912 ) ;
  assign n35351 = n26621 & n35350 ;
  assign n35352 = n5842 ^ n2520 ^ 1'b0 ;
  assign n35353 = n35351 & ~n35352 ;
  assign n35354 = n9244 | n26919 ;
  assign n35355 = n5264 & n32017 ;
  assign n35356 = ~n35354 & n35355 ;
  assign n35357 = n31764 ^ n12120 ^ 1'b0 ;
  assign n35358 = ( n15460 & n19665 ) | ( n15460 & n19706 ) | ( n19665 & n19706 ) ;
  assign n35359 = n10732 & ~n29587 ;
  assign n35360 = ~n6848 & n35359 ;
  assign n35361 = n15434 | n35360 ;
  assign n35362 = n22538 ^ n22427 ^ n17489 ;
  assign n35363 = n10739 & n35362 ;
  assign n35364 = ( n5572 & n9949 ) | ( n5572 & ~n35363 ) | ( n9949 & ~n35363 ) ;
  assign n35365 = n15592 ^ n14222 ^ 1'b0 ;
  assign n35366 = n30093 | n35365 ;
  assign n35367 = n16601 ^ n11429 ^ 1'b0 ;
  assign n35368 = n35367 ^ n17917 ^ 1'b0 ;
  assign n35369 = n24279 | n35368 ;
  assign n35370 = n28522 ^ n18867 ^ n13469 ;
  assign n35371 = n23009 | n35370 ;
  assign n35372 = n24097 ^ n10896 ^ 1'b0 ;
  assign n35373 = n1482 & n4757 ;
  assign n35374 = n18839 & n35373 ;
  assign n35375 = ( n5530 & n13190 ) | ( n5530 & n35374 ) | ( n13190 & n35374 ) ;
  assign n35376 = ( n16964 & n35372 ) | ( n16964 & ~n35375 ) | ( n35372 & ~n35375 ) ;
  assign n35377 = n16650 ^ n15159 ^ n2662 ;
  assign n35378 = ( n2270 & n9534 ) | ( n2270 & ~n35377 ) | ( n9534 & ~n35377 ) ;
  assign n35379 = ( n29893 & ~n29960 ) | ( n29893 & n35378 ) | ( ~n29960 & n35378 ) ;
  assign n35380 = n34077 ^ n19158 ^ n17641 ;
  assign n35381 = ( n21449 & n35379 ) | ( n21449 & n35380 ) | ( n35379 & n35380 ) ;
  assign n35382 = ( n4899 & ~n14765 ) | ( n4899 & n20762 ) | ( ~n14765 & n20762 ) ;
  assign n35383 = n35382 ^ n2684 ^ 1'b0 ;
  assign n35384 = n20117 | n35383 ;
  assign n35385 = ~n2134 & n2843 ;
  assign n35386 = n35385 ^ n13563 ^ 1'b0 ;
  assign n35387 = n20787 ^ n1949 ^ 1'b0 ;
  assign n35388 = ~n35386 & n35387 ;
  assign n35391 = n28157 ^ n24149 ^ n17069 ;
  assign n35389 = n32752 ^ n4049 ^ 1'b0 ;
  assign n35390 = n15209 & n35389 ;
  assign n35392 = n35391 ^ n35390 ^ n17891 ;
  assign n35393 = n16028 & n35392 ;
  assign n35394 = n14325 & n35393 ;
  assign n35395 = n2157 & ~n28607 ;
  assign n35396 = ( ~n1322 & n17004 ) | ( ~n1322 & n19524 ) | ( n17004 & n19524 ) ;
  assign n35397 = ~n20262 & n35396 ;
  assign n35398 = n13049 ^ n11440 ^ n1961 ;
  assign n35399 = n10625 ^ n9652 ^ 1'b0 ;
  assign n35400 = n35398 & n35399 ;
  assign n35401 = n35400 ^ n22658 ^ n9587 ;
  assign n35402 = ( ~n4151 & n15418 ) | ( ~n4151 & n34085 ) | ( n15418 & n34085 ) ;
  assign n35403 = n35402 ^ n15491 ^ 1'b0 ;
  assign n35404 = n8777 ^ n546 ^ 1'b0 ;
  assign n35405 = n9356 | n35404 ;
  assign n35406 = n35405 ^ n12832 ^ n5671 ;
  assign n35407 = ( ~n13859 & n24071 ) | ( ~n13859 & n35406 ) | ( n24071 & n35406 ) ;
  assign n35408 = n5454 ^ n5449 ^ n3352 ;
  assign n35409 = ( n12447 & ~n17012 ) | ( n12447 & n35408 ) | ( ~n17012 & n35408 ) ;
  assign n35410 = n32039 ^ n808 ^ 1'b0 ;
  assign n35411 = n24342 & n34882 ;
  assign n35412 = n30454 ^ n17207 ^ 1'b0 ;
  assign n35413 = n21108 ^ n4782 ^ n1822 ;
  assign n35414 = n13580 ^ n10261 ^ n8311 ;
  assign n35415 = ( n4651 & n15764 ) | ( n4651 & n35414 ) | ( n15764 & n35414 ) ;
  assign n35416 = ( ~n6384 & n35413 ) | ( ~n6384 & n35415 ) | ( n35413 & n35415 ) ;
  assign n35417 = n2036 & ~n27867 ;
  assign n35418 = n35417 ^ n23459 ^ 1'b0 ;
  assign n35419 = ( n16348 & n20724 ) | ( n16348 & ~n35418 ) | ( n20724 & ~n35418 ) ;
  assign n35420 = ( ~n4401 & n14838 ) | ( ~n4401 & n19798 ) | ( n14838 & n19798 ) ;
  assign n35421 = n16829 ^ n1865 ^ 1'b0 ;
  assign n35423 = ~n8719 & n27181 ;
  assign n35424 = ~n12764 & n35423 ;
  assign n35422 = ~n1306 & n33339 ;
  assign n35425 = n35424 ^ n35422 ^ 1'b0 ;
  assign n35426 = ( n19796 & ~n35421 ) | ( n19796 & n35425 ) | ( ~n35421 & n35425 ) ;
  assign n35427 = ( n2594 & ~n7708 ) | ( n2594 & n33951 ) | ( ~n7708 & n33951 ) ;
  assign n35428 = n15862 | n35427 ;
  assign n35429 = n35428 ^ n18041 ^ 1'b0 ;
  assign n35430 = n35426 | n35429 ;
  assign n35431 = n13500 & ~n35336 ;
  assign n35432 = ~n2110 & n28336 ;
  assign n35433 = ( n11303 & ~n16068 ) | ( n11303 & n35432 ) | ( ~n16068 & n35432 ) ;
  assign n35434 = ~n5142 & n14994 ;
  assign n35435 = n7664 & n35434 ;
  assign n35436 = n35435 ^ n23209 ^ n6698 ;
  assign n35437 = n32798 ^ n23965 ^ n19800 ;
  assign n35440 = n16649 ^ n3406 ^ n283 ;
  assign n35441 = n17590 & ~n35440 ;
  assign n35442 = n1163 & n35441 ;
  assign n35438 = ( ~n23332 & n31913 ) | ( ~n23332 & n33381 ) | ( n31913 & n33381 ) ;
  assign n35439 = ~n25463 & n35438 ;
  assign n35443 = n35442 ^ n35439 ^ 1'b0 ;
  assign n35444 = n31669 ^ n12022 ^ n4615 ;
  assign n35445 = n35444 ^ n2511 ^ 1'b0 ;
  assign n35446 = ( ~n493 & n957 ) | ( ~n493 & n35445 ) | ( n957 & n35445 ) ;
  assign n35447 = x210 & ~n13146 ;
  assign n35448 = ~n33103 & n35447 ;
  assign n35449 = ( n12796 & n26843 ) | ( n12796 & n35448 ) | ( n26843 & n35448 ) ;
  assign n35450 = n35446 & n35449 ;
  assign n35451 = n35450 ^ n7423 ^ 1'b0 ;
  assign n35452 = n32314 ^ n21020 ^ n6661 ;
  assign n35453 = n14883 | n35452 ;
  assign n35454 = n35453 ^ n30363 ^ 1'b0 ;
  assign n35455 = n20584 ^ n16705 ^ 1'b0 ;
  assign n35456 = n35227 ^ n19801 ^ n6811 ;
  assign n35457 = n14506 ^ n13663 ^ n5374 ;
  assign n35458 = ( ~n21505 & n27312 ) | ( ~n21505 & n35457 ) | ( n27312 & n35457 ) ;
  assign n35462 = n29896 ^ n8519 ^ 1'b0 ;
  assign n35459 = n14553 & ~n21860 ;
  assign n35460 = ~n21050 & n35459 ;
  assign n35461 = n35460 ^ n13871 ^ 1'b0 ;
  assign n35463 = n35462 ^ n35461 ^ n25836 ;
  assign n35464 = n14868 ^ n9579 ^ 1'b0 ;
  assign n35465 = n27046 & ~n35464 ;
  assign n35466 = n7990 & ~n14639 ;
  assign n35467 = n35466 ^ n15187 ^ 1'b0 ;
  assign n35468 = n35467 ^ n34908 ^ n13819 ;
  assign n35469 = n15850 ^ n11633 ^ n6982 ;
  assign n35470 = n7377 & ~n18471 ;
  assign n35471 = ~n566 & n35470 ;
  assign n35472 = ( n2686 & n13294 ) | ( n2686 & n35471 ) | ( n13294 & n35471 ) ;
  assign n35473 = n2426 | n23605 ;
  assign n35474 = n5551 | n16016 ;
  assign n35475 = ( n12017 & n35473 ) | ( n12017 & n35474 ) | ( n35473 & n35474 ) ;
  assign n35476 = n16125 & n18698 ;
  assign n35477 = n15505 & n35476 ;
  assign n35478 = n18765 ^ n8774 ^ 1'b0 ;
  assign n35479 = ~n35477 & n35478 ;
  assign n35483 = n14474 & ~n17775 ;
  assign n35484 = n35483 ^ n2924 ^ 1'b0 ;
  assign n35485 = n10639 & ~n35484 ;
  assign n35480 = n3637 ^ x55 ^ 1'b0 ;
  assign n35481 = ~n20404 & n35480 ;
  assign n35482 = n35481 ^ n22922 ^ n7560 ;
  assign n35486 = n35485 ^ n35482 ^ n18462 ;
  assign n35487 = n6099 & n7759 ;
  assign n35488 = ~n32876 & n35487 ;
  assign n35489 = n35488 ^ n26416 ^ n742 ;
  assign n35490 = n5592 & ~n35489 ;
  assign n35491 = n35486 & n35490 ;
  assign n35492 = ~n520 & n5897 ;
  assign n35493 = n35492 ^ n19168 ^ 1'b0 ;
  assign n35494 = ( n29101 & n34145 ) | ( n29101 & n35493 ) | ( n34145 & n35493 ) ;
  assign n35495 = n16244 ^ n6566 ^ 1'b0 ;
  assign n35496 = ( n7114 & n18367 ) | ( n7114 & n35495 ) | ( n18367 & n35495 ) ;
  assign n35497 = ~n1280 & n9821 ;
  assign n35498 = n35497 ^ n15626 ^ n3335 ;
  assign n35501 = ( n544 & n12226 ) | ( n544 & n20147 ) | ( n12226 & n20147 ) ;
  assign n35499 = n1049 | n19832 ;
  assign n35500 = n25823 | n35499 ;
  assign n35502 = n35501 ^ n35500 ^ 1'b0 ;
  assign n35503 = n24522 | n35502 ;
  assign n35504 = n18259 ^ n276 ^ 1'b0 ;
  assign n35505 = n29495 ^ n24581 ^ n2649 ;
  assign n35506 = n4728 & ~n34685 ;
  assign n35507 = n22858 ^ n13760 ^ n4921 ;
  assign n35508 = n14594 ^ n3495 ^ 1'b0 ;
  assign n35509 = n23141 ^ n19073 ^ 1'b0 ;
  assign n35511 = n16726 ^ n13636 ^ 1'b0 ;
  assign n35512 = n20779 ^ n17434 ^ 1'b0 ;
  assign n35513 = n35511 | n35512 ;
  assign n35514 = n35513 ^ n18593 ^ 1'b0 ;
  assign n35510 = n12687 & n27604 ;
  assign n35515 = n35514 ^ n35510 ^ 1'b0 ;
  assign n35522 = n2529 & ~n5762 ;
  assign n35523 = n35522 ^ n19111 ^ 1'b0 ;
  assign n35519 = n2428 & n7016 ;
  assign n35520 = ~n12214 & n35519 ;
  assign n35516 = n23217 ^ n9952 ^ n6670 ;
  assign n35517 = n35516 ^ n6077 ^ n4965 ;
  assign n35518 = n13856 & n35517 ;
  assign n35521 = n35520 ^ n35518 ^ 1'b0 ;
  assign n35524 = n35523 ^ n35521 ^ 1'b0 ;
  assign n35528 = n7678 ^ n1299 ^ 1'b0 ;
  assign n35525 = n16513 ^ n14373 ^ n1140 ;
  assign n35526 = ~n26994 & n35525 ;
  assign n35527 = n6248 & n35526 ;
  assign n35529 = n35528 ^ n35527 ^ n4492 ;
  assign n35530 = n32737 ^ n7159 ^ 1'b0 ;
  assign n35532 = n28813 ^ n10251 ^ n7402 ;
  assign n35533 = ~n22618 & n35532 ;
  assign n35534 = n35533 ^ n10106 ^ 1'b0 ;
  assign n35531 = ( n8499 & ~n12677 ) | ( n8499 & n14724 ) | ( ~n12677 & n14724 ) ;
  assign n35535 = n35534 ^ n35531 ^ n30005 ;
  assign n35536 = n29442 ^ n26605 ^ n16979 ;
  assign n35537 = n8023 | n31433 ;
  assign n35538 = n32929 | n35537 ;
  assign n35541 = n30148 ^ n23815 ^ n6875 ;
  assign n35542 = ( n15726 & ~n31724 ) | ( n15726 & n35541 ) | ( ~n31724 & n35541 ) ;
  assign n35539 = ( n1810 & ~n27922 ) | ( n1810 & n29518 ) | ( ~n27922 & n29518 ) ;
  assign n35540 = ~n21236 & n35539 ;
  assign n35543 = n35542 ^ n35540 ^ 1'b0 ;
  assign n35544 = n19557 ^ n10500 ^ 1'b0 ;
  assign n35545 = ( n9120 & n24869 ) | ( n9120 & n35544 ) | ( n24869 & n35544 ) ;
  assign n35546 = n16560 ^ n14487 ^ 1'b0 ;
  assign n35547 = n35546 ^ n16640 ^ n13057 ;
  assign n35548 = ~n9626 & n22471 ;
  assign n35549 = n35548 ^ n1544 ^ 1'b0 ;
  assign n35550 = ( n598 & ~n2103 ) | ( n598 & n5082 ) | ( ~n2103 & n5082 ) ;
  assign n35551 = n35550 ^ n9784 ^ n6197 ;
  assign n35552 = ( ~n3097 & n35549 ) | ( ~n3097 & n35551 ) | ( n35549 & n35551 ) ;
  assign n35553 = ( n30151 & ~n35547 ) | ( n30151 & n35552 ) | ( ~n35547 & n35552 ) ;
  assign n35554 = ~n579 & n8730 ;
  assign n35555 = n21147 & ~n35554 ;
  assign n35556 = ~n10208 & n35555 ;
  assign n35557 = ~n5343 & n24996 ;
  assign n35558 = n35557 ^ n34736 ^ 1'b0 ;
  assign n35559 = n7433 ^ n3363 ^ 1'b0 ;
  assign n35560 = n2791 & n18143 ;
  assign n35561 = n8037 | n35560 ;
  assign n35562 = n8389 & ~n29446 ;
  assign n35563 = n35562 ^ n25650 ^ 1'b0 ;
  assign n35564 = n7159 | n13724 ;
  assign n35565 = n28708 ^ n11618 ^ 1'b0 ;
  assign n35566 = ( n11158 & n16118 ) | ( n11158 & ~n31508 ) | ( n16118 & ~n31508 ) ;
  assign n35567 = n26101 | n35566 ;
  assign n35568 = ( n4245 & n6354 ) | ( n4245 & n27793 ) | ( n6354 & n27793 ) ;
  assign n35569 = ( ~n4291 & n27166 ) | ( ~n4291 & n35568 ) | ( n27166 & n35568 ) ;
  assign n35570 = n20786 ^ n19172 ^ n4460 ;
  assign n35572 = n6916 | n21176 ;
  assign n35573 = n35572 ^ n4198 ^ 1'b0 ;
  assign n35571 = ( ~n6151 & n10190 ) | ( ~n6151 & n17118 ) | ( n10190 & n17118 ) ;
  assign n35574 = n35573 ^ n35571 ^ n810 ;
  assign n35575 = n8079 & n14176 ;
  assign n35576 = n35575 ^ n14988 ^ 1'b0 ;
  assign n35577 = n35576 ^ n27679 ^ 1'b0 ;
  assign n35578 = n16559 & n35577 ;
  assign n35579 = n12785 & n35578 ;
  assign n35580 = n30235 ^ n19913 ^ 1'b0 ;
  assign n35581 = ( n5853 & n27579 ) | ( n5853 & ~n35580 ) | ( n27579 & ~n35580 ) ;
  assign n35582 = n24875 | n35581 ;
  assign n35583 = n35582 ^ n24648 ^ 1'b0 ;
  assign n35584 = n25466 ^ n11173 ^ 1'b0 ;
  assign n35585 = ~n17122 & n35584 ;
  assign n35586 = n16703 | n24735 ;
  assign n35592 = n7144 & n10831 ;
  assign n35590 = n27363 ^ n12835 ^ n6282 ;
  assign n35591 = n35590 ^ n1684 ^ 1'b0 ;
  assign n35587 = n6216 ^ n432 ^ 1'b0 ;
  assign n35588 = n2661 & ~n35587 ;
  assign n35589 = n35588 ^ n4595 ^ n4315 ;
  assign n35593 = n35592 ^ n35591 ^ n35589 ;
  assign n35594 = ~n16200 & n33981 ;
  assign n35595 = n22055 ^ n4908 ^ n1765 ;
  assign n35596 = ~n20246 & n27614 ;
  assign n35597 = ( n9222 & n25494 ) | ( n9222 & n35596 ) | ( n25494 & n35596 ) ;
  assign n35598 = n28063 ^ n25371 ^ n19870 ;
  assign n35599 = n19095 & ~n35598 ;
  assign n35600 = ~n35597 & n35599 ;
  assign n35601 = n33284 ^ n21628 ^ 1'b0 ;
  assign n35602 = n35601 ^ n526 ^ 1'b0 ;
  assign n35603 = n17432 & n35602 ;
  assign n35604 = n26454 ^ n20308 ^ 1'b0 ;
  assign n35605 = ~n8073 & n35604 ;
  assign n35607 = ~n1359 & n21720 ;
  assign n35608 = n35607 ^ n12185 ^ 1'b0 ;
  assign n35609 = n35608 ^ n20807 ^ n8595 ;
  assign n35606 = n3314 & ~n33898 ;
  assign n35610 = n35609 ^ n35606 ^ 1'b0 ;
  assign n35611 = ~n17155 & n28189 ;
  assign n35617 = ( ~n7516 & n9424 ) | ( ~n7516 & n18436 ) | ( n9424 & n18436 ) ;
  assign n35618 = n35617 ^ n13230 ^ 1'b0 ;
  assign n35612 = n5482 ^ n4228 ^ 1'b0 ;
  assign n35613 = ( n1190 & n4711 ) | ( n1190 & n35612 ) | ( n4711 & n35612 ) ;
  assign n35614 = n23742 | n35613 ;
  assign n35615 = n2270 & ~n35614 ;
  assign n35616 = n35615 ^ n34453 ^ n27559 ;
  assign n35619 = n35618 ^ n35616 ^ 1'b0 ;
  assign n35620 = ~n35611 & n35619 ;
  assign n35621 = n1414 & ~n29348 ;
  assign n35622 = n18088 & n35621 ;
  assign n35623 = n20776 ^ n8514 ^ n5320 ;
  assign n35624 = ( n10994 & ~n22896 ) | ( n10994 & n23064 ) | ( ~n22896 & n23064 ) ;
  assign n35625 = n35624 ^ n23026 ^ n10941 ;
  assign n35626 = ( n13807 & n34659 ) | ( n13807 & ~n35625 ) | ( n34659 & ~n35625 ) ;
  assign n35627 = n1888 & n2732 ;
  assign n35628 = n12057 & n35627 ;
  assign n35629 = n28940 ^ n27737 ^ n19689 ;
  assign n35630 = n35629 ^ n19566 ^ n18338 ;
  assign n35631 = n28618 ^ n6526 ^ n3526 ;
  assign n35632 = ( n5408 & n24674 ) | ( n5408 & ~n35631 ) | ( n24674 & ~n35631 ) ;
  assign n35635 = ( n3609 & ~n5303 ) | ( n3609 & n5775 ) | ( ~n5303 & n5775 ) ;
  assign n35636 = ( n4082 & n9295 ) | ( n4082 & n35635 ) | ( n9295 & n35635 ) ;
  assign n35633 = ( n1442 & n8802 ) | ( n1442 & ~n17590 ) | ( n8802 & ~n17590 ) ;
  assign n35634 = ( ~n12838 & n15976 ) | ( ~n12838 & n35633 ) | ( n15976 & n35633 ) ;
  assign n35637 = n35636 ^ n35634 ^ 1'b0 ;
  assign n35638 = ~n23416 & n31952 ;
  assign n35639 = n11296 | n35638 ;
  assign n35640 = n35639 ^ n23403 ^ 1'b0 ;
  assign n35641 = n20329 ^ n8188 ^ n5297 ;
  assign n35642 = n22075 ^ n12857 ^ 1'b0 ;
  assign n35643 = n11304 ^ n1923 ^ 1'b0 ;
  assign n35644 = n35642 & ~n35643 ;
  assign n35645 = ~n19820 & n35644 ;
  assign n35646 = ~n27607 & n35645 ;
  assign n35647 = ( ~n3399 & n7297 ) | ( ~n3399 & n13332 ) | ( n7297 & n13332 ) ;
  assign n35648 = ( ~n350 & n18527 ) | ( ~n350 & n35647 ) | ( n18527 & n35647 ) ;
  assign n35649 = ( n4481 & ~n15087 ) | ( n4481 & n35648 ) | ( ~n15087 & n35648 ) ;
  assign n35650 = n12814 | n25984 ;
  assign n35651 = n7843 ^ n6010 ^ 1'b0 ;
  assign n35652 = n35651 ^ n29446 ^ 1'b0 ;
  assign n35653 = ( ~n9876 & n17700 ) | ( ~n9876 & n35652 ) | ( n17700 & n35652 ) ;
  assign n35654 = ~n7282 & n11044 ;
  assign n35655 = ~n11536 & n35654 ;
  assign n35658 = n8944 ^ n8102 ^ 1'b0 ;
  assign n35659 = n4541 & ~n35658 ;
  assign n35660 = ( n2402 & n8951 ) | ( n2402 & n35659 ) | ( n8951 & n35659 ) ;
  assign n35656 = n32547 ^ n7196 ^ 1'b0 ;
  assign n35657 = n35656 ^ n19089 ^ 1'b0 ;
  assign n35661 = n35660 ^ n35657 ^ 1'b0 ;
  assign n35662 = n7972 ^ n7470 ^ n4283 ;
  assign n35663 = n35662 ^ n31066 ^ 1'b0 ;
  assign n35664 = ( ~n25349 & n28904 ) | ( ~n25349 & n29618 ) | ( n28904 & n29618 ) ;
  assign n35665 = n23046 ^ n11009 ^ n6712 ;
  assign n35666 = n20978 ^ n18712 ^ 1'b0 ;
  assign n35667 = ( n27963 & ~n30269 ) | ( n27963 & n35666 ) | ( ~n30269 & n35666 ) ;
  assign n35668 = n6333 & ~n35667 ;
  assign n35669 = n19354 ^ n15079 ^ n10488 ;
  assign n35670 = n35669 ^ n5111 ^ 1'b0 ;
  assign n35671 = n33896 | n35670 ;
  assign n35672 = n27266 ^ n15201 ^ n12725 ;
  assign n35673 = n21485 ^ n11873 ^ 1'b0 ;
  assign n35674 = ( x236 & n18727 ) | ( x236 & n35673 ) | ( n18727 & n35673 ) ;
  assign n35675 = n7430 & n20752 ;
  assign n35676 = n35675 ^ n23720 ^ 1'b0 ;
  assign n35677 = n7554 & ~n25040 ;
  assign n35678 = n16436 ^ n4774 ^ n1211 ;
  assign n35680 = n15526 ^ x250 ^ 1'b0 ;
  assign n35681 = n19095 & ~n35680 ;
  assign n35679 = n4409 & n6940 ;
  assign n35682 = n35681 ^ n35679 ^ 1'b0 ;
  assign n35683 = n23398 ^ n15164 ^ n5916 ;
  assign n35684 = n32134 ^ n30997 ^ n1558 ;
  assign n35685 = n35684 ^ n505 ^ 1'b0 ;
  assign n35689 = n16409 ^ n8552 ^ n6486 ;
  assign n35687 = n1002 & ~n33983 ;
  assign n35688 = n35687 ^ n8472 ^ 1'b0 ;
  assign n35690 = n35689 ^ n35688 ^ n31788 ;
  assign n35686 = n33697 ^ n6300 ^ 1'b0 ;
  assign n35691 = n35690 ^ n35686 ^ n10069 ;
  assign n35692 = ~n26346 & n35691 ;
  assign n35693 = n14469 & n35692 ;
  assign n35694 = ~n12510 & n25917 ;
  assign n35695 = n8778 & n35694 ;
  assign n35696 = n14695 | n34476 ;
  assign n35697 = n16221 & ~n35696 ;
  assign n35701 = n9192 ^ n3129 ^ 1'b0 ;
  assign n35698 = ( n2242 & ~n10634 ) | ( n2242 & n25609 ) | ( ~n10634 & n25609 ) ;
  assign n35699 = n35698 ^ n35613 ^ n2782 ;
  assign n35700 = ( ~n26695 & n29441 ) | ( ~n26695 & n35699 ) | ( n29441 & n35699 ) ;
  assign n35702 = n35701 ^ n35700 ^ n20657 ;
  assign n35703 = ( n18254 & ~n19611 ) | ( n18254 & n24712 ) | ( ~n19611 & n24712 ) ;
  assign n35704 = n35703 ^ n28642 ^ n13167 ;
  assign n35705 = ( n16500 & n22975 ) | ( n16500 & ~n35704 ) | ( n22975 & ~n35704 ) ;
  assign n35706 = n14131 ^ n1507 ^ 1'b0 ;
  assign n35707 = n27210 & n35706 ;
  assign n35715 = n15552 | n22776 ;
  assign n35716 = n35715 ^ n2152 ^ 1'b0 ;
  assign n35708 = n9418 | n10192 ;
  assign n35709 = n35708 ^ n5863 ^ 1'b0 ;
  assign n35710 = n27998 ^ n8112 ^ 1'b0 ;
  assign n35711 = ( ~n7407 & n19782 ) | ( ~n7407 & n35710 ) | ( n19782 & n35710 ) ;
  assign n35712 = n25537 & n35711 ;
  assign n35713 = ( n6115 & ~n19621 ) | ( n6115 & n35712 ) | ( ~n19621 & n35712 ) ;
  assign n35714 = n35709 & ~n35713 ;
  assign n35717 = n35716 ^ n35714 ^ 1'b0 ;
  assign n35723 = n5342 | n7514 ;
  assign n35724 = n27660 & ~n35723 ;
  assign n35718 = n11788 ^ n5799 ^ n374 ;
  assign n35719 = ~n7862 & n14542 ;
  assign n35720 = ( n28387 & n30951 ) | ( n28387 & n35719 ) | ( n30951 & n35719 ) ;
  assign n35721 = ( n32018 & n35718 ) | ( n32018 & n35720 ) | ( n35718 & n35720 ) ;
  assign n35722 = n35721 ^ n27576 ^ 1'b0 ;
  assign n35725 = n35724 ^ n35722 ^ n29166 ;
  assign n35726 = ( n719 & ~n1984 ) | ( n719 & n8175 ) | ( ~n1984 & n8175 ) ;
  assign n35727 = n35726 ^ n8156 ^ n4592 ;
  assign n35728 = n31497 ^ n18791 ^ n8361 ;
  assign n35729 = ( n5042 & n9507 ) | ( n5042 & ~n20135 ) | ( n9507 & ~n20135 ) ;
  assign n35730 = ( n270 & n6055 ) | ( n270 & n7235 ) | ( n6055 & n7235 ) ;
  assign n35731 = n25768 ^ n1574 ^ n567 ;
  assign n35732 = n35731 ^ n9062 ^ 1'b0 ;
  assign n35733 = n14140 & n35732 ;
  assign n35734 = n24020 & n35733 ;
  assign n35735 = n35734 ^ n4711 ^ 1'b0 ;
  assign n35736 = n27986 | n31316 ;
  assign n35737 = n35736 ^ n13393 ^ 1'b0 ;
  assign n35738 = x238 & ~n17159 ;
  assign n35739 = n35738 ^ n15151 ^ 1'b0 ;
  assign n35740 = n35739 ^ n33788 ^ 1'b0 ;
  assign n35741 = n12177 ^ n1987 ^ 1'b0 ;
  assign n35742 = n35741 ^ n22974 ^ n12983 ;
  assign n35743 = n17476 ^ n5653 ^ x162 ;
  assign n35744 = n7616 & n18860 ;
  assign n35745 = n5818 & n35744 ;
  assign n35746 = n21793 ^ n17821 ^ n2141 ;
  assign n35747 = n35746 ^ n19202 ^ n9775 ;
  assign n35750 = n5812 ^ n433 ^ 1'b0 ;
  assign n35751 = n11886 & n35750 ;
  assign n35748 = n2770 & ~n19178 ;
  assign n35749 = n35748 ^ n23001 ^ 1'b0 ;
  assign n35752 = n35751 ^ n35749 ^ 1'b0 ;
  assign n35753 = n35747 & n35752 ;
  assign n35754 = n12920 ^ n8766 ^ 1'b0 ;
  assign n35755 = n1599 & ~n4602 ;
  assign n35756 = ~n32505 & n35755 ;
  assign n35757 = n18969 & n29227 ;
  assign n35758 = ( n7873 & n35756 ) | ( n7873 & ~n35757 ) | ( n35756 & ~n35757 ) ;
  assign n35759 = ( n2940 & ~n21988 ) | ( n2940 & n29039 ) | ( ~n21988 & n29039 ) ;
  assign n35760 = ~n3598 & n25423 ;
  assign n35761 = ( ~n35292 & n35759 ) | ( ~n35292 & n35760 ) | ( n35759 & n35760 ) ;
  assign n35762 = n13969 ^ n11241 ^ n8361 ;
  assign n35763 = n6485 & ~n35530 ;
  assign n35764 = n35763 ^ n15237 ^ 1'b0 ;
  assign n35765 = ( ~n5069 & n9331 ) | ( ~n5069 & n27175 ) | ( n9331 & n27175 ) ;
  assign n35766 = n509 | n29562 ;
  assign n35767 = ~n7699 & n35005 ;
  assign n35771 = n23518 & n26569 ;
  assign n35768 = ( n10848 & n27863 ) | ( n10848 & n30899 ) | ( n27863 & n30899 ) ;
  assign n35769 = n24943 ^ n3326 ^ 1'b0 ;
  assign n35770 = ~n35768 & n35769 ;
  assign n35772 = n35771 ^ n35770 ^ n23873 ;
  assign n35773 = n2753 & n35525 ;
  assign n35774 = ~n3308 & n35773 ;
  assign n35775 = n8353 & ~n16982 ;
  assign n35776 = n17440 & n35775 ;
  assign n35777 = ( n8880 & n11367 ) | ( n8880 & n18389 ) | ( n11367 & n18389 ) ;
  assign n35778 = n35777 ^ n8180 ^ n2327 ;
  assign n35779 = n14383 & ~n35778 ;
  assign n35780 = n15877 ^ n15764 ^ n1062 ;
  assign n35781 = n25742 ^ n24928 ^ n1246 ;
  assign n35782 = n35781 ^ n13739 ^ x42 ;
  assign n35783 = ( n11836 & ~n20991 ) | ( n11836 & n35782 ) | ( ~n20991 & n35782 ) ;
  assign n35784 = n11513 ^ n10621 ^ 1'b0 ;
  assign n35785 = n11273 & n35784 ;
  assign n35786 = ( ~n35780 & n35783 ) | ( ~n35780 & n35785 ) | ( n35783 & n35785 ) ;
  assign n35787 = n35786 ^ n28584 ^ x159 ;
  assign n35788 = ( n5710 & n13633 ) | ( n5710 & n28574 ) | ( n13633 & n28574 ) ;
  assign n35789 = n5162 & n32911 ;
  assign n35790 = n35789 ^ n29539 ^ n18201 ;
  assign n35791 = n24768 ^ n11831 ^ n2418 ;
  assign n35792 = n35791 ^ n2878 ^ 1'b0 ;
  assign n35793 = ~n2865 & n10620 ;
  assign n35794 = ~n35792 & n35793 ;
  assign n35795 = n32155 ^ n3516 ^ 1'b0 ;
  assign n35796 = n6483 & n35795 ;
  assign n35797 = ~n23434 & n26411 ;
  assign n35798 = n35797 ^ n33642 ^ 1'b0 ;
  assign n35799 = n22062 ^ n20803 ^ 1'b0 ;
  assign n35800 = n13302 | n35799 ;
  assign n35802 = ~n4275 & n9478 ;
  assign n35801 = n29912 ^ n11679 ^ 1'b0 ;
  assign n35803 = n35802 ^ n35801 ^ n2071 ;
  assign n35806 = n15994 ^ x68 ^ 1'b0 ;
  assign n35807 = n10520 | n35806 ;
  assign n35804 = n32372 ^ n8128 ^ n1010 ;
  assign n35805 = n35804 ^ n32271 ^ n7042 ;
  assign n35808 = n35807 ^ n35805 ^ 1'b0 ;
  assign n35809 = n11310 | n22229 ;
  assign n35810 = n3761 & ~n7320 ;
  assign n35811 = n35810 ^ n10320 ^ 1'b0 ;
  assign n35812 = n13190 & n35811 ;
  assign n35813 = n35812 ^ n2538 ^ 1'b0 ;
  assign n35814 = n35813 ^ n20882 ^ n1779 ;
  assign n35815 = ( n3807 & ~n17667 ) | ( n3807 & n30846 ) | ( ~n17667 & n30846 ) ;
  assign n35816 = n3985 | n29316 ;
  assign n35817 = n35816 ^ n18942 ^ 1'b0 ;
  assign n35822 = ~n10120 & n28545 ;
  assign n35823 = n35822 ^ n10103 ^ 1'b0 ;
  assign n35824 = n6548 & n35823 ;
  assign n35818 = n11139 | n19008 ;
  assign n35819 = n35818 ^ n1036 ^ 1'b0 ;
  assign n35820 = n713 & n35819 ;
  assign n35821 = n35820 ^ n34677 ^ n20016 ;
  assign n35825 = n35824 ^ n35821 ^ 1'b0 ;
  assign n35826 = n18483 ^ n14968 ^ 1'b0 ;
  assign n35827 = n10692 & ~n35826 ;
  assign n35828 = n6103 | n27765 ;
  assign n35829 = n35828 ^ n3149 ^ 1'b0 ;
  assign n35830 = n16030 & n35829 ;
  assign n35831 = ~n35827 & n35830 ;
  assign n35832 = n6986 & ~n18392 ;
  assign n35833 = ( n12104 & ~n35212 ) | ( n12104 & n35832 ) | ( ~n35212 & n35832 ) ;
  assign n35834 = ~n19176 & n35833 ;
  assign n35836 = ( ~n15806 & n17544 ) | ( ~n15806 & n20091 ) | ( n17544 & n20091 ) ;
  assign n35835 = n20584 ^ n9148 ^ 1'b0 ;
  assign n35837 = n35836 ^ n35835 ^ n3097 ;
  assign n35839 = ( n10570 & n15494 ) | ( n10570 & ~n22106 ) | ( n15494 & ~n22106 ) ;
  assign n35838 = n358 | n5895 ;
  assign n35840 = n35839 ^ n35838 ^ 1'b0 ;
  assign n35841 = ( n5399 & n21532 ) | ( n5399 & ~n35840 ) | ( n21532 & ~n35840 ) ;
  assign n35842 = ( n11725 & n26987 ) | ( n11725 & ~n35841 ) | ( n26987 & ~n35841 ) ;
  assign n35843 = n10399 & ~n25959 ;
  assign n35844 = n35843 ^ n24166 ^ 1'b0 ;
  assign n35845 = ( n34241 & n35486 ) | ( n34241 & ~n35844 ) | ( n35486 & ~n35844 ) ;
  assign n35852 = n3363 & n5886 ;
  assign n35853 = ~n12688 & n35852 ;
  assign n35854 = n35853 ^ n6463 ^ n1922 ;
  assign n35847 = n2168 ^ n1570 ^ 1'b0 ;
  assign n35848 = n35847 ^ n10706 ^ 1'b0 ;
  assign n35849 = ~n541 & n35848 ;
  assign n35846 = ( n5392 & n9946 ) | ( n5392 & n16712 ) | ( n9946 & n16712 ) ;
  assign n35850 = n35849 ^ n35846 ^ n19144 ;
  assign n35851 = n35709 & ~n35850 ;
  assign n35855 = n35854 ^ n35851 ^ 1'b0 ;
  assign n35856 = n35855 ^ n9854 ^ n1319 ;
  assign n35857 = n24893 ^ x123 ^ 1'b0 ;
  assign n35858 = n10874 & n35857 ;
  assign n35859 = n15112 ^ n3586 ^ 1'b0 ;
  assign n35860 = n23637 & ~n35859 ;
  assign n35861 = ( ~n15958 & n35858 ) | ( ~n15958 & n35860 ) | ( n35858 & n35860 ) ;
  assign n35862 = n29965 ^ n1510 ^ 1'b0 ;
  assign n35863 = n18071 & ~n35862 ;
  assign n35864 = n35527 ^ n13990 ^ n1295 ;
  assign n35865 = n9807 & ~n35864 ;
  assign n35866 = n22302 & n35865 ;
  assign n35867 = n973 | n22747 ;
  assign n35868 = n35867 ^ n27865 ^ 1'b0 ;
  assign n35869 = n15219 | n35868 ;
  assign n35870 = ~n9312 & n11726 ;
  assign n35871 = n23951 & n35870 ;
  assign n35872 = ~n1826 & n5189 ;
  assign n35873 = n7563 | n35872 ;
  assign n35874 = n35873 ^ n5047 ^ 1'b0 ;
  assign n35875 = ( ~n14823 & n20458 ) | ( ~n14823 & n35874 ) | ( n20458 & n35874 ) ;
  assign n35876 = ( ~n11429 & n17156 ) | ( ~n11429 & n19916 ) | ( n17156 & n19916 ) ;
  assign n35877 = ( x17 & ~n5595 ) | ( x17 & n6115 ) | ( ~n5595 & n6115 ) ;
  assign n35878 = n35877 ^ n34400 ^ 1'b0 ;
  assign n35879 = ~n7840 & n31354 ;
  assign n35880 = n35879 ^ n21342 ^ 1'b0 ;
  assign n35881 = ~n1826 & n11552 ;
  assign n35882 = n35881 ^ n8219 ^ 1'b0 ;
  assign n35883 = n24106 ^ n9524 ^ 1'b0 ;
  assign n35884 = n35882 | n35883 ;
  assign n35885 = ~n5599 & n6136 ;
  assign n35886 = n19539 & n35885 ;
  assign n35887 = n14340 & ~n35886 ;
  assign n35888 = n13652 ^ n5036 ^ 1'b0 ;
  assign n35889 = ( n3353 & ~n27985 ) | ( n3353 & n33506 ) | ( ~n27985 & n33506 ) ;
  assign n35890 = ( ~n10472 & n23124 ) | ( ~n10472 & n26171 ) | ( n23124 & n26171 ) ;
  assign n35891 = ~n7502 & n15204 ;
  assign n35892 = n35891 ^ n14685 ^ n13328 ;
  assign n35893 = ~n6557 & n35892 ;
  assign n35894 = ( n2864 & n30461 ) | ( n2864 & ~n35893 ) | ( n30461 & ~n35893 ) ;
  assign n35895 = n9140 ^ n8104 ^ n6902 ;
  assign n35896 = ( n7374 & n35894 ) | ( n7374 & n35895 ) | ( n35894 & n35895 ) ;
  assign n35897 = n34376 ^ n24854 ^ n23070 ;
  assign n35898 = n35897 ^ n14387 ^ 1'b0 ;
  assign n35899 = n15725 | n35898 ;
  assign n35900 = ~n3885 & n34706 ;
  assign n35901 = n1545 & n35900 ;
  assign n35902 = n23756 ^ n8689 ^ 1'b0 ;
  assign n35903 = n29711 & n35902 ;
  assign n35904 = ( ~n489 & n2903 ) | ( ~n489 & n12634 ) | ( n2903 & n12634 ) ;
  assign n35905 = ( ~n3117 & n15222 ) | ( ~n3117 & n35904 ) | ( n15222 & n35904 ) ;
  assign n35906 = n7906 & n35905 ;
  assign n35907 = n4522 & n12003 ;
  assign n35908 = n35907 ^ n10220 ^ 1'b0 ;
  assign n35909 = n1680 & n1770 ;
  assign n35910 = ~n12036 & n35909 ;
  assign n35911 = n35908 & ~n35910 ;
  assign n35914 = n10071 ^ n5399 ^ n2928 ;
  assign n35915 = n8745 & ~n25249 ;
  assign n35916 = ~n35914 & n35915 ;
  assign n35913 = ( n7206 & n7285 ) | ( n7206 & ~n26599 ) | ( n7285 & ~n26599 ) ;
  assign n35917 = n35916 ^ n35913 ^ n16351 ;
  assign n35912 = n26978 ^ n25840 ^ 1'b0 ;
  assign n35918 = n35917 ^ n35912 ^ n489 ;
  assign n35919 = n19052 ^ n15889 ^ n15057 ;
  assign n35920 = n7188 | n35919 ;
  assign n35921 = n9558 ^ n4305 ^ 1'b0 ;
  assign n35922 = ~n19117 & n35921 ;
  assign n35923 = n35922 ^ n7885 ^ n4230 ;
  assign n35925 = n3353 | n16399 ;
  assign n35926 = n35925 ^ n6848 ^ 1'b0 ;
  assign n35924 = n7141 & n13674 ;
  assign n35927 = n35926 ^ n35924 ^ 1'b0 ;
  assign n35928 = ( n35920 & n35923 ) | ( n35920 & n35927 ) | ( n35923 & n35927 ) ;
  assign n35929 = ( n17501 & n29520 ) | ( n17501 & n31784 ) | ( n29520 & n31784 ) ;
  assign n35930 = n2577 & ~n2997 ;
  assign n35931 = n35929 & n35930 ;
  assign n35932 = ( ~n6113 & n16019 ) | ( ~n6113 & n25095 ) | ( n16019 & n25095 ) ;
  assign n35933 = n35932 ^ n15451 ^ 1'b0 ;
  assign n35934 = n1431 & n35933 ;
  assign n35935 = n25575 ^ n6053 ^ 1'b0 ;
  assign n35939 = n22135 ^ n21924 ^ n12943 ;
  assign n35937 = ( n800 & n7660 ) | ( n800 & n27449 ) | ( n7660 & n27449 ) ;
  assign n35936 = ( n2069 & n11086 ) | ( n2069 & n27536 ) | ( n11086 & n27536 ) ;
  assign n35938 = n35937 ^ n35936 ^ n29155 ;
  assign n35940 = n35939 ^ n35938 ^ n13198 ;
  assign n35941 = n34360 ^ n9397 ^ n1224 ;
  assign n35942 = ( n6462 & n18966 ) | ( n6462 & n35941 ) | ( n18966 & n35941 ) ;
  assign n35943 = ( n6028 & n23642 ) | ( n6028 & ~n26992 ) | ( n23642 & ~n26992 ) ;
  assign n35944 = n7904 | n27475 ;
  assign n35945 = n28438 ^ n22032 ^ n8725 ;
  assign n35946 = n27026 ^ n25515 ^ n11956 ;
  assign n35947 = n35946 ^ n12062 ^ n7216 ;
  assign n35948 = ( n35944 & n35945 ) | ( n35944 & ~n35947 ) | ( n35945 & ~n35947 ) ;
  assign n35949 = n32749 ^ n25157 ^ n20207 ;
  assign n35950 = n14175 & ~n32163 ;
  assign n35951 = n35950 ^ n22254 ^ n2759 ;
  assign n35952 = ~n16052 & n35951 ;
  assign n35955 = ( n3144 & n3690 ) | ( n3144 & ~n22296 ) | ( n3690 & ~n22296 ) ;
  assign n35953 = n6525 ^ n6329 ^ n739 ;
  assign n35954 = n8418 | n35953 ;
  assign n35956 = n35955 ^ n35954 ^ 1'b0 ;
  assign n35957 = n11747 & n12626 ;
  assign n35958 = n35957 ^ n22150 ^ 1'b0 ;
  assign n35961 = n13618 ^ n13030 ^ n11974 ;
  assign n35959 = ( n20747 & ~n24041 ) | ( n20747 & n33458 ) | ( ~n24041 & n33458 ) ;
  assign n35960 = n31612 & ~n35959 ;
  assign n35962 = n35961 ^ n35960 ^ 1'b0 ;
  assign n35963 = n836 | n10475 ;
  assign n35964 = n836 & ~n35963 ;
  assign n35965 = n11386 & ~n14392 ;
  assign n35966 = n6902 & n35965 ;
  assign n35967 = ( n9697 & ~n35964 ) | ( n9697 & n35966 ) | ( ~n35964 & n35966 ) ;
  assign n35968 = ( ~n3413 & n3502 ) | ( ~n3413 & n9027 ) | ( n3502 & n9027 ) ;
  assign n35969 = n1633 & ~n35968 ;
  assign n35970 = n22778 ^ n19089 ^ n5874 ;
  assign n35971 = n35970 ^ n9115 ^ 1'b0 ;
  assign n35972 = n2684 | n20535 ;
  assign n35973 = n35972 ^ n24436 ^ 1'b0 ;
  assign n35977 = n12814 | n25756 ;
  assign n35978 = n35977 ^ n27419 ^ 1'b0 ;
  assign n35974 = ~n19344 & n21355 ;
  assign n35975 = ( n24411 & ~n34932 ) | ( n24411 & n35974 ) | ( ~n34932 & n35974 ) ;
  assign n35976 = n35284 & ~n35975 ;
  assign n35979 = n35978 ^ n35976 ^ 1'b0 ;
  assign n35980 = n35979 ^ n25749 ^ n12710 ;
  assign n35981 = ~n13144 & n28096 ;
  assign n35982 = ( ~n12454 & n18830 ) | ( ~n12454 & n20564 ) | ( n18830 & n20564 ) ;
  assign n35987 = n10902 ^ n9177 ^ 1'b0 ;
  assign n35988 = n9062 & ~n35987 ;
  assign n35983 = n13484 & n15645 ;
  assign n35984 = n35983 ^ n844 ^ 1'b0 ;
  assign n35985 = n7696 & n35984 ;
  assign n35986 = n35985 ^ n9319 ^ 1'b0 ;
  assign n35989 = n35988 ^ n35986 ^ 1'b0 ;
  assign n35990 = n20797 ^ n16655 ^ 1'b0 ;
  assign n35991 = n5943 & ~n20450 ;
  assign n35992 = n35991 ^ n5054 ^ 1'b0 ;
  assign n35993 = ( n33795 & n35990 ) | ( n33795 & ~n35992 ) | ( n35990 & ~n35992 ) ;
  assign n35994 = n13405 ^ n5235 ^ 1'b0 ;
  assign n35995 = n2624 & n35994 ;
  assign n35996 = n35995 ^ n14249 ^ n13168 ;
  assign n35997 = ( n14132 & ~n35320 ) | ( n14132 & n35996 ) | ( ~n35320 & n35996 ) ;
  assign n35998 = n8170 | n11004 ;
  assign n35999 = n12493 & ~n35998 ;
  assign n36000 = n18415 | n35999 ;
  assign n36001 = n12766 | n36000 ;
  assign n36002 = x116 & ~n17225 ;
  assign n36003 = n18572 & n36002 ;
  assign n36005 = n19348 | n22539 ;
  assign n36004 = n327 | n11166 ;
  assign n36006 = n36005 ^ n36004 ^ 1'b0 ;
  assign n36007 = n5444 & ~n36006 ;
  assign n36008 = n9591 ^ n9570 ^ n3347 ;
  assign n36009 = ( n4784 & ~n21475 ) | ( n4784 & n36008 ) | ( ~n21475 & n36008 ) ;
  assign n36010 = n36009 ^ n14790 ^ n12681 ;
  assign n36011 = n34411 ^ n29135 ^ n24192 ;
  assign n36012 = ~n25424 & n36011 ;
  assign n36013 = ( n13567 & n19087 ) | ( n13567 & ~n23431 ) | ( n19087 & ~n23431 ) ;
  assign n36014 = n31113 ^ n14653 ^ n4786 ;
  assign n36015 = n33999 | n36014 ;
  assign n36016 = n36015 ^ n12593 ^ 1'b0 ;
  assign n36017 = n1416 & ~n18630 ;
  assign n36018 = ( n36013 & n36016 ) | ( n36013 & n36017 ) | ( n36016 & n36017 ) ;
  assign n36019 = n16730 ^ n7766 ^ 1'b0 ;
  assign n36020 = ~n24966 & n36019 ;
  assign n36021 = n30057 ^ n7960 ^ n2592 ;
  assign n36024 = ( ~x31 & n7036 ) | ( ~x31 & n11296 ) | ( n7036 & n11296 ) ;
  assign n36022 = n4880 ^ n3785 ^ 1'b0 ;
  assign n36023 = ~n30714 & n36022 ;
  assign n36025 = n36024 ^ n36023 ^ 1'b0 ;
  assign n36026 = n36025 ^ n30098 ^ n27632 ;
  assign n36027 = n15673 ^ n10230 ^ n7280 ;
  assign n36028 = n36027 ^ n2142 ^ 1'b0 ;
  assign n36029 = ( n15959 & ~n17975 ) | ( n15959 & n18400 ) | ( ~n17975 & n18400 ) ;
  assign n36030 = n36029 ^ n34001 ^ n33836 ;
  assign n36031 = ~n4994 & n8949 ;
  assign n36032 = n36031 ^ n1904 ^ 1'b0 ;
  assign n36033 = n15567 & n26178 ;
  assign n36034 = n36033 ^ n20379 ^ 1'b0 ;
  assign n36035 = n14391 ^ n12599 ^ 1'b0 ;
  assign n36036 = n30564 & n36035 ;
  assign n36037 = n36036 ^ n30968 ^ n16032 ;
  assign n36038 = n4478 & ~n6237 ;
  assign n36039 = n36038 ^ n358 ^ 1'b0 ;
  assign n36040 = ( n10845 & n21174 ) | ( n10845 & n36039 ) | ( n21174 & n36039 ) ;
  assign n36041 = n21901 ^ n15148 ^ 1'b0 ;
  assign n36042 = ~n5511 & n36041 ;
  assign n36043 = ~n11487 & n36042 ;
  assign n36044 = n5521 ^ n5118 ^ 1'b0 ;
  assign n36045 = n34478 ^ n18836 ^ n8667 ;
  assign n36046 = n3562 | n18995 ;
  assign n36047 = n36045 & ~n36046 ;
  assign n36049 = n2495 | n23303 ;
  assign n36050 = n36049 ^ n332 ^ 1'b0 ;
  assign n36051 = n11445 | n36050 ;
  assign n36048 = n24849 | n27978 ;
  assign n36052 = n36051 ^ n36048 ^ 1'b0 ;
  assign n36053 = ( n3943 & ~n8583 ) | ( n3943 & n28691 ) | ( ~n8583 & n28691 ) ;
  assign n36054 = ~n21007 & n36053 ;
  assign n36055 = n1084 & ~n16334 ;
  assign n36056 = n36055 ^ n2069 ^ 1'b0 ;
  assign n36057 = n36056 ^ n18807 ^ 1'b0 ;
  assign n36058 = n23534 ^ n22781 ^ n17117 ;
  assign n36059 = n36058 ^ n29629 ^ n12075 ;
  assign n36060 = n20301 ^ n9037 ^ n6871 ;
  assign n36061 = n36060 ^ n35255 ^ n15475 ;
  assign n36062 = ( n9582 & ~n18316 ) | ( n9582 & n21922 ) | ( ~n18316 & n21922 ) ;
  assign n36063 = n6304 ^ n4659 ^ n711 ;
  assign n36064 = ~n7330 & n36063 ;
  assign n36065 = ~n14340 & n36064 ;
  assign n36066 = n36065 ^ n14583 ^ n10052 ;
  assign n36067 = n1077 & ~n31268 ;
  assign n36068 = n14593 ^ n8205 ^ 1'b0 ;
  assign n36069 = n34411 | n36068 ;
  assign n36070 = n17843 | n27671 ;
  assign n36071 = n14545 | n36070 ;
  assign n36072 = n25791 & ~n36071 ;
  assign n36073 = n28264 & n36072 ;
  assign n36074 = ( n14576 & ~n15187 ) | ( n14576 & n36073 ) | ( ~n15187 & n36073 ) ;
  assign n36075 = n5192 & n5648 ;
  assign n36076 = n36075 ^ x107 ^ 1'b0 ;
  assign n36077 = n16474 & n30831 ;
  assign n36078 = n36077 ^ n24837 ^ 1'b0 ;
  assign n36079 = n25948 & ~n36078 ;
  assign n36080 = ( n26682 & n36076 ) | ( n26682 & n36079 ) | ( n36076 & n36079 ) ;
  assign n36081 = n29628 ^ n2429 ^ 1'b0 ;
  assign n36082 = n4307 & n36081 ;
  assign n36083 = n36082 ^ n23023 ^ 1'b0 ;
  assign n36084 = n36083 ^ n31818 ^ n12654 ;
  assign n36085 = ~n6218 & n10991 ;
  assign n36086 = n36085 ^ n14607 ^ 1'b0 ;
  assign n36087 = ( ~n1534 & n18317 ) | ( ~n1534 & n36086 ) | ( n18317 & n36086 ) ;
  assign n36088 = ( ~n5175 & n24014 ) | ( ~n5175 & n36087 ) | ( n24014 & n36087 ) ;
  assign n36089 = ( n8564 & n10321 ) | ( n8564 & n11020 ) | ( n10321 & n11020 ) ;
  assign n36090 = n36089 ^ n1761 ^ 1'b0 ;
  assign n36091 = n36088 | n36090 ;
  assign n36092 = n20742 ^ n5857 ^ n5410 ;
  assign n36093 = n9211 ^ n3779 ^ 1'b0 ;
  assign n36094 = n36093 ^ n10778 ^ 1'b0 ;
  assign n36095 = ( ~n18091 & n26851 ) | ( ~n18091 & n36094 ) | ( n26851 & n36094 ) ;
  assign n36096 = ( ~n7438 & n36092 ) | ( ~n7438 & n36095 ) | ( n36092 & n36095 ) ;
  assign n36097 = n30473 | n36096 ;
  assign n36098 = n20677 & ~n36097 ;
  assign n36099 = n20582 ^ n19832 ^ n307 ;
  assign n36100 = n36099 ^ n17283 ^ n5114 ;
  assign n36101 = ( ~n3107 & n8420 ) | ( ~n3107 & n29559 ) | ( n8420 & n29559 ) ;
  assign n36102 = n36101 ^ n25150 ^ x132 ;
  assign n36103 = ( ~n28510 & n36100 ) | ( ~n28510 & n36102 ) | ( n36100 & n36102 ) ;
  assign n36104 = ( n4387 & n18981 ) | ( n4387 & n36103 ) | ( n18981 & n36103 ) ;
  assign n36105 = ( ~n6213 & n12098 ) | ( ~n6213 & n24123 ) | ( n12098 & n24123 ) ;
  assign n36106 = n17204 ^ n6031 ^ n2799 ;
  assign n36107 = ( n3829 & n27247 ) | ( n3829 & ~n36106 ) | ( n27247 & ~n36106 ) ;
  assign n36108 = ( n4686 & ~n11432 ) | ( n4686 & n36107 ) | ( ~n11432 & n36107 ) ;
  assign n36109 = n36108 ^ n17540 ^ n3900 ;
  assign n36110 = ~n14503 & n18735 ;
  assign n36111 = n36110 ^ n23559 ^ 1'b0 ;
  assign n36112 = n26073 & n29928 ;
  assign n36113 = ~n7942 & n36112 ;
  assign n36114 = n5846 & ~n13855 ;
  assign n36115 = n36113 & n36114 ;
  assign n36116 = n19144 ^ x2 ^ 1'b0 ;
  assign n36117 = ( ~n4339 & n23375 ) | ( ~n4339 & n36116 ) | ( n23375 & n36116 ) ;
  assign n36118 = n36117 ^ n15014 ^ 1'b0 ;
  assign n36119 = n5703 & ~n36118 ;
  assign n36120 = n14773 & n25425 ;
  assign n36121 = n17264 & n25534 ;
  assign n36122 = n36121 ^ n19885 ^ 1'b0 ;
  assign n36123 = ~n3326 & n19849 ;
  assign n36124 = ( n9835 & n14501 ) | ( n9835 & n20432 ) | ( n14501 & n20432 ) ;
  assign n36125 = ( n14408 & n19477 ) | ( n14408 & ~n36124 ) | ( n19477 & ~n36124 ) ;
  assign n36126 = n33983 ^ n10739 ^ 1'b0 ;
  assign n36127 = n20934 & ~n36126 ;
  assign n36128 = ( n11991 & n17244 ) | ( n11991 & ~n36127 ) | ( n17244 & ~n36127 ) ;
  assign n36129 = n36128 ^ n19014 ^ n1261 ;
  assign n36130 = n514 & ~n4309 ;
  assign n36131 = n36130 ^ n18008 ^ n13730 ;
  assign n36132 = n6750 & ~n36131 ;
  assign n36133 = n5282 | n20033 ;
  assign n36134 = n10862 | n36133 ;
  assign n36135 = n9282 & ~n23813 ;
  assign n36136 = n30949 & n36135 ;
  assign n36137 = n7634 & ~n13831 ;
  assign n36138 = n15728 ^ n7418 ^ n7344 ;
  assign n36139 = n36138 ^ n19560 ^ 1'b0 ;
  assign n36140 = n8288 & n36139 ;
  assign n36141 = ( n7994 & n10307 ) | ( n7994 & n36140 ) | ( n10307 & n36140 ) ;
  assign n36142 = ( ~n2478 & n14894 ) | ( ~n2478 & n25271 ) | ( n14894 & n25271 ) ;
  assign n36143 = ( n12948 & n36141 ) | ( n12948 & n36142 ) | ( n36141 & n36142 ) ;
  assign n36144 = ( n1164 & n36137 ) | ( n1164 & ~n36143 ) | ( n36137 & ~n36143 ) ;
  assign n36145 = ( n22136 & ~n25448 ) | ( n22136 & n25654 ) | ( ~n25448 & n25654 ) ;
  assign n36146 = ( n8042 & ~n15418 ) | ( n8042 & n31941 ) | ( ~n15418 & n31941 ) ;
  assign n36147 = n27640 ^ n10039 ^ 1'b0 ;
  assign n36148 = ~n29243 & n36147 ;
  assign n36149 = n15492 & n36148 ;
  assign n36150 = n36149 ^ n35070 ^ n28291 ;
  assign n36151 = n31234 ^ n10353 ^ 1'b0 ;
  assign n36152 = n24820 & n36151 ;
  assign n36153 = n18466 ^ n17363 ^ 1'b0 ;
  assign n36154 = n36153 ^ n7658 ^ 1'b0 ;
  assign n36155 = n36152 & ~n36154 ;
  assign n36156 = n15974 & ~n32177 ;
  assign n36157 = n29921 ^ n2501 ^ 1'b0 ;
  assign n36158 = n3962 & n24793 ;
  assign n36159 = n36158 ^ n13320 ^ 1'b0 ;
  assign n36162 = n13411 | n31393 ;
  assign n36160 = n10417 & n30800 ;
  assign n36161 = n36160 ^ n35340 ^ 1'b0 ;
  assign n36163 = n36162 ^ n36161 ^ 1'b0 ;
  assign n36165 = n25061 ^ n16271 ^ n555 ;
  assign n36164 = ( n12304 & n14834 ) | ( n12304 & ~n15013 ) | ( n14834 & ~n15013 ) ;
  assign n36166 = n36165 ^ n36164 ^ n31872 ;
  assign n36168 = n14078 ^ n266 ^ 1'b0 ;
  assign n36169 = ~n8935 & n36168 ;
  assign n36167 = n5702 | n11678 ;
  assign n36170 = n36169 ^ n36167 ^ 1'b0 ;
  assign n36171 = ( ~n11968 & n30609 ) | ( ~n11968 & n36170 ) | ( n30609 & n36170 ) ;
  assign n36172 = n13661 & n18782 ;
  assign n36173 = ~n28103 & n36172 ;
  assign n36174 = n36173 ^ n3869 ^ 1'b0 ;
  assign n36175 = n16386 & n25740 ;
  assign n36176 = n36175 ^ n24767 ^ 1'b0 ;
  assign n36177 = ( ~n3475 & n23034 ) | ( ~n3475 & n36176 ) | ( n23034 & n36176 ) ;
  assign n36178 = n36177 ^ n30377 ^ 1'b0 ;
  assign n36179 = ( ~n5072 & n16458 ) | ( ~n5072 & n30088 ) | ( n16458 & n30088 ) ;
  assign n36180 = n8499 & ~n36179 ;
  assign n36181 = n36180 ^ n12284 ^ 1'b0 ;
  assign n36182 = n1580 & ~n34848 ;
  assign n36183 = ( n23390 & ~n24582 ) | ( n23390 & n36182 ) | ( ~n24582 & n36182 ) ;
  assign n36184 = n5666 & ~n7160 ;
  assign n36185 = n36183 & n36184 ;
  assign n36186 = n12640 | n29304 ;
  assign n36187 = n5118 | n8563 ;
  assign n36188 = ( ~n12340 & n13786 ) | ( ~n12340 & n36187 ) | ( n13786 & n36187 ) ;
  assign n36189 = n7638 | n14422 ;
  assign n36190 = n36189 ^ n9938 ^ n4933 ;
  assign n36191 = n20741 ^ n15663 ^ n11051 ;
  assign n36192 = n18340 | n36191 ;
  assign n36193 = ( n25786 & n36190 ) | ( n25786 & n36192 ) | ( n36190 & n36192 ) ;
  assign n36194 = ~n12559 & n25394 ;
  assign n36195 = n36194 ^ n23805 ^ n23551 ;
  assign n36196 = ( ~n3943 & n12976 ) | ( ~n3943 & n14656 ) | ( n12976 & n14656 ) ;
  assign n36197 = n11728 ^ n4638 ^ n3947 ;
  assign n36198 = n36197 ^ n15475 ^ 1'b0 ;
  assign n36199 = n18348 ^ n5460 ^ 1'b0 ;
  assign n36200 = ~n36198 & n36199 ;
  assign n36201 = ( n481 & n28177 ) | ( n481 & ~n36200 ) | ( n28177 & ~n36200 ) ;
  assign n36202 = n36201 ^ n23246 ^ n13492 ;
  assign n36204 = ( ~n407 & n21021 ) | ( ~n407 & n23261 ) | ( n21021 & n23261 ) ;
  assign n36203 = n35047 ^ n21377 ^ 1'b0 ;
  assign n36205 = n36204 ^ n36203 ^ n19338 ;
  assign n36206 = n19992 ^ n4283 ^ 1'b0 ;
  assign n36207 = ~n11107 & n36206 ;
  assign n36208 = n2633 & n14050 ;
  assign n36209 = x28 & ~n33564 ;
  assign n36210 = ~n36208 & n36209 ;
  assign n36211 = ~n3465 & n10468 ;
  assign n36212 = n36211 ^ n742 ^ 1'b0 ;
  assign n36213 = ( n10395 & n15394 ) | ( n10395 & ~n36212 ) | ( n15394 & ~n36212 ) ;
  assign n36214 = n36213 ^ n10412 ^ n3525 ;
  assign n36216 = n19528 ^ x67 ^ 1'b0 ;
  assign n36217 = n10930 & ~n36216 ;
  assign n36218 = n36217 ^ n15781 ^ n10400 ;
  assign n36219 = n36198 ^ n19356 ^ 1'b0 ;
  assign n36220 = n36218 & ~n36219 ;
  assign n36215 = n17523 ^ n14116 ^ n12345 ;
  assign n36221 = n36220 ^ n36215 ^ n18654 ;
  assign n36222 = n2596 | n12817 ;
  assign n36223 = n19531 ^ n591 ^ 1'b0 ;
  assign n36224 = ~n12678 & n32460 ;
  assign n36225 = n21483 & ~n36224 ;
  assign n36226 = n17814 ^ n6590 ^ 1'b0 ;
  assign n36227 = n35023 ^ n4570 ^ n3514 ;
  assign n36228 = n24667 ^ n16825 ^ 1'b0 ;
  assign n36229 = n36228 ^ n13358 ^ n13158 ;
  assign n36230 = ( n2388 & n16334 ) | ( n2388 & n36229 ) | ( n16334 & n36229 ) ;
  assign n36231 = n9593 & ~n33543 ;
  assign n36232 = n12446 ^ n8288 ^ 1'b0 ;
  assign n36233 = ~n7887 & n36232 ;
  assign n36234 = ( n2120 & n11298 ) | ( n2120 & ~n36233 ) | ( n11298 & ~n36233 ) ;
  assign n36235 = n16969 & ~n19525 ;
  assign n36236 = n36235 ^ n14437 ^ n1924 ;
  assign n36237 = ( n18008 & ~n31708 ) | ( n18008 & n35142 ) | ( ~n31708 & n35142 ) ;
  assign n36238 = n36236 | n36237 ;
  assign n36239 = n36234 & ~n36238 ;
  assign n36240 = n6389 & ~n34258 ;
  assign n36241 = ~n33761 & n33979 ;
  assign n36242 = ~n36240 & n36241 ;
  assign n36243 = n25085 & ~n27759 ;
  assign n36244 = n36243 ^ n8647 ^ 1'b0 ;
  assign n36245 = n16553 ^ n6123 ^ n3750 ;
  assign n36248 = n29668 ^ n28010 ^ n22150 ;
  assign n36246 = n22321 ^ n21373 ^ 1'b0 ;
  assign n36247 = ~n6998 & n36246 ;
  assign n36249 = n36248 ^ n36247 ^ n30809 ;
  assign n36250 = ~n327 & n7547 ;
  assign n36251 = ~n14246 & n36250 ;
  assign n36252 = ~n1531 & n35897 ;
  assign n36253 = n36252 ^ n9263 ^ 1'b0 ;
  assign n36254 = ( n6421 & n11553 ) | ( n6421 & n20062 ) | ( n11553 & n20062 ) ;
  assign n36255 = n36254 ^ n4240 ^ 1'b0 ;
  assign n36256 = n16456 | n36255 ;
  assign n36257 = n36255 & ~n36256 ;
  assign n36258 = n1914 & ~n25396 ;
  assign n36259 = n36258 ^ n13661 ^ 1'b0 ;
  assign n36260 = n36259 ^ n34416 ^ n28225 ;
  assign n36261 = n7824 ^ n6773 ^ 1'b0 ;
  assign n36262 = n4783 | n36261 ;
  assign n36263 = n36262 ^ n8282 ^ 1'b0 ;
  assign n36264 = n36263 ^ n13926 ^ n618 ;
  assign n36265 = n34368 ^ n21199 ^ n20493 ;
  assign n36266 = ~n10699 & n34426 ;
  assign n36267 = n36266 ^ n28774 ^ 1'b0 ;
  assign n36268 = n27222 ^ n11478 ^ n666 ;
  assign n36269 = ( ~n2851 & n6729 ) | ( ~n2851 & n18004 ) | ( n6729 & n18004 ) ;
  assign n36270 = n29879 & ~n36269 ;
  assign n36271 = n17220 ^ n7102 ^ n301 ;
  assign n36272 = ( n2628 & ~n36270 ) | ( n2628 & n36271 ) | ( ~n36270 & n36271 ) ;
  assign n36273 = ( n5799 & n25114 ) | ( n5799 & ~n36272 ) | ( n25114 & ~n36272 ) ;
  assign n36274 = n9271 & ~n10283 ;
  assign n36275 = n3117 & n36274 ;
  assign n36276 = ( n3236 & n3731 ) | ( n3236 & ~n6428 ) | ( n3731 & ~n6428 ) ;
  assign n36277 = ( ~n20382 & n36275 ) | ( ~n20382 & n36276 ) | ( n36275 & n36276 ) ;
  assign n36278 = ( n6582 & n12592 ) | ( n6582 & n36277 ) | ( n12592 & n36277 ) ;
  assign n36279 = n35922 ^ n20945 ^ 1'b0 ;
  assign n36280 = n13794 ^ n3517 ^ 1'b0 ;
  assign n36281 = n36279 | n36280 ;
  assign n36282 = n16529 & ~n36281 ;
  assign n36283 = n1403 | n3564 ;
  assign n36284 = n36283 ^ n24433 ^ x124 ;
  assign n36285 = n23501 ^ n13394 ^ n7954 ;
  assign n36286 = n3036 & n21905 ;
  assign n36287 = n4913 & n36286 ;
  assign n36288 = ( n11881 & n36285 ) | ( n11881 & n36287 ) | ( n36285 & n36287 ) ;
  assign n36289 = ( n523 & n6774 ) | ( n523 & n24570 ) | ( n6774 & n24570 ) ;
  assign n36290 = n8000 & ~n35874 ;
  assign n36292 = n8701 | n18101 ;
  assign n36293 = n36292 ^ n8864 ^ 1'b0 ;
  assign n36291 = n1356 & ~n8579 ;
  assign n36294 = n36293 ^ n36291 ^ 1'b0 ;
  assign n36295 = n36294 ^ n12312 ^ 1'b0 ;
  assign n36296 = n36295 ^ n4978 ^ 1'b0 ;
  assign n36297 = n2990 & ~n18025 ;
  assign n36298 = ( n4057 & n12239 ) | ( n4057 & n22624 ) | ( n12239 & n22624 ) ;
  assign n36299 = n36298 ^ n381 ^ 1'b0 ;
  assign n36300 = ~n4927 & n13210 ;
  assign n36301 = n36300 ^ n13617 ^ 1'b0 ;
  assign n36302 = ( n9491 & ~n16511 ) | ( n9491 & n36301 ) | ( ~n16511 & n36301 ) ;
  assign n36303 = n29317 ^ n12979 ^ n3514 ;
  assign n36304 = n36303 ^ n12122 ^ 1'b0 ;
  assign n36305 = n6413 & n8876 ;
  assign n36306 = ~n36304 & n36305 ;
  assign n36307 = ~n16794 & n26858 ;
  assign n36308 = n19078 & ~n23849 ;
  assign n36309 = ( n4840 & n19626 ) | ( n4840 & ~n36308 ) | ( n19626 & ~n36308 ) ;
  assign n36311 = ( n2740 & n5421 ) | ( n2740 & n14121 ) | ( n5421 & n14121 ) ;
  assign n36312 = ( n10547 & ~n23954 ) | ( n10547 & n36311 ) | ( ~n23954 & n36311 ) ;
  assign n36310 = ( ~n10482 & n16464 ) | ( ~n10482 & n30248 ) | ( n16464 & n30248 ) ;
  assign n36313 = n36312 ^ n36310 ^ n13290 ;
  assign n36314 = ( n20422 & n28674 ) | ( n20422 & n29919 ) | ( n28674 & n29919 ) ;
  assign n36315 = n36314 ^ n17385 ^ 1'b0 ;
  assign n36316 = ( n9924 & n28302 ) | ( n9924 & ~n36315 ) | ( n28302 & ~n36315 ) ;
  assign n36319 = n17807 ^ n2350 ^ n719 ;
  assign n36317 = n33702 ^ n27105 ^ 1'b0 ;
  assign n36318 = n26468 | n36317 ;
  assign n36320 = n36319 ^ n36318 ^ n33449 ;
  assign n36321 = ( n380 & ~n1840 ) | ( n380 & n5939 ) | ( ~n1840 & n5939 ) ;
  assign n36322 = n36321 ^ n11868 ^ n9680 ;
  assign n36323 = ( n15698 & n25248 ) | ( n15698 & ~n30464 ) | ( n25248 & ~n30464 ) ;
  assign n36324 = ~n23985 & n30864 ;
  assign n36325 = n36324 ^ n8538 ^ 1'b0 ;
  assign n36326 = n4612 & ~n18692 ;
  assign n36327 = n8193 ^ n4569 ^ n401 ;
  assign n36328 = n36327 ^ n6077 ^ 1'b0 ;
  assign n36329 = n13555 ^ n7900 ^ n3545 ;
  assign n36330 = ( n11249 & n32516 ) | ( n11249 & n36329 ) | ( n32516 & n36329 ) ;
  assign n36331 = ~n11013 & n35525 ;
  assign n36332 = n32322 & n36331 ;
  assign n36333 = n25772 & ~n36332 ;
  assign n36334 = n4329 ^ n4004 ^ 1'b0 ;
  assign n36335 = ~n29690 & n36203 ;
  assign n36336 = ~n5302 & n36335 ;
  assign n36337 = n2514 & ~n23904 ;
  assign n36338 = n29844 ^ n17753 ^ n14459 ;
  assign n36339 = ( n2763 & n9154 ) | ( n2763 & n10316 ) | ( n9154 & n10316 ) ;
  assign n36340 = ( ~n6668 & n19614 ) | ( ~n6668 & n36339 ) | ( n19614 & n36339 ) ;
  assign n36341 = n36340 ^ n23756 ^ n1173 ;
  assign n36342 = n14954 ^ n7774 ^ 1'b0 ;
  assign n36343 = n36342 ^ n14129 ^ 1'b0 ;
  assign n36344 = ~n20821 & n36343 ;
  assign n36345 = ( ~n36338 & n36341 ) | ( ~n36338 & n36344 ) | ( n36341 & n36344 ) ;
  assign n36346 = ( n1313 & n3804 ) | ( n1313 & ~n8282 ) | ( n3804 & ~n8282 ) ;
  assign n36347 = n36346 ^ n35674 ^ 1'b0 ;
  assign n36348 = n11296 | n18619 ;
  assign n36349 = n36348 ^ n30473 ^ 1'b0 ;
  assign n36350 = n28642 ^ n15641 ^ 1'b0 ;
  assign n36351 = n36350 ^ n22921 ^ n9469 ;
  assign n36352 = n20824 & n36351 ;
  assign n36353 = n31113 ^ n9092 ^ x8 ;
  assign n36354 = n36353 ^ n25067 ^ n2210 ;
  assign n36355 = ( n3867 & n14320 ) | ( n3867 & n36354 ) | ( n14320 & n36354 ) ;
  assign n36356 = n21644 ^ n14697 ^ n14189 ;
  assign n36357 = n1299 | n11824 ;
  assign n36358 = n36357 ^ n18255 ^ 1'b0 ;
  assign n36359 = n30403 ^ n5234 ^ 1'b0 ;
  assign n36360 = n36358 | n36359 ;
  assign n36361 = n17041 ^ n6930 ^ n1064 ;
  assign n36362 = ( n12701 & n30408 ) | ( n12701 & ~n36361 ) | ( n30408 & ~n36361 ) ;
  assign n36363 = n36362 ^ n2572 ^ 1'b0 ;
  assign n36364 = n36360 | n36363 ;
  assign n36365 = n8158 | n14305 ;
  assign n36366 = ( n18703 & n21064 ) | ( n18703 & n36365 ) | ( n21064 & n36365 ) ;
  assign n36367 = n5847 ^ n3738 ^ 1'b0 ;
  assign n36378 = n5728 | n8646 ;
  assign n36379 = n2628 | n36378 ;
  assign n36375 = n761 | n8124 ;
  assign n36376 = n2947 & ~n36375 ;
  assign n36377 = n36376 ^ n8774 ^ 1'b0 ;
  assign n36368 = ( ~n3330 & n21376 ) | ( ~n3330 & n21987 ) | ( n21376 & n21987 ) ;
  assign n36369 = n36368 ^ n30781 ^ 1'b0 ;
  assign n36370 = ( n13984 & n14208 ) | ( n13984 & ~n25153 ) | ( n14208 & ~n25153 ) ;
  assign n36371 = n1556 & n36370 ;
  assign n36372 = ~n11247 & n36371 ;
  assign n36373 = ( n1813 & n12939 ) | ( n1813 & n36372 ) | ( n12939 & n36372 ) ;
  assign n36374 = ( n7714 & n36369 ) | ( n7714 & n36373 ) | ( n36369 & n36373 ) ;
  assign n36380 = n36379 ^ n36377 ^ n36374 ;
  assign n36384 = n1540 & ~n16484 ;
  assign n36385 = ~n18586 & n36384 ;
  assign n36386 = n32526 ^ n9522 ^ 1'b0 ;
  assign n36387 = n36385 | n36386 ;
  assign n36381 = n29502 ^ n14149 ^ n9075 ;
  assign n36382 = n36381 ^ n20559 ^ n11881 ;
  assign n36383 = n10294 & n36382 ;
  assign n36388 = n36387 ^ n36383 ^ 1'b0 ;
  assign n36389 = n19438 & n25637 ;
  assign n36390 = n36389 ^ n26859 ^ 1'b0 ;
  assign n36391 = x87 & n12572 ;
  assign n36392 = n9304 ^ n7396 ^ n5156 ;
  assign n36393 = ( n27389 & n35370 ) | ( n27389 & n36392 ) | ( n35370 & n36392 ) ;
  assign n36394 = n8849 & ~n14991 ;
  assign n36395 = ~n6398 & n8010 ;
  assign n36396 = n36395 ^ n6058 ^ 1'b0 ;
  assign n36397 = ( n26290 & n27212 ) | ( n26290 & n36396 ) | ( n27212 & n36396 ) ;
  assign n36398 = n36397 ^ n33954 ^ 1'b0 ;
  assign n36399 = n19787 & ~n31323 ;
  assign n36400 = n36399 ^ n13222 ^ 1'b0 ;
  assign n36401 = ~n10022 & n36400 ;
  assign n36402 = ( n18056 & n24568 ) | ( n18056 & ~n35281 ) | ( n24568 & ~n35281 ) ;
  assign n36403 = ~n1206 & n2394 ;
  assign n36404 = n17057 & n36403 ;
  assign n36405 = ~n7904 & n22543 ;
  assign n36406 = n36404 & n36405 ;
  assign n36407 = n36406 ^ n31683 ^ n24585 ;
  assign n36408 = n36407 ^ n17237 ^ 1'b0 ;
  assign n36409 = n36402 & n36408 ;
  assign n36410 = ( ~n2537 & n5871 ) | ( ~n2537 & n11266 ) | ( n5871 & n11266 ) ;
  assign n36411 = ( n8419 & n27072 ) | ( n8419 & ~n35117 ) | ( n27072 & ~n35117 ) ;
  assign n36412 = n34236 ^ n13843 ^ 1'b0 ;
  assign n36413 = n36411 & n36412 ;
  assign n36414 = ( ~n29215 & n33312 ) | ( ~n29215 & n36413 ) | ( n33312 & n36413 ) ;
  assign n36415 = n9909 & n11553 ;
  assign n36416 = n35248 & n36415 ;
  assign n36417 = ( n36410 & ~n36414 ) | ( n36410 & n36416 ) | ( ~n36414 & n36416 ) ;
  assign n36418 = n8609 ^ n3902 ^ n2257 ;
  assign n36419 = ( n1088 & n4120 ) | ( n1088 & ~n27949 ) | ( n4120 & ~n27949 ) ;
  assign n36420 = n2777 | n4281 ;
  assign n36421 = n4130 | n36420 ;
  assign n36422 = n5271 & n14394 ;
  assign n36423 = n36422 ^ n20293 ^ n11074 ;
  assign n36424 = n36423 ^ n24630 ^ 1'b0 ;
  assign n36425 = n36421 & n36424 ;
  assign n36426 = n22778 ^ n8684 ^ 1'b0 ;
  assign n36427 = n25837 & ~n36426 ;
  assign n36428 = ~n1494 & n36427 ;
  assign n36429 = n34802 ^ n19957 ^ n5616 ;
  assign n36430 = n29749 ^ n12426 ^ 1'b0 ;
  assign n36431 = n36429 & ~n36430 ;
  assign n36432 = n8092 ^ x140 ^ 1'b0 ;
  assign n36433 = n26975 ^ n19852 ^ n10173 ;
  assign n36434 = n36433 ^ n15917 ^ n10373 ;
  assign n36435 = n36434 ^ n23023 ^ 1'b0 ;
  assign n36436 = n4011 & ~n24380 ;
  assign n36437 = n13211 & n14735 ;
  assign n36438 = n8444 & n36437 ;
  assign n36439 = n6633 & n36438 ;
  assign n36440 = ( ~n19443 & n29261 ) | ( ~n19443 & n30226 ) | ( n29261 & n30226 ) ;
  assign n36441 = n25331 | n30563 ;
  assign n36442 = n36440 & ~n36441 ;
  assign n36443 = n17154 | n23002 ;
  assign n36444 = n22511 & ~n36443 ;
  assign n36445 = n36444 ^ n8007 ^ 1'b0 ;
  assign n36446 = n36445 ^ n20904 ^ n3860 ;
  assign n36447 = n9730 | n10212 ;
  assign n36448 = ~n2914 & n15012 ;
  assign n36449 = ~n1311 & n36448 ;
  assign n36450 = ( n1474 & n35544 ) | ( n1474 & ~n36449 ) | ( n35544 & ~n36449 ) ;
  assign n36451 = n36450 ^ n5869 ^ 1'b0 ;
  assign n36452 = n36451 ^ n33083 ^ n33061 ;
  assign n36453 = n15979 ^ n7224 ^ n5791 ;
  assign n36454 = n6637 & n18946 ;
  assign n36455 = ~n36453 & n36454 ;
  assign n36456 = n36455 ^ n9911 ^ 1'b0 ;
  assign n36457 = n26064 | n36456 ;
  assign n36458 = n36457 ^ n35484 ^ 1'b0 ;
  assign n36459 = n15401 & ~n36458 ;
  assign n36460 = n8627 | n36459 ;
  assign n36461 = ~n20434 & n23235 ;
  assign n36462 = n36461 ^ n4248 ^ 1'b0 ;
  assign n36463 = n23527 | n24867 ;
  assign n36464 = n36463 ^ n29730 ^ 1'b0 ;
  assign n36465 = n18690 & ~n25782 ;
  assign n36466 = n13534 & n36465 ;
  assign n36467 = n20778 & ~n36466 ;
  assign n36468 = ( n2251 & ~n16547 ) | ( n2251 & n28204 ) | ( ~n16547 & n28204 ) ;
  assign n36469 = ( ~n20399 & n32696 ) | ( ~n20399 & n36468 ) | ( n32696 & n36468 ) ;
  assign n36470 = n17231 | n33100 ;
  assign n36471 = n36470 ^ n15623 ^ 1'b0 ;
  assign n36472 = n2638 & n29809 ;
  assign n36473 = ( n1970 & n6388 ) | ( n1970 & ~n36472 ) | ( n6388 & ~n36472 ) ;
  assign n36474 = n30500 ^ n26911 ^ n10582 ;
  assign n36475 = n18509 ^ n5757 ^ 1'b0 ;
  assign n36476 = n12188 | n36475 ;
  assign n36477 = ( n1304 & ~n23867 ) | ( n1304 & n33999 ) | ( ~n23867 & n33999 ) ;
  assign n36478 = ( ~n14049 & n36476 ) | ( ~n14049 & n36477 ) | ( n36476 & n36477 ) ;
  assign n36479 = n36478 ^ n36423 ^ 1'b0 ;
  assign n36480 = ~n10998 & n36479 ;
  assign n36481 = n36042 ^ n10836 ^ 1'b0 ;
  assign n36482 = ~n21525 & n36481 ;
  assign n36483 = n11580 & n20339 ;
  assign n36484 = ~n36482 & n36483 ;
  assign n36485 = n22972 | n26195 ;
  assign n36486 = n2338 | n36485 ;
  assign n36487 = n15850 & ~n32376 ;
  assign n36488 = ( n8968 & n36486 ) | ( n8968 & n36487 ) | ( n36486 & n36487 ) ;
  assign n36491 = n3128 | n4608 ;
  assign n36492 = n36491 ^ n10385 ^ n2139 ;
  assign n36489 = ( n1791 & ~n6507 ) | ( n1791 & n7652 ) | ( ~n6507 & n7652 ) ;
  assign n36490 = ( n16043 & n35159 ) | ( n16043 & n36489 ) | ( n35159 & n36489 ) ;
  assign n36493 = n36492 ^ n36490 ^ n6797 ;
  assign n36494 = n25658 ^ n17403 ^ 1'b0 ;
  assign n36495 = ( n9852 & n16138 ) | ( n9852 & n34766 ) | ( n16138 & n34766 ) ;
  assign n36496 = ~n1195 & n1505 ;
  assign n36497 = ( n12169 & n14375 ) | ( n12169 & n16914 ) | ( n14375 & n16914 ) ;
  assign n36498 = n36496 & n36497 ;
  assign n36499 = n36498 ^ n10998 ^ 1'b0 ;
  assign n36500 = n36495 | n36499 ;
  assign n36501 = n31760 ^ n25564 ^ n9267 ;
  assign n36502 = n4216 & ~n36501 ;
  assign n36503 = n26488 ^ n5815 ^ 1'b0 ;
  assign n36504 = n36503 ^ n16723 ^ n5052 ;
  assign n36505 = n34459 & n36504 ;
  assign n36506 = n1821 | n3140 ;
  assign n36507 = ( n7680 & n10937 ) | ( n7680 & n12759 ) | ( n10937 & n12759 ) ;
  assign n36508 = n36507 ^ n2102 ^ 1'b0 ;
  assign n36509 = n36506 | n36508 ;
  assign n36510 = n6769 & ~n28299 ;
  assign n36511 = n36510 ^ n10112 ^ 1'b0 ;
  assign n36512 = n22169 ^ n10544 ^ n8663 ;
  assign n36513 = n36511 | n36512 ;
  assign n36514 = ( n3898 & n4104 ) | ( n3898 & ~n5799 ) | ( n4104 & ~n5799 ) ;
  assign n36515 = n36514 ^ n29664 ^ n23557 ;
  assign n36516 = ( n5029 & ~n14167 ) | ( n5029 & n14619 ) | ( ~n14167 & n14619 ) ;
  assign n36517 = n15163 & n24182 ;
  assign n36518 = n20700 ^ n18914 ^ 1'b0 ;
  assign n36519 = n9980 ^ n1551 ^ 1'b0 ;
  assign n36520 = n36518 & ~n36519 ;
  assign n36521 = n35872 & n36520 ;
  assign n36522 = ( n13430 & n14557 ) | ( n13430 & ~n36315 ) | ( n14557 & ~n36315 ) ;
  assign n36524 = n17770 ^ n3233 ^ 1'b0 ;
  assign n36525 = n13173 & n36524 ;
  assign n36526 = n36525 ^ n31339 ^ n6322 ;
  assign n36523 = ~n10150 & n12723 ;
  assign n36527 = n36526 ^ n36523 ^ 1'b0 ;
  assign n36528 = n36527 ^ n24772 ^ 1'b0 ;
  assign n36530 = n3655 & n5741 ;
  assign n36531 = n36530 ^ n3450 ^ 1'b0 ;
  assign n36532 = ~n13980 & n36531 ;
  assign n36533 = n36532 ^ n13824 ^ 1'b0 ;
  assign n36529 = ( ~n10005 & n20728 ) | ( ~n10005 & n31785 ) | ( n20728 & n31785 ) ;
  assign n36534 = n36533 ^ n36529 ^ n36295 ;
  assign n36535 = n11635 | n16118 ;
  assign n36536 = n28403 ^ n7131 ^ 1'b0 ;
  assign n36537 = n13130 ^ n4885 ^ 1'b0 ;
  assign n36538 = ( n4466 & n18870 ) | ( n4466 & n33950 ) | ( n18870 & n33950 ) ;
  assign n36539 = n36538 ^ n36531 ^ n15066 ;
  assign n36540 = n15322 | n36539 ;
  assign n36541 = n9182 & ~n36540 ;
  assign n36542 = n36541 ^ n35321 ^ 1'b0 ;
  assign n36543 = ( n6926 & n26660 ) | ( n6926 & n26869 ) | ( n26660 & n26869 ) ;
  assign n36544 = n36543 ^ n35251 ^ n14195 ;
  assign n36545 = ( ~n2881 & n4362 ) | ( ~n2881 & n12045 ) | ( n4362 & n12045 ) ;
  assign n36546 = ( n6297 & ~n22778 ) | ( n6297 & n36545 ) | ( ~n22778 & n36545 ) ;
  assign n36547 = ( n25602 & ~n36518 ) | ( n25602 & n36546 ) | ( ~n36518 & n36546 ) ;
  assign n36548 = n13519 & ~n19267 ;
  assign n36549 = ( n17018 & n17213 ) | ( n17018 & n35009 ) | ( n17213 & n35009 ) ;
  assign n36550 = ~x63 & n519 ;
  assign n36551 = n824 | n36550 ;
  assign n36552 = n36551 ^ n11916 ^ n6596 ;
  assign n36553 = n36552 ^ n24802 ^ 1'b0 ;
  assign n36554 = n28986 & n36553 ;
  assign n36555 = ~n6381 & n36554 ;
  assign n36556 = n36555 ^ n7186 ^ 1'b0 ;
  assign n36557 = n17574 & ~n19786 ;
  assign n36558 = n24065 & n36557 ;
  assign n36560 = ( ~n4827 & n8024 ) | ( ~n4827 & n10885 ) | ( n8024 & n10885 ) ;
  assign n36559 = n16306 & n30634 ;
  assign n36561 = n36560 ^ n36559 ^ 1'b0 ;
  assign n36562 = n11493 ^ n10393 ^ 1'b0 ;
  assign n36563 = n36561 | n36562 ;
  assign n36564 = n10647 ^ n4777 ^ n3667 ;
  assign n36565 = ( n26417 & n28559 ) | ( n26417 & n36564 ) | ( n28559 & n36564 ) ;
  assign n36566 = n23782 & ~n36565 ;
  assign n36567 = n36563 & n36566 ;
  assign n36569 = ~n22886 & n25541 ;
  assign n36568 = n8188 | n21582 ;
  assign n36570 = n36569 ^ n36568 ^ 1'b0 ;
  assign n36571 = ( ~n2374 & n12983 ) | ( ~n2374 & n24257 ) | ( n12983 & n24257 ) ;
  assign n36572 = ( n3979 & n13202 ) | ( n3979 & ~n36571 ) | ( n13202 & ~n36571 ) ;
  assign n36573 = n32749 ^ n7753 ^ 1'b0 ;
  assign n36574 = n36573 ^ n2200 ^ x89 ;
  assign n36575 = n36574 ^ n6434 ^ 1'b0 ;
  assign n36576 = n36575 ^ n11589 ^ n3458 ;
  assign n36577 = n36576 ^ n14193 ^ 1'b0 ;
  assign n36578 = n4580 & n36577 ;
  assign n36579 = n36578 ^ n21160 ^ n5322 ;
  assign n36581 = n16000 ^ n4492 ^ 1'b0 ;
  assign n36580 = ~n1246 & n8056 ;
  assign n36582 = n36581 ^ n36580 ^ n10960 ;
  assign n36587 = n3254 & ~n7211 ;
  assign n36585 = n10892 | n19822 ;
  assign n36586 = n36585 ^ n21228 ^ 1'b0 ;
  assign n36583 = n13679 & n30763 ;
  assign n36584 = x67 & ~n36583 ;
  assign n36588 = n36587 ^ n36586 ^ n36584 ;
  assign n36589 = n30372 ^ n16742 ^ n15136 ;
  assign n36590 = n3331 & ~n19378 ;
  assign n36591 = ( n7102 & ~n31888 ) | ( n7102 & n36590 ) | ( ~n31888 & n36590 ) ;
  assign n36592 = n1990 & ~n18025 ;
  assign n36593 = ( ~n19782 & n23339 ) | ( ~n19782 & n36592 ) | ( n23339 & n36592 ) ;
  assign n36594 = n723 & n19352 ;
  assign n36595 = n1656 & n12844 ;
  assign n36596 = n36595 ^ n13906 ^ 1'b0 ;
  assign n36597 = n29839 & ~n34719 ;
  assign n36598 = n36597 ^ n26366 ^ 1'b0 ;
  assign n36599 = n26101 ^ n19458 ^ x178 ;
  assign n36600 = n5416 | n13694 ;
  assign n36601 = n6101 & n36600 ;
  assign n36602 = n5853 & ~n13583 ;
  assign n36603 = n36602 ^ n654 ^ 1'b0 ;
  assign n36604 = ( ~n730 & n1682 ) | ( ~n730 & n36603 ) | ( n1682 & n36603 ) ;
  assign n36605 = n36604 ^ n9424 ^ 1'b0 ;
  assign n36606 = n36601 | n36605 ;
  assign n36607 = n36606 ^ n27514 ^ n19053 ;
  assign n36608 = ( n8773 & n10538 ) | ( n8773 & ~n35321 ) | ( n10538 & ~n35321 ) ;
  assign n36609 = ( ~n3659 & n14972 ) | ( ~n3659 & n36608 ) | ( n14972 & n36608 ) ;
  assign n36610 = n19019 | n27812 ;
  assign n36611 = n980 | n36610 ;
  assign n36612 = ( n1458 & n13246 ) | ( n1458 & n22073 ) | ( n13246 & n22073 ) ;
  assign n36613 = n36612 ^ n4913 ^ 1'b0 ;
  assign n36614 = n19811 ^ n10567 ^ 1'b0 ;
  assign n36615 = n36614 ^ n20663 ^ n14075 ;
  assign n36616 = n17105 & ~n36615 ;
  assign n36617 = n36616 ^ n21698 ^ 1'b0 ;
  assign n36618 = n33385 ^ n13718 ^ 1'b0 ;
  assign n36619 = n19820 & ~n36618 ;
  assign n36620 = n23235 & ~n34724 ;
  assign n36621 = ~n36619 & n36620 ;
  assign n36622 = n19106 | n36621 ;
  assign n36623 = n36622 ^ n11379 ^ 1'b0 ;
  assign n36624 = ~n29335 & n32818 ;
  assign n36625 = n11406 & ~n20854 ;
  assign n36626 = ( ~n9662 & n28417 ) | ( ~n9662 & n36625 ) | ( n28417 & n36625 ) ;
  assign n36627 = n3202 | n4564 ;
  assign n36628 = n11484 & ~n36627 ;
  assign n36629 = n36628 ^ n10162 ^ 1'b0 ;
  assign n36630 = n1657 & n18628 ;
  assign n36631 = n22659 ^ n14920 ^ n3368 ;
  assign n36632 = n21572 | n36631 ;
  assign n36633 = n28063 ^ n21531 ^ n5232 ;
  assign n36634 = n36632 & ~n36633 ;
  assign n36635 = n36634 ^ n7399 ^ 1'b0 ;
  assign n36637 = n28336 ^ n22572 ^ 1'b0 ;
  assign n36638 = ( x32 & ~n22663 ) | ( x32 & n36637 ) | ( ~n22663 & n36637 ) ;
  assign n36636 = n13693 | n26236 ;
  assign n36639 = n36638 ^ n36636 ^ 1'b0 ;
  assign n36640 = n8386 & ~n23997 ;
  assign n36641 = n36640 ^ n5378 ^ 1'b0 ;
  assign n36642 = ( n9375 & n9576 ) | ( n9375 & n20706 ) | ( n9576 & n20706 ) ;
  assign n36643 = ( n2145 & ~n23834 ) | ( n2145 & n31866 ) | ( ~n23834 & n31866 ) ;
  assign n36646 = n16480 | n36124 ;
  assign n36647 = n16680 & ~n36646 ;
  assign n36644 = n948 & n23711 ;
  assign n36645 = n36644 ^ n6883 ^ 1'b0 ;
  assign n36648 = n36647 ^ n36645 ^ 1'b0 ;
  assign n36649 = n17331 ^ n6734 ^ n3828 ;
  assign n36650 = n36649 ^ n12729 ^ n4478 ;
  assign n36651 = n5732 & n36650 ;
  assign n36652 = n36651 ^ n14740 ^ 1'b0 ;
  assign n36654 = n19295 ^ n8931 ^ 1'b0 ;
  assign n36653 = n2809 | n6439 ;
  assign n36655 = n36654 ^ n36653 ^ 1'b0 ;
  assign n36656 = ( ~n4430 & n15311 ) | ( ~n4430 & n18008 ) | ( n15311 & n18008 ) ;
  assign n36657 = n36656 ^ n9074 ^ 1'b0 ;
  assign n36658 = ( ~n4676 & n7164 ) | ( ~n4676 & n12619 ) | ( n7164 & n12619 ) ;
  assign n36659 = n20818 ^ n19631 ^ n10969 ;
  assign n36660 = n36659 ^ n843 ^ 1'b0 ;
  assign n36661 = n36658 | n36660 ;
  assign n36662 = n36661 ^ n22943 ^ n6778 ;
  assign n36663 = n26335 ^ n7677 ^ x68 ;
  assign n36664 = n36663 ^ n33757 ^ 1'b0 ;
  assign n36665 = n12080 ^ n7790 ^ n5171 ;
  assign n36666 = n5183 ^ n3290 ^ 1'b0 ;
  assign n36667 = n6744 | n36666 ;
  assign n36668 = n36667 ^ n15057 ^ 1'b0 ;
  assign n36669 = n36665 | n36668 ;
  assign n36670 = n23575 ^ n19725 ^ n1794 ;
  assign n36671 = n8855 ^ n7077 ^ n4268 ;
  assign n36672 = n36671 ^ n17981 ^ 1'b0 ;
  assign n36673 = n36670 & n36672 ;
  assign n36674 = n5321 & n16960 ;
  assign n36675 = ~n23476 & n36674 ;
  assign n36676 = n18402 ^ n3630 ^ 1'b0 ;
  assign n36677 = n32832 & ~n36676 ;
  assign n36678 = n26963 ^ n22687 ^ 1'b0 ;
  assign n36679 = n3771 | n27835 ;
  assign n36680 = n36679 ^ n13112 ^ 1'b0 ;
  assign n36681 = ~n22361 & n36680 ;
  assign n36682 = ( n3849 & n30275 ) | ( n3849 & n35532 ) | ( n30275 & n35532 ) ;
  assign n36683 = n3941 ^ n3828 ^ 1'b0 ;
  assign n36687 = ( n5075 & n6101 ) | ( n5075 & n11810 ) | ( n6101 & n11810 ) ;
  assign n36684 = n25650 ^ n18525 ^ n14215 ;
  assign n36685 = n26534 & ~n36684 ;
  assign n36686 = ~n5617 & n36685 ;
  assign n36688 = n36687 ^ n36686 ^ 1'b0 ;
  assign n36691 = n4281 | n4644 ;
  assign n36689 = n31493 ^ n8926 ^ 1'b0 ;
  assign n36690 = n22254 | n36689 ;
  assign n36692 = n36691 ^ n36690 ^ n25881 ;
  assign n36693 = ( n1573 & n18617 ) | ( n1573 & n27530 ) | ( n18617 & n27530 ) ;
  assign n36694 = n2540 & n36693 ;
  assign n36695 = ( ~n6474 & n17743 ) | ( ~n6474 & n32751 ) | ( n17743 & n32751 ) ;
  assign n36696 = ( n11033 & ~n11659 ) | ( n11033 & n25746 ) | ( ~n11659 & n25746 ) ;
  assign n36697 = n24395 ^ n14522 ^ 1'b0 ;
  assign n36698 = n13816 & n36697 ;
  assign n36699 = ~n11625 & n20399 ;
  assign n36700 = n23412 & n36699 ;
  assign n36701 = n4024 | n36700 ;
  assign n36702 = n2295 & ~n36701 ;
  assign n36703 = n5620 & n9064 ;
  assign n36704 = n3819 | n36703 ;
  assign n36705 = n29394 & ~n36704 ;
  assign n36706 = n18869 ^ n7517 ^ 1'b0 ;
  assign n36707 = ~n13829 & n36706 ;
  assign n36708 = n26073 & ~n27154 ;
  assign n36709 = n36708 ^ n7403 ^ 1'b0 ;
  assign n36710 = ( n4681 & n6709 ) | ( n4681 & n26679 ) | ( n6709 & n26679 ) ;
  assign n36711 = n36710 ^ n30997 ^ n7364 ;
  assign n36712 = n31323 ^ n14826 ^ 1'b0 ;
  assign n36713 = n7216 & n36712 ;
  assign n36714 = n5433 | n36713 ;
  assign n36715 = ( x145 & n982 ) | ( x145 & n36714 ) | ( n982 & n36714 ) ;
  assign n36716 = x155 & ~n5860 ;
  assign n36717 = ( n22355 & n26026 ) | ( n22355 & n36716 ) | ( n26026 & n36716 ) ;
  assign n36718 = n36717 ^ n12145 ^ 1'b0 ;
  assign n36719 = n1193 | n6655 ;
  assign n36720 = n36719 ^ n20893 ^ 1'b0 ;
  assign n36721 = ( n8424 & n30146 ) | ( n8424 & ~n36720 ) | ( n30146 & ~n36720 ) ;
  assign n36723 = n1086 & n2230 ;
  assign n36724 = n11706 & n36723 ;
  assign n36722 = n11000 & ~n19367 ;
  assign n36725 = n36724 ^ n36722 ^ 1'b0 ;
  assign n36726 = n19631 ^ n11708 ^ 1'b0 ;
  assign n36727 = ~n4398 & n14291 ;
  assign n36728 = n36727 ^ n29584 ^ 1'b0 ;
  assign n36729 = n8060 ^ n4997 ^ 1'b0 ;
  assign n36730 = n13111 ^ n9193 ^ 1'b0 ;
  assign n36731 = ( ~n8928 & n36729 ) | ( ~n8928 & n36730 ) | ( n36729 & n36730 ) ;
  assign n36732 = ( n2432 & n23001 ) | ( n2432 & n36731 ) | ( n23001 & n36731 ) ;
  assign n36733 = n13895 ^ n13502 ^ 1'b0 ;
  assign n36734 = n28751 ^ n8580 ^ 1'b0 ;
  assign n36735 = n36733 & ~n36734 ;
  assign n36736 = n13155 & n35320 ;
  assign n36737 = n36736 ^ n34241 ^ 1'b0 ;
  assign n36738 = n36737 ^ n31778 ^ n7611 ;
  assign n36739 = ( n20772 & ~n31033 ) | ( n20772 & n36738 ) | ( ~n31033 & n36738 ) ;
  assign n36740 = n23688 & n33730 ;
  assign n36741 = ~n5354 & n36740 ;
  assign n36742 = n29548 ^ n19588 ^ n18156 ;
  assign n36743 = n30795 ^ n21666 ^ n4560 ;
  assign n36749 = n10491 & n28191 ;
  assign n36744 = n8533 | n27970 ;
  assign n36745 = n36744 ^ n17873 ^ n11011 ;
  assign n36746 = ~n7914 & n36745 ;
  assign n36747 = n36746 ^ n812 ^ x170 ;
  assign n36748 = n36747 ^ n24079 ^ n23358 ;
  assign n36750 = n36749 ^ n36748 ^ n6168 ;
  assign n36751 = n7055 & n9625 ;
  assign n36752 = n36751 ^ n7080 ^ 1'b0 ;
  assign n36753 = n36752 ^ n24441 ^ n11114 ;
  assign n36754 = ( n10287 & n11810 ) | ( n10287 & n14767 ) | ( n11810 & n14767 ) ;
  assign n36755 = ( n32861 & n36753 ) | ( n32861 & ~n36754 ) | ( n36753 & ~n36754 ) ;
  assign n36756 = ~n2804 & n5204 ;
  assign n36757 = ~n11678 & n15833 ;
  assign n36758 = ~n36756 & n36757 ;
  assign n36759 = n16639 ^ n7146 ^ n1872 ;
  assign n36760 = ( n3765 & n9298 ) | ( n3765 & n36759 ) | ( n9298 & n36759 ) ;
  assign n36761 = n20773 | n36760 ;
  assign n36762 = n36758 & ~n36761 ;
  assign n36763 = n20646 | n36762 ;
  assign n36764 = n16245 & ~n36763 ;
  assign n36765 = n10778 ^ n6424 ^ 1'b0 ;
  assign n36766 = n10659 | n27180 ;
  assign n36767 = n8178 & ~n36766 ;
  assign n36768 = n9621 ^ n1971 ^ 1'b0 ;
  assign n36769 = n23164 & n36768 ;
  assign n36770 = ( n5747 & n18217 ) | ( n5747 & ~n21917 ) | ( n18217 & ~n21917 ) ;
  assign n36771 = ~n2799 & n19949 ;
  assign n36772 = n36771 ^ n18014 ^ 1'b0 ;
  assign n36773 = n36772 ^ n17444 ^ n13529 ;
  assign n36774 = n36440 ^ n3436 ^ 1'b0 ;
  assign n36775 = ~n27477 & n36774 ;
  assign n36777 = ( n7395 & n12418 ) | ( n7395 & n21340 ) | ( n12418 & n21340 ) ;
  assign n36776 = n554 & n5568 ;
  assign n36778 = n36777 ^ n36776 ^ 1'b0 ;
  assign n36779 = n36342 ^ n7258 ^ n3388 ;
  assign n36780 = n17716 ^ n7279 ^ 1'b0 ;
  assign n36781 = n18624 | n36780 ;
  assign n36782 = n36779 & n36781 ;
  assign n36783 = n36396 ^ n25484 ^ n16725 ;
  assign n36784 = n29904 | n36783 ;
  assign n36785 = n36784 ^ n32638 ^ n23642 ;
  assign n36791 = n5981 & n20213 ;
  assign n36792 = ~n5913 & n36791 ;
  assign n36786 = n2131 & ~n29378 ;
  assign n36787 = n36786 ^ n12921 ^ 1'b0 ;
  assign n36788 = n36787 ^ n9738 ^ n3839 ;
  assign n36789 = ~x48 & n36788 ;
  assign n36790 = n36789 ^ n33510 ^ n7093 ;
  assign n36793 = n36792 ^ n36790 ^ n27715 ;
  assign n36795 = n12607 ^ n3450 ^ n1830 ;
  assign n36794 = n2904 & ~n17713 ;
  assign n36796 = n36795 ^ n36794 ^ 1'b0 ;
  assign n36797 = ( n751 & n6114 ) | ( n751 & n23882 ) | ( n6114 & n23882 ) ;
  assign n36798 = n13838 | n24166 ;
  assign n36799 = n36797 | n36798 ;
  assign n36800 = n23951 & ~n36525 ;
  assign n36801 = ~n933 & n4555 ;
  assign n36802 = n35112 & n36801 ;
  assign n36803 = n36802 ^ n3087 ^ 1'b0 ;
  assign n36804 = n7313 & n36803 ;
  assign n36805 = ~n17673 & n27389 ;
  assign n36806 = n4641 | n36805 ;
  assign n36810 = n34272 ^ n1896 ^ n1091 ;
  assign n36807 = ( n2569 & ~n7541 ) | ( n2569 & n19715 ) | ( ~n7541 & n19715 ) ;
  assign n36808 = ( n20291 & n27610 ) | ( n20291 & n28087 ) | ( n27610 & n28087 ) ;
  assign n36809 = ( n19481 & ~n36807 ) | ( n19481 & n36808 ) | ( ~n36807 & n36808 ) ;
  assign n36811 = n36810 ^ n36809 ^ n4929 ;
  assign n36812 = ~n24449 & n33883 ;
  assign n36813 = n1241 & ~n19800 ;
  assign n36814 = ( n1618 & ~n10052 ) | ( n1618 & n21075 ) | ( ~n10052 & n21075 ) ;
  assign n36815 = ~n28721 & n36814 ;
  assign n36816 = n36815 ^ n19576 ^ 1'b0 ;
  assign n36817 = n2936 & ~n4223 ;
  assign n36818 = n5750 & n36817 ;
  assign n36819 = ( n2659 & n12321 ) | ( n2659 & ~n36818 ) | ( n12321 & ~n36818 ) ;
  assign n36820 = n36819 ^ n26707 ^ n5968 ;
  assign n36825 = n19812 | n24342 ;
  assign n36821 = n32565 ^ n11485 ^ n4100 ;
  assign n36822 = n20739 & n36821 ;
  assign n36823 = n2364 & n36822 ;
  assign n36824 = ( ~n17288 & n24793 ) | ( ~n17288 & n36823 ) | ( n24793 & n36823 ) ;
  assign n36826 = n36825 ^ n36824 ^ n6930 ;
  assign n36829 = ( n5177 & n11598 ) | ( n5177 & ~n18916 ) | ( n11598 & ~n18916 ) ;
  assign n36827 = ~n26965 & n32496 ;
  assign n36828 = ~n29743 & n36827 ;
  assign n36830 = n36829 ^ n36828 ^ 1'b0 ;
  assign n36831 = n15908 ^ n8051 ^ n6734 ;
  assign n36832 = x5 & n36831 ;
  assign n36833 = ( n34279 & ~n35234 ) | ( n34279 & n36832 ) | ( ~n35234 & n36832 ) ;
  assign n36834 = ~n11205 & n13166 ;
  assign n36835 = n582 & n36834 ;
  assign n36836 = n36835 ^ n17319 ^ n5512 ;
  assign n36837 = n2261 | n36836 ;
  assign n36838 = n12769 ^ n7868 ^ 1'b0 ;
  assign n36839 = n13292 & n36838 ;
  assign n36840 = n12686 & ~n36839 ;
  assign n36841 = n36840 ^ n34702 ^ n6406 ;
  assign n36842 = ~n13824 & n15526 ;
  assign n36843 = n2246 | n22687 ;
  assign n36844 = n36843 ^ n12804 ^ 1'b0 ;
  assign n36845 = n36844 ^ n21843 ^ 1'b0 ;
  assign n36846 = n29557 & ~n36845 ;
  assign n36848 = n32069 ^ n16109 ^ n8734 ;
  assign n36847 = ( n2149 & n24402 ) | ( n2149 & ~n27904 ) | ( n24402 & ~n27904 ) ;
  assign n36849 = n36848 ^ n36847 ^ n31474 ;
  assign n36850 = ( n16962 & ~n36846 ) | ( n16962 & n36849 ) | ( ~n36846 & n36849 ) ;
  assign n36851 = ( n9010 & n13114 ) | ( n9010 & n18993 ) | ( n13114 & n18993 ) ;
  assign n36852 = n36851 ^ n35829 ^ n1408 ;
  assign n36853 = n9599 ^ n4634 ^ n3573 ;
  assign n36854 = ( ~n10881 & n12860 ) | ( ~n10881 & n36853 ) | ( n12860 & n36853 ) ;
  assign n36855 = ~n29746 & n31633 ;
  assign n36856 = ( ~n8472 & n36854 ) | ( ~n8472 & n36855 ) | ( n36854 & n36855 ) ;
  assign n36857 = n16538 ^ n10571 ^ n3257 ;
  assign n36858 = n21325 & ~n36857 ;
  assign n36859 = n2315 | n12286 ;
  assign n36860 = n36859 ^ n1088 ^ 1'b0 ;
  assign n36861 = ( ~n6197 & n7677 ) | ( ~n6197 & n8799 ) | ( n7677 & n8799 ) ;
  assign n36862 = ~n36860 & n36861 ;
  assign n36863 = n36862 ^ n1489 ^ 1'b0 ;
  assign n36864 = ~n2824 & n6181 ;
  assign n36865 = ~n7110 & n36864 ;
  assign n36866 = n30564 ^ n2265 ^ n337 ;
  assign n36867 = ( ~n8191 & n16601 ) | ( ~n8191 & n36866 ) | ( n16601 & n36866 ) ;
  assign n36868 = n28416 ^ n21799 ^ n7902 ;
  assign n36869 = ~n26933 & n36868 ;
  assign n36870 = n8274 & n36869 ;
  assign n36871 = n36867 | n36870 ;
  assign n36872 = n11001 | n20315 ;
  assign n36873 = ( n20106 & ~n34635 ) | ( n20106 & n36872 ) | ( ~n34635 & n36872 ) ;
  assign n36874 = ~n4990 & n18345 ;
  assign n36875 = n34258 ^ n20454 ^ 1'b0 ;
  assign n36876 = n14139 | n20008 ;
  assign n36877 = n36876 ^ n1322 ^ 1'b0 ;
  assign n36878 = n17396 & n36877 ;
  assign n36879 = n15692 & n36878 ;
  assign n36882 = n12570 ^ n10846 ^ n502 ;
  assign n36880 = n11441 & ~n13396 ;
  assign n36881 = ( n3954 & n10627 ) | ( n3954 & n36880 ) | ( n10627 & n36880 ) ;
  assign n36883 = n36882 ^ n36881 ^ 1'b0 ;
  assign n36884 = n4139 & ~n31043 ;
  assign n36885 = ~n9548 & n36884 ;
  assign n36888 = n6027 & n11755 ;
  assign n36889 = n36888 ^ n21258 ^ 1'b0 ;
  assign n36886 = n34786 ^ n34237 ^ 1'b0 ;
  assign n36887 = ( n8276 & n36587 ) | ( n8276 & n36886 ) | ( n36587 & n36886 ) ;
  assign n36890 = n36889 ^ n36887 ^ 1'b0 ;
  assign n36891 = n12751 & ~n36890 ;
  assign n36892 = n34417 ^ n13010 ^ 1'b0 ;
  assign n36893 = n23403 ^ n10267 ^ 1'b0 ;
  assign n36894 = n3587 | n36893 ;
  assign n36895 = n7313 & n29214 ;
  assign n36896 = n36895 ^ n16526 ^ 1'b0 ;
  assign n36897 = ( ~n4651 & n16570 ) | ( ~n4651 & n36896 ) | ( n16570 & n36896 ) ;
  assign n36898 = ( ~n27169 & n36894 ) | ( ~n27169 & n36897 ) | ( n36894 & n36897 ) ;
  assign n36899 = n27214 ^ n25612 ^ n8267 ;
  assign n36900 = n16435 ^ n1966 ^ x108 ;
  assign n36901 = n17110 ^ n16478 ^ 1'b0 ;
  assign n36902 = n17795 & ~n36901 ;
  assign n36903 = ( ~n26493 & n36900 ) | ( ~n26493 & n36902 ) | ( n36900 & n36902 ) ;
  assign n36904 = x62 & n25250 ;
  assign n36905 = n12916 & n36904 ;
  assign n36906 = n36905 ^ n9167 ^ n6735 ;
  assign n36907 = n36906 ^ n24674 ^ 1'b0 ;
  assign n36908 = n11232 | n36907 ;
  assign n36909 = ~n13212 & n24627 ;
  assign n36910 = n5569 & n9179 ;
  assign n36911 = n36910 ^ n22366 ^ n6780 ;
  assign n36912 = n30809 ^ n21330 ^ n6450 ;
  assign n36913 = n7120 ^ n6849 ^ 1'b0 ;
  assign n36914 = n22218 ^ n16580 ^ 1'b0 ;
  assign n36917 = n29317 ^ n2569 ^ 1'b0 ;
  assign n36918 = n15821 & n36917 ;
  assign n36915 = n24514 ^ n5305 ^ n4034 ;
  assign n36916 = n36915 ^ n31124 ^ 1'b0 ;
  assign n36919 = n36918 ^ n36916 ^ 1'b0 ;
  assign n36920 = ~n36914 & n36919 ;
  assign n36921 = n5778 ^ n1710 ^ 1'b0 ;
  assign n36922 = n2716 & ~n3543 ;
  assign n36923 = n30861 & n36922 ;
  assign n36924 = n36143 ^ n15603 ^ n12475 ;
  assign n36925 = n23559 ^ n15316 ^ n10177 ;
  assign n36928 = n11178 | n25514 ;
  assign n36926 = ( n3186 & n3623 ) | ( n3186 & ~n11218 ) | ( n3623 & ~n11218 ) ;
  assign n36927 = n22087 | n36926 ;
  assign n36929 = n36928 ^ n36927 ^ n8637 ;
  assign n36930 = ( ~n11507 & n22732 ) | ( ~n11507 & n25818 ) | ( n22732 & n25818 ) ;
  assign n36931 = ( x24 & n5723 ) | ( x24 & n15859 ) | ( n5723 & n15859 ) ;
  assign n36932 = n36931 ^ n33143 ^ 1'b0 ;
  assign n36933 = ~n1091 & n19376 ;
  assign n36934 = n13183 & n36933 ;
  assign n36935 = n36934 ^ n26926 ^ 1'b0 ;
  assign n36936 = n16578 & n36935 ;
  assign n36937 = ( n8726 & n9063 ) | ( n8726 & n26848 ) | ( n9063 & n26848 ) ;
  assign n36938 = ~n1153 & n16137 ;
  assign n36939 = ( n15831 & ~n21160 ) | ( n15831 & n29897 ) | ( ~n21160 & n29897 ) ;
  assign n36940 = n20056 ^ n19898 ^ 1'b0 ;
  assign n36941 = n16478 & n36940 ;
  assign n36942 = n32409 ^ n9949 ^ 1'b0 ;
  assign n36943 = n36942 ^ n36137 ^ n22050 ;
  assign n36944 = n17513 ^ x72 ^ 1'b0 ;
  assign n36945 = n36943 & n36944 ;
  assign n36946 = ( n3808 & ~n11517 ) | ( n3808 & n12275 ) | ( ~n11517 & n12275 ) ;
  assign n36947 = n36946 ^ n11375 ^ n10813 ;
  assign n36948 = n29378 ^ n18865 ^ n2770 ;
  assign n36949 = ( n2467 & n36947 ) | ( n2467 & ~n36948 ) | ( n36947 & ~n36948 ) ;
  assign n36950 = n36949 ^ n29957 ^ 1'b0 ;
  assign n36951 = n3722 ^ n3527 ^ n2790 ;
  assign n36952 = n19157 ^ n11634 ^ n10946 ;
  assign n36953 = n9017 ^ n3568 ^ 1'b0 ;
  assign n36954 = ( n36951 & ~n36952 ) | ( n36951 & n36953 ) | ( ~n36952 & n36953 ) ;
  assign n36955 = n1010 & n15434 ;
  assign n36956 = n7772 ^ n2924 ^ 1'b0 ;
  assign n36957 = ~n1682 & n36956 ;
  assign n36958 = ~n4990 & n36957 ;
  assign n36959 = ~n36955 & n36958 ;
  assign n36960 = n14266 & n22111 ;
  assign n36961 = ( n2471 & ~n5616 ) | ( n2471 & n21850 ) | ( ~n5616 & n21850 ) ;
  assign n36962 = n16557 | n36961 ;
  assign n36963 = n36960 & ~n36962 ;
  assign n36964 = n8304 ^ n558 ^ 1'b0 ;
  assign n36965 = ~n9885 & n36964 ;
  assign n36966 = n4975 & ~n11525 ;
  assign n36967 = n36966 ^ n16060 ^ 1'b0 ;
  assign n36968 = ( ~n3364 & n12549 ) | ( ~n3364 & n36967 ) | ( n12549 & n36967 ) ;
  assign n36969 = ( n4376 & ~n25537 ) | ( n4376 & n36968 ) | ( ~n25537 & n36968 ) ;
  assign n36970 = n20047 ^ n16141 ^ n10363 ;
  assign n36971 = ( ~n17463 & n32542 ) | ( ~n17463 & n36970 ) | ( n32542 & n36970 ) ;
  assign n36972 = n31152 ^ n10423 ^ 1'b0 ;
  assign n36973 = ( n29041 & ~n30553 ) | ( n29041 & n36972 ) | ( ~n30553 & n36972 ) ;
  assign n36974 = ~n1549 & n10223 ;
  assign n36975 = ~n14013 & n36974 ;
  assign n36976 = ( ~n3580 & n34659 ) | ( ~n3580 & n36975 ) | ( n34659 & n36975 ) ;
  assign n36977 = n36976 ^ n30111 ^ n19056 ;
  assign n36978 = n12770 & n16691 ;
  assign n36979 = n3807 & n36978 ;
  assign n36980 = n36979 ^ n31307 ^ 1'b0 ;
  assign n36981 = n16300 ^ n15735 ^ 1'b0 ;
  assign n36982 = n34197 & ~n36981 ;
  assign n36983 = n36982 ^ n14778 ^ n14523 ;
  assign n36984 = n13703 | n36983 ;
  assign n36985 = ( n963 & ~n17547 ) | ( n963 & n20240 ) | ( ~n17547 & n20240 ) ;
  assign n36987 = n4391 & n5433 ;
  assign n36988 = n11632 & n36987 ;
  assign n36986 = ( ~n12772 & n18350 ) | ( ~n12772 & n21340 ) | ( n18350 & n21340 ) ;
  assign n36989 = n36988 ^ n36986 ^ n11848 ;
  assign n36990 = ( n6209 & n11458 ) | ( n6209 & ~n12097 ) | ( n11458 & ~n12097 ) ;
  assign n36991 = ( n12783 & ~n17374 ) | ( n12783 & n36990 ) | ( ~n17374 & n36990 ) ;
  assign n36992 = n17777 & ~n36991 ;
  assign n36993 = ~n14106 & n36992 ;
  assign n36994 = n23930 & ~n36993 ;
  assign n36995 = n36994 ^ n12455 ^ 1'b0 ;
  assign n36996 = n22424 ^ n22119 ^ n1177 ;
  assign n36997 = ( n9212 & n23886 ) | ( n9212 & ~n26402 ) | ( n23886 & ~n26402 ) ;
  assign n36998 = n29444 ^ n15864 ^ n358 ;
  assign n36999 = n5348 & ~n36998 ;
  assign n37000 = n15316 ^ n15079 ^ 1'b0 ;
  assign n37001 = ~n17973 & n20695 ;
  assign n37002 = n5731 & ~n7073 ;
  assign n37003 = n37002 ^ n30022 ^ 1'b0 ;
  assign n37004 = n31170 ^ n11264 ^ 1'b0 ;
  assign n37005 = n10330 ^ n513 ^ 1'b0 ;
  assign n37006 = n9482 & n37005 ;
  assign n37007 = ( n7576 & ~n11240 ) | ( n7576 & n37006 ) | ( ~n11240 & n37006 ) ;
  assign n37008 = n29858 | n37007 ;
  assign n37009 = ~n37004 & n37008 ;
  assign n37010 = n2816 | n37009 ;
  assign n37011 = x47 | n37010 ;
  assign n37012 = ( n5714 & n7178 ) | ( n5714 & n13909 ) | ( n7178 & n13909 ) ;
  assign n37013 = n33344 ^ n20685 ^ n5981 ;
  assign n37014 = n12618 | n37013 ;
  assign n37015 = n37012 & ~n37014 ;
  assign n37016 = n7300 | n19894 ;
  assign n37017 = n30569 ^ n2539 ^ 1'b0 ;
  assign n37018 = n9740 & n37017 ;
  assign n37019 = ( n14698 & ~n26251 ) | ( n14698 & n37018 ) | ( ~n26251 & n37018 ) ;
  assign n37020 = ( n758 & ~n1131 ) | ( n758 & n24520 ) | ( ~n1131 & n24520 ) ;
  assign n37021 = n6193 ^ n5573 ^ n1587 ;
  assign n37022 = n3999 & ~n37021 ;
  assign n37023 = n37022 ^ n15825 ^ n657 ;
  assign n37024 = ( ~n2247 & n6947 ) | ( ~n2247 & n24407 ) | ( n6947 & n24407 ) ;
  assign n37025 = n37024 ^ n6312 ^ 1'b0 ;
  assign n37026 = n12679 & ~n37025 ;
  assign n37027 = n35326 ^ n10844 ^ n7907 ;
  assign n37028 = ~n16338 & n25233 ;
  assign n37029 = ~n37027 & n37028 ;
  assign n37030 = n18344 | n22196 ;
  assign n37031 = n25028 & ~n37030 ;
  assign n37032 = ( n498 & ~n3717 ) | ( n498 & n18563 ) | ( ~n3717 & n18563 ) ;
  assign n37033 = ( ~n5064 & n21753 ) | ( ~n5064 & n37032 ) | ( n21753 & n37032 ) ;
  assign n37034 = ( n2489 & n12253 ) | ( n2489 & n24169 ) | ( n12253 & n24169 ) ;
  assign n37035 = ( n10844 & ~n17511 ) | ( n10844 & n20610 ) | ( ~n17511 & n20610 ) ;
  assign n37036 = n36821 ^ n9146 ^ 1'b0 ;
  assign n37037 = n37035 & ~n37036 ;
  assign n37038 = ( n14685 & n37034 ) | ( n14685 & ~n37037 ) | ( n37034 & ~n37037 ) ;
  assign n37039 = n8272 ^ n1136 ^ n793 ;
  assign n37040 = ( n11728 & n12422 ) | ( n11728 & ~n37039 ) | ( n12422 & ~n37039 ) ;
  assign n37041 = n23422 & ~n34177 ;
  assign n37042 = n37040 & ~n37041 ;
  assign n37043 = n37042 ^ n29280 ^ 1'b0 ;
  assign n37044 = n19053 | n37043 ;
  assign n37045 = n22495 | n37044 ;
  assign n37046 = n11592 ^ n7842 ^ 1'b0 ;
  assign n37047 = n13694 | n37046 ;
  assign n37048 = n23549 ^ n14499 ^ 1'b0 ;
  assign n37049 = n4358 | n35316 ;
  assign n37050 = n34553 | n37049 ;
  assign n37051 = n37050 ^ n18544 ^ n2461 ;
  assign n37052 = n37051 ^ n12493 ^ 1'b0 ;
  assign n37053 = ~n37048 & n37052 ;
  assign n37054 = n2651 | n30395 ;
  assign n37055 = n37054 ^ n25336 ^ n5218 ;
  assign n37056 = n34266 ^ n20423 ^ 1'b0 ;
  assign n37057 = ( ~n772 & n11215 ) | ( ~n772 & n14632 ) | ( n11215 & n14632 ) ;
  assign n37058 = ( n18436 & ~n36234 ) | ( n18436 & n37057 ) | ( ~n36234 & n37057 ) ;
  assign n37059 = n6388 | n12674 ;
  assign n37060 = n35258 | n37059 ;
  assign n37061 = n37060 ^ n30941 ^ n29729 ;
  assign n37062 = ( n3787 & n16179 ) | ( n3787 & n35829 ) | ( n16179 & n35829 ) ;
  assign n37063 = n26695 | n37062 ;
  assign n37064 = n2376 & n10886 ;
  assign n37065 = n1638 & n17278 ;
  assign n37066 = n37065 ^ n10897 ^ 1'b0 ;
  assign n37067 = n595 & ~n32425 ;
  assign n37068 = n37067 ^ n31589 ^ 1'b0 ;
  assign n37069 = n37066 & n37068 ;
  assign n37070 = n33163 ^ n24413 ^ 1'b0 ;
  assign n37071 = ~n8677 & n24273 ;
  assign n37072 = n37071 ^ n23863 ^ 1'b0 ;
  assign n37073 = n22720 | n23104 ;
  assign n37074 = n20143 ^ n11137 ^ 1'b0 ;
  assign n37075 = n37074 ^ n26484 ^ 1'b0 ;
  assign n37076 = n8539 & ~n9505 ;
  assign n37077 = ~n5715 & n9482 ;
  assign n37078 = n37077 ^ n15395 ^ 1'b0 ;
  assign n37079 = ( ~n7346 & n25630 ) | ( ~n7346 & n37078 ) | ( n25630 & n37078 ) ;
  assign n37080 = n14516 ^ n13728 ^ 1'b0 ;
  assign n37081 = n23503 & n37080 ;
  assign n37082 = ( n24901 & ~n37079 ) | ( n24901 & n37081 ) | ( ~n37079 & n37081 ) ;
  assign n37083 = ( n4329 & ~n21279 ) | ( n4329 & n25667 ) | ( ~n21279 & n25667 ) ;
  assign n37084 = n21263 & ~n37083 ;
  assign n37085 = n18807 & ~n27084 ;
  assign n37086 = ~n12063 & n37085 ;
  assign n37087 = n15359 & n28720 ;
  assign n37088 = n37087 ^ n10249 ^ 1'b0 ;
  assign n37093 = ( ~n10765 & n11190 ) | ( ~n10765 & n14410 ) | ( n11190 & n14410 ) ;
  assign n37089 = n11821 | n18747 ;
  assign n37090 = ( n4219 & n5264 ) | ( n4219 & n28927 ) | ( n5264 & n28927 ) ;
  assign n37091 = n25149 & ~n37090 ;
  assign n37092 = n37089 & n37091 ;
  assign n37094 = n37093 ^ n37092 ^ n13611 ;
  assign n37095 = ( n3787 & ~n4384 ) | ( n3787 & n12032 ) | ( ~n4384 & n12032 ) ;
  assign n37096 = n5587 | n8216 ;
  assign n37097 = n5904 & ~n37096 ;
  assign n37098 = ( n26378 & n37095 ) | ( n26378 & ~n37097 ) | ( n37095 & ~n37097 ) ;
  assign n37099 = n16015 ^ n1427 ^ 1'b0 ;
  assign n37100 = ( n7385 & ~n17181 ) | ( n7385 & n29987 ) | ( ~n17181 & n29987 ) ;
  assign n37101 = ~n5281 & n30214 ;
  assign n37102 = n17780 & n37101 ;
  assign n37103 = n16593 & ~n36165 ;
  assign n37104 = ( n2111 & n4337 ) | ( n2111 & ~n37103 ) | ( n4337 & ~n37103 ) ;
  assign n37105 = n37104 ^ n33062 ^ n23087 ;
  assign n37106 = n13499 | n18033 ;
  assign n37108 = n5869 & n7211 ;
  assign n37107 = n15498 ^ n14195 ^ n5363 ;
  assign n37109 = n37108 ^ n37107 ^ n6899 ;
  assign n37110 = n37104 ^ n1897 ^ 1'b0 ;
  assign n37111 = ~n2580 & n37110 ;
  assign n37112 = ~n22795 & n34232 ;
  assign n37113 = ( n2215 & n6784 ) | ( n2215 & n18174 ) | ( n6784 & n18174 ) ;
  assign n37114 = n37113 ^ n25686 ^ n1195 ;
  assign n37115 = ( n2425 & n5227 ) | ( n2425 & ~n12415 ) | ( n5227 & ~n12415 ) ;
  assign n37116 = ( n3689 & n4826 ) | ( n3689 & n37115 ) | ( n4826 & n37115 ) ;
  assign n37117 = ( n3547 & n29634 ) | ( n3547 & n33566 ) | ( n29634 & n33566 ) ;
  assign n37118 = n23906 ^ n10921 ^ n4412 ;
  assign n37119 = n11329 & n37118 ;
  assign n37120 = n23895 & n37119 ;
  assign n37121 = n25524 ^ n19187 ^ 1'b0 ;
  assign n37122 = ~n7901 & n24517 ;
  assign n37126 = n11774 ^ n9009 ^ 1'b0 ;
  assign n37127 = n24003 & n37126 ;
  assign n37128 = n37127 ^ n16844 ^ n7075 ;
  assign n37123 = n2681 & n5769 ;
  assign n37124 = ( ~n23549 & n30474 ) | ( ~n23549 & n37123 ) | ( n30474 & n37123 ) ;
  assign n37125 = n2317 & n37124 ;
  assign n37129 = n37128 ^ n37125 ^ 1'b0 ;
  assign n37130 = ~n5043 & n9305 ;
  assign n37131 = n5142 & n37130 ;
  assign n37132 = n37131 ^ n17463 ^ n8787 ;
  assign n37133 = ~n14102 & n37132 ;
  assign n37134 = ( x246 & ~n8968 ) | ( x246 & n33945 ) | ( ~n8968 & n33945 ) ;
  assign n37135 = ( n5370 & ~n18312 ) | ( n5370 & n37134 ) | ( ~n18312 & n37134 ) ;
  assign n37137 = n13127 | n16635 ;
  assign n37136 = n29088 ^ n3701 ^ n773 ;
  assign n37138 = n37137 ^ n37136 ^ n19183 ;
  assign n37142 = ( n5365 & ~n15971 ) | ( n5365 & n16051 ) | ( ~n15971 & n16051 ) ;
  assign n37139 = n19142 ^ n10155 ^ n3811 ;
  assign n37140 = n30384 & ~n37139 ;
  assign n37141 = ~n18376 & n37140 ;
  assign n37143 = n37142 ^ n37141 ^ n4237 ;
  assign n37144 = n22863 ^ n8955 ^ n7186 ;
  assign n37145 = n28354 & ~n37144 ;
  assign n37146 = n37145 ^ n34959 ^ 1'b0 ;
  assign n37147 = ~n2980 & n17274 ;
  assign n37148 = ~n2690 & n37147 ;
  assign n37149 = n28278 ^ n4755 ^ 1'b0 ;
  assign n37150 = n32981 & ~n37149 ;
  assign n37151 = ( n11588 & n24965 ) | ( n11588 & n37150 ) | ( n24965 & n37150 ) ;
  assign n37152 = ( ~n695 & n13850 ) | ( ~n695 & n15958 ) | ( n13850 & n15958 ) ;
  assign n37153 = ( n11084 & ~n16105 ) | ( n11084 & n37152 ) | ( ~n16105 & n37152 ) ;
  assign n37155 = n8035 | n13360 ;
  assign n37154 = n23650 ^ n21074 ^ 1'b0 ;
  assign n37156 = n37155 ^ n37154 ^ n30421 ;
  assign n37157 = n8112 | n26673 ;
  assign n37166 = n8596 ^ n3645 ^ 1'b0 ;
  assign n37167 = n27234 & n37166 ;
  assign n37160 = n21470 ^ n4769 ^ 1'b0 ;
  assign n37161 = n6873 | n37160 ;
  assign n37162 = n7783 & n25674 ;
  assign n37163 = n37161 & n37162 ;
  assign n37158 = n20419 ^ n10344 ^ 1'b0 ;
  assign n37159 = ~n6973 & n37158 ;
  assign n37164 = n37163 ^ n37159 ^ n20476 ;
  assign n37165 = n14300 & n37164 ;
  assign n37168 = n37167 ^ n37165 ^ 1'b0 ;
  assign n37169 = n11413 & ~n37168 ;
  assign n37170 = n8567 & n37169 ;
  assign n37171 = n11477 & ~n14724 ;
  assign n37172 = ( n586 & ~n10139 ) | ( n586 & n37171 ) | ( ~n10139 & n37171 ) ;
  assign n37173 = ( ~n443 & n17147 ) | ( ~n443 & n37172 ) | ( n17147 & n37172 ) ;
  assign n37174 = n37173 ^ n35175 ^ 1'b0 ;
  assign n37175 = n497 & n33653 ;
  assign n37176 = n37175 ^ n27904 ^ 1'b0 ;
  assign n37177 = n31331 & n37176 ;
  assign n37178 = n37174 & n37177 ;
  assign n37179 = n21526 & n27324 ;
  assign n37180 = ( n2049 & n11558 ) | ( n2049 & n35392 ) | ( n11558 & n35392 ) ;
  assign n37181 = n24953 ^ n13249 ^ 1'b0 ;
  assign n37182 = n34932 ^ n14677 ^ n9643 ;
  assign n37183 = ( n4043 & n37181 ) | ( n4043 & n37182 ) | ( n37181 & n37182 ) ;
  assign n37184 = n6074 ^ n5752 ^ 1'b0 ;
  assign n37185 = n18981 & ~n37184 ;
  assign n37186 = ( ~n9740 & n11730 ) | ( ~n9740 & n21353 ) | ( n11730 & n21353 ) ;
  assign n37187 = n4585 & n36489 ;
  assign n37188 = n37186 & n37187 ;
  assign n37189 = ( n5145 & n9840 ) | ( n5145 & ~n30930 ) | ( n9840 & ~n30930 ) ;
  assign n37195 = n16469 & n21544 ;
  assign n37196 = ~n12700 & n37195 ;
  assign n37190 = n8297 | n11040 ;
  assign n37191 = n37190 ^ n11967 ^ 1'b0 ;
  assign n37192 = n16176 ^ n12653 ^ n6219 ;
  assign n37193 = n37192 ^ n34130 ^ n24012 ;
  assign n37194 = ~n37191 & n37193 ;
  assign n37197 = n37196 ^ n37194 ^ n18882 ;
  assign n37198 = n21615 ^ n7309 ^ 1'b0 ;
  assign n37199 = n37198 ^ n29743 ^ n15910 ;
  assign n37200 = ~n447 & n9622 ;
  assign n37201 = n37200 ^ n1545 ^ 1'b0 ;
  assign n37202 = ~n2956 & n37201 ;
  assign n37203 = ~n26093 & n28957 ;
  assign n37204 = n37203 ^ n3342 ^ 1'b0 ;
  assign n37205 = n17461 & ~n24506 ;
  assign n37206 = n37205 ^ n10843 ^ 1'b0 ;
  assign n37207 = n7663 & ~n10488 ;
  assign n37208 = n7160 & n37207 ;
  assign n37209 = n14581 ^ n10236 ^ 1'b0 ;
  assign n37210 = n18157 | n37209 ;
  assign n37211 = n25978 & n37210 ;
  assign n37212 = n12522 & n16367 ;
  assign n37213 = n8507 & n37212 ;
  assign n37214 = ( n37208 & ~n37211 ) | ( n37208 & n37213 ) | ( ~n37211 & n37213 ) ;
  assign n37215 = ( n11068 & n31896 ) | ( n11068 & n32771 ) | ( n31896 & n32771 ) ;
  assign n37216 = n30121 ^ n29781 ^ 1'b0 ;
  assign n37217 = n9730 ^ n8550 ^ n317 ;
  assign n37218 = n20742 & n37217 ;
  assign n37219 = n37218 ^ n1666 ^ 1'b0 ;
  assign n37220 = n12916 ^ n7180 ^ n1319 ;
  assign n37221 = ( n17369 & ~n37219 ) | ( n17369 & n37220 ) | ( ~n37219 & n37220 ) ;
  assign n37222 = ( n6691 & ~n13586 ) | ( n6691 & n33387 ) | ( ~n13586 & n33387 ) ;
  assign n37223 = ( n1690 & n6659 ) | ( n1690 & ~n24855 ) | ( n6659 & ~n24855 ) ;
  assign n37224 = n37222 & ~n37223 ;
  assign n37225 = n37224 ^ n11514 ^ 1'b0 ;
  assign n37226 = n23816 ^ n5245 ^ 1'b0 ;
  assign n37227 = n23440 ^ n22903 ^ n5867 ;
  assign n37228 = ~n33402 & n37227 ;
  assign n37229 = n18279 ^ n11057 ^ n3584 ;
  assign n37230 = n37229 ^ n8922 ^ n3446 ;
  assign n37231 = ~n690 & n15467 ;
  assign n37232 = n17594 & ~n30182 ;
  assign n37233 = n24026 & n37232 ;
  assign n37234 = ~n1448 & n23620 ;
  assign n37235 = n35346 & n37234 ;
  assign n37236 = ( n1790 & ~n37233 ) | ( n1790 & n37235 ) | ( ~n37233 & n37235 ) ;
  assign n37238 = ( n4421 & n6652 ) | ( n4421 & n23034 ) | ( n6652 & n23034 ) ;
  assign n37237 = n3736 & n5645 ;
  assign n37239 = n37238 ^ n37237 ^ n33715 ;
  assign n37240 = ( n19725 & n27862 ) | ( n19725 & ~n37239 ) | ( n27862 & ~n37239 ) ;
  assign n37241 = ( n21843 & n31393 ) | ( n21843 & n32018 ) | ( n31393 & n32018 ) ;
  assign n37242 = n13847 & n24085 ;
  assign n37244 = ( n3216 & n12608 ) | ( n3216 & n22008 ) | ( n12608 & n22008 ) ;
  assign n37243 = n24067 ^ n8320 ^ 1'b0 ;
  assign n37245 = n37244 ^ n37243 ^ n18193 ;
  assign n37246 = n1831 & ~n19363 ;
  assign n37247 = ~n14007 & n37246 ;
  assign n37248 = n36581 ^ n27063 ^ 1'b0 ;
  assign n37249 = n25332 & ~n37248 ;
  assign n37250 = n11593 ^ n7836 ^ 1'b0 ;
  assign n37251 = n27289 ^ n23542 ^ n12470 ;
  assign n37252 = n18840 | n30625 ;
  assign n37253 = n5014 & ~n37252 ;
  assign n37254 = n5516 & n7987 ;
  assign n37255 = n17139 & n37254 ;
  assign n37256 = ~n18272 & n37255 ;
  assign n37257 = n12757 | n37256 ;
  assign n37258 = n1998 & ~n37257 ;
  assign n37259 = ( n19600 & ~n37253 ) | ( n19600 & n37258 ) | ( ~n37253 & n37258 ) ;
  assign n37260 = ~n36758 & n37259 ;
  assign n37261 = n37260 ^ n8659 ^ 1'b0 ;
  assign n37262 = n8682 & ~n37261 ;
  assign n37263 = ( ~n25609 & n37251 ) | ( ~n25609 & n37262 ) | ( n37251 & n37262 ) ;
  assign n37264 = n33638 ^ n7971 ^ n761 ;
  assign n37265 = n37264 ^ n24493 ^ 1'b0 ;
  assign n37266 = n4271 & n7163 ;
  assign n37267 = n12178 & n37266 ;
  assign n37268 = n37267 ^ n15636 ^ 1'b0 ;
  assign n37269 = n15554 & n37268 ;
  assign n37270 = n37269 ^ n5996 ^ 1'b0 ;
  assign n37275 = n5799 & ~n9104 ;
  assign n37276 = n13226 & n37275 ;
  assign n37271 = n26271 ^ n13169 ^ 1'b0 ;
  assign n37272 = ~n4315 & n37271 ;
  assign n37273 = ( n30558 & n34300 ) | ( n30558 & ~n37272 ) | ( n34300 & ~n37272 ) ;
  assign n37274 = ~n24107 & n37273 ;
  assign n37277 = n37276 ^ n37274 ^ 1'b0 ;
  assign n37278 = n23959 ^ n18192 ^ n13020 ;
  assign n37279 = ( n899 & n7073 ) | ( n899 & n28677 ) | ( n7073 & n28677 ) ;
  assign n37280 = ( ~n16145 & n31732 ) | ( ~n16145 & n37279 ) | ( n31732 & n37279 ) ;
  assign n37281 = n18727 ^ n12870 ^ n1733 ;
  assign n37282 = ~n5726 & n10635 ;
  assign n37283 = n37282 ^ n4196 ^ 1'b0 ;
  assign n37284 = n19820 ^ n13249 ^ 1'b0 ;
  assign n37285 = n37284 ^ n20975 ^ 1'b0 ;
  assign n37286 = ~n7423 & n29475 ;
  assign n37287 = ( n4277 & n16063 ) | ( n4277 & n30166 ) | ( n16063 & n30166 ) ;
  assign n37288 = n33288 ^ n31197 ^ n19095 ;
  assign n37289 = n20791 | n21742 ;
  assign n37290 = n7548 | n37289 ;
  assign n37291 = n17322 & ~n37290 ;
  assign n37293 = n15035 ^ n9406 ^ 1'b0 ;
  assign n37294 = n10086 | n37293 ;
  assign n37295 = ( n9940 & n33499 ) | ( n9940 & n37294 ) | ( n33499 & n37294 ) ;
  assign n37292 = n11210 | n14941 ;
  assign n37296 = n37295 ^ n37292 ^ 1'b0 ;
  assign n37297 = n13195 ^ n7911 ^ n7230 ;
  assign n37298 = n37297 ^ n22077 ^ n14639 ;
  assign n37299 = n37298 ^ n20433 ^ n407 ;
  assign n37302 = n24341 ^ n2003 ^ n737 ;
  assign n37300 = n3406 & n17787 ;
  assign n37301 = ( n2931 & n32427 ) | ( n2931 & ~n37300 ) | ( n32427 & ~n37300 ) ;
  assign n37303 = n37302 ^ n37301 ^ n9790 ;
  assign n37304 = n28060 ^ n7561 ^ 1'b0 ;
  assign n37305 = n37304 ^ n18524 ^ n9156 ;
  assign n37306 = ( n14451 & n27832 ) | ( n14451 & n37305 ) | ( n27832 & n37305 ) ;
  assign n37307 = n37306 ^ n22107 ^ 1'b0 ;
  assign n37308 = n18459 ^ n1226 ^ 1'b0 ;
  assign n37309 = n27275 & n37308 ;
  assign n37312 = ( n5475 & n18036 ) | ( n5475 & n34720 ) | ( n18036 & n34720 ) ;
  assign n37310 = n17443 ^ n5699 ^ 1'b0 ;
  assign n37311 = n8328 & ~n37310 ;
  assign n37313 = n37312 ^ n37311 ^ 1'b0 ;
  assign n37314 = n6752 | n37313 ;
  assign n37315 = n13657 & n30375 ;
  assign n37316 = n37314 & n37315 ;
  assign n37317 = n30562 ^ n24318 ^ 1'b0 ;
  assign n37318 = n22662 ^ n17295 ^ n1896 ;
  assign n37324 = ~n1216 & n15660 ;
  assign n37325 = ( ~n9624 & n14180 ) | ( ~n9624 & n37324 ) | ( n14180 & n37324 ) ;
  assign n37326 = n37325 ^ n7725 ^ 1'b0 ;
  assign n37327 = ~n17451 & n37326 ;
  assign n37328 = n12725 & n37327 ;
  assign n37319 = n7576 | n25816 ;
  assign n37320 = n21676 ^ n13244 ^ n8853 ;
  assign n37321 = ~n37319 & n37320 ;
  assign n37322 = n7478 & n37321 ;
  assign n37323 = n23855 & ~n37322 ;
  assign n37329 = n37328 ^ n37323 ^ n9654 ;
  assign n37331 = ( n1769 & n15914 ) | ( n1769 & n25973 ) | ( n15914 & n25973 ) ;
  assign n37330 = n13664 & n32318 ;
  assign n37332 = n37331 ^ n37330 ^ n13209 ;
  assign n37333 = n1949 & ~n21919 ;
  assign n37334 = ~n9234 & n22138 ;
  assign n37335 = ~n6860 & n37334 ;
  assign n37336 = n35363 ^ n23243 ^ 1'b0 ;
  assign n37337 = ~n37335 & n37336 ;
  assign n37338 = n20339 ^ n12352 ^ n11919 ;
  assign n37339 = ( n8124 & n26100 ) | ( n8124 & ~n37338 ) | ( n26100 & ~n37338 ) ;
  assign n37340 = ( n5542 & n10662 ) | ( n5542 & ~n37339 ) | ( n10662 & ~n37339 ) ;
  assign n37341 = ( n9644 & n24905 ) | ( n9644 & ~n37340 ) | ( n24905 & ~n37340 ) ;
  assign n37342 = n6297 & ~n30927 ;
  assign n37343 = n37342 ^ n2469 ^ 1'b0 ;
  assign n37344 = n37343 ^ n10693 ^ n848 ;
  assign n37345 = n18524 & n21111 ;
  assign n37346 = ( ~n7638 & n27161 ) | ( ~n7638 & n37345 ) | ( n27161 & n37345 ) ;
  assign n37347 = n16940 ^ n3465 ^ 1'b0 ;
  assign n37348 = ( n3146 & ~n12188 ) | ( n3146 & n12817 ) | ( ~n12188 & n12817 ) ;
  assign n37349 = n14898 & n37348 ;
  assign n37350 = n37349 ^ n18316 ^ 1'b0 ;
  assign n37361 = ( n941 & n15318 ) | ( n941 & n27510 ) | ( n15318 & n27510 ) ;
  assign n37355 = n6413 ^ n3905 ^ 1'b0 ;
  assign n37356 = n3206 | n37355 ;
  assign n37352 = ~n8290 & n10689 ;
  assign n37353 = n37352 ^ n5574 ^ 1'b0 ;
  assign n37351 = ~n1538 & n6001 ;
  assign n37354 = n37353 ^ n37351 ^ 1'b0 ;
  assign n37357 = n37356 ^ n37354 ^ n7182 ;
  assign n37358 = n31310 & n37357 ;
  assign n37359 = n37358 ^ n22818 ^ 1'b0 ;
  assign n37360 = ~n5239 & n37359 ;
  assign n37362 = n37361 ^ n37360 ^ 1'b0 ;
  assign n37363 = n26363 ^ n18213 ^ 1'b0 ;
  assign n37364 = n2780 & ~n36637 ;
  assign n37365 = ~n2600 & n37364 ;
  assign n37366 = ~n37363 & n37365 ;
  assign n37367 = ( ~n3880 & n9266 ) | ( ~n3880 & n14682 ) | ( n9266 & n14682 ) ;
  assign n37368 = n16257 ^ n12062 ^ n2567 ;
  assign n37370 = n29198 & ~n35473 ;
  assign n37369 = ~n8663 & n25959 ;
  assign n37371 = n37370 ^ n37369 ^ 1'b0 ;
  assign n37372 = n25642 ^ n15079 ^ n3364 ;
  assign n37373 = n3636 & ~n37372 ;
  assign n37375 = n16353 ^ n15215 ^ 1'b0 ;
  assign n37376 = ( n2860 & n34885 ) | ( n2860 & ~n37375 ) | ( n34885 & ~n37375 ) ;
  assign n37374 = n29077 & ~n36360 ;
  assign n37377 = n37376 ^ n37374 ^ 1'b0 ;
  assign n37378 = n37377 ^ n9917 ^ 1'b0 ;
  assign n37379 = n37373 & n37378 ;
  assign n37380 = n13450 ^ n9993 ^ 1'b0 ;
  assign n37381 = n16317 ^ n11028 ^ n2365 ;
  assign n37387 = n24067 & ~n31123 ;
  assign n37388 = n37387 ^ n19588 ^ 1'b0 ;
  assign n37384 = n14315 ^ n1289 ^ 1'b0 ;
  assign n37385 = n14922 | n37384 ;
  assign n37386 = x181 | n37385 ;
  assign n37382 = n10629 ^ n672 ^ 1'b0 ;
  assign n37383 = n19112 | n37382 ;
  assign n37389 = n37388 ^ n37386 ^ n37383 ;
  assign n37390 = n37389 ^ n16086 ^ n14183 ;
  assign n37391 = n18101 ^ n9108 ^ n945 ;
  assign n37392 = n576 | n37391 ;
  assign n37393 = n2648 | n37392 ;
  assign n37394 = ~n36306 & n37393 ;
  assign n37395 = n35306 ^ n34562 ^ 1'b0 ;
  assign n37396 = n4213 & ~n27872 ;
  assign n37397 = n37396 ^ n1358 ^ 1'b0 ;
  assign n37398 = n7439 & n9751 ;
  assign n37399 = n1521 & n37398 ;
  assign n37400 = n29858 ^ n6668 ^ 1'b0 ;
  assign n37401 = n5768 | n37400 ;
  assign n37402 = n31444 & ~n33075 ;
  assign n37403 = ~n9568 & n34265 ;
  assign n37404 = ( ~n6355 & n12429 ) | ( ~n6355 & n19524 ) | ( n12429 & n19524 ) ;
  assign n37405 = n37404 ^ n13432 ^ 1'b0 ;
  assign n37406 = n2597 | n20203 ;
  assign n37407 = n2980 & ~n37406 ;
  assign n37408 = ~n11346 & n34009 ;
  assign n37409 = n3435 & ~n19931 ;
  assign n37410 = n37409 ^ n17985 ^ 1'b0 ;
  assign n37411 = ~n2605 & n22512 ;
  assign n37412 = n8647 & n37411 ;
  assign n37413 = ( n32670 & n37410 ) | ( n32670 & ~n37412 ) | ( n37410 & ~n37412 ) ;
  assign n37414 = ( n26847 & n27623 ) | ( n26847 & ~n28886 ) | ( n27623 & ~n28886 ) ;
  assign n37415 = n18141 ^ n4243 ^ 1'b0 ;
  assign n37416 = ~n1727 & n3404 ;
  assign n37417 = n37415 & ~n37416 ;
  assign n37418 = n25425 ^ n22502 ^ n10446 ;
  assign n37421 = n33157 ^ n20587 ^ n19355 ;
  assign n37419 = n16950 ^ n16511 ^ n2987 ;
  assign n37420 = n37419 ^ n31739 ^ 1'b0 ;
  assign n37422 = n37421 ^ n37420 ^ n5128 ;
  assign n37423 = n36918 ^ n12266 ^ n8538 ;
  assign n37424 = n6077 | n9515 ;
  assign n37425 = n37424 ^ n22809 ^ 1'b0 ;
  assign n37426 = n4295 & n37425 ;
  assign n37427 = ~n37423 & n37426 ;
  assign n37429 = n1429 | n14553 ;
  assign n37428 = ( x23 & n4082 ) | ( x23 & n6328 ) | ( n4082 & n6328 ) ;
  assign n37430 = n37429 ^ n37428 ^ n20641 ;
  assign n37431 = n37430 ^ n16528 ^ 1'b0 ;
  assign n37432 = n24428 ^ n5432 ^ n4563 ;
  assign n37436 = n5514 ^ n3428 ^ n2243 ;
  assign n37433 = ( n15827 & n19503 ) | ( n15827 & ~n34642 ) | ( n19503 & ~n34642 ) ;
  assign n37434 = ( n4023 & n13021 ) | ( n4023 & ~n37433 ) | ( n13021 & ~n37433 ) ;
  assign n37435 = n37434 ^ n21352 ^ 1'b0 ;
  assign n37437 = n37436 ^ n37435 ^ n19848 ;
  assign n37438 = ~n12014 & n21725 ;
  assign n37439 = n28940 & n37438 ;
  assign n37440 = ( n12207 & n24364 ) | ( n12207 & ~n37439 ) | ( n24364 & ~n37439 ) ;
  assign n37441 = n37440 ^ n25795 ^ n6370 ;
  assign n37444 = n34931 ^ n4325 ^ n1692 ;
  assign n37442 = n10309 ^ n7514 ^ 1'b0 ;
  assign n37443 = n24378 | n37442 ;
  assign n37445 = n37444 ^ n37443 ^ 1'b0 ;
  assign n37446 = ~n9810 & n37445 ;
  assign n37447 = ~n16983 & n36499 ;
  assign n37448 = ( n24016 & n36397 ) | ( n24016 & ~n37447 ) | ( n36397 & ~n37447 ) ;
  assign n37449 = n15090 ^ n9761 ^ 1'b0 ;
  assign n37450 = n37449 ^ n24578 ^ n24049 ;
  assign n37451 = n37450 ^ n4917 ^ n2739 ;
  assign n37452 = ( n6457 & n15906 ) | ( n6457 & n37451 ) | ( n15906 & n37451 ) ;
  assign n37453 = n18188 & n34123 ;
  assign n37457 = n26584 ^ n3154 ^ 1'b0 ;
  assign n37454 = ( x134 & n20590 ) | ( x134 & n32883 ) | ( n20590 & n32883 ) ;
  assign n37455 = ( ~n1104 & n25678 ) | ( ~n1104 & n37454 ) | ( n25678 & n37454 ) ;
  assign n37456 = n37455 ^ n11161 ^ 1'b0 ;
  assign n37458 = n37457 ^ n37456 ^ n2899 ;
  assign n37459 = ( ~n26783 & n30012 ) | ( ~n26783 & n37458 ) | ( n30012 & n37458 ) ;
  assign n37460 = n29434 ^ n12215 ^ 1'b0 ;
  assign n37461 = n4300 & n37460 ;
  assign n37462 = n24285 ^ n23577 ^ n20747 ;
  assign n37463 = n27175 ^ n18987 ^ 1'b0 ;
  assign n37464 = n37462 & ~n37463 ;
  assign n37465 = ~n37362 & n37464 ;
  assign n37466 = n32892 & n37465 ;
  assign n37467 = ( n2707 & ~n9356 ) | ( n2707 & n28753 ) | ( ~n9356 & n28753 ) ;
  assign n37468 = n18548 & n26918 ;
  assign n37469 = ~n2405 & n37468 ;
  assign n37470 = ~n4520 & n37469 ;
  assign n37471 = n13504 ^ n9299 ^ 1'b0 ;
  assign n37472 = n4864 & ~n6999 ;
  assign n37473 = n18085 ^ n3214 ^ n2438 ;
  assign n37474 = ( ~n18846 & n37472 ) | ( ~n18846 & n37473 ) | ( n37472 & n37473 ) ;
  assign n37475 = ( n32790 & n36541 ) | ( n32790 & n37474 ) | ( n36541 & n37474 ) ;
  assign n37477 = n16113 ^ n15235 ^ n10418 ;
  assign n37478 = ~n16317 & n37477 ;
  assign n37479 = n37478 ^ n14023 ^ 1'b0 ;
  assign n37476 = ( n17404 & ~n18376 ) | ( n17404 & n35532 ) | ( ~n18376 & n35532 ) ;
  assign n37480 = n37479 ^ n37476 ^ n13031 ;
  assign n37481 = n23141 ^ n19770 ^ 1'b0 ;
  assign n37482 = n736 & n37481 ;
  assign n37483 = n20936 ^ n12366 ^ 1'b0 ;
  assign n37484 = n18139 | n37483 ;
  assign n37485 = ( ~n5426 & n6999 ) | ( ~n5426 & n9175 ) | ( n6999 & n9175 ) ;
  assign n37486 = n25607 ^ n24621 ^ n20395 ;
  assign n37487 = n37485 & n37486 ;
  assign n37488 = ~n7174 & n37487 ;
  assign n37489 = n18061 ^ n6181 ^ 1'b0 ;
  assign n37490 = ( n1693 & n25251 ) | ( n1693 & n33276 ) | ( n25251 & n33276 ) ;
  assign n37491 = n37490 ^ n12451 ^ n5832 ;
  assign n37492 = ( n2330 & n37489 ) | ( n2330 & ~n37491 ) | ( n37489 & ~n37491 ) ;
  assign n37493 = n8243 & n20174 ;
  assign n37494 = n37493 ^ n4582 ^ n1233 ;
  assign n37495 = ( n12247 & ~n16475 ) | ( n12247 & n16855 ) | ( ~n16475 & n16855 ) ;
  assign n37496 = n37495 ^ n32143 ^ n9819 ;
  assign n37497 = n37496 ^ n8881 ^ 1'b0 ;
  assign n37499 = ( n1745 & ~n7354 ) | ( n1745 & n9412 ) | ( ~n7354 & n9412 ) ;
  assign n37498 = n23946 & n29840 ;
  assign n37500 = n37499 ^ n37498 ^ 1'b0 ;
  assign n37501 = n25715 ^ n24809 ^ n523 ;
  assign n37502 = n37501 ^ n29317 ^ n27214 ;
  assign n37503 = n37502 ^ n3672 ^ 1'b0 ;
  assign n37504 = ( n11798 & n18345 ) | ( n11798 & n37503 ) | ( n18345 & n37503 ) ;
  assign n37505 = n628 | n31377 ;
  assign n37506 = n37505 ^ n20108 ^ n745 ;
  assign n37507 = n16790 ^ n11649 ^ n5924 ;
  assign n37508 = n37507 ^ n34080 ^ n17164 ;
  assign n37509 = n24748 ^ n4162 ^ n3845 ;
  assign n37510 = n37509 ^ n13271 ^ n11766 ;
  assign n37511 = n15544 ^ n3140 ^ 1'b0 ;
  assign n37512 = ~n35426 & n37511 ;
  assign n37513 = n22108 & n37353 ;
  assign n37514 = n37513 ^ n23192 ^ n3833 ;
  assign n37515 = ( ~n7560 & n24373 ) | ( ~n7560 & n37514 ) | ( n24373 & n37514 ) ;
  assign n37516 = n24016 | n37515 ;
  assign n37517 = n10043 ^ n4078 ^ 1'b0 ;
  assign n37518 = n37517 ^ n34381 ^ n25746 ;
  assign n37519 = n35280 & n37518 ;
  assign n37520 = ~n5810 & n7857 ;
  assign n37521 = n37520 ^ n6543 ^ 1'b0 ;
  assign n37522 = n36603 & ~n37521 ;
  assign n37523 = ( n19966 & n36517 ) | ( n19966 & n37522 ) | ( n36517 & n37522 ) ;
  assign n37524 = ~n12340 & n23823 ;
  assign n37525 = n37524 ^ n24862 ^ n8352 ;
  assign n37526 = ( ~n17183 & n20797 ) | ( ~n17183 & n37525 ) | ( n20797 & n37525 ) ;
  assign n37527 = n15232 | n19823 ;
  assign n37529 = n36853 ^ n10959 ^ 1'b0 ;
  assign n37530 = n5044 & ~n37529 ;
  assign n37528 = n15531 ^ n6443 ^ n3759 ;
  assign n37531 = n37530 ^ n37528 ^ n1598 ;
  assign n37532 = ( n11677 & n19586 ) | ( n11677 & n28510 ) | ( n19586 & n28510 ) ;
  assign n37533 = n3373 | n3785 ;
  assign n37534 = n37532 | n37533 ;
  assign n37535 = n4438 ^ n1133 ^ x207 ;
  assign n37536 = ~n24457 & n37535 ;
  assign n37537 = n17811 | n23838 ;
  assign n37538 = n31212 | n37537 ;
  assign n37539 = n37538 ^ n32943 ^ n32338 ;
  assign n37541 = ( n3208 & ~n9482 ) | ( n3208 & n23635 ) | ( ~n9482 & n23635 ) ;
  assign n37540 = n10811 & ~n19714 ;
  assign n37542 = n37541 ^ n37540 ^ 1'b0 ;
  assign n37543 = ( n6431 & ~n24441 ) | ( n6431 & n32737 ) | ( ~n24441 & n32737 ) ;
  assign n37544 = n37543 ^ n17155 ^ n2577 ;
  assign n37545 = n35402 ^ n32392 ^ n14512 ;
  assign n37546 = n37545 ^ n16257 ^ n14385 ;
  assign n37547 = ~n1897 & n34568 ;
  assign n37548 = n35095 ^ n16691 ^ n13035 ;
  assign n37549 = n5738 & n12493 ;
  assign n37550 = n37549 ^ n8040 ^ 1'b0 ;
  assign n37551 = n4166 ^ n513 ^ 1'b0 ;
  assign n37552 = ~n21111 & n37551 ;
  assign n37553 = n6180 | n14342 ;
  assign n37554 = n18257 ^ n16811 ^ n2177 ;
  assign n37555 = ( n902 & ~n7605 ) | ( n902 & n8494 ) | ( ~n7605 & n8494 ) ;
  assign n37556 = n37554 & n37555 ;
  assign n37557 = ~n25250 & n37556 ;
  assign n37558 = n37553 & n37557 ;
  assign n37559 = n14537 ^ n1838 ^ 1'b0 ;
  assign n37560 = n37559 ^ n30170 ^ n15230 ;
  assign n37562 = ( ~n2331 & n26164 ) | ( ~n2331 & n29066 ) | ( n26164 & n29066 ) ;
  assign n37563 = ( n2592 & ~n9635 ) | ( n2592 & n37562 ) | ( ~n9635 & n37562 ) ;
  assign n37561 = ( ~n5620 & n15728 ) | ( ~n5620 & n17983 ) | ( n15728 & n17983 ) ;
  assign n37564 = n37563 ^ n37561 ^ n12603 ;
  assign n37565 = n14580 ^ n6946 ^ n5928 ;
  assign n37566 = n17167 ^ n12239 ^ 1'b0 ;
  assign n37567 = n37565 | n37566 ;
  assign n37568 = n20332 ^ n5600 ^ 1'b0 ;
  assign n37571 = n25232 ^ n14823 ^ 1'b0 ;
  assign n37572 = ~n4484 & n37571 ;
  assign n37569 = n8802 & ~n21234 ;
  assign n37570 = ~n26164 & n37569 ;
  assign n37573 = n37572 ^ n37570 ^ n35932 ;
  assign n37575 = n9328 | n16039 ;
  assign n37576 = n37575 ^ n35827 ^ 1'b0 ;
  assign n37577 = n14545 & n37576 ;
  assign n37578 = ~n8034 & n37577 ;
  assign n37579 = n37578 ^ n5333 ^ 1'b0 ;
  assign n37574 = n5643 & ~n23327 ;
  assign n37580 = n37579 ^ n37574 ^ 1'b0 ;
  assign n37581 = ( n11814 & n12186 ) | ( n11814 & n17582 ) | ( n12186 & n17582 ) ;
  assign n37582 = n30635 ^ n4271 ^ 1'b0 ;
  assign n37583 = n270 | n37223 ;
  assign n37584 = n9078 | n37583 ;
  assign n37585 = ~n6789 & n37584 ;
  assign n37586 = ~n9940 & n37585 ;
  assign n37587 = n37586 ^ n4090 ^ 1'b0 ;
  assign n37588 = n10287 ^ n3245 ^ n1643 ;
  assign n37589 = n30768 ^ n10501 ^ 1'b0 ;
  assign n37590 = n37588 & n37589 ;
  assign n37591 = n36590 ^ n17870 ^ 1'b0 ;
  assign n37592 = n29232 | n37591 ;
  assign n37593 = n20533 ^ n15685 ^ n10412 ;
  assign n37594 = ~n2064 & n5403 ;
  assign n37595 = n37593 & n37594 ;
  assign n37596 = n26816 ^ n13543 ^ n2999 ;
  assign n37597 = n37596 ^ n36573 ^ 1'b0 ;
  assign n37598 = ( n5404 & n7327 ) | ( n5404 & n18555 ) | ( n7327 & n18555 ) ;
  assign n37599 = n6092 & n17578 ;
  assign n37602 = n28824 & n33932 ;
  assign n37600 = n7047 & ~n28900 ;
  assign n37601 = n37600 ^ n6662 ^ 1'b0 ;
  assign n37603 = n37602 ^ n37601 ^ n8810 ;
  assign n37604 = n37603 ^ n27875 ^ 1'b0 ;
  assign n37605 = ( n5409 & n16870 ) | ( n5409 & ~n21585 ) | ( n16870 & ~n21585 ) ;
  assign n37608 = n8985 ^ n2887 ^ 1'b0 ;
  assign n37607 = n25988 ^ n12080 ^ 1'b0 ;
  assign n37606 = ( n9380 & n12018 ) | ( n9380 & n16859 ) | ( n12018 & n16859 ) ;
  assign n37609 = n37608 ^ n37607 ^ n37606 ;
  assign n37610 = n2329 | n2643 ;
  assign n37611 = n37610 ^ n20610 ^ 1'b0 ;
  assign n37612 = ~n2624 & n28041 ;
  assign n37618 = ( n6488 & n13192 ) | ( n6488 & ~n31123 ) | ( n13192 & ~n31123 ) ;
  assign n37619 = ( n2076 & n16856 ) | ( n2076 & ~n37618 ) | ( n16856 & ~n37618 ) ;
  assign n37620 = n27061 ^ n5104 ^ 1'b0 ;
  assign n37621 = n37619 & ~n37620 ;
  assign n37622 = n37621 ^ n15636 ^ 1'b0 ;
  assign n37613 = ( n5631 & n11212 ) | ( n5631 & n12914 ) | ( n11212 & n12914 ) ;
  assign n37614 = n1600 & n9414 ;
  assign n37615 = n37613 & n37614 ;
  assign n37616 = ( n295 & n20151 ) | ( n295 & ~n37615 ) | ( n20151 & ~n37615 ) ;
  assign n37617 = n9533 | n37616 ;
  assign n37623 = n37622 ^ n37617 ^ 1'b0 ;
  assign n37624 = n27701 ^ n12855 ^ x110 ;
  assign n37625 = n5189 ^ n1583 ^ 1'b0 ;
  assign n37626 = ( n4268 & n12286 ) | ( n4268 & n37625 ) | ( n12286 & n37625 ) ;
  assign n37627 = n25247 ^ n22770 ^ 1'b0 ;
  assign n37629 = ( ~n1050 & n2118 ) | ( ~n1050 & n6304 ) | ( n2118 & n6304 ) ;
  assign n37630 = n37629 ^ n15723 ^ n5670 ;
  assign n37628 = ~n690 & n8028 ;
  assign n37631 = n37630 ^ n37628 ^ n11400 ;
  assign n37638 = n9195 ^ n5482 ^ n3675 ;
  assign n37634 = n10288 ^ n9166 ^ 1'b0 ;
  assign n37635 = n1692 | n37634 ;
  assign n37636 = n24382 ^ n3911 ^ 1'b0 ;
  assign n37637 = ~n37635 & n37636 ;
  assign n37639 = n37638 ^ n37637 ^ n2975 ;
  assign n37632 = ( n3373 & n13863 ) | ( n3373 & ~n20265 ) | ( n13863 & ~n20265 ) ;
  assign n37633 = n37632 ^ n6640 ^ n2863 ;
  assign n37640 = n37639 ^ n37633 ^ 1'b0 ;
  assign n37641 = n16743 ^ n6313 ^ 1'b0 ;
  assign n37642 = n37640 & ~n37641 ;
  assign n37649 = n26893 ^ n24373 ^ n1028 ;
  assign n37650 = n37649 ^ n7381 ^ 1'b0 ;
  assign n37645 = n1396 & n13137 ;
  assign n37646 = ~n21854 & n37645 ;
  assign n37647 = ~n28423 & n37646 ;
  assign n37648 = ~n26260 & n37647 ;
  assign n37643 = ( n4297 & n20886 ) | ( n4297 & n32012 ) | ( n20886 & n32012 ) ;
  assign n37644 = ( ~n3203 & n33655 ) | ( ~n3203 & n37643 ) | ( n33655 & n37643 ) ;
  assign n37651 = n37650 ^ n37648 ^ n37644 ;
  assign n37652 = n17772 | n26958 ;
  assign n37653 = n28568 | n37652 ;
  assign n37654 = ( ~n13764 & n14778 ) | ( ~n13764 & n29632 ) | ( n14778 & n29632 ) ;
  assign n37655 = n37654 ^ n36728 ^ n12603 ;
  assign n37656 = n15494 & n31289 ;
  assign n37657 = n37656 ^ n26820 ^ 1'b0 ;
  assign n37658 = n37657 ^ n36293 ^ 1'b0 ;
  assign n37659 = n518 & ~n11784 ;
  assign n37660 = n37659 ^ n8319 ^ 1'b0 ;
  assign n37661 = n14946 & n37660 ;
  assign n37662 = n37661 ^ n17472 ^ 1'b0 ;
  assign n37663 = n37662 ^ n23503 ^ n22627 ;
  assign n37664 = n10048 | n37663 ;
  assign n37665 = n31770 & n34064 ;
  assign n37666 = n37665 ^ n19259 ^ 1'b0 ;
  assign n37667 = n28512 ^ n3881 ^ 1'b0 ;
  assign n37668 = ( n10075 & ~n17225 ) | ( n10075 & n37667 ) | ( ~n17225 & n37667 ) ;
  assign n37669 = n22846 | n37668 ;
  assign n37670 = n10290 & n37669 ;
  assign n37671 = n37670 ^ n16327 ^ 1'b0 ;
  assign n37672 = n3535 & ~n17178 ;
  assign n37686 = ~n12920 & n26845 ;
  assign n37678 = ( n1400 & n13082 ) | ( n1400 & n25280 ) | ( n13082 & n25280 ) ;
  assign n37679 = n20778 ^ n19820 ^ n1990 ;
  assign n37680 = ~n14485 & n31756 ;
  assign n37681 = ~n37679 & n37680 ;
  assign n37682 = ( n6948 & ~n21823 ) | ( n6948 & n37681 ) | ( ~n21823 & n37681 ) ;
  assign n37683 = ( ~n10411 & n37678 ) | ( ~n10411 & n37682 ) | ( n37678 & n37682 ) ;
  assign n37684 = n6229 | n37683 ;
  assign n37685 = n37684 ^ n23093 ^ 1'b0 ;
  assign n37687 = n37686 ^ n37685 ^ n23904 ;
  assign n37673 = n6064 ^ n5537 ^ 1'b0 ;
  assign n37674 = n11357 & n19512 ;
  assign n37675 = n37673 & n37674 ;
  assign n37676 = n3126 | n37675 ;
  assign n37677 = n29284 & ~n37676 ;
  assign n37688 = n37687 ^ n37677 ^ n14967 ;
  assign n37689 = n37688 ^ n6095 ^ 1'b0 ;
  assign n37690 = n7415 & n12515 ;
  assign n37691 = n2357 | n16256 ;
  assign n37692 = n37691 ^ n13087 ^ 1'b0 ;
  assign n37693 = ~n17410 & n23482 ;
  assign n37694 = ( ~n12854 & n37692 ) | ( ~n12854 & n37693 ) | ( n37692 & n37693 ) ;
  assign n37695 = n8836 & n23576 ;
  assign n37696 = n37694 & ~n37695 ;
  assign n37697 = ( n25619 & n37690 ) | ( n25619 & n37696 ) | ( n37690 & n37696 ) ;
  assign n37698 = n36927 ^ n14278 ^ 1'b0 ;
  assign n37699 = ~n6569 & n37698 ;
  assign n37700 = n1874 | n12767 ;
  assign n37701 = n37700 ^ n4706 ^ 1'b0 ;
  assign n37702 = n34725 ^ n23711 ^ 1'b0 ;
  assign n37703 = ~n37701 & n37702 ;
  assign n37704 = ( n1670 & n15137 ) | ( n1670 & ~n21287 ) | ( n15137 & ~n21287 ) ;
  assign n37705 = n37704 ^ n5866 ^ n458 ;
  assign n37706 = n37705 ^ n5786 ^ 1'b0 ;
  assign n37707 = n31222 ^ n15738 ^ 1'b0 ;
  assign n37708 = n2863 & ~n37707 ;
  assign n37709 = n15900 & n31328 ;
  assign n37710 = ( n37706 & ~n37708 ) | ( n37706 & n37709 ) | ( ~n37708 & n37709 ) ;
  assign n37711 = n32818 ^ n17160 ^ 1'b0 ;
  assign n37712 = n16563 & ~n32440 ;
  assign n37713 = n37712 ^ n8336 ^ 1'b0 ;
  assign n37714 = ( ~n36738 & n37711 ) | ( ~n36738 & n37713 ) | ( n37711 & n37713 ) ;
  assign n37715 = n18504 & ~n20276 ;
  assign n37716 = n19525 & n37715 ;
  assign n37717 = n19675 ^ n4374 ^ n3963 ;
  assign n37718 = n7259 & n12262 ;
  assign n37719 = ~n37717 & n37718 ;
  assign n37720 = ~n20186 & n21830 ;
  assign n37721 = n37720 ^ n28122 ^ 1'b0 ;
  assign n37722 = n23899 & n37721 ;
  assign n37723 = n37722 ^ n16454 ^ n6706 ;
  assign n37724 = n31902 & n37723 ;
  assign n37725 = n32972 ^ n6477 ^ n3838 ;
  assign n37726 = n372 & ~n2179 ;
  assign n37727 = n37726 ^ n16145 ^ n7662 ;
  assign n37728 = n13288 & n37727 ;
  assign n37729 = ~n6909 & n37728 ;
  assign n37730 = ( n1183 & ~n34863 ) | ( n1183 & n37729 ) | ( ~n34863 & n37729 ) ;
  assign n37731 = ~n25651 & n37730 ;
  assign n37732 = n21406 ^ n1826 ^ n1446 ;
  assign n37733 = n12845 | n14941 ;
  assign n37734 = n37733 ^ n9754 ^ 1'b0 ;
  assign n37735 = ( x5 & ~n11838 ) | ( x5 & n23628 ) | ( ~n11838 & n23628 ) ;
  assign n37736 = ( ~n13385 & n33664 ) | ( ~n13385 & n37735 ) | ( n33664 & n37735 ) ;
  assign n37737 = n37736 ^ n22817 ^ 1'b0 ;
  assign n37738 = n37734 & ~n37737 ;
  assign n37739 = n21133 | n37738 ;
  assign n37740 = n20649 ^ n20135 ^ 1'b0 ;
  assign n37741 = ~n7247 & n37740 ;
  assign n37744 = n24013 ^ n9071 ^ 1'b0 ;
  assign n37745 = n25657 ^ n17449 ^ 1'b0 ;
  assign n37746 = n37744 & ~n37745 ;
  assign n37742 = n9256 ^ n7468 ^ n4642 ;
  assign n37743 = ~n8290 & n37742 ;
  assign n37747 = n37746 ^ n37743 ^ 1'b0 ;
  assign n37749 = n5232 ^ n2946 ^ n1670 ;
  assign n37748 = n2106 & n10939 ;
  assign n37750 = n37749 ^ n37748 ^ n25658 ;
  assign n37752 = ( ~n9292 & n9991 ) | ( ~n9292 & n19095 ) | ( n9991 & n19095 ) ;
  assign n37751 = ( n258 & n16308 ) | ( n258 & ~n27989 ) | ( n16308 & ~n27989 ) ;
  assign n37753 = n37752 ^ n37751 ^ n6127 ;
  assign n37754 = ( n20944 & n28173 ) | ( n20944 & ~n37753 ) | ( n28173 & ~n37753 ) ;
  assign n37755 = ~n37678 & n37754 ;
  assign n37756 = n7070 & n37755 ;
  assign n37757 = n37756 ^ n9736 ^ 1'b0 ;
  assign n37758 = n6947 & ~n16703 ;
  assign n37759 = ~n2693 & n37758 ;
  assign n37760 = n37759 ^ n18944 ^ n15913 ;
  assign n37761 = ( ~n1988 & n17549 ) | ( ~n1988 & n37760 ) | ( n17549 & n37760 ) ;
  assign n37762 = n37761 ^ n31415 ^ 1'b0 ;
  assign n37763 = ~n1570 & n37762 ;
  assign n37765 = ( n11319 & n15217 ) | ( n11319 & ~n18998 ) | ( n15217 & ~n18998 ) ;
  assign n37764 = n11717 ^ n9512 ^ 1'b0 ;
  assign n37766 = n37765 ^ n37764 ^ n17653 ;
  assign n37767 = n37766 ^ n8178 ^ 1'b0 ;
  assign n37768 = n32763 ^ n28790 ^ n5889 ;
  assign n37769 = ~n7836 & n37768 ;
  assign n37770 = n37769 ^ n26824 ^ n13321 ;
  assign n37771 = n21789 ^ n13312 ^ n6165 ;
  assign n37772 = ~n15401 & n37771 ;
  assign n37773 = ~n10475 & n20849 ;
  assign n37774 = ~n4939 & n37773 ;
  assign n37775 = n16640 & ~n33246 ;
  assign n37776 = n23823 ^ n18336 ^ 1'b0 ;
  assign n37777 = ~n37775 & n37776 ;
  assign n37778 = n17220 ^ n11022 ^ 1'b0 ;
  assign n37779 = n25042 & n37778 ;
  assign n37780 = n35426 ^ n27555 ^ n23375 ;
  assign n37781 = n3111 & n32565 ;
  assign n37782 = n19418 ^ n7333 ^ 1'b0 ;
  assign n37783 = n2510 | n37782 ;
  assign n37784 = n5921 | n37783 ;
  assign n37785 = ( n678 & n34598 ) | ( n678 & n37784 ) | ( n34598 & n37784 ) ;
  assign n37786 = n37785 ^ n32072 ^ n934 ;
  assign n37787 = n10154 & n19128 ;
  assign n37788 = n10723 & ~n37787 ;
  assign n37789 = n36808 & n37788 ;
  assign n37790 = n12295 ^ n5650 ^ 1'b0 ;
  assign n37791 = n22670 ^ n9621 ^ 1'b0 ;
  assign n37792 = n37790 | n37791 ;
  assign n37793 = n19629 | n37792 ;
  assign n37794 = n37793 ^ n18620 ^ 1'b0 ;
  assign n37795 = n6061 & ~n12132 ;
  assign n37796 = n37795 ^ n34346 ^ n7958 ;
  assign n37797 = n37796 ^ n18237 ^ x230 ;
  assign n37798 = n9892 | n31058 ;
  assign n37799 = n37798 ^ n22736 ^ 1'b0 ;
  assign n37800 = n5703 | n20887 ;
  assign n37801 = ( n23848 & n24972 ) | ( n23848 & n37800 ) | ( n24972 & n37800 ) ;
  assign n37802 = n37801 ^ n34538 ^ 1'b0 ;
  assign n37803 = n37802 ^ n13954 ^ 1'b0 ;
  assign n37804 = n1555 & n13286 ;
  assign n37805 = n37804 ^ n12766 ^ 1'b0 ;
  assign n37806 = n32601 | n37805 ;
  assign n37807 = n17260 & ~n37806 ;
  assign n37808 = ( n1140 & n4339 ) | ( n1140 & n21740 ) | ( n4339 & n21740 ) ;
  assign n37809 = n37808 ^ n2217 ^ 1'b0 ;
  assign n37810 = ~n14214 & n37809 ;
  assign n37811 = n22658 ^ n1545 ^ 1'b0 ;
  assign n37812 = n26310 & n37811 ;
  assign n37813 = n7009 & n17622 ;
  assign n37815 = ( n481 & n15517 ) | ( n481 & n28774 ) | ( n15517 & n28774 ) ;
  assign n37814 = n17807 ^ n10943 ^ 1'b0 ;
  assign n37816 = n37815 ^ n37814 ^ 1'b0 ;
  assign n37817 = x253 & n37816 ;
  assign n37818 = ( n6472 & n34917 ) | ( n6472 & ~n37817 ) | ( n34917 & ~n37817 ) ;
  assign n37819 = n37818 ^ n18993 ^ 1'b0 ;
  assign n37820 = n37813 & n37819 ;
  assign n37821 = n32496 ^ n16839 ^ 1'b0 ;
  assign n37822 = n25096 ^ n16367 ^ 1'b0 ;
  assign n37823 = n2732 & ~n37822 ;
  assign n37824 = n37823 ^ n13656 ^ n5786 ;
  assign n37825 = n24492 & n37824 ;
  assign n37826 = ( ~n15083 & n29904 ) | ( ~n15083 & n37825 ) | ( n29904 & n37825 ) ;
  assign n37828 = n4228 ^ n1226 ^ 1'b0 ;
  assign n37827 = n3642 & ~n10318 ;
  assign n37829 = n37828 ^ n37827 ^ n8601 ;
  assign n37830 = ( n2128 & ~n6776 ) | ( n2128 & n16753 ) | ( ~n6776 & n16753 ) ;
  assign n37831 = ( n713 & n37829 ) | ( n713 & ~n37830 ) | ( n37829 & ~n37830 ) ;
  assign n37832 = n37831 ^ n26515 ^ n16292 ;
  assign n37833 = n16354 ^ n8522 ^ 1'b0 ;
  assign n37834 = n28908 ^ n13932 ^ 1'b0 ;
  assign n37835 = ~n19310 & n37834 ;
  assign n37836 = n9349 & n13723 ;
  assign n37837 = n37836 ^ n32028 ^ 1'b0 ;
  assign n37838 = ~n6020 & n6432 ;
  assign n37839 = n37838 ^ n20013 ^ 1'b0 ;
  assign n37840 = ( ~n2014 & n10067 ) | ( ~n2014 & n37839 ) | ( n10067 & n37839 ) ;
  assign n37841 = n37840 ^ n767 ^ 1'b0 ;
  assign n37842 = n26312 & ~n37841 ;
  assign n37843 = n7262 ^ n896 ^ 1'b0 ;
  assign n37844 = n37404 | n37843 ;
  assign n37845 = n29634 ^ n5046 ^ 1'b0 ;
  assign n37846 = n9656 | n37845 ;
  assign n37847 = n37846 ^ n6255 ^ 1'b0 ;
  assign n37848 = ~n6712 & n16040 ;
  assign n37849 = n37848 ^ n13168 ^ 1'b0 ;
  assign n37850 = n20450 ^ n9080 ^ 1'b0 ;
  assign n37851 = ( n9611 & n17966 ) | ( n9611 & n37850 ) | ( n17966 & n37850 ) ;
  assign n37854 = n10712 ^ n7897 ^ 1'b0 ;
  assign n37852 = n35988 ^ n7480 ^ 1'b0 ;
  assign n37853 = n4313 | n37852 ;
  assign n37855 = n37854 ^ n37853 ^ n33217 ;
  assign n37856 = ~n10223 & n16658 ;
  assign n37857 = ( n33564 & ~n37276 ) | ( n33564 & n37856 ) | ( ~n37276 & n37856 ) ;
  assign n37858 = n20200 ^ n1781 ^ 1'b0 ;
  assign n37859 = n514 | n37858 ;
  assign n37860 = n6948 | n37859 ;
  assign n37861 = ~n7858 & n25250 ;
  assign n37862 = n37861 ^ n34562 ^ n11746 ;
  assign n37863 = n37862 ^ n14108 ^ 1'b0 ;
  assign n37864 = n28303 ^ n8654 ^ n7645 ;
  assign n37865 = ( n6342 & n8869 ) | ( n6342 & ~n22658 ) | ( n8869 & ~n22658 ) ;
  assign n37866 = n15147 ^ n9114 ^ n4348 ;
  assign n37867 = ( n3948 & n29062 ) | ( n3948 & ~n37866 ) | ( n29062 & ~n37866 ) ;
  assign n37868 = ( n4217 & ~n7734 ) | ( n4217 & n15234 ) | ( ~n7734 & n15234 ) ;
  assign n37869 = n8196 | n37868 ;
  assign n37870 = n33373 & ~n37869 ;
  assign n37871 = n31200 ^ n9864 ^ 1'b0 ;
  assign n37872 = n32244 & ~n37871 ;
  assign n37873 = x206 & ~n20754 ;
  assign n37874 = n37873 ^ n17313 ^ 1'b0 ;
  assign n37875 = ( n9609 & n13702 ) | ( n9609 & ~n18677 ) | ( n13702 & ~n18677 ) ;
  assign n37876 = n37875 ^ n8828 ^ 1'b0 ;
  assign n37877 = ( n12162 & n19421 ) | ( n12162 & n37876 ) | ( n19421 & n37876 ) ;
  assign n37878 = n34017 ^ n22517 ^ 1'b0 ;
  assign n37879 = n19811 ^ n9017 ^ n7403 ;
  assign n37880 = n37879 ^ n33074 ^ n7721 ;
  assign n37881 = ( n20169 & n37878 ) | ( n20169 & ~n37880 ) | ( n37878 & ~n37880 ) ;
  assign n37882 = n7333 | n10638 ;
  assign n37883 = n37882 ^ n15733 ^ 1'b0 ;
  assign n37884 = n16601 & ~n37883 ;
  assign n37885 = ~n29081 & n37884 ;
  assign n37886 = ~n883 & n6828 ;
  assign n37887 = ( n20625 & ~n20939 ) | ( n20625 & n25946 ) | ( ~n20939 & n25946 ) ;
  assign n37888 = ( n7845 & n12700 ) | ( n7845 & n27210 ) | ( n12700 & n27210 ) ;
  assign n37889 = ( n3668 & n37887 ) | ( n3668 & n37888 ) | ( n37887 & n37888 ) ;
  assign n37890 = ~n2947 & n15843 ;
  assign n37891 = ~n10212 & n37890 ;
  assign n37892 = n26630 & n37891 ;
  assign n37893 = ( n8982 & n24537 ) | ( n8982 & n29666 ) | ( n24537 & n29666 ) ;
  assign n37894 = ( n27675 & n31328 ) | ( n27675 & ~n37893 ) | ( n31328 & ~n37893 ) ;
  assign n37895 = ( ~n5140 & n6503 ) | ( ~n5140 & n11883 ) | ( n6503 & n11883 ) ;
  assign n37896 = n37895 ^ n24563 ^ n5929 ;
  assign n37897 = n37896 ^ n16174 ^ n7989 ;
  assign n37898 = n37897 ^ n22063 ^ 1'b0 ;
  assign n37900 = n18403 | n29431 ;
  assign n37899 = ( n7334 & n28912 ) | ( n7334 & n33244 ) | ( n28912 & n33244 ) ;
  assign n37901 = n37900 ^ n37899 ^ n8625 ;
  assign n37902 = n1786 | n9156 ;
  assign n37903 = n9505 | n37902 ;
  assign n37904 = n37903 ^ n27985 ^ n8834 ;
  assign n37905 = n37324 ^ n33782 ^ n14912 ;
  assign n37906 = ~n11762 & n13256 ;
  assign n37907 = n37906 ^ n23683 ^ n20701 ;
  assign n37908 = ~n3951 & n29619 ;
  assign n37909 = n37907 & n37908 ;
  assign n37910 = ~n37905 & n37909 ;
  assign n37911 = n4379 | n25580 ;
  assign n37912 = n37911 ^ n11915 ^ 1'b0 ;
  assign n37913 = n16634 ^ n508 ^ 1'b0 ;
  assign n37914 = n7351 | n37913 ;
  assign n37915 = n37914 ^ n20136 ^ 1'b0 ;
  assign n37916 = n9492 & n26992 ;
  assign n37917 = n13618 & n37916 ;
  assign n37918 = ( n6423 & n20639 ) | ( n6423 & ~n37917 ) | ( n20639 & ~n37917 ) ;
  assign n37919 = n37918 ^ n32705 ^ n3520 ;
  assign n37920 = n23331 & n27371 ;
  assign n37921 = ~n14455 & n16042 ;
  assign n37922 = ~n37920 & n37921 ;
  assign n37923 = ( n6928 & ~n16484 ) | ( n6928 & n37922 ) | ( ~n16484 & n37922 ) ;
  assign n37924 = n37923 ^ n20318 ^ n16082 ;
  assign n37925 = ( n9955 & n20807 ) | ( n9955 & ~n24013 ) | ( n20807 & ~n24013 ) ;
  assign n37926 = n37925 ^ n17183 ^ 1'b0 ;
  assign n37927 = n37926 ^ n6671 ^ 1'b0 ;
  assign n37928 = n8583 & n12339 ;
  assign n37929 = n30379 ^ n4626 ^ n2158 ;
  assign n37930 = n37929 ^ n8253 ^ 1'b0 ;
  assign n37931 = n37930 ^ n37522 ^ n9084 ;
  assign n37932 = n37338 ^ n5140 ^ 1'b0 ;
  assign n37933 = n37932 ^ n10967 ^ 1'b0 ;
  assign n37934 = n18885 ^ n18386 ^ 1'b0 ;
  assign n37935 = n14019 & n37934 ;
  assign n37936 = n31243 ^ n30498 ^ 1'b0 ;
  assign n37937 = n6033 ^ n2860 ^ n2648 ;
  assign n37938 = n37937 ^ n3748 ^ 1'b0 ;
  assign n37939 = n31177 | n37938 ;
  assign n37940 = n3253 & ~n37939 ;
  assign n37941 = n7903 & ~n37940 ;
  assign n37942 = ( n14007 & ~n16513 ) | ( n14007 & n29741 ) | ( ~n16513 & n29741 ) ;
  assign n37944 = ( n4210 & ~n8092 ) | ( n4210 & n14197 ) | ( ~n8092 & n14197 ) ;
  assign n37945 = n18723 ^ n5385 ^ 1'b0 ;
  assign n37946 = n37944 & n37945 ;
  assign n37943 = n19306 ^ n10137 ^ 1'b0 ;
  assign n37947 = n37946 ^ n37943 ^ n29173 ;
  assign n37948 = n37947 ^ n23025 ^ n1664 ;
  assign n37950 = n3293 & n15337 ;
  assign n37949 = n2467 & ~n15529 ;
  assign n37951 = n37950 ^ n37949 ^ 1'b0 ;
  assign n37952 = n37951 ^ n12763 ^ n3353 ;
  assign n37954 = n23929 ^ n9285 ^ 1'b0 ;
  assign n37955 = n28518 | n37954 ;
  assign n37953 = n31344 ^ n20335 ^ n352 ;
  assign n37956 = n37955 ^ n37953 ^ 1'b0 ;
  assign n37957 = n12755 & n12821 ;
  assign n37958 = n17690 ^ n10139 ^ 1'b0 ;
  assign n37959 = n3380 & n37958 ;
  assign n37960 = n28707 ^ n14504 ^ 1'b0 ;
  assign n37961 = ( n1313 & n1600 ) | ( n1313 & n5404 ) | ( n1600 & n5404 ) ;
  assign n37962 = ( n683 & ~n14406 ) | ( n683 & n37961 ) | ( ~n14406 & n37961 ) ;
  assign n37963 = n6992 | n26479 ;
  assign n37964 = n37963 ^ n5163 ^ 1'b0 ;
  assign n37965 = n37964 ^ n29004 ^ n5164 ;
  assign n37966 = ~n16068 & n22272 ;
  assign n37967 = n24924 & n37966 ;
  assign n37968 = n28496 & n37967 ;
  assign n37970 = n23868 ^ n15142 ^ 1'b0 ;
  assign n37971 = n9483 & ~n37970 ;
  assign n37972 = ( n1684 & n8841 ) | ( n1684 & n37971 ) | ( n8841 & n37971 ) ;
  assign n37969 = n21694 & n22882 ;
  assign n37973 = n37972 ^ n37969 ^ 1'b0 ;
  assign n37974 = n8701 & ~n37973 ;
  assign n37975 = n8638 | n14590 ;
  assign n37976 = n24458 ^ n21339 ^ 1'b0 ;
  assign n37977 = n6327 & ~n37976 ;
  assign n37979 = n6315 | n24576 ;
  assign n37978 = n4624 | n34400 ;
  assign n37980 = n37979 ^ n37978 ^ 1'b0 ;
  assign n37981 = ~n11051 & n20650 ;
  assign n37982 = n37980 & n37981 ;
  assign n37983 = ( ~n2935 & n15142 ) | ( ~n2935 & n32283 ) | ( n15142 & n32283 ) ;
  assign n37987 = n18345 ^ n5224 ^ x41 ;
  assign n37985 = n6654 & n11681 ;
  assign n37984 = n22395 ^ n20460 ^ n488 ;
  assign n37986 = n37985 ^ n37984 ^ n29975 ;
  assign n37988 = n37987 ^ n37986 ^ n22443 ;
  assign n37989 = n2432 | n17482 ;
  assign n37990 = n37989 ^ n7550 ^ n3311 ;
  assign n37992 = n8907 ^ n5430 ^ 1'b0 ;
  assign n37993 = n5458 | n37992 ;
  assign n37991 = ~n3500 & n9936 ;
  assign n37994 = n37993 ^ n37991 ^ 1'b0 ;
  assign n37995 = ~n3773 & n23796 ;
  assign n37996 = n25729 | n37995 ;
  assign n37997 = n19189 & ~n37996 ;
  assign n37998 = n37997 ^ n2312 ^ 1'b0 ;
  assign n38000 = n6014 & ~n20872 ;
  assign n38001 = n15595 & n38000 ;
  assign n38002 = n38001 ^ n27784 ^ n25294 ;
  assign n37999 = n22086 ^ n10620 ^ n394 ;
  assign n38003 = n38002 ^ n37999 ^ 1'b0 ;
  assign n38004 = n35681 ^ n32753 ^ n29669 ;
  assign n38005 = n18197 ^ n9139 ^ n5472 ;
  assign n38006 = n38005 ^ n26671 ^ 1'b0 ;
  assign n38007 = n22439 & ~n38006 ;
  assign n38008 = n11779 ^ x45 ^ 1'b0 ;
  assign n38009 = n22574 & ~n38008 ;
  assign n38010 = n38009 ^ n12830 ^ 1'b0 ;
  assign n38011 = n4601 & n38010 ;
  assign n38012 = ~n387 & n15059 ;
  assign n38013 = n26449 ^ n25641 ^ 1'b0 ;
  assign n38014 = n4217 | n38013 ;
  assign n38015 = n38014 ^ n23304 ^ n19659 ;
  assign n38016 = n21485 ^ n5882 ^ n3952 ;
  assign n38017 = n29649 & ~n38016 ;
  assign n38020 = ( n1671 & n3817 ) | ( n1671 & n23861 ) | ( n3817 & n23861 ) ;
  assign n38021 = n34412 ^ n12717 ^ n2305 ;
  assign n38022 = ( n26874 & n38020 ) | ( n26874 & ~n38021 ) | ( n38020 & ~n38021 ) ;
  assign n38018 = ( ~n18893 & n22472 ) | ( ~n18893 & n24297 ) | ( n22472 & n24297 ) ;
  assign n38019 = n34832 | n38018 ;
  assign n38023 = n38022 ^ n38019 ^ 1'b0 ;
  assign n38024 = n18526 & n23518 ;
  assign n38025 = n6061 | n38024 ;
  assign n38026 = n38025 ^ n17451 ^ 1'b0 ;
  assign n38027 = n22286 ^ n384 ^ x217 ;
  assign n38028 = ( n18621 & n23946 ) | ( n18621 & n38027 ) | ( n23946 & n38027 ) ;
  assign n38029 = ( n426 & n10334 ) | ( n426 & ~n33100 ) | ( n10334 & ~n33100 ) ;
  assign n38030 = n19014 ^ n16615 ^ 1'b0 ;
  assign n38039 = n31727 ^ n29813 ^ n28173 ;
  assign n38040 = ~n12200 & n38039 ;
  assign n38041 = n38040 ^ n617 ^ 1'b0 ;
  assign n38033 = ( n18810 & n23088 ) | ( n18810 & n27316 ) | ( n23088 & n27316 ) ;
  assign n38034 = ( ~n16336 & n30047 ) | ( ~n16336 & n38033 ) | ( n30047 & n38033 ) ;
  assign n38032 = ~n10201 & n26363 ;
  assign n38031 = n30843 | n32090 ;
  assign n38035 = n38034 ^ n38032 ^ n38031 ;
  assign n38036 = ( n20729 & n29039 ) | ( n20729 & n38035 ) | ( n29039 & n38035 ) ;
  assign n38037 = n7188 | n38036 ;
  assign n38038 = n36240 | n38037 ;
  assign n38042 = n38041 ^ n38038 ^ n615 ;
  assign n38043 = n31094 ^ n6678 ^ 1'b0 ;
  assign n38044 = ( n18693 & n18804 ) | ( n18693 & ~n38043 ) | ( n18804 & ~n38043 ) ;
  assign n38045 = n8792 & ~n19242 ;
  assign n38046 = ( n4526 & ~n5722 ) | ( n4526 & n20357 ) | ( ~n5722 & n20357 ) ;
  assign n38047 = ( n1131 & ~n32267 ) | ( n1131 & n37113 ) | ( ~n32267 & n37113 ) ;
  assign n38049 = n744 | n7069 ;
  assign n38050 = n38049 ^ n23144 ^ 1'b0 ;
  assign n38051 = n4853 & n38050 ;
  assign n38048 = ~n12609 & n37570 ;
  assign n38052 = n38051 ^ n38048 ^ n4593 ;
  assign n38053 = n11289 & n30046 ;
  assign n38054 = n2973 & n38053 ;
  assign n38055 = n38054 ^ n27843 ^ 1'b0 ;
  assign n38056 = n21911 ^ n2716 ^ 1'b0 ;
  assign n38057 = ( n12238 & n17780 ) | ( n12238 & ~n38056 ) | ( n17780 & ~n38056 ) ;
  assign n38058 = n6386 & ~n16037 ;
  assign n38059 = n38058 ^ n28687 ^ 1'b0 ;
  assign n38060 = ( n626 & ~n22639 ) | ( n626 & n37013 ) | ( ~n22639 & n37013 ) ;
  assign n38061 = n6678 & n15877 ;
  assign n38062 = n33564 & n38061 ;
  assign n38063 = n13072 ^ n529 ^ 1'b0 ;
  assign n38064 = n20973 ^ n13985 ^ n11058 ;
  assign n38065 = ( ~n38062 & n38063 ) | ( ~n38062 & n38064 ) | ( n38063 & n38064 ) ;
  assign n38066 = n32304 ^ n25442 ^ n13888 ;
  assign n38067 = n37808 ^ n7993 ^ n1233 ;
  assign n38068 = ( ~n12521 & n30045 ) | ( ~n12521 & n38067 ) | ( n30045 & n38067 ) ;
  assign n38069 = n32158 ^ n31794 ^ 1'b0 ;
  assign n38070 = n2728 | n3557 ;
  assign n38071 = n9232 & ~n38070 ;
  assign n38072 = n30207 ^ n24545 ^ 1'b0 ;
  assign n38073 = n12350 ^ n2317 ^ 1'b0 ;
  assign n38074 = n16019 | n38073 ;
  assign n38075 = n25114 ^ n23356 ^ 1'b0 ;
  assign n38076 = n854 & n38075 ;
  assign n38077 = n38076 ^ n29656 ^ n27426 ;
  assign n38079 = ( n2048 & n5669 ) | ( n2048 & n18127 ) | ( n5669 & n18127 ) ;
  assign n38078 = ( n5417 & n5778 ) | ( n5417 & n21303 ) | ( n5778 & n21303 ) ;
  assign n38080 = n38079 ^ n38078 ^ n31185 ;
  assign n38081 = n5732 | n27093 ;
  assign n38082 = n38081 ^ n16864 ^ 1'b0 ;
  assign n38083 = n18159 ^ n3611 ^ 1'b0 ;
  assign n38084 = n5782 ^ n1098 ^ 1'b0 ;
  assign n38085 = n675 & n38084 ;
  assign n38086 = ~n38083 & n38085 ;
  assign n38087 = n38086 ^ n34035 ^ n8394 ;
  assign n38088 = n30997 ^ n24817 ^ 1'b0 ;
  assign n38089 = ( n16710 & n29502 ) | ( n16710 & ~n38088 ) | ( n29502 & ~n38088 ) ;
  assign n38090 = ~n22178 & n38089 ;
  assign n38091 = n38090 ^ n18389 ^ 1'b0 ;
  assign n38092 = n3489 & ~n17621 ;
  assign n38093 = n26793 ^ n25419 ^ n6691 ;
  assign n38094 = n16983 ^ n2545 ^ 1'b0 ;
  assign n38095 = n10016 & n38094 ;
  assign n38096 = n11536 ^ n8083 ^ 1'b0 ;
  assign n38097 = n9647 & ~n38096 ;
  assign n38098 = n31271 ^ n12532 ^ n11006 ;
  assign n38099 = n19991 ^ n4914 ^ 1'b0 ;
  assign n38100 = ( ~n2474 & n38098 ) | ( ~n2474 & n38099 ) | ( n38098 & n38099 ) ;
  assign n38101 = n28055 ^ n27457 ^ 1'b0 ;
  assign n38102 = n35501 ^ n28348 ^ n11048 ;
  assign n38103 = ( n7411 & ~n16317 ) | ( n7411 & n38102 ) | ( ~n16317 & n38102 ) ;
  assign n38104 = ( n7209 & n10896 ) | ( n7209 & ~n38103 ) | ( n10896 & ~n38103 ) ;
  assign n38105 = n17343 ^ n9119 ^ 1'b0 ;
  assign n38106 = ( n12522 & n20423 ) | ( n12522 & ~n38105 ) | ( n20423 & ~n38105 ) ;
  assign n38107 = ( n3771 & n19045 ) | ( n3771 & n38106 ) | ( n19045 & n38106 ) ;
  assign n38108 = n4336 | n9790 ;
  assign n38109 = n38108 ^ n14228 ^ 1'b0 ;
  assign n38110 = n22668 & ~n32350 ;
  assign n38111 = ~x127 & n38110 ;
  assign n38112 = n9720 & n15262 ;
  assign n38113 = ~n25280 & n38112 ;
  assign n38114 = n27029 & n38113 ;
  assign n38115 = ( ~n1523 & n3439 ) | ( ~n1523 & n5727 ) | ( n3439 & n5727 ) ;
  assign n38116 = n7972 & ~n38115 ;
  assign n38117 = n38116 ^ n19576 ^ 1'b0 ;
  assign n38118 = n36254 ^ n34749 ^ n10856 ;
  assign n38119 = ~n31732 & n38118 ;
  assign n38120 = n38117 & n38119 ;
  assign n38121 = n32517 ^ n21139 ^ n13220 ;
  assign n38122 = ( n3955 & n26611 ) | ( n3955 & ~n38121 ) | ( n26611 & ~n38121 ) ;
  assign n38123 = n10179 | n20310 ;
  assign n38124 = n28983 ^ n2579 ^ 1'b0 ;
  assign n38125 = n8652 | n38124 ;
  assign n38126 = ( n1863 & ~n10336 ) | ( n1863 & n19494 ) | ( ~n10336 & n19494 ) ;
  assign n38127 = n25791 ^ n21049 ^ n11927 ;
  assign n38128 = n38127 ^ n24526 ^ 1'b0 ;
  assign n38129 = n18548 ^ n4328 ^ 1'b0 ;
  assign n38130 = ~n4123 & n38129 ;
  assign n38131 = ~n5590 & n21651 ;
  assign n38132 = ( n5873 & n37243 ) | ( n5873 & ~n38131 ) | ( n37243 & ~n38131 ) ;
  assign n38133 = ( n416 & n23138 ) | ( n416 & ~n38132 ) | ( n23138 & ~n38132 ) ;
  assign n38134 = n16282 & ~n38133 ;
  assign n38140 = n478 & ~n34642 ;
  assign n38139 = n19179 & n34843 ;
  assign n38138 = ( n10702 & ~n11507 ) | ( n10702 & n12592 ) | ( ~n11507 & n12592 ) ;
  assign n38141 = n38140 ^ n38139 ^ n38138 ;
  assign n38135 = ( n10285 & n24869 ) | ( n10285 & n36756 ) | ( n24869 & n36756 ) ;
  assign n38136 = n1606 | n38135 ;
  assign n38137 = ( ~n21707 & n30116 ) | ( ~n21707 & n38136 ) | ( n30116 & n38136 ) ;
  assign n38142 = n38141 ^ n38137 ^ 1'b0 ;
  assign n38143 = n26206 ^ n12151 ^ 1'b0 ;
  assign n38144 = ( n3593 & n22936 ) | ( n3593 & n38143 ) | ( n22936 & n38143 ) ;
  assign n38145 = n1974 & n19901 ;
  assign n38146 = ~n11375 & n38145 ;
  assign n38147 = n38146 ^ n34571 ^ 1'b0 ;
  assign n38148 = n5149 & n38147 ;
  assign n38149 = n38148 ^ n24938 ^ n5042 ;
  assign n38150 = n7424 | n21956 ;
  assign n38151 = n17981 | n38150 ;
  assign n38152 = n27273 ^ n24893 ^ 1'b0 ;
  assign n38153 = ~n9980 & n38152 ;
  assign n38154 = n38153 ^ n13388 ^ 1'b0 ;
  assign n38155 = ( n3234 & ~n38151 ) | ( n3234 & n38154 ) | ( ~n38151 & n38154 ) ;
  assign n38163 = n25584 ^ n603 ^ 1'b0 ;
  assign n38161 = n6562 | n21893 ;
  assign n38162 = n38161 ^ n16737 ^ 1'b0 ;
  assign n38158 = ~n6666 & n9497 ;
  assign n38159 = ~n12140 & n38158 ;
  assign n38160 = ( n19658 & ~n25940 ) | ( n19658 & n38159 ) | ( ~n25940 & n38159 ) ;
  assign n38164 = n38163 ^ n38162 ^ n38160 ;
  assign n38156 = n14095 & ~n23474 ;
  assign n38157 = n38156 ^ n23680 ^ n4145 ;
  assign n38165 = n38164 ^ n38157 ^ n352 ;
  assign n38166 = n14261 | n27270 ;
  assign n38167 = n11226 & ~n32027 ;
  assign n38168 = n38167 ^ n24953 ^ 1'b0 ;
  assign n38170 = ( ~n5816 & n10027 ) | ( ~n5816 & n10679 ) | ( n10027 & n10679 ) ;
  assign n38169 = n11286 | n22339 ;
  assign n38171 = n38170 ^ n38169 ^ 1'b0 ;
  assign n38172 = n12402 & n31566 ;
  assign n38173 = n38172 ^ n4576 ^ 1'b0 ;
  assign n38174 = n18259 & n24568 ;
  assign n38175 = ( n18072 & n18241 ) | ( n18072 & n19298 ) | ( n18241 & n19298 ) ;
  assign n38179 = n6785 & n7600 ;
  assign n38180 = n38179 ^ n5118 ^ 1'b0 ;
  assign n38181 = ( ~n10713 & n28915 ) | ( ~n10713 & n38180 ) | ( n28915 & n38180 ) ;
  assign n38178 = n2398 & ~n27410 ;
  assign n38176 = n3823 | n32042 ;
  assign n38177 = n38176 ^ n15258 ^ 1'b0 ;
  assign n38182 = n38181 ^ n38178 ^ n38177 ;
  assign n38183 = n17704 | n36823 ;
  assign n38184 = ( n15594 & ~n37696 ) | ( n15594 & n38183 ) | ( ~n37696 & n38183 ) ;
  assign n38186 = n25391 ^ n9758 ^ n7356 ;
  assign n38185 = n3546 | n19458 ;
  assign n38187 = n38186 ^ n38185 ^ 1'b0 ;
  assign n38188 = n10356 ^ n9591 ^ n701 ;
  assign n38189 = ( n1732 & ~n5382 ) | ( n1732 & n10060 ) | ( ~n5382 & n10060 ) ;
  assign n38190 = n38189 ^ n28543 ^ 1'b0 ;
  assign n38191 = n38188 & n38190 ;
  assign n38192 = n13870 ^ n7471 ^ 1'b0 ;
  assign n38193 = n930 & n7550 ;
  assign n38194 = n14515 & ~n26192 ;
  assign n38195 = n38189 ^ n14139 ^ n10696 ;
  assign n38196 = ~n8954 & n32499 ;
  assign n38197 = n17261 ^ n4649 ^ 1'b0 ;
  assign n38198 = n23744 | n38197 ;
  assign n38199 = ( n1611 & n9234 ) | ( n1611 & n12500 ) | ( n9234 & n12500 ) ;
  assign n38200 = ( n16064 & n32535 ) | ( n16064 & n38199 ) | ( n32535 & n38199 ) ;
  assign n38201 = n28780 ^ n22972 ^ 1'b0 ;
  assign n38202 = ~n9547 & n38201 ;
  assign n38203 = ( n24834 & n33524 ) | ( n24834 & ~n38202 ) | ( n33524 & ~n38202 ) ;
  assign n38204 = n38203 ^ n33109 ^ n27894 ;
  assign n38205 = ( ~n1274 & n3844 ) | ( ~n1274 & n26719 ) | ( n3844 & n26719 ) ;
  assign n38206 = ~n28702 & n38205 ;
  assign n38207 = n38206 ^ n29524 ^ 1'b0 ;
  assign n38208 = n15846 ^ n2569 ^ 1'b0 ;
  assign n38209 = ( ~n15246 & n38207 ) | ( ~n15246 & n38208 ) | ( n38207 & n38208 ) ;
  assign n38210 = ( n10007 & ~n29084 ) | ( n10007 & n30285 ) | ( ~n29084 & n30285 ) ;
  assign n38211 = ( n3083 & ~n11240 ) | ( n3083 & n38210 ) | ( ~n11240 & n38210 ) ;
  assign n38212 = n38211 ^ n1229 ^ 1'b0 ;
  assign n38213 = n38212 ^ n27052 ^ n14725 ;
  assign n38214 = n38213 ^ n22406 ^ 1'b0 ;
  assign n38215 = n21344 ^ n17504 ^ n8188 ;
  assign n38216 = ( ~n18363 & n25515 ) | ( ~n18363 & n38215 ) | ( n25515 & n38215 ) ;
  assign n38217 = n38216 ^ n18863 ^ n2533 ;
  assign n38218 = n2632 & n8135 ;
  assign n38219 = n256 & n7471 ;
  assign n38220 = n38218 & n38219 ;
  assign n38221 = n29199 ^ n24810 ^ 1'b0 ;
  assign n38222 = n31415 | n38221 ;
  assign n38225 = n8224 ^ n8045 ^ 1'b0 ;
  assign n38223 = ~n15866 & n29729 ;
  assign n38224 = ~n4521 & n38223 ;
  assign n38226 = n38225 ^ n38224 ^ n36631 ;
  assign n38227 = ( x80 & n638 ) | ( x80 & ~n33671 ) | ( n638 & ~n33671 ) ;
  assign n38228 = ( n4412 & n14803 ) | ( n4412 & ~n18131 ) | ( n14803 & ~n18131 ) ;
  assign n38229 = ( n7977 & n11404 ) | ( n7977 & ~n19545 ) | ( n11404 & ~n19545 ) ;
  assign n38230 = ( n1135 & ~n18988 ) | ( n1135 & n38229 ) | ( ~n18988 & n38229 ) ;
  assign n38231 = n38230 ^ n38028 ^ 1'b0 ;
  assign n38232 = n22618 ^ n11592 ^ n7850 ;
  assign n38233 = n14188 & ~n38232 ;
  assign n38234 = n29997 ^ n28971 ^ n7788 ;
  assign n38235 = n25423 ^ n20566 ^ 1'b0 ;
  assign n38236 = n29224 & ~n38235 ;
  assign n38237 = n11633 ^ n6767 ^ n6584 ;
  assign n38238 = n2977 & ~n20705 ;
  assign n38239 = n4446 & ~n22942 ;
  assign n38240 = n38239 ^ n9551 ^ 1'b0 ;
  assign n38241 = n38240 ^ n16181 ^ n10424 ;
  assign n38242 = n38241 ^ n7824 ^ n7239 ;
  assign n38243 = ( ~n6916 & n38238 ) | ( ~n6916 & n38242 ) | ( n38238 & n38242 ) ;
  assign n38244 = n38243 ^ n21499 ^ 1'b0 ;
  assign n38245 = n38237 & ~n38244 ;
  assign n38246 = n12127 & n19319 ;
  assign n38247 = n38246 ^ n6302 ^ 1'b0 ;
  assign n38248 = ( ~n1452 & n2841 ) | ( ~n1452 & n4951 ) | ( n2841 & n4951 ) ;
  assign n38249 = n38248 ^ n7027 ^ 1'b0 ;
  assign n38250 = n7746 & n38249 ;
  assign n38251 = ( n8103 & n26628 ) | ( n8103 & n38250 ) | ( n26628 & n38250 ) ;
  assign n38252 = ( n2179 & n10604 ) | ( n2179 & n18804 ) | ( n10604 & n18804 ) ;
  assign n38253 = n6127 ^ n2736 ^ 1'b0 ;
  assign n38254 = ( n3878 & n20450 ) | ( n3878 & n38253 ) | ( n20450 & n38253 ) ;
  assign n38255 = n20707 ^ n17369 ^ n2707 ;
  assign n38256 = ( n2117 & n3371 ) | ( n2117 & ~n29544 ) | ( n3371 & ~n29544 ) ;
  assign n38257 = n6992 | n27989 ;
  assign n38258 = n38256 & ~n38257 ;
  assign n38259 = n38255 & ~n38258 ;
  assign n38260 = n13168 & n38259 ;
  assign n38261 = n17964 ^ n4639 ^ n1823 ;
  assign n38262 = ( n7856 & ~n32646 ) | ( n7856 & n34462 ) | ( ~n32646 & n34462 ) ;
  assign n38263 = ( n12178 & ~n19163 ) | ( n12178 & n28661 ) | ( ~n19163 & n28661 ) ;
  assign n38264 = n14189 ^ n4011 ^ 1'b0 ;
  assign n38265 = ( n557 & n8040 ) | ( n557 & ~n31655 ) | ( n8040 & ~n31655 ) ;
  assign n38266 = n38265 ^ n14418 ^ 1'b0 ;
  assign n38267 = n25307 & n38266 ;
  assign n38268 = n15931 & n30776 ;
  assign n38269 = n38268 ^ n10845 ^ 1'b0 ;
  assign n38270 = n10506 & n33782 ;
  assign n38271 = ( ~n438 & n9177 ) | ( ~n438 & n21793 ) | ( n9177 & n21793 ) ;
  assign n38272 = ~n10196 & n38271 ;
  assign n38273 = ( ~n3552 & n24457 ) | ( ~n3552 & n38272 ) | ( n24457 & n38272 ) ;
  assign n38274 = n24093 ^ n23434 ^ n18778 ;
  assign n38275 = ~n14901 & n37107 ;
  assign n38276 = n38275 ^ n14348 ^ n9639 ;
  assign n38277 = n38276 ^ n35332 ^ n2475 ;
  assign n38278 = n2209 & n12820 ;
  assign n38279 = ~n3914 & n38278 ;
  assign n38280 = ~n25497 & n37219 ;
  assign n38281 = ~n3358 & n9509 ;
  assign n38282 = n38281 ^ n10854 ^ 1'b0 ;
  assign n38283 = ~n2199 & n4896 ;
  assign n38284 = ~n18169 & n38283 ;
  assign n38285 = n38284 ^ n11451 ^ 1'b0 ;
  assign n38286 = n38282 & n38285 ;
  assign n38287 = n34600 ^ n18748 ^ 1'b0 ;
  assign n38288 = n36368 ^ n17152 ^ n13087 ;
  assign n38289 = n38288 ^ n19295 ^ n10254 ;
  assign n38290 = n12924 ^ n8887 ^ 1'b0 ;
  assign n38291 = n3044 & n38290 ;
  assign n38292 = ( n15074 & ~n32853 ) | ( n15074 & n38291 ) | ( ~n32853 & n38291 ) ;
  assign n38293 = n38292 ^ n27489 ^ 1'b0 ;
  assign n38294 = n38289 | n38293 ;
  assign n38295 = ( n3864 & ~n6180 ) | ( n3864 & n12661 ) | ( ~n6180 & n12661 ) ;
  assign n38296 = n30261 ^ n1863 ^ n1848 ;
  assign n38297 = ~n22339 & n35480 ;
  assign n38298 = n38297 ^ n5554 ^ 1'b0 ;
  assign n38299 = ~n31942 & n38298 ;
  assign n38300 = ( ~n4340 & n19176 ) | ( ~n4340 & n35551 ) | ( n19176 & n35551 ) ;
  assign n38301 = ( n7019 & ~n16393 ) | ( n7019 & n25605 ) | ( ~n16393 & n25605 ) ;
  assign n38302 = ~n6728 & n37798 ;
  assign n38303 = n15648 & n38302 ;
  assign n38304 = n2859 & n15022 ;
  assign n38305 = n22210 ^ n802 ^ 1'b0 ;
  assign n38306 = ~n9005 & n38305 ;
  assign n38307 = ( ~n1644 & n28480 ) | ( ~n1644 & n38306 ) | ( n28480 & n38306 ) ;
  assign n38308 = n6420 & ~n25554 ;
  assign n38309 = ~n7382 & n38308 ;
  assign n38310 = ( n9898 & ~n13594 ) | ( n9898 & n15467 ) | ( ~n13594 & n15467 ) ;
  assign n38311 = n22032 | n38310 ;
  assign n38312 = n38311 ^ n24734 ^ 1'b0 ;
  assign n38313 = n34638 ^ n8403 ^ n3430 ;
  assign n38314 = n2993 & ~n5904 ;
  assign n38315 = n5795 ^ n1525 ^ 1'b0 ;
  assign n38319 = n25781 ^ n7387 ^ n6876 ;
  assign n38320 = n15772 ^ n4819 ^ 1'b0 ;
  assign n38321 = n38319 & ~n38320 ;
  assign n38318 = n18676 ^ n5914 ^ 1'b0 ;
  assign n38316 = n1691 | n38146 ;
  assign n38317 = n21973 & ~n38316 ;
  assign n38322 = n38321 ^ n38318 ^ n38317 ;
  assign n38323 = n32142 ^ n22102 ^ n8149 ;
  assign n38324 = n4564 ^ n4552 ^ n800 ;
  assign n38327 = n22152 ^ n17244 ^ n12764 ;
  assign n38328 = n38327 ^ n31227 ^ 1'b0 ;
  assign n38329 = n30613 & ~n38328 ;
  assign n38325 = n27270 | n37759 ;
  assign n38326 = n38325 ^ n18130 ^ 1'b0 ;
  assign n38330 = n38329 ^ n38326 ^ n34074 ;
  assign n38331 = ( n4674 & n11794 ) | ( n4674 & n36946 ) | ( n11794 & n36946 ) ;
  assign n38332 = n38242 & n38331 ;
  assign n38333 = n5749 ^ n2986 ^ 1'b0 ;
  assign n38334 = n2095 & n26904 ;
  assign n38335 = ( x46 & ~n2751 ) | ( x46 & n9873 ) | ( ~n2751 & n9873 ) ;
  assign n38336 = ( n31483 & n38334 ) | ( n31483 & ~n38335 ) | ( n38334 & ~n38335 ) ;
  assign n38337 = ( n18599 & n19786 ) | ( n18599 & n38336 ) | ( n19786 & n38336 ) ;
  assign n38338 = n21772 ^ n14572 ^ n6625 ;
  assign n38339 = ~n10627 & n20485 ;
  assign n38340 = ~n38338 & n38339 ;
  assign n38341 = n24288 ^ n21585 ^ 1'b0 ;
  assign n38342 = n36808 ^ n20047 ^ n3863 ;
  assign n38343 = n38342 ^ n33028 ^ 1'b0 ;
  assign n38344 = n6493 & n38343 ;
  assign n38345 = ( ~n10170 & n14552 ) | ( ~n10170 & n18215 ) | ( n14552 & n18215 ) ;
  assign n38346 = n38345 ^ n22010 ^ n5114 ;
  assign n38347 = ( n19142 & ~n28081 ) | ( n19142 & n30987 ) | ( ~n28081 & n30987 ) ;
  assign n38348 = ( ~n25208 & n31372 ) | ( ~n25208 & n38347 ) | ( n31372 & n38347 ) ;
  assign n38349 = n17077 ^ n1721 ^ n963 ;
  assign n38350 = n16766 & n38349 ;
  assign n38351 = n38350 ^ n14499 ^ 1'b0 ;
  assign n38352 = ( n2943 & n14841 ) | ( n2943 & n38351 ) | ( n14841 & n38351 ) ;
  assign n38353 = n38352 ^ n10138 ^ n5909 ;
  assign n38356 = ~n26730 & n36926 ;
  assign n38357 = n11582 & n38356 ;
  assign n38354 = n3867 ^ n1827 ^ x123 ;
  assign n38355 = ~n30259 & n38354 ;
  assign n38358 = n38357 ^ n38355 ^ 1'b0 ;
  assign n38359 = ~n11884 & n35406 ;
  assign n38360 = n18968 | n21033 ;
  assign n38361 = n38360 ^ n1276 ^ 1'b0 ;
  assign n38362 = n5906 & n26334 ;
  assign n38363 = n31435 ^ n30509 ^ n5076 ;
  assign n38364 = n19746 ^ n5224 ^ 1'b0 ;
  assign n38365 = n19051 | n38364 ;
  assign n38367 = ~n2826 & n9670 ;
  assign n38368 = ~n31339 & n38367 ;
  assign n38366 = n9216 & n28542 ;
  assign n38369 = n38368 ^ n38366 ^ 1'b0 ;
  assign n38370 = n38365 & n38369 ;
  assign n38371 = ( n19635 & ~n38363 ) | ( n19635 & n38370 ) | ( ~n38363 & n38370 ) ;
  assign n38372 = ~n3174 & n21904 ;
  assign n38373 = n19626 & n38372 ;
  assign n38374 = n38373 ^ n6491 ^ 1'b0 ;
  assign n38375 = n38374 ^ n22354 ^ 1'b0 ;
  assign n38376 = n10896 | n38375 ;
  assign n38377 = n38376 ^ n22505 ^ n9121 ;
  assign n38384 = n893 & n9490 ;
  assign n38380 = n30415 ^ n20318 ^ n11273 ;
  assign n38381 = ~n3969 & n38380 ;
  assign n38382 = n24698 & n38381 ;
  assign n38383 = ( n25396 & n35609 ) | ( n25396 & n38382 ) | ( n35609 & n38382 ) ;
  assign n38378 = n7354 & ~n23859 ;
  assign n38379 = n38378 ^ n22545 ^ 1'b0 ;
  assign n38385 = n38384 ^ n38383 ^ n38379 ;
  assign n38386 = n24008 ^ n16720 ^ 1'b0 ;
  assign n38387 = n38386 ^ n18284 ^ n6848 ;
  assign n38388 = n19518 ^ n15037 ^ n6986 ;
  assign n38389 = n15708 ^ n4327 ^ 1'b0 ;
  assign n38390 = n38388 | n38389 ;
  assign n38391 = n20766 ^ n16877 ^ n2574 ;
  assign n38392 = n35252 ^ n7843 ^ 1'b0 ;
  assign n38393 = ( n7317 & n13661 ) | ( n7317 & ~n38392 ) | ( n13661 & ~n38392 ) ;
  assign n38394 = n32456 ^ n19357 ^ 1'b0 ;
  assign n38395 = n36983 ^ n8201 ^ 1'b0 ;
  assign n38396 = n23376 & n38395 ;
  assign n38397 = n8456 & n38396 ;
  assign n38398 = ~n29640 & n38397 ;
  assign n38399 = n16140 & n37434 ;
  assign n38400 = n38399 ^ n27033 ^ 1'b0 ;
  assign n38401 = n38400 ^ n15246 ^ 1'b0 ;
  assign n38402 = ( x236 & n5622 ) | ( x236 & n38401 ) | ( n5622 & n38401 ) ;
  assign n38403 = n37258 ^ n5996 ^ 1'b0 ;
  assign n38404 = ~n2769 & n16832 ;
  assign n38405 = n38404 ^ n4350 ^ 1'b0 ;
  assign n38406 = ~n7405 & n38405 ;
  assign n38407 = n38406 ^ n8260 ^ 1'b0 ;
  assign n38408 = ~n19202 & n38407 ;
  assign n38409 = ( n2012 & ~n10165 ) | ( n2012 & n13344 ) | ( ~n10165 & n13344 ) ;
  assign n38410 = ( n494 & n8686 ) | ( n494 & ~n8888 ) | ( n8686 & ~n8888 ) ;
  assign n38411 = ( n13493 & n21001 ) | ( n13493 & n38410 ) | ( n21001 & n38410 ) ;
  assign n38412 = n18410 | n38272 ;
  assign n38413 = n38412 ^ n21181 ^ n12160 ;
  assign n38414 = ( ~n18077 & n26742 ) | ( ~n18077 & n38413 ) | ( n26742 & n38413 ) ;
  assign n38415 = n2712 & ~n12461 ;
  assign n38416 = ~n346 & n38415 ;
  assign n38418 = n30251 ^ n20130 ^ n12788 ;
  assign n38417 = n10233 | n23196 ;
  assign n38419 = n38418 ^ n38417 ^ 1'b0 ;
  assign n38420 = ( ~n24834 & n38416 ) | ( ~n24834 & n38419 ) | ( n38416 & n38419 ) ;
  assign n38421 = n33856 ^ n22906 ^ 1'b0 ;
  assign n38422 = n11762 ^ x130 ^ 1'b0 ;
  assign n38423 = n345 & n2100 ;
  assign n38424 = ~n7470 & n38423 ;
  assign n38425 = n18843 ^ n8180 ^ 1'b0 ;
  assign n38426 = n38425 ^ n2590 ^ 1'b0 ;
  assign n38427 = n1537 & ~n38426 ;
  assign n38429 = n26220 ^ n22243 ^ n19068 ;
  assign n38428 = n25888 ^ n7686 ^ n6990 ;
  assign n38430 = n38429 ^ n38428 ^ 1'b0 ;
  assign n38431 = ~n15856 & n38430 ;
  assign n38432 = ( n38424 & n38427 ) | ( n38424 & ~n38431 ) | ( n38427 & ~n38431 ) ;
  assign n38434 = n25565 ^ n14269 ^ 1'b0 ;
  assign n38433 = n12593 & n17874 ;
  assign n38435 = n38434 ^ n38433 ^ n16330 ;
  assign n38436 = n817 & ~n28204 ;
  assign n38437 = ~n33923 & n35135 ;
  assign n38438 = ~n4720 & n11178 ;
  assign n38439 = n26645 ^ n12740 ^ 1'b0 ;
  assign n38440 = n14670 & ~n38439 ;
  assign n38441 = n11674 & ~n17520 ;
  assign n38442 = n38441 ^ n15467 ^ 1'b0 ;
  assign n38443 = ( n3983 & n31165 ) | ( n3983 & ~n38442 ) | ( n31165 & ~n38442 ) ;
  assign n38444 = ( ~n811 & n38440 ) | ( ~n811 & n38443 ) | ( n38440 & n38443 ) ;
  assign n38445 = ( n7500 & ~n38438 ) | ( n7500 & n38444 ) | ( ~n38438 & n38444 ) ;
  assign n38446 = n38445 ^ n24603 ^ n2204 ;
  assign n38447 = n19718 & ~n27302 ;
  assign n38448 = n38447 ^ n7189 ^ 1'b0 ;
  assign n38449 = n18473 ^ n14290 ^ 1'b0 ;
  assign n38450 = ~n14960 & n38449 ;
  assign n38451 = n38450 ^ n20013 ^ n3549 ;
  assign n38452 = n27465 ^ n8508 ^ n7638 ;
  assign n38453 = n38452 ^ n38283 ^ n1876 ;
  assign n38454 = n38453 ^ n14870 ^ n14625 ;
  assign n38455 = n9072 & ~n12244 ;
  assign n38456 = n14992 | n38455 ;
  assign n38457 = n26720 ^ n15153 ^ 1'b0 ;
  assign n38458 = n20369 ^ n2791 ^ n640 ;
  assign n38459 = n38458 ^ n1640 ^ 1'b0 ;
  assign n38460 = n33973 ^ n30727 ^ n18441 ;
  assign n38461 = n38460 ^ n21524 ^ x205 ;
  assign n38462 = ( n2913 & ~n17824 ) | ( n2913 & n19117 ) | ( ~n17824 & n19117 ) ;
  assign n38463 = n38462 ^ n3476 ^ n911 ;
  assign n38464 = n4654 & n13451 ;
  assign n38465 = n29972 & n38464 ;
  assign n38466 = n31591 ^ n31177 ^ n4746 ;
  assign n38467 = n27758 ^ n13823 ^ 1'b0 ;
  assign n38468 = ~n38466 & n38467 ;
  assign n38469 = n1867 & n11515 ;
  assign n38470 = n38469 ^ n13664 ^ 1'b0 ;
  assign n38471 = ~n5054 & n7268 ;
  assign n38472 = n38471 ^ n19829 ^ 1'b0 ;
  assign n38473 = n15148 ^ n8682 ^ n937 ;
  assign n38474 = n25939 ^ n10712 ^ 1'b0 ;
  assign n38475 = n3775 & ~n38474 ;
  assign n38476 = ( n12339 & n23892 ) | ( n12339 & n38475 ) | ( n23892 & n38475 ) ;
  assign n38477 = ~n31977 & n38476 ;
  assign n38478 = n21290 ^ n3522 ^ 1'b0 ;
  assign n38479 = n7620 | n38478 ;
  assign n38480 = n38479 ^ n13126 ^ 1'b0 ;
  assign n38481 = n38477 & n38480 ;
  assign n38482 = ( n14396 & n30844 ) | ( n14396 & n38481 ) | ( n30844 & n38481 ) ;
  assign n38483 = n38482 ^ n8881 ^ n6849 ;
  assign n38484 = n9140 & n26812 ;
  assign n38485 = n5069 & n38484 ;
  assign n38486 = n38485 ^ n23826 ^ 1'b0 ;
  assign n38487 = ~n19639 & n38486 ;
  assign n38488 = n38487 ^ n4245 ^ 1'b0 ;
  assign n38489 = n25188 & ~n38488 ;
  assign n38490 = n14880 | n31633 ;
  assign n38491 = n25833 ^ n24188 ^ n14330 ;
  assign n38492 = n3699 | n5541 ;
  assign n38493 = n38492 ^ n4950 ^ 1'b0 ;
  assign n38494 = n18252 & ~n38493 ;
  assign n38495 = n10671 ^ n8970 ^ n2847 ;
  assign n38496 = ~n6134 & n38495 ;
  assign n38497 = n38494 & n38496 ;
  assign n38498 = n1974 & ~n32459 ;
  assign n38499 = n38498 ^ n3111 ^ 1'b0 ;
  assign n38500 = ( ~n16501 & n27779 ) | ( ~n16501 & n38499 ) | ( n27779 & n38499 ) ;
  assign n38501 = ( n4726 & n22853 ) | ( n4726 & n38500 ) | ( n22853 & n38500 ) ;
  assign n38502 = n36130 ^ n8718 ^ 1'b0 ;
  assign n38503 = ~n38501 & n38502 ;
  assign n38504 = ( n4846 & ~n13836 ) | ( n4846 & n25318 ) | ( ~n13836 & n25318 ) ;
  assign n38505 = ~n6615 & n38504 ;
  assign n38506 = n38505 ^ n35872 ^ 1'b0 ;
  assign n38507 = ( n6434 & n9213 ) | ( n6434 & ~n38506 ) | ( n9213 & ~n38506 ) ;
  assign n38509 = n15573 ^ n6677 ^ 1'b0 ;
  assign n38510 = n10426 & n38509 ;
  assign n38508 = ( n16497 & n19348 ) | ( n16497 & n25512 ) | ( n19348 & n25512 ) ;
  assign n38511 = n38510 ^ n38508 ^ 1'b0 ;
  assign n38512 = ( ~n14098 & n37357 ) | ( ~n14098 & n38511 ) | ( n37357 & n38511 ) ;
  assign n38513 = ( n27188 & n27600 ) | ( n27188 & n36056 ) | ( n27600 & n36056 ) ;
  assign n38514 = ( n1232 & ~n11848 ) | ( n1232 & n14113 ) | ( ~n11848 & n14113 ) ;
  assign n38515 = n38514 ^ n8398 ^ n3674 ;
  assign n38516 = n38515 ^ n28546 ^ n12042 ;
  assign n38517 = ( n11554 & n38513 ) | ( n11554 & n38516 ) | ( n38513 & n38516 ) ;
  assign n38518 = n32226 ^ n28545 ^ n1714 ;
  assign n38519 = n6831 & n38518 ;
  assign n38520 = n8094 & n38519 ;
  assign n38521 = n18999 & ~n32405 ;
  assign n38522 = ( n5842 & ~n27399 ) | ( n5842 & n32734 ) | ( ~n27399 & n32734 ) ;
  assign n38523 = n5272 & n25867 ;
  assign n38524 = n38522 & n38523 ;
  assign n38525 = n27420 & ~n37370 ;
  assign n38527 = ~n3606 & n6528 ;
  assign n38528 = n38527 ^ n6469 ^ 1'b0 ;
  assign n38529 = ( ~n12684 & n29913 ) | ( ~n12684 & n38528 ) | ( n29913 & n38528 ) ;
  assign n38530 = n38529 ^ n33883 ^ 1'b0 ;
  assign n38526 = n1054 & n25824 ;
  assign n38531 = n38530 ^ n38526 ^ n33958 ;
  assign n38532 = n21487 ^ n9084 ^ 1'b0 ;
  assign n38533 = n19095 | n38532 ;
  assign n38534 = n4053 & ~n14980 ;
  assign n38535 = ~n38533 & n38534 ;
  assign n38536 = n38535 ^ n17713 ^ n9664 ;
  assign n38537 = n18120 ^ n11509 ^ n3567 ;
  assign n38538 = ( n14908 & n38536 ) | ( n14908 & n38537 ) | ( n38536 & n38537 ) ;
  assign n38539 = ( ~n10263 & n15739 ) | ( ~n10263 & n21788 ) | ( n15739 & n21788 ) ;
  assign n38540 = n20371 | n38539 ;
  assign n38541 = n21403 ^ n11253 ^ n1523 ;
  assign n38542 = n37619 ^ n8984 ^ n966 ;
  assign n38543 = x103 & ~n10673 ;
  assign n38544 = n17041 ^ n8457 ^ n4824 ;
  assign n38545 = n312 & ~n905 ;
  assign n38546 = n38545 ^ n16317 ^ 1'b0 ;
  assign n38547 = n38546 ^ n38140 ^ n5714 ;
  assign n38548 = n1261 & ~n34508 ;
  assign n38549 = n24555 & n38548 ;
  assign n38550 = n24192 ^ n7586 ^ n1295 ;
  assign n38551 = ( n9576 & n20724 ) | ( n9576 & ~n20753 ) | ( n20724 & ~n20753 ) ;
  assign n38552 = n7482 & n10547 ;
  assign n38553 = ( n19361 & n21890 ) | ( n19361 & n38552 ) | ( n21890 & n38552 ) ;
  assign n38556 = ~n2288 & n9593 ;
  assign n38557 = n38556 ^ n13760 ^ 1'b0 ;
  assign n38554 = n14875 & n17012 ;
  assign n38555 = n24488 & n38554 ;
  assign n38558 = n38557 ^ n38555 ^ n14370 ;
  assign n38559 = n38558 ^ n31937 ^ n2146 ;
  assign n38560 = n26599 ^ n13039 ^ 1'b0 ;
  assign n38561 = n12540 ^ n9041 ^ 1'b0 ;
  assign n38562 = n15008 | n38561 ;
  assign n38563 = n38562 ^ n16529 ^ 1'b0 ;
  assign n38564 = n9277 & n38563 ;
  assign n38565 = n13129 ^ n536 ^ 1'b0 ;
  assign n38566 = n11086 & n38565 ;
  assign n38567 = n14451 ^ n4415 ^ 1'b0 ;
  assign n38568 = n20537 & n38567 ;
  assign n38570 = n21448 ^ n11757 ^ n5500 ;
  assign n38571 = n38570 ^ n37613 ^ n6370 ;
  assign n38572 = ( n2864 & ~n9021 ) | ( n2864 & n38571 ) | ( ~n9021 & n38571 ) ;
  assign n38569 = n18598 & n35612 ;
  assign n38573 = n38572 ^ n38569 ^ 1'b0 ;
  assign n38574 = n2717 ^ n1394 ^ 1'b0 ;
  assign n38575 = n38574 ^ n29611 ^ n325 ;
  assign n38576 = n38575 ^ n2594 ^ 1'b0 ;
  assign n38577 = n23536 ^ n12606 ^ n2002 ;
  assign n38581 = ~n1905 & n18467 ;
  assign n38578 = n8372 & n10760 ;
  assign n38579 = n38450 & ~n38578 ;
  assign n38580 = n38579 ^ n15845 ^ 1'b0 ;
  assign n38582 = n38581 ^ n38580 ^ n5171 ;
  assign n38583 = n37089 ^ n32273 ^ n24308 ;
  assign n38584 = ( n2610 & n9340 ) | ( n2610 & ~n11360 ) | ( n9340 & ~n11360 ) ;
  assign n38585 = n38584 ^ n23600 ^ 1'b0 ;
  assign n38586 = n13869 & n23164 ;
  assign n38587 = n5408 & ~n29931 ;
  assign n38588 = n38586 & n38587 ;
  assign n38589 = ( n17013 & n21582 ) | ( n17013 & n22670 ) | ( n21582 & n22670 ) ;
  assign n38590 = n28587 & n38589 ;
  assign n38591 = n37353 ^ n14613 ^ 1'b0 ;
  assign n38592 = ~n12697 & n38591 ;
  assign n38593 = ( n32734 & ~n38537 ) | ( n32734 & n38592 ) | ( ~n38537 & n38592 ) ;
  assign n38594 = ~n17584 & n22361 ;
  assign n38595 = n38594 ^ n16481 ^ x228 ;
  assign n38596 = ( n2338 & n5729 ) | ( n2338 & ~n13725 ) | ( n5729 & ~n13725 ) ;
  assign n38597 = n21917 & n23897 ;
  assign n38598 = n18722 | n22068 ;
  assign n38599 = n38598 ^ n703 ^ 1'b0 ;
  assign n38600 = n26424 & ~n34446 ;
  assign n38601 = n38599 & n38600 ;
  assign n38602 = n6026 | n38601 ;
  assign n38603 = ( n12485 & ~n23039 ) | ( n12485 & n29976 ) | ( ~n23039 & n29976 ) ;
  assign n38604 = n38603 ^ n8510 ^ n3965 ;
  assign n38605 = ( n1050 & ~n18462 ) | ( n1050 & n38604 ) | ( ~n18462 & n38604 ) ;
  assign n38606 = n13340 & n17936 ;
  assign n38607 = n38606 ^ n21078 ^ n19497 ;
  assign n38608 = ( ~n1760 & n10062 ) | ( ~n1760 & n15484 ) | ( n10062 & n15484 ) ;
  assign n38609 = ( ~n576 & n33458 ) | ( ~n576 & n38608 ) | ( n33458 & n38608 ) ;
  assign n38610 = n425 & ~n23267 ;
  assign n38611 = n38610 ^ n31152 ^ 1'b0 ;
  assign n38612 = ( n5806 & n21346 ) | ( n5806 & ~n38611 ) | ( n21346 & ~n38611 ) ;
  assign n38613 = n38612 ^ n35525 ^ n32251 ;
  assign n38614 = n21196 ^ x245 ^ 1'b0 ;
  assign n38615 = n19558 | n38614 ;
  assign n38616 = ( n4556 & n18429 ) | ( n4556 & ~n38615 ) | ( n18429 & ~n38615 ) ;
  assign n38617 = n19600 ^ n2657 ^ 1'b0 ;
  assign n38618 = ~n18746 & n38617 ;
  assign n38619 = n38618 ^ n2988 ^ 1'b0 ;
  assign n38620 = ~n35442 & n38619 ;
  assign n38621 = n15106 ^ n5064 ^ 1'b0 ;
  assign n38622 = ~n811 & n38621 ;
  assign n38623 = n10318 & ~n11823 ;
  assign n38624 = ~n15689 & n38623 ;
  assign n38625 = n38622 & ~n38624 ;
  assign n38626 = n38625 ^ n14956 ^ 1'b0 ;
  assign n38627 = n1747 | n29004 ;
  assign n38628 = n16971 ^ n13672 ^ 1'b0 ;
  assign n38629 = n13312 & n38628 ;
  assign n38630 = n38629 ^ n21170 ^ n8648 ;
  assign n38631 = ( ~n16047 & n18255 ) | ( ~n16047 & n38630 ) | ( n18255 & n38630 ) ;
  assign n38632 = n15575 ^ n2735 ^ 1'b0 ;
  assign n38633 = n753 & ~n38632 ;
  assign n38634 = ~n38631 & n38633 ;
  assign n38635 = ~n33572 & n38634 ;
  assign n38636 = n15494 & ~n38635 ;
  assign n38637 = n23112 ^ n20246 ^ 1'b0 ;
  assign n38638 = n33315 ^ n31603 ^ n395 ;
  assign n38639 = ( n2773 & n24373 ) | ( n2773 & n38638 ) | ( n24373 & n38638 ) ;
  assign n38640 = ( n37203 & n38637 ) | ( n37203 & n38639 ) | ( n38637 & n38639 ) ;
  assign n38641 = n38336 ^ n13097 ^ n6362 ;
  assign n38642 = n14847 ^ n7892 ^ 1'b0 ;
  assign n38643 = ~n9669 & n16587 ;
  assign n38644 = n36218 & n38643 ;
  assign n38645 = n38644 ^ n30248 ^ 1'b0 ;
  assign n38646 = n38002 ^ n26236 ^ 1'b0 ;
  assign n38647 = ~n24083 & n38646 ;
  assign n38648 = n14312 & ~n20582 ;
  assign n38649 = n5999 | n38648 ;
  assign n38650 = n6376 | n38649 ;
  assign n38651 = n12670 ^ n12122 ^ n6328 ;
  assign n38652 = n27756 ^ n10327 ^ 1'b0 ;
  assign n38653 = n38651 & ~n38652 ;
  assign n38654 = n21724 ^ n7535 ^ 1'b0 ;
  assign n38655 = n5433 ^ n2602 ^ 1'b0 ;
  assign n38656 = n38655 ^ n26322 ^ n6347 ;
  assign n38657 = n13792 ^ n10136 ^ 1'b0 ;
  assign n38659 = ( x99 & n3999 ) | ( x99 & ~n10550 ) | ( n3999 & ~n10550 ) ;
  assign n38658 = n2809 | n4635 ;
  assign n38660 = n38659 ^ n38658 ^ 1'b0 ;
  assign n38663 = n26767 | n30045 ;
  assign n38661 = ~n18654 & n25835 ;
  assign n38662 = n38661 ^ n11188 ^ n4359 ;
  assign n38664 = n38663 ^ n38662 ^ n6815 ;
  assign n38665 = n4434 & ~n38664 ;
  assign n38666 = n34107 ^ n21047 ^ n7072 ;
  assign n38667 = n38666 ^ n29966 ^ n6311 ;
  assign n38668 = n12601 & ~n12909 ;
  assign n38669 = ( n1010 & n19480 ) | ( n1010 & ~n29939 ) | ( n19480 & ~n29939 ) ;
  assign n38670 = ( ~n2220 & n4532 ) | ( ~n2220 & n35747 ) | ( n4532 & n35747 ) ;
  assign n38671 = n38670 ^ n33954 ^ 1'b0 ;
  assign n38672 = n4349 | n25396 ;
  assign n38673 = n38672 ^ n4348 ^ 1'b0 ;
  assign n38674 = n1508 & n38673 ;
  assign n38675 = n38674 ^ n36076 ^ 1'b0 ;
  assign n38676 = n28352 ^ n27719 ^ n16376 ;
  assign n38677 = n7737 ^ n5996 ^ n3838 ;
  assign n38678 = n38677 ^ n11995 ^ n1160 ;
  assign n38682 = n3743 ^ n1644 ^ 1'b0 ;
  assign n38683 = n17467 & n38682 ;
  assign n38684 = n5424 & n38683 ;
  assign n38679 = n2187 & n17061 ;
  assign n38680 = n22843 ^ n3379 ^ 1'b0 ;
  assign n38681 = n38679 & ~n38680 ;
  assign n38685 = n38684 ^ n38681 ^ n16846 ;
  assign n38686 = ( n5835 & ~n12017 ) | ( n5835 & n32988 ) | ( ~n12017 & n32988 ) ;
  assign n38687 = x80 & ~n13063 ;
  assign n38688 = ~n33681 & n38687 ;
  assign n38689 = n38688 ^ n18345 ^ n11016 ;
  assign n38690 = ~n34959 & n38689 ;
  assign n38692 = n8132 ^ n4821 ^ 1'b0 ;
  assign n38693 = n38608 & ~n38692 ;
  assign n38691 = n36531 ^ n20516 ^ 1'b0 ;
  assign n38694 = n38693 ^ n38691 ^ n17321 ;
  assign n38695 = n38694 ^ n20368 ^ 1'b0 ;
  assign n38696 = n27101 | n38695 ;
  assign n38697 = n19391 ^ n11708 ^ n5123 ;
  assign n38698 = ~n16613 & n20975 ;
  assign n38699 = ~n38697 & n38698 ;
  assign n38700 = n2863 & n21556 ;
  assign n38701 = n26257 ^ n17396 ^ n10057 ;
  assign n38702 = n24996 ^ n3552 ^ 1'b0 ;
  assign n38703 = n7163 & ~n38702 ;
  assign n38704 = ~n18187 & n38703 ;
  assign n38705 = n38704 ^ n9217 ^ 1'b0 ;
  assign n38706 = n14415 | n38705 ;
  assign n38707 = n5973 | n17035 ;
  assign n38708 = n38707 ^ n26618 ^ n4197 ;
  assign n38712 = n26591 ^ n16954 ^ n1099 ;
  assign n38709 = n18151 ^ n17415 ^ n9756 ;
  assign n38710 = n1558 & ~n38709 ;
  assign n38711 = ~n11237 & n38710 ;
  assign n38713 = n38712 ^ n38711 ^ n26703 ;
  assign n38714 = ( n12146 & n25578 ) | ( n12146 & ~n38713 ) | ( n25578 & ~n38713 ) ;
  assign n38715 = n38714 ^ n27683 ^ n24266 ;
  assign n38716 = ( n6850 & ~n23192 ) | ( n6850 & n29963 ) | ( ~n23192 & n29963 ) ;
  assign n38717 = ( ~n16376 & n23516 ) | ( ~n16376 & n32453 ) | ( n23516 & n32453 ) ;
  assign n38718 = ( ~n12311 & n23324 ) | ( ~n12311 & n38717 ) | ( n23324 & n38717 ) ;
  assign n38719 = n3136 & n38718 ;
  assign n38720 = n35078 ^ n26275 ^ 1'b0 ;
  assign n38721 = ( x167 & n15605 ) | ( x167 & n38720 ) | ( n15605 & n38720 ) ;
  assign n38724 = ( n3002 & n5002 ) | ( n3002 & ~n18047 ) | ( n5002 & ~n18047 ) ;
  assign n38722 = n3886 & ~n10669 ;
  assign n38723 = ~n10355 & n38722 ;
  assign n38725 = n38724 ^ n38723 ^ n2845 ;
  assign n38726 = ( n1189 & n35456 ) | ( n1189 & ~n38725 ) | ( n35456 & ~n38725 ) ;
  assign n38727 = n4547 & ~n17588 ;
  assign n38728 = n38727 ^ n9711 ^ n9235 ;
  assign n38729 = n35531 ^ n23614 ^ 1'b0 ;
  assign n38730 = n19405 | n27376 ;
  assign n38731 = n38730 ^ n24976 ^ 1'b0 ;
  assign n38732 = n19360 | n38731 ;
  assign n38733 = ( n27776 & n38729 ) | ( n27776 & n38732 ) | ( n38729 & n38732 ) ;
  assign n38736 = n8299 ^ n6350 ^ n4042 ;
  assign n38737 = n38736 ^ n25052 ^ n9013 ;
  assign n38734 = n13638 | n22690 ;
  assign n38735 = n38734 ^ n9478 ^ 1'b0 ;
  assign n38738 = n38737 ^ n38735 ^ n33885 ;
  assign n38739 = n9655 & ~n13335 ;
  assign n38740 = n38739 ^ n29454 ^ 1'b0 ;
  assign n38741 = n11885 & n23095 ;
  assign n38742 = ( n1637 & n19552 ) | ( n1637 & n20987 ) | ( n19552 & n20987 ) ;
  assign n38743 = n11901 ^ n4501 ^ n971 ;
  assign n38746 = n8257 | n21082 ;
  assign n38747 = n15458 | n38746 ;
  assign n38744 = ( n3892 & ~n11037 ) | ( n3892 & n17761 ) | ( ~n11037 & n17761 ) ;
  assign n38745 = ( ~n3124 & n4309 ) | ( ~n3124 & n38744 ) | ( n4309 & n38744 ) ;
  assign n38748 = n38747 ^ n38745 ^ n16548 ;
  assign n38749 = n1032 & ~n37086 ;
  assign n38750 = n31307 | n37419 ;
  assign n38751 = n9279 | n15050 ;
  assign n38752 = n38751 ^ n33383 ^ n2701 ;
  assign n38753 = n38752 ^ n16494 ^ 1'b0 ;
  assign n38754 = n38753 ^ n34298 ^ 1'b0 ;
  assign n38755 = ( x1 & n6570 ) | ( x1 & ~n7747 ) | ( n6570 & ~n7747 ) ;
  assign n38756 = ( n25448 & ~n37607 ) | ( n25448 & n38755 ) | ( ~n37607 & n38755 ) ;
  assign n38757 = n1334 | n3211 ;
  assign n38758 = n13149 & n22382 ;
  assign n38759 = ( n25970 & n38757 ) | ( n25970 & ~n38758 ) | ( n38757 & ~n38758 ) ;
  assign n38760 = n38759 ^ n17750 ^ n10400 ;
  assign n38761 = n37559 ^ n21757 ^ 1'b0 ;
  assign n38762 = n25412 & ~n38761 ;
  assign n38763 = ~n1447 & n23677 ;
  assign n38764 = n38763 ^ n16359 ^ 1'b0 ;
  assign n38765 = n3935 & n38764 ;
  assign n38766 = ~n12487 & n22933 ;
  assign n38767 = n38766 ^ n9520 ^ 1'b0 ;
  assign n38768 = n16568 ^ n11525 ^ 1'b0 ;
  assign n38769 = ( n910 & ~n13335 ) | ( n910 & n13926 ) | ( ~n13335 & n13926 ) ;
  assign n38770 = n38769 ^ n17167 ^ n12623 ;
  assign n38771 = n38770 ^ n14698 ^ 1'b0 ;
  assign n38772 = x203 & ~n10269 ;
  assign n38773 = n38772 ^ n35286 ^ 1'b0 ;
  assign n38774 = n38773 ^ n3896 ^ 1'b0 ;
  assign n38776 = n22702 ^ n14305 ^ 1'b0 ;
  assign n38775 = n8806 & n9454 ;
  assign n38777 = n38776 ^ n38775 ^ n2242 ;
  assign n38778 = n13226 ^ n10870 ^ 1'b0 ;
  assign n38779 = ~n8637 & n38778 ;
  assign n38780 = ( n3160 & ~n35858 ) | ( n3160 & n38779 ) | ( ~n35858 & n38779 ) ;
  assign n38781 = ( n676 & n26374 ) | ( n676 & n38780 ) | ( n26374 & n38780 ) ;
  assign n38782 = ( n816 & n28141 ) | ( n816 & ~n38781 ) | ( n28141 & ~n38781 ) ;
  assign n38783 = ( n6817 & ~n13216 ) | ( n6817 & n38782 ) | ( ~n13216 & n38782 ) ;
  assign n38787 = n10174 | n34400 ;
  assign n38788 = n38787 ^ n29727 ^ 1'b0 ;
  assign n38784 = ( n6851 & ~n7485 ) | ( n6851 & n13278 ) | ( ~n7485 & n13278 ) ;
  assign n38785 = n16353 & ~n38784 ;
  assign n38786 = ~n10774 & n38785 ;
  assign n38789 = n38788 ^ n38786 ^ n26520 ;
  assign n38790 = n2230 & n7428 ;
  assign n38791 = ~n26763 & n38790 ;
  assign n38793 = ( n1288 & n3468 ) | ( n1288 & n4626 ) | ( n3468 & n4626 ) ;
  assign n38794 = n2829 | n37449 ;
  assign n38795 = n38793 & ~n38794 ;
  assign n38792 = n5556 | n11898 ;
  assign n38796 = n38795 ^ n38792 ^ 1'b0 ;
  assign n38797 = n6537 & ~n21309 ;
  assign n38798 = n4307 ^ n2401 ^ 1'b0 ;
  assign n38799 = ( n8861 & n31323 ) | ( n8861 & n38798 ) | ( n31323 & n38798 ) ;
  assign n38800 = n38799 ^ n16306 ^ 1'b0 ;
  assign n38801 = n36839 ^ n7407 ^ n7274 ;
  assign n38802 = ( n4615 & n17062 ) | ( n4615 & n38801 ) | ( n17062 & n38801 ) ;
  assign n38803 = n19860 | n38802 ;
  assign n38804 = n14730 & ~n38803 ;
  assign n38805 = n1544 & n38804 ;
  assign n38806 = ( ~n1384 & n13665 ) | ( ~n1384 & n31200 ) | ( n13665 & n31200 ) ;
  assign n38809 = n28044 | n33960 ;
  assign n38810 = n5755 & ~n38809 ;
  assign n38811 = ~n7700 & n12712 ;
  assign n38812 = ( n4397 & n38810 ) | ( n4397 & ~n38811 ) | ( n38810 & ~n38811 ) ;
  assign n38807 = n15906 | n28777 ;
  assign n38808 = n2934 & n38807 ;
  assign n38813 = n38812 ^ n38808 ^ 1'b0 ;
  assign n38814 = n24943 | n31083 ;
  assign n38815 = n38814 ^ n13168 ^ 1'b0 ;
  assign n38816 = n11450 & n29843 ;
  assign n38817 = ( n25248 & ~n29747 ) | ( n25248 & n32482 ) | ( ~n29747 & n32482 ) ;
  assign n38818 = n8955 & ~n9392 ;
  assign n38819 = n38818 ^ n33966 ^ 1'b0 ;
  assign n38820 = n38819 ^ n27078 ^ n3762 ;
  assign n38821 = n16268 ^ n3083 ^ 1'b0 ;
  assign n38822 = ~n23604 & n38821 ;
  assign n38823 = n38578 ^ n1644 ^ x42 ;
  assign n38824 = n23232 & n30811 ;
  assign n38825 = n20807 & n38824 ;
  assign n38826 = n24645 ^ n1330 ^ 1'b0 ;
  assign n38827 = n38124 & n38826 ;
  assign n38828 = n11994 ^ n5847 ^ n5619 ;
  assign n38829 = ( n22942 & ~n24248 ) | ( n22942 & n38828 ) | ( ~n24248 & n38828 ) ;
  assign n38832 = n6543 ^ n1230 ^ n1153 ;
  assign n38830 = n8856 ^ n8063 ^ 1'b0 ;
  assign n38831 = n23824 & n38830 ;
  assign n38833 = n38832 ^ n38831 ^ 1'b0 ;
  assign n38834 = n30843 ^ n30433 ^ n15246 ;
  assign n38835 = n31461 ^ n6226 ^ 1'b0 ;
  assign n38836 = n38835 ^ n15828 ^ 1'b0 ;
  assign n38837 = ~n38834 & n38836 ;
  assign n38838 = n32302 ^ n6983 ^ n5961 ;
  assign n38839 = n38838 ^ n3459 ^ 1'b0 ;
  assign n38840 = n15804 ^ n5156 ^ 1'b0 ;
  assign n38841 = ~n6650 & n6813 ;
  assign n38842 = ~n12441 & n38841 ;
  assign n38843 = ~n929 & n34071 ;
  assign n38844 = ~n17407 & n29112 ;
  assign n38845 = n38844 ^ n6337 ^ 1'b0 ;
  assign n38846 = n25442 ^ n23070 ^ n10506 ;
  assign n38847 = n22687 ^ n6328 ^ 1'b0 ;
  assign n38848 = n38846 & ~n38847 ;
  assign n38849 = n29261 ^ n2898 ^ 1'b0 ;
  assign n38850 = n38848 & ~n38849 ;
  assign n38851 = n38850 ^ n16237 ^ n2036 ;
  assign n38853 = n9948 & ~n24509 ;
  assign n38854 = n5623 & n38853 ;
  assign n38852 = n8484 | n12083 ;
  assign n38855 = n38854 ^ n38852 ^ 1'b0 ;
  assign n38856 = n1482 & ~n34029 ;
  assign n38857 = n8341 & n38856 ;
  assign n38858 = n31243 ^ n24659 ^ n8384 ;
  assign n38859 = n17274 ^ n11541 ^ n2353 ;
  assign n38865 = n9739 ^ n6483 ^ n6267 ;
  assign n38864 = ~n10155 & n27275 ;
  assign n38866 = n38865 ^ n38864 ^ 1'b0 ;
  assign n38867 = n18986 & ~n38866 ;
  assign n38860 = n29045 ^ n2898 ^ 1'b0 ;
  assign n38861 = n24120 | n38860 ;
  assign n38862 = n9833 & ~n38861 ;
  assign n38863 = ~n28016 & n38862 ;
  assign n38868 = n38867 ^ n38863 ^ n6946 ;
  assign n38869 = ~n38859 & n38868 ;
  assign n38870 = ~n38858 & n38869 ;
  assign n38871 = n4356 | n15798 ;
  assign n38872 = n11261 & ~n38871 ;
  assign n38873 = n38872 ^ n17540 ^ n3235 ;
  assign n38874 = ~n36897 & n38873 ;
  assign n38875 = n7364 ^ n4621 ^ 1'b0 ;
  assign n38876 = ~n12621 & n38875 ;
  assign n38877 = n8341 | n38876 ;
  assign n38878 = n35611 ^ n33614 ^ n8649 ;
  assign n38880 = n6806 & ~n10561 ;
  assign n38879 = n22633 ^ n19523 ^ n3065 ;
  assign n38881 = n38880 ^ n38879 ^ n15157 ;
  assign n38882 = n22977 ^ n6157 ^ 1'b0 ;
  assign n38883 = n10042 | n36934 ;
  assign n38884 = n38883 ^ n23414 ^ 1'b0 ;
  assign n38885 = n14516 ^ n9052 ^ n2085 ;
  assign n38886 = n38885 ^ n10343 ^ n6164 ;
  assign n38887 = n38886 ^ n28494 ^ 1'b0 ;
  assign n38888 = n6499 & n38887 ;
  assign n38889 = n38888 ^ n28886 ^ 1'b0 ;
  assign n38890 = ( n10214 & n19995 ) | ( n10214 & ~n38889 ) | ( n19995 & ~n38889 ) ;
  assign n38891 = ( ~n2500 & n18623 ) | ( ~n2500 & n37507 ) | ( n18623 & n37507 ) ;
  assign n38892 = n10606 ^ n8796 ^ 1'b0 ;
  assign n38893 = n14046 & n38892 ;
  assign n38894 = n26983 ^ n16072 ^ n2512 ;
  assign n38895 = n20117 | n38894 ;
  assign n38896 = n38895 ^ n33401 ^ 1'b0 ;
  assign n38897 = n6913 | n14172 ;
  assign n38898 = n38897 ^ n30963 ^ 1'b0 ;
  assign n38899 = ( n38893 & n38896 ) | ( n38893 & n38898 ) | ( n38896 & n38898 ) ;
  assign n38900 = ( n4336 & ~n8768 ) | ( n4336 & n30301 ) | ( ~n8768 & n30301 ) ;
  assign n38901 = n15505 & n17322 ;
  assign n38902 = n11076 ^ n2424 ^ 1'b0 ;
  assign n38903 = n3430 & n38902 ;
  assign n38904 = ~n9118 & n38903 ;
  assign n38905 = ( n4115 & n27081 ) | ( n4115 & ~n38904 ) | ( n27081 & ~n38904 ) ;
  assign n38906 = n37331 ^ n1740 ^ 1'b0 ;
  assign n38907 = n3716 | n30160 ;
  assign n38908 = n38906 | n38907 ;
  assign n38909 = n20422 ^ n19918 ^ n16066 ;
  assign n38910 = ( ~n3151 & n7874 ) | ( ~n3151 & n21517 ) | ( n7874 & n21517 ) ;
  assign n38911 = n38909 & n38910 ;
  assign n38912 = n29921 & n38911 ;
  assign n38913 = ~n8468 & n20037 ;
  assign n38914 = n1573 & n38913 ;
  assign n38915 = n38914 ^ n23047 ^ n9361 ;
  assign n38916 = ( n12414 & n31389 ) | ( n12414 & ~n38915 ) | ( n31389 & ~n38915 ) ;
  assign n38917 = ( ~x58 & n2085 ) | ( ~x58 & n17735 ) | ( n2085 & n17735 ) ;
  assign n38918 = n34235 ^ n4569 ^ 1'b0 ;
  assign n38919 = n38918 ^ n32533 ^ n19393 ;
  assign n38920 = n38919 ^ n38405 ^ n28495 ;
  assign n38921 = ~n3626 & n17845 ;
  assign n38922 = n16236 & n38921 ;
  assign n38923 = ( ~n4542 & n18487 ) | ( ~n4542 & n37840 ) | ( n18487 & n37840 ) ;
  assign n38924 = n24110 ^ n20841 ^ n8326 ;
  assign n38925 = ~n9427 & n31417 ;
  assign n38926 = n2272 & n38925 ;
  assign n38930 = n5671 ^ n3069 ^ n1293 ;
  assign n38927 = n3704 & ~n5864 ;
  assign n38928 = ~n19844 & n38927 ;
  assign n38929 = n38928 ^ n19112 ^ n5155 ;
  assign n38931 = n38930 ^ n38929 ^ n25486 ;
  assign n38932 = ~n1524 & n38931 ;
  assign n38933 = ~n13848 & n38932 ;
  assign n38934 = n3588 | n15277 ;
  assign n38935 = n38933 & ~n38934 ;
  assign n38936 = n8181 & ~n25921 ;
  assign n38937 = ( n17787 & n38935 ) | ( n17787 & ~n38936 ) | ( n38935 & ~n38936 ) ;
  assign n38938 = n26039 & n26076 ;
  assign n38939 = ( n736 & n22577 ) | ( n736 & n25984 ) | ( n22577 & n25984 ) ;
  assign n38940 = n38939 ^ n35006 ^ n12908 ;
  assign n38941 = n4645 & n37507 ;
  assign n38942 = ~n8286 & n38941 ;
  assign n38943 = n15855 & ~n20106 ;
  assign n38944 = n31963 & n38943 ;
  assign n38945 = n12573 & n30148 ;
  assign n38946 = n38945 ^ n6875 ^ 1'b0 ;
  assign n38947 = n31120 ^ n18392 ^ n5549 ;
  assign n38948 = ( n5548 & n25948 ) | ( n5548 & n38947 ) | ( n25948 & n38947 ) ;
  assign n38949 = n38948 ^ n6299 ^ 1'b0 ;
  assign n38950 = n24967 & ~n38949 ;
  assign n38951 = ( n4179 & ~n38946 ) | ( n4179 & n38950 ) | ( ~n38946 & n38950 ) ;
  assign n38952 = n18701 | n38951 ;
  assign n38953 = n22646 ^ n12694 ^ n3484 ;
  assign n38954 = n17246 ^ n14992 ^ n5742 ;
  assign n38955 = n7683 ^ n4920 ^ 1'b0 ;
  assign n38956 = ~n17391 & n38955 ;
  assign n38957 = ( ~n13390 & n22138 ) | ( ~n13390 & n33992 ) | ( n22138 & n33992 ) ;
  assign n38958 = n36574 ^ n603 ^ 1'b0 ;
  assign n38959 = ~n38957 & n38958 ;
  assign n38960 = n9115 & ~n12744 ;
  assign n38961 = n38960 ^ n27125 ^ 1'b0 ;
  assign n38963 = n15134 & n22621 ;
  assign n38964 = n26045 & n38963 ;
  assign n38962 = n585 & ~n17107 ;
  assign n38965 = n38964 ^ n38962 ^ 1'b0 ;
  assign n38966 = n3536 & ~n25585 ;
  assign n38967 = ( n16497 & ~n36991 ) | ( n16497 & n38966 ) | ( ~n36991 & n38966 ) ;
  assign n38968 = n25316 ^ n12213 ^ n2192 ;
  assign n38969 = n1899 & ~n12290 ;
  assign n38970 = n24822 & n38969 ;
  assign n38971 = n24293 ^ n10597 ^ 1'b0 ;
  assign n38972 = n7907 & ~n38971 ;
  assign n38973 = ~n26003 & n26266 ;
  assign n38974 = n38973 ^ n1390 ^ 1'b0 ;
  assign n38975 = ( ~x72 & n10461 ) | ( ~x72 & n18221 ) | ( n10461 & n18221 ) ;
  assign n38976 = n38975 ^ n32995 ^ 1'b0 ;
  assign n38977 = ~n22393 & n38976 ;
  assign n38978 = n2376 ^ n1876 ^ 1'b0 ;
  assign n38979 = n4771 & ~n38978 ;
  assign n38980 = n38979 ^ n18377 ^ 1'b0 ;
  assign n38981 = n29553 ^ n17079 ^ n4495 ;
  assign n38982 = n38980 & n38981 ;
  assign n38984 = n12427 | n14707 ;
  assign n38985 = n38984 ^ n13142 ^ 1'b0 ;
  assign n38983 = n4920 | n6856 ;
  assign n38986 = n38985 ^ n38983 ^ x153 ;
  assign n38987 = n38986 ^ n34822 ^ n517 ;
  assign n38988 = n12618 | n21761 ;
  assign n38989 = n38988 ^ n31895 ^ 1'b0 ;
  assign n38990 = n38989 ^ n16656 ^ n329 ;
  assign n38991 = n38990 ^ n11114 ^ n7434 ;
  assign n38992 = ( n3530 & ~n29896 ) | ( n3530 & n35895 ) | ( ~n29896 & n35895 ) ;
  assign n38993 = n36137 ^ n22591 ^ n8592 ;
  assign n38994 = n38993 ^ n25406 ^ n6289 ;
  assign n38997 = n2064 | n16423 ;
  assign n38995 = x242 & ~n32089 ;
  assign n38996 = n38995 ^ n6492 ^ 1'b0 ;
  assign n38998 = n38997 ^ n38996 ^ n16272 ;
  assign n38999 = x146 & n32646 ;
  assign n39000 = n9066 & n10094 ;
  assign n39001 = n2993 & n39000 ;
  assign n39002 = n39001 ^ n37765 ^ 1'b0 ;
  assign n39003 = n12848 & ~n39002 ;
  assign n39004 = n11094 ^ n6998 ^ n2838 ;
  assign n39005 = n29271 | n39004 ;
  assign n39006 = ~n3494 & n6963 ;
  assign n39007 = n39006 ^ x42 ^ 1'b0 ;
  assign n39008 = n39007 ^ n24108 ^ 1'b0 ;
  assign n39009 = n9977 & n39008 ;
  assign n39010 = ( ~n15304 & n19712 ) | ( ~n15304 & n28818 ) | ( n19712 & n28818 ) ;
  assign n39011 = n27842 ^ n9205 ^ n4191 ;
  assign n39012 = ( ~n10155 & n18823 ) | ( ~n10155 & n26477 ) | ( n18823 & n26477 ) ;
  assign n39013 = ~n39011 & n39012 ;
  assign n39014 = n4535 ^ n3945 ^ n2110 ;
  assign n39015 = n39014 ^ n13987 ^ 1'b0 ;
  assign n39016 = ~n31266 & n39015 ;
  assign n39017 = n37705 ^ n36346 ^ 1'b0 ;
  assign n39018 = n18508 ^ n10876 ^ n397 ;
  assign n39019 = n39018 ^ n33315 ^ n20117 ;
  assign n39020 = ( ~n4469 & n10801 ) | ( ~n4469 & n24251 ) | ( n10801 & n24251 ) ;
  assign n39021 = ( n7497 & n28067 ) | ( n7497 & ~n39020 ) | ( n28067 & ~n39020 ) ;
  assign n39022 = ( n497 & ~n8357 ) | ( n497 & n19674 ) | ( ~n8357 & n19674 ) ;
  assign n39023 = n39022 ^ n14432 ^ n6620 ;
  assign n39024 = n10115 | n39023 ;
  assign n39025 = n10822 ^ n9642 ^ 1'b0 ;
  assign n39026 = n39025 ^ n1427 ^ 1'b0 ;
  assign n39027 = ~n279 & n6399 ;
  assign n39031 = n29965 ^ n29674 ^ 1'b0 ;
  assign n39032 = n7463 & ~n39031 ;
  assign n39029 = n2301 & ~n3148 ;
  assign n39030 = n39029 ^ n23574 ^ 1'b0 ;
  assign n39028 = ( n18308 & n22106 ) | ( n18308 & ~n24057 ) | ( n22106 & ~n24057 ) ;
  assign n39033 = n39032 ^ n39030 ^ n39028 ;
  assign n39035 = ( n1760 & n4807 ) | ( n1760 & n7843 ) | ( n4807 & n7843 ) ;
  assign n39034 = n7354 ^ n7116 ^ n1200 ;
  assign n39036 = n39035 ^ n39034 ^ n24413 ;
  assign n39037 = ( ~n15974 & n19117 ) | ( ~n15974 & n39036 ) | ( n19117 & n39036 ) ;
  assign n39038 = n39037 ^ n20709 ^ 1'b0 ;
  assign n39039 = n39033 & ~n39038 ;
  assign n39040 = n9677 | n16487 ;
  assign n39041 = n39040 ^ n17864 ^ 1'b0 ;
  assign n39042 = n39041 ^ n727 ^ 1'b0 ;
  assign n39043 = n19602 | n39042 ;
  assign n39044 = n20109 | n31594 ;
  assign n39045 = n5960 | n19111 ;
  assign n39046 = n13469 & ~n39045 ;
  assign n39047 = n27446 | n39046 ;
  assign n39048 = n39044 | n39047 ;
  assign n39049 = ( n11777 & n23072 ) | ( n11777 & n35099 ) | ( n23072 & n35099 ) ;
  assign n39050 = n31826 ^ n23888 ^ n5864 ;
  assign n39051 = n39050 ^ n19918 ^ n6915 ;
  assign n39052 = n39051 ^ n9260 ^ 1'b0 ;
  assign n39053 = ( n17858 & ~n18483 ) | ( n17858 & n30375 ) | ( ~n18483 & n30375 ) ;
  assign n39054 = n26498 ^ n23586 ^ 1'b0 ;
  assign n39055 = ( n9486 & n17129 ) | ( n9486 & ~n39054 ) | ( n17129 & ~n39054 ) ;
  assign n39056 = n29304 ^ n1877 ^ 1'b0 ;
  assign n39057 = n10060 ^ n7896 ^ 1'b0 ;
  assign n39058 = n27983 | n39057 ;
  assign n39059 = ~n16752 & n27206 ;
  assign n39060 = n39059 ^ n13405 ^ 1'b0 ;
  assign n39061 = n26128 | n28798 ;
  assign n39062 = n39061 ^ n19774 ^ 1'b0 ;
  assign n39063 = n22148 ^ n13900 ^ 1'b0 ;
  assign n39064 = n29597 | n29691 ;
  assign n39065 = n39064 ^ n1916 ^ 1'b0 ;
  assign n39066 = n39065 ^ n13665 ^ n10659 ;
  assign n39067 = ~n5006 & n29946 ;
  assign n39068 = n1049 & n39067 ;
  assign n39069 = n36197 & ~n39068 ;
  assign n39070 = n37432 ^ n16465 ^ 1'b0 ;
  assign n39071 = ~n17078 & n39070 ;
  assign n39072 = n36120 ^ n12542 ^ 1'b0 ;
  assign n39073 = n6025 & n39072 ;
  assign n39074 = ( n1547 & n27746 ) | ( n1547 & ~n30963 ) | ( n27746 & ~n30963 ) ;
  assign n39075 = ( n362 & ~n3200 ) | ( n362 & n5753 ) | ( ~n3200 & n5753 ) ;
  assign n39076 = n39075 ^ n34625 ^ n23074 ;
  assign n39077 = n526 & ~n13192 ;
  assign n39078 = ~n11640 & n39077 ;
  assign n39079 = n39078 ^ n13649 ^ n4375 ;
  assign n39080 = n14961 & ~n39079 ;
  assign n39081 = n32098 ^ n14580 ^ 1'b0 ;
  assign n39082 = ~n8701 & n8891 ;
  assign n39083 = n39082 ^ n8955 ^ 1'b0 ;
  assign n39084 = ( n21639 & n31991 ) | ( n21639 & n39083 ) | ( n31991 & n39083 ) ;
  assign n39085 = n12813 ^ n2036 ^ 1'b0 ;
  assign n39086 = n2274 & n20709 ;
  assign n39087 = n16395 & n39086 ;
  assign n39088 = n11816 | n28006 ;
  assign n39089 = n28006 & ~n39088 ;
  assign n39090 = n13198 | n36835 ;
  assign n39091 = n11351 & ~n33294 ;
  assign n39092 = ( n13654 & n21116 ) | ( n13654 & ~n39091 ) | ( n21116 & ~n39091 ) ;
  assign n39093 = n9177 ^ n9056 ^ n8002 ;
  assign n39094 = n17635 & n39093 ;
  assign n39095 = n19717 ^ n13581 ^ n1967 ;
  assign n39096 = ( n10415 & n11526 ) | ( n10415 & ~n21462 ) | ( n11526 & ~n21462 ) ;
  assign n39097 = n39096 ^ n5994 ^ 1'b0 ;
  assign n39098 = n20291 | n39097 ;
  assign n39099 = n28303 ^ n12469 ^ n9852 ;
  assign n39100 = n39099 ^ n6926 ^ n979 ;
  assign n39101 = n39100 ^ n36724 ^ n4506 ;
  assign n39102 = n17405 & n28957 ;
  assign n39103 = n39101 & n39102 ;
  assign n39104 = n12216 & ~n13085 ;
  assign n39105 = n39104 ^ n9125 ^ 1'b0 ;
  assign n39106 = n39105 ^ n33284 ^ 1'b0 ;
  assign n39107 = n17710 & ~n39106 ;
  assign n39108 = ( n17880 & n23965 ) | ( n17880 & ~n32150 ) | ( n23965 & ~n32150 ) ;
  assign n39109 = ( n6903 & n7355 ) | ( n6903 & ~n7719 ) | ( n7355 & ~n7719 ) ;
  assign n39110 = n39109 ^ n2097 ^ 1'b0 ;
  assign n39111 = n29231 & n36829 ;
  assign n39112 = n4566 & n39111 ;
  assign n39113 = n39112 ^ n18498 ^ n3784 ;
  assign n39114 = n12136 ^ n10395 ^ 1'b0 ;
  assign n39115 = n5218 | n39114 ;
  assign n39116 = n39115 ^ n5468 ^ 1'b0 ;
  assign n39117 = n36169 ^ n10112 ^ 1'b0 ;
  assign n39118 = ~n16163 & n39117 ;
  assign n39119 = n5855 & ~n7025 ;
  assign n39120 = ~n3746 & n4426 ;
  assign n39121 = n39120 ^ n8792 ^ 1'b0 ;
  assign n39125 = n37201 ^ n8508 ^ n2155 ;
  assign n39122 = n28640 ^ n6151 ^ 1'b0 ;
  assign n39123 = n32479 & n39122 ;
  assign n39124 = n39123 ^ n24169 ^ n4801 ;
  assign n39126 = n39125 ^ n39124 ^ 1'b0 ;
  assign n39127 = n39121 | n39126 ;
  assign n39128 = n39127 ^ n5769 ^ 1'b0 ;
  assign n39131 = n10561 ^ n5068 ^ 1'b0 ;
  assign n39129 = ~n2575 & n17839 ;
  assign n39130 = n39129 ^ n7539 ^ 1'b0 ;
  assign n39132 = n39131 ^ n39130 ^ n4612 ;
  assign n39133 = ( n29546 & n34154 ) | ( n29546 & n39132 ) | ( n34154 & n39132 ) ;
  assign n39134 = n21888 & ~n39133 ;
  assign n39135 = ( ~n667 & n19009 ) | ( ~n667 & n24546 ) | ( n19009 & n24546 ) ;
  assign n39136 = ( ~n4572 & n38694 ) | ( ~n4572 & n39135 ) | ( n38694 & n39135 ) ;
  assign n39139 = n30101 ^ n16327 ^ n5708 ;
  assign n39137 = n31879 ^ n7627 ^ n3877 ;
  assign n39138 = ( n1901 & ~n4720 ) | ( n1901 & n39137 ) | ( ~n4720 & n39137 ) ;
  assign n39140 = n39139 ^ n39138 ^ n13722 ;
  assign n39141 = n39140 ^ n35501 ^ n30127 ;
  assign n39142 = n36538 ^ n20207 ^ n7572 ;
  assign n39143 = n20214 & n29044 ;
  assign n39144 = n19770 ^ n10928 ^ 1'b0 ;
  assign n39145 = n11730 ^ n7788 ^ 1'b0 ;
  assign n39146 = n39144 | n39145 ;
  assign n39147 = n39146 ^ n8074 ^ 1'b0 ;
  assign n39148 = ~n13949 & n39147 ;
  assign n39150 = ( ~n8632 & n15780 ) | ( ~n8632 & n34125 ) | ( n15780 & n34125 ) ;
  assign n39149 = ~n13353 & n13806 ;
  assign n39151 = n39150 ^ n39149 ^ 1'b0 ;
  assign n39152 = ( ~n11218 & n15831 ) | ( ~n11218 & n39151 ) | ( n15831 & n39151 ) ;
  assign n39153 = ( n6041 & n21790 ) | ( n6041 & ~n28552 ) | ( n21790 & ~n28552 ) ;
  assign n39154 = n7798 & ~n11009 ;
  assign n39155 = n39154 ^ n22944 ^ 1'b0 ;
  assign n39156 = n9873 | n39155 ;
  assign n39157 = ( n7863 & n10379 ) | ( n7863 & n39156 ) | ( n10379 & n39156 ) ;
  assign n39163 = ~n1224 & n5326 ;
  assign n39164 = ~n2963 & n39163 ;
  assign n39160 = ( ~n3333 & n6045 ) | ( ~n3333 & n8256 ) | ( n6045 & n8256 ) ;
  assign n39158 = ( n3439 & ~n6100 ) | ( n3439 & n6575 ) | ( ~n6100 & n6575 ) ;
  assign n39159 = ~n5295 & n39158 ;
  assign n39161 = n39160 ^ n39159 ^ 1'b0 ;
  assign n39162 = n5752 & ~n39161 ;
  assign n39165 = n39164 ^ n39162 ^ n3653 ;
  assign n39166 = ( n9201 & n21661 ) | ( n9201 & n39165 ) | ( n21661 & n39165 ) ;
  assign n39169 = n14469 ^ n7195 ^ n4488 ;
  assign n39170 = n39169 ^ n16306 ^ 1'b0 ;
  assign n39171 = ~n12703 & n39170 ;
  assign n39167 = ( x7 & n1545 ) | ( x7 & ~n12742 ) | ( n1545 & ~n12742 ) ;
  assign n39168 = n1289 | n39167 ;
  assign n39172 = n39171 ^ n39168 ^ 1'b0 ;
  assign n39173 = n39172 ^ n36684 ^ 1'b0 ;
  assign n39174 = n4584 | n39173 ;
  assign n39176 = n14939 ^ n6149 ^ 1'b0 ;
  assign n39175 = n7004 & n7347 ;
  assign n39177 = n39176 ^ n39175 ^ 1'b0 ;
  assign n39178 = ( n1461 & ~n7411 ) | ( n1461 & n33826 ) | ( ~n7411 & n33826 ) ;
  assign n39179 = n36137 ^ n12885 ^ n6727 ;
  assign n39180 = n7842 | n39179 ;
  assign n39183 = n7786 & n10405 ;
  assign n39181 = ~n28867 & n29471 ;
  assign n39182 = n39181 ^ n37694 ^ n11167 ;
  assign n39184 = n39183 ^ n39182 ^ 1'b0 ;
  assign n39185 = ( n2737 & ~n25836 ) | ( n2737 & n29454 ) | ( ~n25836 & n29454 ) ;
  assign n39186 = n17299 & ~n28661 ;
  assign n39187 = n2706 & ~n6160 ;
  assign n39188 = n8779 & n39187 ;
  assign n39189 = n13148 | n39188 ;
  assign n39190 = n39189 ^ n16074 ^ n12303 ;
  assign n39191 = ~n2360 & n39190 ;
  assign n39192 = n39109 ^ n15186 ^ n5300 ;
  assign n39193 = ( n8288 & ~n12640 ) | ( n8288 & n33188 ) | ( ~n12640 & n33188 ) ;
  assign n39194 = n37191 ^ n2625 ^ 1'b0 ;
  assign n39195 = n1629 | n9823 ;
  assign n39196 = n26724 & ~n39195 ;
  assign n39197 = n13323 ^ n10690 ^ 1'b0 ;
  assign n39198 = n17214 & n39197 ;
  assign n39199 = x128 & ~n27664 ;
  assign n39200 = ~n12667 & n39199 ;
  assign n39201 = n1897 | n39200 ;
  assign n39202 = n39198 | n39201 ;
  assign n39203 = n2525 & n21481 ;
  assign n39204 = n39203 ^ n12231 ^ 1'b0 ;
  assign n39205 = ( n14150 & n20926 ) | ( n14150 & n39204 ) | ( n20926 & n39204 ) ;
  assign n39206 = n38705 ^ n38452 ^ n1186 ;
  assign n39207 = ( ~n35674 & n39205 ) | ( ~n35674 & n39206 ) | ( n39205 & n39206 ) ;
  assign n39208 = n22951 ^ n9580 ^ n7558 ;
  assign n39209 = ( ~n22876 & n23965 ) | ( ~n22876 & n39208 ) | ( n23965 & n39208 ) ;
  assign n39210 = n33272 & ~n39209 ;
  assign n39215 = n24166 ^ n22638 ^ n6300 ;
  assign n39216 = ( ~n12109 & n36514 ) | ( ~n12109 & n39215 ) | ( n36514 & n39215 ) ;
  assign n39211 = n16397 ^ n7843 ^ x114 ;
  assign n39212 = ~n10820 & n12515 ;
  assign n39213 = ( ~n8250 & n22962 ) | ( ~n8250 & n35227 ) | ( n22962 & n35227 ) ;
  assign n39214 = ( n39211 & n39212 ) | ( n39211 & n39213 ) | ( n39212 & n39213 ) ;
  assign n39217 = n39216 ^ n39214 ^ n2791 ;
  assign n39218 = ( n15976 & n24379 ) | ( n15976 & ~n39217 ) | ( n24379 & ~n39217 ) ;
  assign n39219 = n11638 & n24676 ;
  assign n39220 = n32601 ^ n3520 ^ 1'b0 ;
  assign n39221 = n12792 & ~n39220 ;
  assign n39222 = n30570 & ~n33442 ;
  assign n39223 = n25912 & ~n29243 ;
  assign n39224 = n11846 & n39223 ;
  assign n39225 = n29914 | n39224 ;
  assign n39226 = n39225 ^ n26039 ^ 1'b0 ;
  assign n39227 = n15562 ^ n12772 ^ n3322 ;
  assign n39228 = ( n5444 & n7362 ) | ( n5444 & n39227 ) | ( n7362 & n39227 ) ;
  assign n39229 = ~n5710 & n39228 ;
  assign n39234 = ( n4818 & ~n5943 ) | ( n4818 & n7491 ) | ( ~n5943 & n7491 ) ;
  assign n39230 = n1395 | n30899 ;
  assign n39231 = n39230 ^ n4714 ^ 1'b0 ;
  assign n39232 = n39231 ^ n8198 ^ n2495 ;
  assign n39233 = ( n11994 & ~n17998 ) | ( n11994 & n39232 ) | ( ~n17998 & n39232 ) ;
  assign n39235 = n39234 ^ n39233 ^ n2171 ;
  assign n39236 = ( n529 & n10931 ) | ( n529 & ~n30749 ) | ( n10931 & ~n30749 ) ;
  assign n39237 = n26059 | n39236 ;
  assign n39238 = n39237 ^ n1891 ^ 1'b0 ;
  assign n39239 = n39238 ^ n38782 ^ 1'b0 ;
  assign n39240 = n37168 ^ n34806 ^ n26222 ;
  assign n39241 = n8691 & n34453 ;
  assign n39242 = ( n22134 & n22861 ) | ( n22134 & ~n39241 ) | ( n22861 & ~n39241 ) ;
  assign n39243 = ( n1011 & ~n9816 ) | ( n1011 & n39242 ) | ( ~n9816 & n39242 ) ;
  assign n39244 = ~n5645 & n25643 ;
  assign n39245 = n39244 ^ n5197 ^ 1'b0 ;
  assign n39246 = n13134 & ~n15338 ;
  assign n39247 = n27109 & n39246 ;
  assign n39248 = n7110 & ~n35481 ;
  assign n39249 = n5245 & n39248 ;
  assign n39250 = n39249 ^ n12471 ^ 1'b0 ;
  assign n39251 = n20976 ^ n19263 ^ n9468 ;
  assign n39252 = n36583 ^ n9479 ^ 1'b0 ;
  assign n39253 = n10336 ^ n5562 ^ 1'b0 ;
  assign n39254 = n8947 & ~n39253 ;
  assign n39255 = ~n26773 & n39254 ;
  assign n39256 = n16684 & n39255 ;
  assign n39257 = n29820 ^ n20594 ^ n11733 ;
  assign n39258 = ( n13461 & ~n27072 ) | ( n13461 & n39257 ) | ( ~n27072 & n39257 ) ;
  assign n39259 = n39258 ^ n35741 ^ 1'b0 ;
  assign n39260 = n31982 ^ n11997 ^ n6051 ;
  assign n39261 = ( n4376 & ~n17069 ) | ( n4376 & n39260 ) | ( ~n17069 & n39260 ) ;
  assign n39262 = ( n25740 & ~n38493 ) | ( n25740 & n39261 ) | ( ~n38493 & n39261 ) ;
  assign n39263 = ~n15444 & n21428 ;
  assign n39264 = n39263 ^ n12682 ^ 1'b0 ;
  assign n39265 = n39264 ^ n21367 ^ n1633 ;
  assign n39268 = n15422 ^ n2637 ^ n2191 ;
  assign n39266 = n31180 ^ n21049 ^ n9290 ;
  assign n39267 = n5046 & n39266 ;
  assign n39269 = n39268 ^ n39267 ^ 1'b0 ;
  assign n39270 = n39269 ^ n24517 ^ 1'b0 ;
  assign n39271 = n24453 & ~n39270 ;
  assign n39272 = n29575 ^ n12943 ^ 1'b0 ;
  assign n39273 = n5271 | n39272 ;
  assign n39274 = n39273 ^ n20190 ^ n18481 ;
  assign n39275 = n8147 & n39274 ;
  assign n39276 = n39275 ^ n3604 ^ 1'b0 ;
  assign n39277 = ~n23617 & n27408 ;
  assign n39278 = n39277 ^ n15914 ^ 1'b0 ;
  assign n39279 = ~n16602 & n39278 ;
  assign n39280 = n39279 ^ n23112 ^ n5383 ;
  assign n39281 = n8995 ^ n4660 ^ 1'b0 ;
  assign n39282 = n4783 | n39281 ;
  assign n39283 = n9385 & ~n26070 ;
  assign n39284 = ~n16730 & n39283 ;
  assign n39285 = n4339 | n34355 ;
  assign n39286 = n39284 & ~n39285 ;
  assign n39287 = n10795 | n29711 ;
  assign n39288 = n14663 ^ x200 ^ 1'b0 ;
  assign n39289 = n36094 | n39288 ;
  assign n39290 = n15508 | n39289 ;
  assign n39291 = n39290 ^ n20464 ^ n5809 ;
  assign n39292 = n29164 ^ n4533 ^ 1'b0 ;
  assign n39293 = n7627 & ~n39292 ;
  assign n39294 = ~n10782 & n16290 ;
  assign n39295 = n32312 ^ n19811 ^ n9968 ;
  assign n39296 = n1184 ^ n736 ^ x34 ;
  assign n39297 = n23512 ^ n23331 ^ n15687 ;
  assign n39298 = n39296 & n39297 ;
  assign n39299 = n39295 & n39298 ;
  assign n39300 = ( n5028 & ~n39294 ) | ( n5028 & n39299 ) | ( ~n39294 & n39299 ) ;
  assign n39301 = ~n852 & n4477 ;
  assign n39302 = ( n7445 & ~n31529 ) | ( n7445 & n39301 ) | ( ~n31529 & n39301 ) ;
  assign n39304 = n1643 & n5259 ;
  assign n39305 = n28721 & n39304 ;
  assign n39306 = n39305 ^ n20253 ^ n509 ;
  assign n39303 = ~n1274 & n25735 ;
  assign n39307 = n39306 ^ n39303 ^ 1'b0 ;
  assign n39308 = n27372 ^ n26148 ^ 1'b0 ;
  assign n39309 = n38062 | n39308 ;
  assign n39310 = n3440 | n21480 ;
  assign n39311 = ( n13913 & ~n20200 ) | ( n13913 & n39310 ) | ( ~n20200 & n39310 ) ;
  assign n39312 = n15014 & ~n19566 ;
  assign n39313 = n10687 & n18894 ;
  assign n39314 = n39313 ^ n31193 ^ 1'b0 ;
  assign n39315 = n39314 ^ n38357 ^ n19831 ;
  assign n39316 = n3160 & n39315 ;
  assign n39317 = ( n18843 & n23465 ) | ( n18843 & ~n24772 ) | ( n23465 & ~n24772 ) ;
  assign n39318 = n8090 ^ n6679 ^ n1881 ;
  assign n39319 = n39318 ^ n19026 ^ n8842 ;
  assign n39320 = ~n13353 & n39319 ;
  assign n39321 = n34515 & n39320 ;
  assign n39322 = n39321 ^ n2592 ^ 1'b0 ;
  assign n39323 = n39322 ^ n25063 ^ n18235 ;
  assign n39324 = ~n13041 & n39323 ;
  assign n39325 = ~n34456 & n39324 ;
  assign n39326 = n8561 & n14136 ;
  assign n39327 = n38521 ^ n3151 ^ 1'b0 ;
  assign n39328 = n8489 ^ n4221 ^ n1531 ;
  assign n39329 = n39328 ^ n35841 ^ n5044 ;
  assign n39330 = n29103 ^ n26919 ^ 1'b0 ;
  assign n39335 = ( n6440 & n15431 ) | ( n6440 & ~n36304 ) | ( n15431 & ~n36304 ) ;
  assign n39332 = n9523 ^ n494 ^ 1'b0 ;
  assign n39331 = n35566 ^ n30372 ^ 1'b0 ;
  assign n39333 = n39332 ^ n39331 ^ n933 ;
  assign n39334 = n35304 & ~n39333 ;
  assign n39336 = n39335 ^ n39334 ^ 1'b0 ;
  assign n39337 = n39336 ^ n10108 ^ n9431 ;
  assign n39342 = ~n2250 & n11802 ;
  assign n39338 = ~n4399 & n9548 ;
  assign n39339 = n39338 ^ n4243 ^ 1'b0 ;
  assign n39340 = n14071 ^ n12063 ^ n4422 ;
  assign n39341 = ( n11912 & n39339 ) | ( n11912 & n39340 ) | ( n39339 & n39340 ) ;
  assign n39343 = n39342 ^ n39341 ^ n20062 ;
  assign n39344 = n13063 | n17112 ;
  assign n39345 = n2997 & ~n20549 ;
  assign n39346 = ~n2193 & n25585 ;
  assign n39347 = n24544 & n39346 ;
  assign n39348 = n13381 & n15263 ;
  assign n39349 = n15211 ^ n13693 ^ n2948 ;
  assign n39350 = ( n15029 & n23729 ) | ( n15029 & n39349 ) | ( n23729 & n39349 ) ;
  assign n39351 = ( n301 & n21101 ) | ( n301 & n24220 ) | ( n21101 & n24220 ) ;
  assign n39352 = ~n15130 & n37535 ;
  assign n39353 = ( n18464 & n34736 ) | ( n18464 & n39352 ) | ( n34736 & n39352 ) ;
  assign n39354 = n4580 & ~n36541 ;
  assign n39355 = n18860 ^ n1666 ^ 1'b0 ;
  assign n39356 = ~n1890 & n39355 ;
  assign n39357 = n11607 ^ n729 ^ x132 ;
  assign n39358 = n36191 & ~n39357 ;
  assign n39359 = n28936 & n39358 ;
  assign n39360 = n10310 & n15454 ;
  assign n39361 = n4024 & n39360 ;
  assign n39362 = n30329 ^ n26638 ^ 1'b0 ;
  assign n39363 = n933 & n39362 ;
  assign n39364 = n32687 & n39363 ;
  assign n39365 = n4348 & ~n7088 ;
  assign n39366 = ~n12394 & n39365 ;
  assign n39367 = n39366 ^ n2779 ^ 1'b0 ;
  assign n39368 = n39367 ^ x8 ^ 1'b0 ;
  assign n39369 = x145 | n32444 ;
  assign n39370 = ( n36612 & ~n37181 ) | ( n36612 & n39369 ) | ( ~n37181 & n39369 ) ;
  assign n39371 = n36645 ^ n21310 ^ n10779 ;
  assign n39372 = n8150 ^ n7452 ^ 1'b0 ;
  assign n39373 = ( n2190 & n33356 ) | ( n2190 & n39372 ) | ( n33356 & n39372 ) ;
  assign n39374 = ( n3492 & ~n9295 ) | ( n3492 & n28589 ) | ( ~n9295 & n28589 ) ;
  assign n39375 = n4158 & n21257 ;
  assign n39376 = n19813 & n28722 ;
  assign n39377 = n39376 ^ n11960 ^ 1'b0 ;
  assign n39378 = n2365 & n13161 ;
  assign n39379 = ~n28546 & n39378 ;
  assign n39380 = n6051 & n39379 ;
  assign n39381 = n19341 | n36011 ;
  assign n39382 = ( n15050 & n18996 ) | ( n15050 & ~n21110 ) | ( n18996 & ~n21110 ) ;
  assign n39383 = ( n25003 & ~n33955 ) | ( n25003 & n39382 ) | ( ~n33955 & n39382 ) ;
  assign n39384 = n6010 | n10236 ;
  assign n39385 = n31282 ^ n4187 ^ x249 ;
  assign n39386 = ( n12073 & ~n35330 ) | ( n12073 & n39385 ) | ( ~n35330 & n39385 ) ;
  assign n39387 = ~n27995 & n30221 ;
  assign n39388 = ( ~n502 & n11413 ) | ( ~n502 & n14063 ) | ( n11413 & n14063 ) ;
  assign n39389 = n39388 ^ n30198 ^ 1'b0 ;
  assign n39390 = n37808 ^ n18926 ^ 1'b0 ;
  assign n39391 = ~n2062 & n9180 ;
  assign n39392 = ~n5085 & n39391 ;
  assign n39395 = ( n7155 & n8695 ) | ( n7155 & n13201 ) | ( n8695 & n13201 ) ;
  assign n39393 = n38298 ^ n12968 ^ 1'b0 ;
  assign n39394 = n22359 & ~n39393 ;
  assign n39396 = n39395 ^ n39394 ^ 1'b0 ;
  assign n39397 = n14086 & ~n37152 ;
  assign n39398 = ( n9317 & ~n14347 ) | ( n9317 & n39397 ) | ( ~n14347 & n39397 ) ;
  assign n39399 = n31576 ^ n10636 ^ 1'b0 ;
  assign n39400 = n39399 ^ n24998 ^ n10952 ;
  assign n39401 = n31786 ^ n28461 ^ 1'b0 ;
  assign n39402 = n9318 ^ n4374 ^ 1'b0 ;
  assign n39403 = ( ~n1469 & n10716 ) | ( ~n1469 & n15825 ) | ( n10716 & n15825 ) ;
  assign n39404 = ( n6753 & n39402 ) | ( n6753 & ~n39403 ) | ( n39402 & ~n39403 ) ;
  assign n39405 = n12493 & ~n39404 ;
  assign n39406 = n4938 & ~n39405 ;
  assign n39407 = n39401 & n39406 ;
  assign n39408 = n10613 ^ n3507 ^ 1'b0 ;
  assign n39409 = n39408 ^ n21039 ^ n17472 ;
  assign n39410 = n39409 ^ n1396 ^ 1'b0 ;
  assign n39411 = ~n13436 & n39410 ;
  assign n39412 = n15313 ^ n8436 ^ 1'b0 ;
  assign n39413 = n30801 & ~n39412 ;
  assign n39417 = n19164 & n28627 ;
  assign n39418 = n39417 ^ n2029 ^ 1'b0 ;
  assign n39414 = ( n5385 & n14136 ) | ( n5385 & n30721 ) | ( n14136 & n30721 ) ;
  assign n39415 = n39414 ^ n38536 ^ n2603 ;
  assign n39416 = n9101 & ~n39415 ;
  assign n39419 = n39418 ^ n39416 ^ 1'b0 ;
  assign n39420 = n10293 & n10340 ;
  assign n39421 = n39420 ^ n25305 ^ n2727 ;
  assign n39422 = n13682 & n18894 ;
  assign n39423 = n28228 ^ n13986 ^ 1'b0 ;
  assign n39424 = n39422 & n39423 ;
  assign n39425 = ~n1776 & n8812 ;
  assign n39426 = ~n39424 & n39425 ;
  assign n39427 = ( n19466 & ~n31022 ) | ( n19466 & n39426 ) | ( ~n31022 & n39426 ) ;
  assign n39428 = n13935 ^ n7535 ^ n3346 ;
  assign n39432 = n12870 | n16349 ;
  assign n39430 = ~n868 & n12543 ;
  assign n39429 = ~n11366 & n13346 ;
  assign n39431 = n39430 ^ n39429 ^ 1'b0 ;
  assign n39433 = n39432 ^ n39431 ^ n17069 ;
  assign n39437 = n24775 ^ n22477 ^ n10385 ;
  assign n39438 = n39437 ^ n27875 ^ n14561 ;
  assign n39434 = n1396 | n26798 ;
  assign n39435 = ( n7354 & n16000 ) | ( n7354 & ~n39434 ) | ( n16000 & ~n39434 ) ;
  assign n39436 = ( n4999 & n8954 ) | ( n4999 & ~n39435 ) | ( n8954 & ~n39435 ) ;
  assign n39439 = n39438 ^ n39436 ^ n35432 ;
  assign n39440 = ( n2455 & n2501 ) | ( n2455 & ~n12121 ) | ( n2501 & ~n12121 ) ;
  assign n39441 = ( n24338 & n26234 ) | ( n24338 & ~n39440 ) | ( n26234 & ~n39440 ) ;
  assign n39442 = n39441 ^ n8324 ^ n2238 ;
  assign n39443 = n287 & n26620 ;
  assign n39444 = n39443 ^ n15913 ^ 1'b0 ;
  assign n39445 = n26286 | n37107 ;
  assign n39446 = n36108 & ~n39445 ;
  assign n39448 = ( n14706 & n19928 ) | ( n14706 & ~n21848 ) | ( n19928 & ~n21848 ) ;
  assign n39447 = n32102 ^ n21307 ^ n10236 ;
  assign n39449 = n39448 ^ n39447 ^ 1'b0 ;
  assign n39450 = x56 & n22820 ;
  assign n39451 = n39450 ^ x201 ^ 1'b0 ;
  assign n39452 = ( ~n32704 & n38253 ) | ( ~n32704 & n39451 ) | ( n38253 & n39451 ) ;
  assign n39453 = n29227 ^ n21885 ^ 1'b0 ;
  assign n39454 = n13563 & ~n14583 ;
  assign n39455 = n39454 ^ n24133 ^ 1'b0 ;
  assign n39459 = ~n11816 & n26739 ;
  assign n39460 = n39459 ^ n35617 ^ n308 ;
  assign n39456 = n3300 & ~n37294 ;
  assign n39457 = ~n6399 & n39456 ;
  assign n39458 = n23221 | n39457 ;
  assign n39461 = n39460 ^ n39458 ^ 1'b0 ;
  assign n39462 = n10858 | n36298 ;
  assign n39463 = ( n3489 & n9005 ) | ( n3489 & n10673 ) | ( n9005 & n10673 ) ;
  assign n39464 = ~n21485 & n39463 ;
  assign n39465 = n10689 & n12723 ;
  assign n39466 = n39464 & n39465 ;
  assign n39467 = ( n33354 & n37746 ) | ( n33354 & n39065 ) | ( n37746 & n39065 ) ;
  assign n39469 = ( n2348 & ~n7076 ) | ( n2348 & n21570 ) | ( ~n7076 & n21570 ) ;
  assign n39468 = ( n8062 & n14168 ) | ( n8062 & n15016 ) | ( n14168 & n15016 ) ;
  assign n39470 = n39469 ^ n39468 ^ n19521 ;
  assign n39471 = n29920 ^ n18838 ^ n2799 ;
  assign n39472 = n39471 ^ n12717 ^ 1'b0 ;
  assign n39473 = n12623 | n39472 ;
  assign n39474 = n464 & ~n39473 ;
  assign n39475 = ~n31888 & n39474 ;
  assign n39476 = n33758 ^ n22130 ^ n19357 ;
  assign n39477 = ~n10693 & n39476 ;
  assign n39478 = n39475 & n39477 ;
  assign n39479 = n39470 & ~n39478 ;
  assign n39481 = n31271 ^ n11633 ^ 1'b0 ;
  assign n39482 = n6057 & ~n39481 ;
  assign n39480 = n32226 ^ n28563 ^ n15744 ;
  assign n39483 = n39482 ^ n39480 ^ n1694 ;
  assign n39484 = n7169 | n26392 ;
  assign n39485 = n9078 | n39484 ;
  assign n39486 = ( n5180 & n12013 ) | ( n5180 & n12082 ) | ( n12013 & n12082 ) ;
  assign n39487 = n20669 ^ n12944 ^ 1'b0 ;
  assign n39488 = n39486 & ~n39487 ;
  assign n39489 = ( n10069 & n39485 ) | ( n10069 & ~n39488 ) | ( n39485 & ~n39488 ) ;
  assign n39490 = ( ~n3606 & n12630 ) | ( ~n3606 & n38211 ) | ( n12630 & n38211 ) ;
  assign n39491 = n5665 & n7423 ;
  assign n39492 = n39491 ^ n1465 ^ 1'b0 ;
  assign n39493 = n39492 ^ n10848 ^ n1010 ;
  assign n39494 = n39493 ^ n9192 ^ 1'b0 ;
  assign n39496 = ( n13048 & n19139 ) | ( n13048 & ~n27389 ) | ( n19139 & ~n27389 ) ;
  assign n39495 = n18009 ^ n8985 ^ n5590 ;
  assign n39497 = n39496 ^ n39495 ^ n12532 ;
  assign n39498 = n39406 ^ n8091 ^ n6626 ;
  assign n39499 = n6968 ^ x180 ^ x168 ;
  assign n39500 = n8011 | n39499 ;
  assign n39501 = n27580 & ~n39500 ;
  assign n39502 = n32001 ^ n10613 ^ 1'b0 ;
  assign n39504 = n10949 ^ n9572 ^ 1'b0 ;
  assign n39505 = n36039 & ~n39504 ;
  assign n39503 = n1638 & n23895 ;
  assign n39506 = n39505 ^ n39503 ^ 1'b0 ;
  assign n39507 = n2908 & ~n3181 ;
  assign n39508 = n33490 ^ n27919 ^ n5263 ;
  assign n39509 = ( ~n2903 & n10967 ) | ( ~n2903 & n15201 ) | ( n10967 & n15201 ) ;
  assign n39510 = ( n4191 & ~n11189 ) | ( n4191 & n36275 ) | ( ~n11189 & n36275 ) ;
  assign n39511 = n39509 | n39510 ;
  assign n39512 = n7073 & ~n21676 ;
  assign n39513 = n15263 & ~n16024 ;
  assign n39514 = ~n11276 & n39513 ;
  assign n39515 = n39514 ^ n29385 ^ n10966 ;
  assign n39516 = ( n11609 & n29085 ) | ( n11609 & n39515 ) | ( n29085 & n39515 ) ;
  assign n39517 = n25792 & n27613 ;
  assign n39523 = ( x43 & n2001 ) | ( x43 & n9387 ) | ( n2001 & n9387 ) ;
  assign n39519 = n12350 & n22210 ;
  assign n39520 = ( n9635 & n16734 ) | ( n9635 & ~n17360 ) | ( n16734 & ~n17360 ) ;
  assign n39521 = n39520 ^ n18463 ^ n3394 ;
  assign n39522 = ( n10506 & ~n39519 ) | ( n10506 & n39521 ) | ( ~n39519 & n39521 ) ;
  assign n39518 = ( n8669 & ~n27779 ) | ( n8669 & n28031 ) | ( ~n27779 & n28031 ) ;
  assign n39524 = n39523 ^ n39522 ^ n39518 ;
  assign n39525 = n11937 & n39524 ;
  assign n39526 = n39525 ^ n13924 ^ 1'b0 ;
  assign n39527 = ( ~n4003 & n14934 ) | ( ~n4003 & n34382 ) | ( n14934 & n34382 ) ;
  assign n39528 = n9765 & n30875 ;
  assign n39529 = n24403 & ~n32884 ;
  assign n39530 = n6632 & n39529 ;
  assign n39531 = n39530 ^ n5713 ^ n1474 ;
  assign n39532 = ~n13267 & n28598 ;
  assign n39533 = n39532 ^ n28021 ^ 1'b0 ;
  assign n39534 = n21781 ^ n15065 ^ n2329 ;
  assign n39535 = n26155 ^ n22304 ^ n6693 ;
  assign n39536 = n39535 ^ n32048 ^ n24427 ;
  assign n39537 = n12096 & n14123 ;
  assign n39540 = n8954 | n13468 ;
  assign n39538 = n9338 & ~n18992 ;
  assign n39539 = n7119 & n39538 ;
  assign n39541 = n39540 ^ n39539 ^ n4262 ;
  assign n39542 = ( n17622 & n26342 ) | ( n17622 & ~n39541 ) | ( n26342 & ~n39541 ) ;
  assign n39546 = ~n295 & n24388 ;
  assign n39544 = n10834 ^ n8158 ^ 1'b0 ;
  assign n39543 = ~n12684 & n32193 ;
  assign n39545 = n39544 ^ n39543 ^ 1'b0 ;
  assign n39547 = n39546 ^ n39545 ^ n5298 ;
  assign n39548 = n34678 ^ n1662 ^ 1'b0 ;
  assign n39549 = ~n22591 & n39548 ;
  assign n39550 = n20079 ^ n1518 ^ 1'b0 ;
  assign n39551 = ~n7309 & n39550 ;
  assign n39552 = ~n33739 & n39551 ;
  assign n39553 = n14900 & n39552 ;
  assign n39554 = n2251 & ~n16964 ;
  assign n39555 = n17013 & n39554 ;
  assign n39556 = n31228 | n39555 ;
  assign n39557 = n13138 ^ n11250 ^ 1'b0 ;
  assign n39558 = n29486 | n39557 ;
  assign n39559 = n39558 ^ n38711 ^ n8070 ;
  assign n39560 = n15182 & n17075 ;
  assign n39561 = n39560 ^ n20528 ^ 1'b0 ;
  assign n39562 = n39561 ^ n31328 ^ n8592 ;
  assign n39563 = n16123 ^ n4920 ^ 1'b0 ;
  assign n39564 = n6542 & n39563 ;
  assign n39565 = ( ~n16911 & n28365 ) | ( ~n16911 & n39564 ) | ( n28365 & n39564 ) ;
  assign n39566 = n20766 ^ n16812 ^ n2881 ;
  assign n39567 = n39566 ^ n21711 ^ 1'b0 ;
  assign n39568 = n39567 ^ n9591 ^ 1'b0 ;
  assign n39569 = n4354 & n19209 ;
  assign n39570 = n16939 & n39569 ;
  assign n39571 = n13211 & n32093 ;
  assign n39572 = n39570 & n39571 ;
  assign n39573 = ( n39565 & ~n39568 ) | ( n39565 & n39572 ) | ( ~n39568 & n39572 ) ;
  assign n39575 = ( ~n16719 & n23320 ) | ( ~n16719 & n32343 ) | ( n23320 & n32343 ) ;
  assign n39574 = n26380 ^ n12318 ^ n6761 ;
  assign n39576 = n39575 ^ n39574 ^ n23647 ;
  assign n39577 = n9437 ^ n3813 ^ n932 ;
  assign n39578 = n6111 & ~n9908 ;
  assign n39579 = n39578 ^ n19629 ^ n12513 ;
  assign n39580 = ( ~n19604 & n30669 ) | ( ~n19604 & n39579 ) | ( n30669 & n39579 ) ;
  assign n39581 = ( n12147 & ~n39577 ) | ( n12147 & n39580 ) | ( ~n39577 & n39580 ) ;
  assign n39582 = n39581 ^ n23397 ^ n16179 ;
  assign n39583 = ~n793 & n859 ;
  assign n39584 = ~n460 & n39583 ;
  assign n39585 = n9609 | n20621 ;
  assign n39586 = n39584 | n39585 ;
  assign n39587 = n36802 ^ n28458 ^ 1'b0 ;
  assign n39588 = n26275 & ~n39587 ;
  assign n39589 = n31571 ^ n1408 ^ 1'b0 ;
  assign n39590 = ~n21873 & n39589 ;
  assign n39591 = n9805 & n39590 ;
  assign n39592 = ~n3399 & n39591 ;
  assign n39593 = ( ~n715 & n24376 ) | ( ~n715 & n39592 ) | ( n24376 & n39592 ) ;
  assign n39594 = n1900 & n7851 ;
  assign n39595 = n39594 ^ n37258 ^ n4506 ;
  assign n39596 = ( ~n1644 & n23484 ) | ( ~n1644 & n32975 ) | ( n23484 & n32975 ) ;
  assign n39597 = n7741 & ~n23099 ;
  assign n39598 = n3125 & n39597 ;
  assign n39599 = ( n7326 & n9555 ) | ( n7326 & n39598 ) | ( n9555 & n39598 ) ;
  assign n39600 = ( n13291 & ~n18300 ) | ( n13291 & n39599 ) | ( ~n18300 & n39599 ) ;
  assign n39601 = n32680 ^ n18209 ^ 1'b0 ;
  assign n39602 = n4095 & n13275 ;
  assign n39603 = ~n39601 & n39602 ;
  assign n39605 = n317 & n2984 ;
  assign n39606 = n39605 ^ n8293 ^ 1'b0 ;
  assign n39604 = ~n17052 & n20930 ;
  assign n39607 = n39606 ^ n39604 ^ 1'b0 ;
  assign n39608 = n19742 & n27029 ;
  assign n39620 = n4391 & n28011 ;
  assign n39621 = n9756 & n39620 ;
  assign n39617 = ( ~n2739 & n4865 ) | ( ~n2739 & n5301 ) | ( n4865 & n5301 ) ;
  assign n39618 = ~n5536 & n39617 ;
  assign n39619 = ( n11013 & n13325 ) | ( n11013 & ~n39618 ) | ( n13325 & ~n39618 ) ;
  assign n39609 = n13654 & ~n19602 ;
  assign n39610 = n39609 ^ n28152 ^ 1'b0 ;
  assign n39614 = n4300 & ~n18841 ;
  assign n39611 = ~n2295 & n6727 ;
  assign n39612 = n39611 ^ n8371 ^ 1'b0 ;
  assign n39613 = n16000 | n39612 ;
  assign n39615 = n39614 ^ n39613 ^ n34195 ;
  assign n39616 = ( n26236 & n39610 ) | ( n26236 & n39615 ) | ( n39610 & n39615 ) ;
  assign n39622 = n39621 ^ n39619 ^ n39616 ;
  assign n39623 = n23023 ^ n9064 ^ n7308 ;
  assign n39624 = ~n3015 & n12361 ;
  assign n39625 = n39624 ^ n781 ^ 1'b0 ;
  assign n39626 = n2661 & n20916 ;
  assign n39627 = ~n1113 & n39626 ;
  assign n39628 = n23355 | n39627 ;
  assign n39629 = n39628 ^ n21111 ^ 1'b0 ;
  assign n39630 = n686 & ~n24785 ;
  assign n39631 = ( n902 & n29056 ) | ( n902 & n39630 ) | ( n29056 & n39630 ) ;
  assign n39632 = n3176 & ~n27676 ;
  assign n39633 = n2349 & ~n2824 ;
  assign n39634 = ~n2653 & n39633 ;
  assign n39635 = n29062 & n39634 ;
  assign n39636 = n10154 ^ n7722 ^ 1'b0 ;
  assign n39637 = ~n39635 & n39636 ;
  assign n39638 = n39637 ^ n10552 ^ 1'b0 ;
  assign n39639 = n13372 ^ n5427 ^ 1'b0 ;
  assign n39640 = n5284 & n34602 ;
  assign n39641 = n544 | n28371 ;
  assign n39642 = n16950 & ~n34894 ;
  assign n39643 = ~n39641 & n39642 ;
  assign n39645 = n25228 ^ n9090 ^ n7789 ;
  assign n39644 = n7586 & n27141 ;
  assign n39646 = n39645 ^ n39644 ^ 1'b0 ;
  assign n39647 = ( n17023 & n17604 ) | ( n17023 & ~n29696 ) | ( n17604 & ~n29696 ) ;
  assign n39648 = ( ~n5355 & n8170 ) | ( ~n5355 & n39647 ) | ( n8170 & n39647 ) ;
  assign n39649 = n12650 ^ n4572 ^ n2162 ;
  assign n39650 = n8883 & ~n39649 ;
  assign n39651 = n39648 & n39650 ;
  assign n39652 = n27135 ^ n5878 ^ 1'b0 ;
  assign n39653 = n2326 & ~n39652 ;
  assign n39654 = n28121 & n39653 ;
  assign n39655 = ~n14297 & n39654 ;
  assign n39656 = ( n6765 & n10485 ) | ( n6765 & n16752 ) | ( n10485 & n16752 ) ;
  assign n39657 = n39656 ^ n4332 ^ 1'b0 ;
  assign n39658 = ( n10832 & n39655 ) | ( n10832 & n39657 ) | ( n39655 & n39657 ) ;
  assign n39659 = n11926 ^ n8088 ^ 1'b0 ;
  assign n39660 = n39659 ^ n39535 ^ n19580 ;
  assign n39661 = n10525 & n19045 ;
  assign n39662 = ~n35711 & n39661 ;
  assign n39663 = n39662 ^ n28132 ^ x10 ;
  assign n39664 = n4187 & n6204 ;
  assign n39665 = ~n20840 & n39664 ;
  assign n39666 = n27669 ^ n840 ^ 1'b0 ;
  assign n39667 = n3747 & ~n39666 ;
  assign n39668 = ( ~n37984 & n39665 ) | ( ~n37984 & n39667 ) | ( n39665 & n39667 ) ;
  assign n39669 = n21600 ^ n10107 ^ n534 ;
  assign n39670 = n38896 ^ n6042 ^ 1'b0 ;
  assign n39671 = n31603 | n39670 ;
  assign n39672 = n29581 ^ n17313 ^ 1'b0 ;
  assign n39673 = ~n33791 & n39672 ;
  assign n39674 = n21785 ^ n11627 ^ n6477 ;
  assign n39675 = ( n16812 & ~n35770 ) | ( n16812 & n39674 ) | ( ~n35770 & n39674 ) ;
  assign n39676 = n22554 ^ n16702 ^ n6739 ;
  assign n39677 = n17780 ^ n13713 ^ n2979 ;
  assign n39678 = ~n39676 & n39677 ;
  assign n39679 = n39678 ^ n31252 ^ n19170 ;
  assign n39680 = n33937 ^ n11572 ^ n6146 ;
  assign n39681 = n32586 ^ n27040 ^ n15694 ;
  assign n39682 = n30509 ^ n1310 ^ 1'b0 ;
  assign n39683 = n1144 & n28076 ;
  assign n39684 = n20491 ^ n10840 ^ 1'b0 ;
  assign n39685 = n39684 ^ n858 ^ 1'b0 ;
  assign n39686 = ( n11314 & n22664 ) | ( n11314 & ~n39685 ) | ( n22664 & ~n39685 ) ;
  assign n39687 = n39686 ^ n36129 ^ 1'b0 ;
  assign n39688 = n29736 ^ n19732 ^ 1'b0 ;
  assign n39689 = ~n6151 & n39688 ;
  assign n39690 = ( ~n13590 & n15427 ) | ( ~n13590 & n18386 ) | ( n15427 & n18386 ) ;
  assign n39691 = n32638 ^ n24040 ^ 1'b0 ;
  assign n39692 = n17850 ^ n3747 ^ x118 ;
  assign n39693 = n22511 ^ n6167 ^ 1'b0 ;
  assign n39694 = n39692 & n39693 ;
  assign n39695 = n39694 ^ n18153 ^ 1'b0 ;
  assign n39696 = n39691 & ~n39695 ;
  assign n39697 = n5791 ^ n4523 ^ 1'b0 ;
  assign n39698 = ( ~n509 & n14433 ) | ( ~n509 & n39697 ) | ( n14433 & n39697 ) ;
  assign n39699 = n1677 & n39231 ;
  assign n39700 = n39699 ^ n16438 ^ 1'b0 ;
  assign n39701 = n34274 ^ n7671 ^ 1'b0 ;
  assign n39702 = n39700 & n39701 ;
  assign n39703 = n2712 & ~n6425 ;
  assign n39704 = n39703 ^ n5495 ^ 1'b0 ;
  assign n39705 = n39704 ^ x192 ^ 1'b0 ;
  assign n39706 = n21943 ^ n1261 ^ 1'b0 ;
  assign n39707 = ~n8212 & n39706 ;
  assign n39708 = ~n32878 & n39707 ;
  assign n39709 = n39708 ^ n36754 ^ n34571 ;
  assign n39710 = ( n17082 & n18450 ) | ( n17082 & n27634 ) | ( n18450 & n27634 ) ;
  assign n39711 = n39710 ^ n35028 ^ 1'b0 ;
  assign n39712 = n8200 ^ n7397 ^ 1'b0 ;
  assign n39713 = n39437 & n39712 ;
  assign n39714 = n19281 & n39713 ;
  assign n39715 = n23570 ^ n16357 ^ 1'b0 ;
  assign n39716 = ( ~n6712 & n23235 ) | ( ~n6712 & n39715 ) | ( n23235 & n39715 ) ;
  assign n39717 = n1749 & n39716 ;
  assign n39718 = ~n6877 & n17851 ;
  assign n39719 = n39718 ^ n4213 ^ 1'b0 ;
  assign n39720 = n9422 ^ n7314 ^ n2592 ;
  assign n39721 = n39720 ^ n36096 ^ 1'b0 ;
  assign n39722 = n37802 | n39721 ;
  assign n39723 = n39722 ^ n2880 ^ 1'b0 ;
  assign n39724 = n32825 & ~n39723 ;
  assign n39725 = n4538 & n29332 ;
  assign n39726 = n10563 & n24580 ;
  assign n39727 = n6073 & n20385 ;
  assign n39728 = n39290 & n39727 ;
  assign n39729 = n39728 ^ n7181 ^ 1'b0 ;
  assign n39730 = n9252 & n11777 ;
  assign n39731 = ~n23313 & n39730 ;
  assign n39732 = n39731 ^ n1561 ^ n1347 ;
  assign n39733 = n26485 ^ x121 ^ 1'b0 ;
  assign n39734 = ( n18258 & ~n25198 ) | ( n18258 & n39733 ) | ( ~n25198 & n39733 ) ;
  assign n39735 = ( n28815 & ~n37555 ) | ( n28815 & n37685 ) | ( ~n37555 & n37685 ) ;
  assign n39736 = n3362 ^ n2967 ^ 1'b0 ;
  assign n39737 = ~n33411 & n39736 ;
  assign n39738 = n23990 ^ n3902 ^ 1'b0 ;
  assign n39739 = n15243 & ~n39738 ;
  assign n39740 = ~n22696 & n39739 ;
  assign n39741 = n39740 ^ n6932 ^ 1'b0 ;
  assign n39742 = ( n27938 & n29287 ) | ( n27938 & ~n30329 ) | ( n29287 & ~n30329 ) ;
  assign n39743 = n39742 ^ n3612 ^ 1'b0 ;
  assign n39744 = ( n9951 & ~n26691 ) | ( n9951 & n28057 ) | ( ~n26691 & n28057 ) ;
  assign n39745 = n39744 ^ n15368 ^ 1'b0 ;
  assign n39746 = n3228 & n23928 ;
  assign n39747 = n39746 ^ n16219 ^ 1'b0 ;
  assign n39748 = n28021 ^ n21616 ^ n14037 ;
  assign n39749 = ( n1548 & n15148 ) | ( n1548 & n39748 ) | ( n15148 & n39748 ) ;
  assign n39750 = ( n2553 & n6551 ) | ( n2553 & ~n22006 ) | ( n6551 & ~n22006 ) ;
  assign n39751 = n4646 & n28102 ;
  assign n39752 = n39750 & ~n39751 ;
  assign n39753 = ~n26204 & n39752 ;
  assign n39754 = ~n1953 & n4660 ;
  assign n39755 = n39754 ^ n22578 ^ 1'b0 ;
  assign n39756 = n5204 & ~n39755 ;
  assign n39757 = ( n7783 & n24725 ) | ( n7783 & ~n39756 ) | ( n24725 & ~n39756 ) ;
  assign n39758 = ( ~n2300 & n13271 ) | ( ~n2300 & n24937 ) | ( n13271 & n24937 ) ;
  assign n39759 = n39758 ^ n20596 ^ n16708 ;
  assign n39760 = ( n1923 & ~n12975 ) | ( n1923 & n39759 ) | ( ~n12975 & n39759 ) ;
  assign n39761 = n7518 ^ n1934 ^ 1'b0 ;
  assign n39762 = n14001 & ~n39761 ;
  assign n39763 = n39762 ^ n28027 ^ n19125 ;
  assign n39764 = n39763 ^ n35427 ^ 1'b0 ;
  assign n39765 = n38049 ^ n9175 ^ 1'b0 ;
  assign n39766 = n5570 ^ n4463 ^ 1'b0 ;
  assign n39767 = n19009 ^ n10890 ^ n8034 ;
  assign n39768 = ( n12085 & n39766 ) | ( n12085 & ~n39767 ) | ( n39766 & ~n39767 ) ;
  assign n39769 = n38250 ^ n32579 ^ n16530 ;
  assign n39770 = n29098 | n30359 ;
  assign n39771 = n39770 ^ n1693 ^ 1'b0 ;
  assign n39772 = ( n1924 & n5961 ) | ( n1924 & n26561 ) | ( n5961 & n26561 ) ;
  assign n39773 = ( n1046 & n2988 ) | ( n1046 & n11588 ) | ( n2988 & n11588 ) ;
  assign n39777 = n622 ^ x161 ^ 1'b0 ;
  assign n39778 = n39777 ^ n11540 ^ 1'b0 ;
  assign n39779 = n28892 | n39778 ;
  assign n39775 = n9298 & ~n17416 ;
  assign n39776 = n39775 ^ n36049 ^ 1'b0 ;
  assign n39780 = n39779 ^ n39776 ^ 1'b0 ;
  assign n39774 = n15163 ^ n4354 ^ 1'b0 ;
  assign n39781 = n39780 ^ n39774 ^ n15681 ;
  assign n39782 = n34136 ^ n5557 ^ n2658 ;
  assign n39783 = ( n3262 & n8665 ) | ( n3262 & ~n39782 ) | ( n8665 & ~n39782 ) ;
  assign n39784 = ( n4435 & n19003 ) | ( n4435 & n23185 ) | ( n19003 & n23185 ) ;
  assign n39785 = n9832 ^ n7576 ^ 1'b0 ;
  assign n39786 = n5357 & n39785 ;
  assign n39787 = n3182 ^ n1790 ^ n676 ;
  assign n39788 = ~n16208 & n22666 ;
  assign n39789 = n13209 & n39788 ;
  assign n39790 = ( n4245 & n39787 ) | ( n4245 & ~n39789 ) | ( n39787 & ~n39789 ) ;
  assign n39791 = n6339 & n39790 ;
  assign n39792 = n27032 ^ n11845 ^ 1'b0 ;
  assign n39793 = n19859 & ~n39792 ;
  assign n39794 = n19013 ^ n3828 ^ 1'b0 ;
  assign n39795 = n459 & n11954 ;
  assign n39796 = n39795 ^ n772 ^ 1'b0 ;
  assign n39797 = n21794 ^ n13949 ^ n1652 ;
  assign n39798 = n15979 & n39797 ;
  assign n39799 = ~n12522 & n39798 ;
  assign n39800 = ( n39794 & n39796 ) | ( n39794 & n39799 ) | ( n39796 & n39799 ) ;
  assign n39801 = ( x104 & n9832 ) | ( x104 & ~n39800 ) | ( n9832 & ~n39800 ) ;
  assign n39802 = ~n7578 & n32610 ;
  assign n39803 = n39802 ^ n15609 ^ 1'b0 ;
  assign n39804 = ( n5091 & n7558 ) | ( n5091 & n39803 ) | ( n7558 & n39803 ) ;
  assign n39805 = n22993 ^ n2560 ^ 1'b0 ;
  assign n39806 = ~n32223 & n39805 ;
  assign n39807 = ( ~n8946 & n30976 ) | ( ~n8946 & n39806 ) | ( n30976 & n39806 ) ;
  assign n39808 = n13203 & n31998 ;
  assign n39809 = n39808 ^ n2051 ^ 1'b0 ;
  assign n39810 = n39809 ^ n9599 ^ 1'b0 ;
  assign n39811 = ( n6305 & ~n10926 ) | ( n6305 & n37955 ) | ( ~n10926 & n37955 ) ;
  assign n39812 = ( n2732 & n8248 ) | ( n2732 & ~n13504 ) | ( n8248 & ~n13504 ) ;
  assign n39813 = n39812 ^ n37109 ^ 1'b0 ;
  assign n39814 = n14102 ^ n4333 ^ 1'b0 ;
  assign n39815 = n2924 | n39814 ;
  assign n39816 = n6933 & n30483 ;
  assign n39817 = n39815 & n39816 ;
  assign n39818 = n2804 | n18511 ;
  assign n39819 = n39818 ^ n6870 ^ 1'b0 ;
  assign n39820 = n24085 ^ n13956 ^ 1'b0 ;
  assign n39821 = ~n39819 & n39820 ;
  assign n39822 = ( n14603 & n23113 ) | ( n14603 & ~n27599 ) | ( n23113 & ~n27599 ) ;
  assign n39823 = n34828 ^ n14600 ^ 1'b0 ;
  assign n39824 = n3821 & ~n22434 ;
  assign n39825 = n39824 ^ n9807 ^ 1'b0 ;
  assign n39826 = n32341 & ~n39825 ;
  assign n39827 = n7217 | n10842 ;
  assign n39828 = n35280 & ~n39827 ;
  assign n39829 = n39828 ^ n39572 ^ n29450 ;
  assign n39830 = n12634 & n21562 ;
  assign n39831 = n5895 & n39830 ;
  assign n39832 = n39831 ^ n11854 ^ n6553 ;
  assign n39833 = n28801 ^ n24402 ^ 1'b0 ;
  assign n39834 = n6994 & ~n7992 ;
  assign n39835 = n10420 ^ n4694 ^ 1'b0 ;
  assign n39836 = n3471 & n39835 ;
  assign n39838 = n4043 ^ n3510 ^ 1'b0 ;
  assign n39839 = n24137 & ~n39838 ;
  assign n39837 = n15203 ^ n8408 ^ n7558 ;
  assign n39840 = n39839 ^ n39837 ^ 1'b0 ;
  assign n39841 = ( ~n737 & n2875 ) | ( ~n737 & n11428 ) | ( n2875 & n11428 ) ;
  assign n39842 = n393 & n622 ;
  assign n39843 = n39842 ^ n17178 ^ 1'b0 ;
  assign n39844 = ( n1995 & n30577 ) | ( n1995 & n39843 ) | ( n30577 & n39843 ) ;
  assign n39845 = n27912 ^ n21321 ^ n1404 ;
  assign n39846 = n39845 ^ n34653 ^ n21063 ;
  assign n39847 = n23604 ^ n3647 ^ 1'b0 ;
  assign n39848 = n9350 & n25503 ;
  assign n39849 = n39848 ^ n19529 ^ 1'b0 ;
  assign n39850 = n23280 ^ n13315 ^ n4747 ;
  assign n39851 = n2681 | n28380 ;
  assign n39852 = n39850 | n39851 ;
  assign n39853 = n35414 ^ n14625 ^ n9840 ;
  assign n39854 = n2025 & n22781 ;
  assign n39855 = ~n39853 & n39854 ;
  assign n39856 = n24666 ^ n10602 ^ 1'b0 ;
  assign n39857 = ~n39855 & n39856 ;
  assign n39858 = n24697 ^ n13258 ^ n3217 ;
  assign n39859 = ( ~n3634 & n27058 ) | ( ~n3634 & n39858 ) | ( n27058 & n39858 ) ;
  assign n39860 = n38419 ^ n38212 ^ n25385 ;
  assign n39861 = n24130 ^ n3217 ^ 1'b0 ;
  assign n39862 = n23239 ^ n20122 ^ 1'b0 ;
  assign n39863 = ~n39861 & n39862 ;
  assign n39866 = n23310 ^ n501 ^ 1'b0 ;
  assign n39864 = n6479 ^ n1445 ^ 1'b0 ;
  assign n39865 = n10095 & n39864 ;
  assign n39867 = n39866 ^ n39865 ^ n7707 ;
  assign n39868 = ( n7645 & ~n39863 ) | ( n7645 & n39867 ) | ( ~n39863 & n39867 ) ;
  assign n39869 = n20767 & ~n21312 ;
  assign n39870 = n945 ^ n897 ^ 1'b0 ;
  assign n39871 = ~n36975 & n39870 ;
  assign n39872 = n30178 & n39871 ;
  assign n39873 = n39872 ^ n1042 ^ 1'b0 ;
  assign n39874 = n28617 ^ n10944 ^ 1'b0 ;
  assign n39875 = n27248 ^ n23724 ^ n6460 ;
  assign n39876 = n8327 & n14202 ;
  assign n39877 = n1105 & n39876 ;
  assign n39878 = ( n9018 & n17425 ) | ( n9018 & n39877 ) | ( n17425 & n39877 ) ;
  assign n39879 = n38292 ^ n11901 ^ 1'b0 ;
  assign n39880 = ( n6005 & n8416 ) | ( n6005 & n16722 ) | ( n8416 & n16722 ) ;
  assign n39882 = n24806 ^ n6362 ^ 1'b0 ;
  assign n39883 = n39882 ^ n19782 ^ n2541 ;
  assign n39881 = ~n534 & n8672 ;
  assign n39884 = n39883 ^ n39881 ^ 1'b0 ;
  assign n39885 = n6433 ^ n6364 ^ 1'b0 ;
  assign n39886 = n17549 & n39885 ;
  assign n39887 = n38779 ^ n11033 ^ 1'b0 ;
  assign n39888 = ( n39884 & n39886 ) | ( n39884 & n39887 ) | ( n39886 & n39887 ) ;
  assign n39889 = n33688 ^ n25514 ^ n13336 ;
  assign n39890 = n35792 & n39889 ;
  assign n39894 = ( x59 & n8654 ) | ( x59 & n9378 ) | ( n8654 & n9378 ) ;
  assign n39891 = n16519 ^ n5026 ^ 1'b0 ;
  assign n39892 = n39891 ^ n33510 ^ n2920 ;
  assign n39893 = ( n25699 & n38638 ) | ( n25699 & n39892 ) | ( n38638 & n39892 ) ;
  assign n39895 = n39894 ^ n39893 ^ n3214 ;
  assign n39896 = n2492 & ~n13831 ;
  assign n39897 = n4033 & ~n32964 ;
  assign n39898 = n39896 & n39897 ;
  assign n39899 = n4949 & ~n34894 ;
  assign n39900 = n716 & n39899 ;
  assign n39901 = ~n4615 & n20112 ;
  assign n39902 = n358 | n27354 ;
  assign n39903 = n39901 & ~n39902 ;
  assign n39904 = n11736 | n23951 ;
  assign n39905 = ( n5750 & n24185 ) | ( n5750 & ~n39904 ) | ( n24185 & ~n39904 ) ;
  assign n39906 = n37356 ^ n28774 ^ n6601 ;
  assign n39907 = ( n18977 & ~n19310 ) | ( n18977 & n39906 ) | ( ~n19310 & n39906 ) ;
  assign n39908 = n39176 ^ n23997 ^ n3491 ;
  assign n39909 = n39908 ^ n4465 ^ 1'b0 ;
  assign n39910 = ( ~n15391 & n31444 ) | ( ~n15391 & n39909 ) | ( n31444 & n39909 ) ;
  assign n39911 = n29887 & ~n31161 ;
  assign n39912 = n15000 ^ n9879 ^ n4632 ;
  assign n39913 = n39912 ^ n31578 ^ n4158 ;
  assign n39914 = ( n26163 & n33854 ) | ( n26163 & ~n39913 ) | ( n33854 & ~n39913 ) ;
  assign n39915 = n18558 ^ n12751 ^ n4533 ;
  assign n39916 = n14104 | n39915 ;
  assign n39917 = n39916 ^ n14518 ^ 1'b0 ;
  assign n39918 = n7699 | n13163 ;
  assign n39919 = n36124 & ~n39918 ;
  assign n39920 = n39919 ^ n35756 ^ n4519 ;
  assign n39921 = ( n8451 & n9353 ) | ( n8451 & ~n21694 ) | ( n9353 & ~n21694 ) ;
  assign n39922 = n7279 & n27845 ;
  assign n39923 = n29353 ^ n24823 ^ n7344 ;
  assign n39924 = n12467 & n26143 ;
  assign n39925 = n39924 ^ n2727 ^ 1'b0 ;
  assign n39926 = n29182 ^ n6961 ^ 1'b0 ;
  assign n39927 = n39925 | n39926 ;
  assign n39928 = n31721 | n32483 ;
  assign n39929 = n6494 & ~n39928 ;
  assign n39930 = n23960 ^ n14348 ^ 1'b0 ;
  assign n39931 = ~n31975 & n39930 ;
  assign n39932 = n39931 ^ n8064 ^ 1'b0 ;
  assign n39933 = x31 & ~n8413 ;
  assign n39934 = ( n19957 & n21428 ) | ( n19957 & n39933 ) | ( n21428 & n39933 ) ;
  assign n39935 = ~n3924 & n39934 ;
  assign n39936 = n39935 ^ n27784 ^ 1'b0 ;
  assign n39937 = n39936 ^ n3885 ^ n3458 ;
  assign n39938 = ~n9575 & n26280 ;
  assign n39939 = ( n15109 & n17807 ) | ( n15109 & ~n19391 ) | ( n17807 & ~n19391 ) ;
  assign n39940 = n39939 ^ n17033 ^ 1'b0 ;
  assign n39941 = n858 & ~n39940 ;
  assign n39942 = ( ~n17156 & n24748 ) | ( ~n17156 & n39941 ) | ( n24748 & n39941 ) ;
  assign n39943 = ( n39937 & ~n39938 ) | ( n39937 & n39942 ) | ( ~n39938 & n39942 ) ;
  assign n39944 = n4652 ^ n4475 ^ 1'b0 ;
  assign n39945 = n23501 & ~n39944 ;
  assign n39946 = n39945 ^ n16457 ^ 1'b0 ;
  assign n39947 = ~n23577 & n32492 ;
  assign n39948 = ( n4640 & n5711 ) | ( n4640 & n39947 ) | ( n5711 & n39947 ) ;
  assign n39949 = n15147 ^ n14708 ^ n6127 ;
  assign n39950 = n2838 | n5226 ;
  assign n39951 = n39950 ^ n18579 ^ 1'b0 ;
  assign n39952 = n25912 ^ n10426 ^ 1'b0 ;
  assign n39953 = ~n2250 & n39952 ;
  assign n39954 = n39953 ^ n18033 ^ n16051 ;
  assign n39955 = n39171 ^ n33555 ^ n1271 ;
  assign n39956 = ~n25338 & n37464 ;
  assign n39957 = n19655 | n24849 ;
  assign n39958 = n4368 | n39957 ;
  assign n39959 = n8600 ^ n3537 ^ 1'b0 ;
  assign n39960 = ( n1561 & ~n5709 ) | ( n1561 & n39959 ) | ( ~n5709 & n39959 ) ;
  assign n39961 = n39960 ^ n23465 ^ n19832 ;
  assign n39962 = ~n1086 & n39961 ;
  assign n39963 = ( n6455 & ~n27844 ) | ( n6455 & n30536 ) | ( ~n27844 & n30536 ) ;
  assign n39964 = n33985 ^ n8403 ^ n3468 ;
  assign n39965 = n26843 ^ n4090 ^ 1'b0 ;
  assign n39966 = n7818 & n37541 ;
  assign n39967 = n39966 ^ n9010 ^ 1'b0 ;
  assign n39968 = n39965 & n39967 ;
  assign n39969 = n29761 ^ n9151 ^ n3515 ;
  assign n39970 = ( n20587 & ~n36518 ) | ( n20587 & n39969 ) | ( ~n36518 & n39969 ) ;
  assign n39971 = ~n12971 & n16342 ;
  assign n39972 = n39971 ^ n1282 ^ 1'b0 ;
  assign n39973 = n21082 | n39972 ;
  assign n39974 = n39686 ^ n14926 ^ n9072 ;
  assign n39975 = n39974 ^ n28192 ^ 1'b0 ;
  assign n39976 = ( n317 & n9821 ) | ( n317 & ~n9832 ) | ( n9821 & ~n9832 ) ;
  assign n39977 = n707 & n913 ;
  assign n39978 = ( n28453 & n39976 ) | ( n28453 & ~n39977 ) | ( n39976 & ~n39977 ) ;
  assign n39980 = ( n12042 & n24250 ) | ( n12042 & ~n37937 ) | ( n24250 & ~n37937 ) ;
  assign n39979 = n26485 ^ n6916 ^ n768 ;
  assign n39981 = n39980 ^ n39979 ^ 1'b0 ;
  assign n39982 = n15411 & ~n17607 ;
  assign n39983 = n17496 ^ n8371 ^ 1'b0 ;
  assign n39984 = n39983 ^ n10653 ^ 1'b0 ;
  assign n39985 = n7426 & n39984 ;
  assign n39986 = n18204 & ~n21501 ;
  assign n39987 = n36789 & n39986 ;
  assign n39988 = n23895 & ~n38083 ;
  assign n39989 = n22047 | n29166 ;
  assign n39990 = n39989 ^ n11730 ^ n1015 ;
  assign n39991 = n39990 ^ n39521 ^ n10831 ;
  assign n39994 = n29787 ^ n12641 ^ 1'b0 ;
  assign n39992 = n1951 | n15906 ;
  assign n39993 = n39992 ^ n26911 ^ 1'b0 ;
  assign n39995 = n39994 ^ n39993 ^ n8379 ;
  assign n39996 = n8447 | n32734 ;
  assign n39997 = n39996 ^ n700 ^ 1'b0 ;
  assign n39998 = n3776 ^ n2311 ^ 1'b0 ;
  assign n39999 = n34432 ^ n11735 ^ n3472 ;
  assign n40000 = n5902 ^ n260 ^ 1'b0 ;
  assign n40001 = x192 & ~n40000 ;
  assign n40002 = n40001 ^ n8422 ^ 1'b0 ;
  assign n40003 = n2939 & ~n27600 ;
  assign n40004 = n40003 ^ n19402 ^ 1'b0 ;
  assign n40005 = ~n6481 & n12374 ;
  assign n40006 = n40005 ^ n6004 ^ 1'b0 ;
  assign n40007 = n32670 | n40006 ;
  assign n40008 = ( n3939 & n6648 ) | ( n3939 & ~n10343 ) | ( n6648 & ~n10343 ) ;
  assign n40011 = n1489 & ~n2950 ;
  assign n40009 = ~n4779 & n9693 ;
  assign n40010 = n40009 ^ n11509 ^ n11011 ;
  assign n40012 = n40011 ^ n40010 ^ n13177 ;
  assign n40013 = n40012 ^ n5708 ^ 1'b0 ;
  assign n40014 = n38757 ^ n7590 ^ n1775 ;
  assign n40015 = ( n1189 & ~n40013 ) | ( n1189 & n40014 ) | ( ~n40013 & n40014 ) ;
  assign n40016 = n36902 ^ n35765 ^ n14112 ;
  assign n40017 = ~n18937 & n27002 ;
  assign n40018 = n40017 ^ n21913 ^ 1'b0 ;
  assign n40019 = n16098 & ~n30850 ;
  assign n40020 = n26241 & ~n40019 ;
  assign n40021 = n40020 ^ n20444 ^ 1'b0 ;
  assign n40022 = n15065 & n40021 ;
  assign n40033 = n14933 & n20430 ;
  assign n40027 = ~n10432 & n18070 ;
  assign n40029 = n34720 ^ n28826 ^ n1473 ;
  assign n40028 = n1951 & n10277 ;
  assign n40030 = n40029 ^ n40028 ^ 1'b0 ;
  assign n40031 = n5799 & n40030 ;
  assign n40032 = ( n32294 & ~n40027 ) | ( n32294 & n40031 ) | ( ~n40027 & n40031 ) ;
  assign n40023 = ~n18627 & n27749 ;
  assign n40024 = n27900 ^ n1208 ^ 1'b0 ;
  assign n40025 = n12739 & n40024 ;
  assign n40026 = ( n32299 & n40023 ) | ( n32299 & n40025 ) | ( n40023 & n40025 ) ;
  assign n40034 = n40033 ^ n40032 ^ n40026 ;
  assign n40035 = n12586 ^ n2661 ^ 1'b0 ;
  assign n40036 = n25877 ^ n3281 ^ 1'b0 ;
  assign n40037 = ~n19568 & n40036 ;
  assign n40039 = n7215 ^ n5634 ^ n463 ;
  assign n40040 = n40039 ^ n10751 ^ n3787 ;
  assign n40038 = n36860 ^ n3552 ^ 1'b0 ;
  assign n40041 = n40040 ^ n40038 ^ n38230 ;
  assign n40042 = ( n1171 & ~n40037 ) | ( n1171 & n40041 ) | ( ~n40037 & n40041 ) ;
  assign n40043 = n37399 ^ n34170 ^ n1854 ;
  assign n40044 = n40043 ^ n2205 ^ 1'b0 ;
  assign n40045 = n40042 & n40044 ;
  assign n40046 = ( n1353 & n2398 ) | ( n1353 & ~n4713 ) | ( n2398 & ~n4713 ) ;
  assign n40047 = n663 & n8168 ;
  assign n40048 = n2036 & n40047 ;
  assign n40049 = n40048 ^ n12277 ^ 1'b0 ;
  assign n40050 = ( n15614 & ~n40046 ) | ( n15614 & n40049 ) | ( ~n40046 & n40049 ) ;
  assign n40051 = n37679 ^ n8455 ^ n5783 ;
  assign n40052 = ( n11976 & ~n38886 ) | ( n11976 & n40051 ) | ( ~n38886 & n40051 ) ;
  assign n40053 = n1260 | n14512 ;
  assign n40054 = n15510 | n40053 ;
  assign n40056 = n9876 ^ n9558 ^ 1'b0 ;
  assign n40057 = n460 & ~n40056 ;
  assign n40055 = n33415 ^ n20471 ^ n525 ;
  assign n40058 = n40057 ^ n40055 ^ 1'b0 ;
  assign n40059 = n16241 | n40058 ;
  assign n40060 = n8617 & ~n40059 ;
  assign n40061 = n31343 ^ n28787 ^ n3061 ;
  assign n40062 = n40061 ^ n26858 ^ 1'b0 ;
  assign n40063 = ( n12239 & ~n20772 ) | ( n12239 & n33395 ) | ( ~n20772 & n33395 ) ;
  assign n40064 = n40063 ^ n18257 ^ 1'b0 ;
  assign n40065 = n7844 & n39759 ;
  assign n40066 = ~n40064 & n40065 ;
  assign n40067 = n23373 ^ n13033 ^ 1'b0 ;
  assign n40068 = n32223 ^ n26038 ^ n19768 ;
  assign n40069 = ~n8023 & n19628 ;
  assign n40070 = n14446 & n15864 ;
  assign n40071 = ( n21071 & n40069 ) | ( n21071 & ~n40070 ) | ( n40069 & ~n40070 ) ;
  assign n40072 = n9234 | n15095 ;
  assign n40073 = n21485 | n29465 ;
  assign n40074 = n40073 ^ n39099 ^ 1'b0 ;
  assign n40075 = n35765 ^ n5354 ^ 1'b0 ;
  assign n40076 = n23508 ^ n9926 ^ n3083 ;
  assign n40077 = n32472 ^ n19672 ^ 1'b0 ;
  assign n40078 = n14127 ^ n11443 ^ n2126 ;
  assign n40079 = n15960 & ~n22509 ;
  assign n40080 = ~n7776 & n40079 ;
  assign n40081 = ( x149 & n13175 ) | ( x149 & n40080 ) | ( n13175 & n40080 ) ;
  assign n40082 = n11595 ^ n11322 ^ n7500 ;
  assign n40083 = n40082 ^ n20117 ^ 1'b0 ;
  assign n40084 = ( n3397 & ~n3644 ) | ( n3397 & n19591 ) | ( ~n3644 & n19591 ) ;
  assign n40085 = ( n19450 & n22438 ) | ( n19450 & ~n26767 ) | ( n22438 & ~n26767 ) ;
  assign n40090 = n26488 ^ n6219 ^ n1272 ;
  assign n40086 = ~n5176 & n33751 ;
  assign n40087 = n18333 & n40086 ;
  assign n40088 = n40087 ^ n23327 ^ n15751 ;
  assign n40089 = n26763 & ~n40088 ;
  assign n40091 = n40090 ^ n40089 ^ n9543 ;
  assign n40092 = ( n448 & ~n1943 ) | ( n448 & n10052 ) | ( ~n1943 & n10052 ) ;
  assign n40093 = n32898 ^ n28991 ^ n9801 ;
  assign n40094 = n35438 & n40093 ;
  assign n40095 = n40094 ^ n38406 ^ 1'b0 ;
  assign n40096 = ~n23756 & n40095 ;
  assign n40097 = n12040 & n40096 ;
  assign n40098 = ( n26013 & ~n40092 ) | ( n26013 & n40097 ) | ( ~n40092 & n40097 ) ;
  assign n40101 = n9369 ^ n6236 ^ n4376 ;
  assign n40099 = n35294 ^ n16483 ^ 1'b0 ;
  assign n40100 = n40051 | n40099 ;
  assign n40102 = n40101 ^ n40100 ^ n1089 ;
  assign n40103 = n26113 ^ n10388 ^ 1'b0 ;
  assign n40104 = n40103 ^ n14916 ^ 1'b0 ;
  assign n40105 = n27108 | n40104 ;
  assign n40106 = n40105 ^ n24347 ^ n9656 ;
  assign n40107 = ( n3349 & n12247 ) | ( n3349 & ~n25486 ) | ( n12247 & ~n25486 ) ;
  assign n40108 = n40107 ^ n9980 ^ 1'b0 ;
  assign n40109 = n11215 ^ n7595 ^ 1'b0 ;
  assign n40110 = n37742 & ~n40109 ;
  assign n40111 = ( n627 & n5734 ) | ( n627 & n14620 ) | ( n5734 & n14620 ) ;
  assign n40112 = n7454 ^ n6835 ^ n3124 ;
  assign n40113 = ~n22164 & n40112 ;
  assign n40114 = ( ~n34943 & n40111 ) | ( ~n34943 & n40113 ) | ( n40111 & n40113 ) ;
  assign n40115 = n38035 ^ n28860 ^ n18463 ;
  assign n40116 = n8946 | n12889 ;
  assign n40117 = n40116 ^ n23844 ^ n15556 ;
  assign n40118 = n39012 ^ n19107 ^ n9801 ;
  assign n40119 = n14545 & n16049 ;
  assign n40120 = n40119 ^ n10384 ^ 1'b0 ;
  assign n40121 = n9689 & n40120 ;
  assign n40122 = n40121 ^ n32027 ^ n1284 ;
  assign n40123 = n14593 | n18159 ;
  assign n40124 = ( n1362 & n21822 ) | ( n1362 & ~n30055 ) | ( n21822 & ~n30055 ) ;
  assign n40125 = ( ~n12324 & n40123 ) | ( ~n12324 & n40124 ) | ( n40123 & n40124 ) ;
  assign n40126 = n40125 ^ n4595 ^ 1'b0 ;
  assign n40127 = n5953 & n9586 ;
  assign n40128 = n40127 ^ x84 ^ 1'b0 ;
  assign n40129 = ( n29095 & n32285 ) | ( n29095 & n40128 ) | ( n32285 & n40128 ) ;
  assign n40131 = ( n1011 & n4593 ) | ( n1011 & n9844 ) | ( n4593 & n9844 ) ;
  assign n40130 = n258 & ~n5911 ;
  assign n40132 = n40131 ^ n40130 ^ n26461 ;
  assign n40133 = n7285 ^ n6424 ^ n1640 ;
  assign n40137 = n3333 & n9623 ;
  assign n40138 = n40137 ^ n33748 ^ 1'b0 ;
  assign n40134 = ~n14451 & n40112 ;
  assign n40135 = n17853 & n40134 ;
  assign n40136 = n24543 | n40135 ;
  assign n40139 = n40138 ^ n40136 ^ n5256 ;
  assign n40143 = n20008 ^ n1046 ^ 1'b0 ;
  assign n40144 = n1004 & n40143 ;
  assign n40140 = x212 & n13017 ;
  assign n40141 = ~n4111 & n10570 ;
  assign n40142 = ( x74 & n40140 ) | ( x74 & n40141 ) | ( n40140 & n40141 ) ;
  assign n40145 = n40144 ^ n40142 ^ n18969 ;
  assign n40146 = n2905 & ~n3703 ;
  assign n40147 = n29526 | n40146 ;
  assign n40148 = n40147 ^ n4050 ^ 1'b0 ;
  assign n40149 = n34409 ^ n24924 ^ 1'b0 ;
  assign n40150 = ~n40148 & n40149 ;
  assign n40151 = n35720 ^ n3879 ^ 1'b0 ;
  assign n40152 = n33438 ^ n9513 ^ n6275 ;
  assign n40153 = n21365 | n37830 ;
  assign n40154 = n25973 | n40153 ;
  assign n40155 = n20367 ^ n6748 ^ n4121 ;
  assign n40156 = ~n24131 & n40155 ;
  assign n40157 = n40154 & n40156 ;
  assign n40158 = n27848 ^ n787 ^ 1'b0 ;
  assign n40159 = n18730 ^ n17792 ^ 1'b0 ;
  assign n40160 = n40158 & n40159 ;
  assign n40161 = n33715 ^ n17737 ^ n8677 ;
  assign n40162 = n40161 ^ n34145 ^ 1'b0 ;
  assign n40163 = n1710 & n8264 ;
  assign n40164 = n40163 ^ n9271 ^ 1'b0 ;
  assign n40165 = ( ~n11679 & n13271 ) | ( ~n11679 & n16884 ) | ( n13271 & n16884 ) ;
  assign n40166 = n40165 ^ n19451 ^ n5003 ;
  assign n40167 = ~n40164 & n40166 ;
  assign n40169 = n7238 & ~n26715 ;
  assign n40170 = n40169 ^ n20081 ^ 1'b0 ;
  assign n40168 = n287 | n16032 ;
  assign n40171 = n40170 ^ n40168 ^ n7172 ;
  assign n40172 = n19080 | n26352 ;
  assign n40173 = n40172 ^ n17225 ^ 1'b0 ;
  assign n40174 = ( n10254 & ~n16593 ) | ( n10254 & n25584 ) | ( ~n16593 & n25584 ) ;
  assign n40175 = ( n13722 & n14497 ) | ( n13722 & n40174 ) | ( n14497 & n40174 ) ;
  assign n40176 = n33910 ^ n3223 ^ 1'b0 ;
  assign n40177 = n16125 & n40176 ;
  assign n40181 = ( n3047 & ~n11730 ) | ( n3047 & n12485 ) | ( ~n11730 & n12485 ) ;
  assign n40178 = ( n5724 & ~n10833 ) | ( n5724 & n21298 ) | ( ~n10833 & n21298 ) ;
  assign n40179 = ( n8686 & n11316 ) | ( n8686 & ~n40178 ) | ( n11316 & ~n40178 ) ;
  assign n40180 = ~n15016 & n40179 ;
  assign n40182 = n40181 ^ n40180 ^ 1'b0 ;
  assign n40183 = n10297 ^ n9275 ^ n1298 ;
  assign n40184 = n35922 & n40183 ;
  assign n40185 = ~n14777 & n37086 ;
  assign n40186 = x239 & ~n2024 ;
  assign n40187 = n40186 ^ n12906 ^ 1'b0 ;
  assign n40188 = ( n17560 & n23612 ) | ( n17560 & ~n40187 ) | ( n23612 & ~n40187 ) ;
  assign n40189 = n20808 ^ n7820 ^ n2973 ;
  assign n40190 = n14873 & n17874 ;
  assign n40191 = n1971 & n40190 ;
  assign n40192 = n24934 | n40191 ;
  assign n40193 = n35010 ^ n31497 ^ n10870 ;
  assign n40194 = ( ~n40189 & n40192 ) | ( ~n40189 & n40193 ) | ( n40192 & n40193 ) ;
  assign n40195 = n13194 ^ n5885 ^ 1'b0 ;
  assign n40196 = ( n12175 & n25288 ) | ( n12175 & n40195 ) | ( n25288 & n40195 ) ;
  assign n40197 = n40196 ^ n27237 ^ n26339 ;
  assign n40198 = n28494 ^ n3560 ^ 1'b0 ;
  assign n40199 = n20571 | n40198 ;
  assign n40200 = ( n7553 & n16910 ) | ( n7553 & ~n40199 ) | ( n16910 & ~n40199 ) ;
  assign n40201 = ( n7057 & n9402 ) | ( n7057 & n38210 ) | ( n9402 & n38210 ) ;
  assign n40202 = ( n15770 & n16560 ) | ( n15770 & n16935 ) | ( n16560 & n16935 ) ;
  assign n40203 = ( n20114 & n40201 ) | ( n20114 & ~n40202 ) | ( n40201 & ~n40202 ) ;
  assign n40204 = n23681 ^ n9050 ^ n2123 ;
  assign n40205 = n40204 ^ n24565 ^ x236 ;
  assign n40206 = n14772 | n25444 ;
  assign n40207 = n40206 ^ n29921 ^ 1'b0 ;
  assign n40208 = n6026 & ~n40207 ;
  assign n40209 = ~n40205 & n40208 ;
  assign n40210 = n1301 | n40209 ;
  assign n40211 = n40203 & ~n40210 ;
  assign n40212 = n14100 ^ n8024 ^ n7830 ;
  assign n40213 = n7439 & ~n40212 ;
  assign n40214 = n40213 ^ n16145 ^ 1'b0 ;
  assign n40215 = n5469 | n22106 ;
  assign n40216 = ( n3224 & n8887 ) | ( n3224 & n22809 ) | ( n8887 & n22809 ) ;
  assign n40217 = n40216 ^ n21211 ^ 1'b0 ;
  assign n40218 = n16632 | n40217 ;
  assign n40219 = n38311 ^ n16414 ^ n14606 ;
  assign n40220 = ( n32964 & n40218 ) | ( n32964 & n40219 ) | ( n40218 & n40219 ) ;
  assign n40223 = ~n9455 & n25486 ;
  assign n40222 = n6488 | n6517 ;
  assign n40221 = n614 & n36953 ;
  assign n40224 = n40223 ^ n40222 ^ n40221 ;
  assign n40225 = n14987 ^ n3796 ^ 1'b0 ;
  assign n40226 = x211 & ~n40225 ;
  assign n40227 = n15347 | n18363 ;
  assign n40228 = n12536 & ~n40227 ;
  assign n40229 = n14552 & n40228 ;
  assign n40230 = ( n8876 & ~n14544 ) | ( n8876 & n40229 ) | ( ~n14544 & n40229 ) ;
  assign n40231 = n40230 ^ n16887 ^ 1'b0 ;
  assign n40232 = ~n22059 & n40231 ;
  assign n40233 = ( ~n6031 & n6157 ) | ( ~n6031 & n12063 ) | ( n6157 & n12063 ) ;
  assign n40234 = n40233 ^ n39203 ^ 1'b0 ;
  assign n40235 = n40234 ^ n31400 ^ 1'b0 ;
  assign n40236 = n25845 & ~n29714 ;
  assign n40237 = n34709 ^ n13134 ^ 1'b0 ;
  assign n40238 = n20984 ^ n10800 ^ 1'b0 ;
  assign n40239 = n13163 | n37654 ;
  assign n40240 = n14555 & ~n40239 ;
  assign n40241 = n29243 ^ n13755 ^ 1'b0 ;
  assign n40242 = ( n35382 & n40240 ) | ( n35382 & ~n40241 ) | ( n40240 & ~n40241 ) ;
  assign n40243 = n29198 | n40242 ;
  assign n40244 = ~n28232 & n35003 ;
  assign n40245 = ~n7118 & n28238 ;
  assign n40246 = n17673 ^ n2727 ^ 1'b0 ;
  assign n40247 = n40246 ^ n4311 ^ 1'b0 ;
  assign n40248 = n18867 & n40247 ;
  assign n40249 = n9956 | n27154 ;
  assign n40250 = n40249 ^ n21096 ^ 1'b0 ;
  assign n40251 = n33262 ^ n24975 ^ n11686 ;
  assign n40252 = n37608 & ~n40251 ;
  assign n40253 = ( n27078 & ~n27459 ) | ( n27078 & n34246 ) | ( ~n27459 & n34246 ) ;
  assign n40254 = ( ~n3497 & n15269 ) | ( ~n3497 & n40253 ) | ( n15269 & n40253 ) ;
  assign n40257 = n40039 ^ n36379 ^ n5076 ;
  assign n40258 = ~n2591 & n6113 ;
  assign n40259 = n40257 & n40258 ;
  assign n40255 = n16990 ^ n10697 ^ 1'b0 ;
  assign n40256 = n17391 & n40255 ;
  assign n40260 = n40259 ^ n40256 ^ n28228 ;
  assign n40261 = n37432 ^ n8299 ^ 1'b0 ;
  assign n40262 = n3967 & ~n22891 ;
  assign n40263 = ~n7244 & n40262 ;
  assign n40264 = ~n5725 & n26405 ;
  assign n40265 = n13764 & n40264 ;
  assign n40266 = n40265 ^ n14465 ^ 1'b0 ;
  assign n40267 = n38413 ^ n23988 ^ 1'b0 ;
  assign n40268 = n10472 & n40267 ;
  assign n40269 = ( ~n4293 & n8369 ) | ( ~n4293 & n39993 ) | ( n8369 & n39993 ) ;
  assign n40270 = ( ~n826 & n27763 ) | ( ~n826 & n32543 ) | ( n27763 & n32543 ) ;
  assign n40271 = n11494 ^ n9365 ^ n1325 ;
  assign n40272 = ( n11425 & n14861 ) | ( n11425 & ~n40271 ) | ( n14861 & ~n40271 ) ;
  assign n40273 = n40272 ^ n16205 ^ 1'b0 ;
  assign n40274 = n25841 ^ n22320 ^ n1235 ;
  assign n40275 = n40274 ^ n7577 ^ 1'b0 ;
  assign n40276 = n13674 & n40275 ;
  assign n40277 = n10607 | n14741 ;
  assign n40278 = n40277 ^ n10571 ^ 1'b0 ;
  assign n40279 = n1050 | n27758 ;
  assign n40280 = n40278 & ~n40279 ;
  assign n40281 = n35719 ^ n35673 ^ n2183 ;
  assign n40282 = n10268 | n40281 ;
  assign n40283 = n39677 ^ n29587 ^ n19661 ;
  assign n40284 = ~n596 & n18445 ;
  assign n40285 = ~n775 & n40284 ;
  assign n40286 = n40146 ^ n10722 ^ 1'b0 ;
  assign n40287 = ~n40285 & n40286 ;
  assign n40288 = ( ~n12965 & n30315 ) | ( ~n12965 & n40287 ) | ( n30315 & n40287 ) ;
  assign n40289 = n13958 ^ n1293 ^ 1'b0 ;
  assign n40291 = n31180 & ~n40011 ;
  assign n40290 = n10558 | n24512 ;
  assign n40292 = n40291 ^ n40290 ^ 1'b0 ;
  assign n40293 = n40292 ^ x38 ^ 1'b0 ;
  assign n40294 = ( n40288 & ~n40289 ) | ( n40288 & n40293 ) | ( ~n40289 & n40293 ) ;
  assign n40295 = n37660 ^ n11117 ^ n4488 ;
  assign n40296 = n20214 & n29930 ;
  assign n40297 = n40296 ^ n26589 ^ 1'b0 ;
  assign n40298 = n10725 & ~n40297 ;
  assign n40299 = n40298 ^ n18191 ^ n11107 ;
  assign n40300 = n20232 & n24048 ;
  assign n40301 = n4776 | n5867 ;
  assign n40302 = n40301 ^ n3972 ^ 1'b0 ;
  assign n40303 = n15286 & n20608 ;
  assign n40304 = n17987 & n40303 ;
  assign n40305 = n37887 ^ n30217 ^ n2696 ;
  assign n40306 = n40305 ^ n38388 ^ n26171 ;
  assign n40307 = n40306 ^ n4488 ^ 1'b0 ;
  assign n40308 = n40304 | n40307 ;
  assign n40309 = n11406 ^ n8062 ^ 1'b0 ;
  assign n40310 = n2615 & n40309 ;
  assign n40311 = n40310 ^ n8319 ^ 1'b0 ;
  assign n40312 = n518 | n23694 ;
  assign n40313 = n40311 & ~n40312 ;
  assign n40314 = ( n18491 & n37361 ) | ( n18491 & ~n40313 ) | ( n37361 & ~n40313 ) ;
  assign n40315 = n33001 ^ n14193 ^ n4783 ;
  assign n40320 = n12735 | n14358 ;
  assign n40321 = n2443 | n40320 ;
  assign n40316 = n1388 & n8508 ;
  assign n40317 = ( ~n20540 & n29020 ) | ( ~n20540 & n30373 ) | ( n29020 & n30373 ) ;
  assign n40318 = n40316 & ~n40317 ;
  assign n40319 = ( n7704 & n19711 ) | ( n7704 & n40318 ) | ( n19711 & n40318 ) ;
  assign n40322 = n40321 ^ n40319 ^ n34417 ;
  assign n40323 = n22297 ^ n9132 ^ x85 ;
  assign n40324 = ( n22742 & ~n32372 ) | ( n22742 & n40323 ) | ( ~n32372 & n40323 ) ;
  assign n40325 = ( n10842 & n35454 ) | ( n10842 & n40324 ) | ( n35454 & n40324 ) ;
  assign n40326 = n2053 | n12046 ;
  assign n40327 = n1997 & ~n5818 ;
  assign n40328 = ~n17797 & n40327 ;
  assign n40329 = ( ~n25364 & n28356 ) | ( ~n25364 & n37272 ) | ( n28356 & n37272 ) ;
  assign n40330 = ~n20355 & n36813 ;
  assign n40331 = n17104 & ~n19584 ;
  assign n40332 = n1667 | n40331 ;
  assign n40333 = n24188 & ~n40332 ;
  assign n40334 = ( n4414 & n18850 ) | ( n4414 & n40333 ) | ( n18850 & n40333 ) ;
  assign n40335 = n12783 | n27184 ;
  assign n40336 = n1390 & ~n34863 ;
  assign n40337 = ~n17912 & n40336 ;
  assign n40338 = ( ~n5017 & n9724 ) | ( ~n5017 & n26115 ) | ( n9724 & n26115 ) ;
  assign n40339 = ~n20073 & n40338 ;
  assign n40340 = n40337 & n40339 ;
  assign n40341 = n18494 ^ n950 ^ n500 ;
  assign n40342 = ( n13384 & n15567 ) | ( n13384 & n40341 ) | ( n15567 & n40341 ) ;
  assign n40343 = n39382 ^ n9584 ^ n7727 ;
  assign n40344 = ( n33349 & n40342 ) | ( n33349 & ~n40343 ) | ( n40342 & ~n40343 ) ;
  assign n40345 = n11296 & n20484 ;
  assign n40346 = n40345 ^ n13838 ^ n1382 ;
  assign n40348 = n14108 ^ n9616 ^ n3692 ;
  assign n40347 = ~n11594 & n31822 ;
  assign n40349 = n40348 ^ n40347 ^ n9837 ;
  assign n40350 = n25466 ^ n19725 ^ 1'b0 ;
  assign n40351 = n30345 ^ n24811 ^ n21395 ;
  assign n40352 = n18728 | n40351 ;
  assign n40353 = n3432 & n15301 ;
  assign n40354 = ( n11431 & n15917 ) | ( n11431 & ~n40353 ) | ( n15917 & ~n40353 ) ;
  assign n40355 = n15899 ^ n3666 ^ 1'b0 ;
  assign n40356 = n29227 ^ n16460 ^ 1'b0 ;
  assign n40357 = ~n2922 & n40356 ;
  assign n40358 = n32039 ^ n21638 ^ 1'b0 ;
  assign n40359 = n40357 & ~n40358 ;
  assign n40360 = n7120 | n13481 ;
  assign n40361 = n40360 ^ n11467 ^ 1'b0 ;
  assign n40363 = ( n9784 & n14740 ) | ( n9784 & ~n25959 ) | ( n14740 & ~n25959 ) ;
  assign n40362 = n22128 | n33123 ;
  assign n40364 = n40363 ^ n40362 ^ 1'b0 ;
  assign n40365 = n35629 | n40364 ;
  assign n40366 = n40365 ^ n17490 ^ 1'b0 ;
  assign n40371 = n1703 & n10867 ;
  assign n40372 = n7948 & n40371 ;
  assign n40373 = n40372 ^ n5546 ^ n3814 ;
  assign n40369 = ( ~n15617 & n18298 ) | ( ~n15617 & n24843 ) | ( n18298 & n24843 ) ;
  assign n40370 = n40369 ^ n530 ^ 1'b0 ;
  assign n40367 = ~n18385 & n36182 ;
  assign n40368 = n40367 ^ n37244 ^ 1'b0 ;
  assign n40374 = n40373 ^ n40370 ^ n40368 ;
  assign n40375 = ( n6905 & n23669 ) | ( n6905 & n28500 ) | ( n23669 & n28500 ) ;
  assign n40376 = ( n32815 & n35846 ) | ( n32815 & n40375 ) | ( n35846 & n40375 ) ;
  assign n40377 = ( x77 & n14824 ) | ( x77 & ~n16244 ) | ( n14824 & ~n16244 ) ;
  assign n40378 = n7867 & ~n40377 ;
  assign n40379 = n13279 ^ n9944 ^ 1'b0 ;
  assign n40380 = x186 & n22662 ;
  assign n40381 = n40380 ^ n16188 ^ 1'b0 ;
  assign n40382 = n40381 ^ n14670 ^ 1'b0 ;
  assign n40383 = n20864 ^ n17955 ^ 1'b0 ;
  assign n40384 = n40382 & n40383 ;
  assign n40385 = n17567 ^ n10073 ^ n5256 ;
  assign n40386 = ~n1213 & n40385 ;
  assign n40387 = n18477 ^ n15508 ^ 1'b0 ;
  assign n40388 = n27456 & ~n34753 ;
  assign n40389 = n40388 ^ n39691 ^ n21485 ;
  assign n40390 = ( n28564 & ~n29060 ) | ( n28564 & n38205 ) | ( ~n29060 & n38205 ) ;
  assign n40393 = n22921 ^ n15378 ^ n4734 ;
  assign n40392 = ( n8128 & ~n9443 ) | ( n8128 & n10425 ) | ( ~n9443 & n10425 ) ;
  assign n40391 = n25769 ^ n13510 ^ 1'b0 ;
  assign n40394 = n40393 ^ n40392 ^ n40391 ;
  assign n40395 = ( ~n4975 & n15077 ) | ( ~n4975 & n37113 ) | ( n15077 & n37113 ) ;
  assign n40396 = n40395 ^ n38033 ^ 1'b0 ;
  assign n40397 = n40396 ^ n30633 ^ n12353 ;
  assign n40398 = ~n13125 & n27337 ;
  assign n40399 = n40398 ^ n37856 ^ 1'b0 ;
  assign n40400 = n27544 ^ n15610 ^ 1'b0 ;
  assign n40401 = ~n25143 & n40400 ;
  assign n40402 = n17195 ^ n12063 ^ 1'b0 ;
  assign n40403 = n40402 ^ n21289 ^ n16336 ;
  assign n40404 = n30342 ^ n27623 ^ n16046 ;
  assign n40405 = n33043 ^ n9571 ^ 1'b0 ;
  assign n40406 = n40405 ^ n29267 ^ n6863 ;
  assign n40407 = n16933 ^ n1156 ^ 1'b0 ;
  assign n40408 = n10921 & ~n40407 ;
  assign n40409 = n15446 ^ n8373 ^ 1'b0 ;
  assign n40410 = ~n14506 & n40409 ;
  assign n40411 = n5268 & n7974 ;
  assign n40412 = n13791 & n40411 ;
  assign n40413 = n40412 ^ n38447 ^ n7993 ;
  assign n40414 = ( n40408 & n40410 ) | ( n40408 & n40413 ) | ( n40410 & n40413 ) ;
  assign n40420 = n2848 & ~n9724 ;
  assign n40421 = n5470 ^ n5339 ^ 1'b0 ;
  assign n40422 = n16160 & n40421 ;
  assign n40423 = ~n13719 & n40422 ;
  assign n40424 = ~n40420 & n40423 ;
  assign n40415 = n22162 ^ n21448 ^ n18398 ;
  assign n40416 = n35493 ^ n4407 ^ 1'b0 ;
  assign n40417 = n40415 | n40416 ;
  assign n40418 = n40417 ^ n39399 ^ n38283 ;
  assign n40419 = n14414 | n40418 ;
  assign n40425 = n40424 ^ n40419 ^ 1'b0 ;
  assign n40426 = ( n9017 & ~n14373 ) | ( n9017 & n19807 ) | ( ~n14373 & n19807 ) ;
  assign n40427 = n40426 ^ n21986 ^ n16192 ;
  assign n40428 = n40427 ^ n16097 ^ 1'b0 ;
  assign n40429 = n4075 | n8999 ;
  assign n40430 = n40429 ^ n28815 ^ 1'b0 ;
  assign n40431 = n20409 ^ n3922 ^ 1'b0 ;
  assign n40432 = n11975 ^ n10363 ^ n1896 ;
  assign n40433 = n40432 ^ n18421 ^ 1'b0 ;
  assign n40434 = ( n12019 & ~n40431 ) | ( n12019 & n40433 ) | ( ~n40431 & n40433 ) ;
  assign n40435 = n9154 ^ n5186 ^ 1'b0 ;
  assign n40436 = n40435 ^ n37469 ^ n4196 ;
  assign n40437 = n2933 | n30982 ;
  assign n40441 = n16225 & n26992 ;
  assign n40442 = ~n16832 & n40441 ;
  assign n40439 = n12616 ^ n12216 ^ n7650 ;
  assign n40440 = n26443 & ~n40439 ;
  assign n40443 = n40442 ^ n40440 ^ 1'b0 ;
  assign n40444 = n40443 ^ n14728 ^ 1'b0 ;
  assign n40438 = ~n7306 & n27964 ;
  assign n40445 = n40444 ^ n40438 ^ 1'b0 ;
  assign n40446 = n17356 ^ n16635 ^ x253 ;
  assign n40447 = n40446 ^ n26789 ^ n12852 ;
  assign n40448 = n7445 | n35061 ;
  assign n40449 = n40448 ^ n14041 ^ 1'b0 ;
  assign n40450 = ( n16274 & ~n27200 ) | ( n16274 & n40449 ) | ( ~n27200 & n40449 ) ;
  assign n40451 = n40450 ^ n25266 ^ 1'b0 ;
  assign n40452 = ( n6065 & n8260 ) | ( n6065 & n18337 ) | ( n8260 & n18337 ) ;
  assign n40453 = ( x191 & ~n443 ) | ( x191 & n15552 ) | ( ~n443 & n15552 ) ;
  assign n40454 = ( n7591 & n34938 ) | ( n7591 & ~n40453 ) | ( n34938 & ~n40453 ) ;
  assign n40455 = n40454 ^ n16232 ^ 1'b0 ;
  assign n40456 = n13368 & ~n30375 ;
  assign n40457 = n8553 & ~n28924 ;
  assign n40458 = n6247 & ~n25112 ;
  assign n40459 = n16076 | n17024 ;
  assign n40460 = n40459 ^ n11675 ^ 1'b0 ;
  assign n40461 = ~n40458 & n40460 ;
  assign n40463 = n7792 & n17731 ;
  assign n40462 = n3947 | n5072 ;
  assign n40464 = n40463 ^ n40462 ^ n7779 ;
  assign n40465 = n1940 | n7424 ;
  assign n40466 = n40465 ^ n26596 ^ 1'b0 ;
  assign n40467 = n40464 | n40466 ;
  assign n40468 = n30846 ^ n25930 ^ n17803 ;
  assign n40469 = ( ~n3287 & n7887 ) | ( ~n3287 & n38750 ) | ( n7887 & n38750 ) ;
  assign n40470 = n21196 & ~n38016 ;
  assign n40471 = n26469 ^ n7680 ^ 1'b0 ;
  assign n40472 = ( n8297 & ~n16200 ) | ( n8297 & n30354 ) | ( ~n16200 & n30354 ) ;
  assign n40473 = ( n6831 & ~n12852 ) | ( n6831 & n20884 ) | ( ~n12852 & n20884 ) ;
  assign n40474 = n40473 ^ n28877 ^ 1'b0 ;
  assign n40475 = n40472 & n40474 ;
  assign n40476 = ( ~n11249 & n14100 ) | ( ~n11249 & n21945 ) | ( n14100 & n21945 ) ;
  assign n40477 = n33387 ^ n7098 ^ n6315 ;
  assign n40478 = n31037 ^ n21269 ^ n10490 ;
  assign n40479 = n40478 ^ n16367 ^ 1'b0 ;
  assign n40480 = ( ~n5715 & n40477 ) | ( ~n5715 & n40479 ) | ( n40477 & n40479 ) ;
  assign n40481 = n8929 ^ n2522 ^ n560 ;
  assign n40482 = n8213 ^ n5953 ^ 1'b0 ;
  assign n40483 = ~n40481 & n40482 ;
  assign n40484 = n30078 & ~n40483 ;
  assign n40485 = n297 | n8871 ;
  assign n40486 = n40485 ^ n39437 ^ 1'b0 ;
  assign n40487 = n16013 | n17440 ;
  assign n40488 = n40487 ^ n31130 ^ 1'b0 ;
  assign n40489 = n3509 & n12919 ;
  assign n40490 = n25158 ^ n10450 ^ 1'b0 ;
  assign n40491 = n40489 & n40490 ;
  assign n40492 = ( ~n7261 & n12895 ) | ( ~n7261 & n17421 ) | ( n12895 & n17421 ) ;
  assign n40493 = n40492 ^ n21529 ^ 1'b0 ;
  assign n40494 = ( n5218 & n8813 ) | ( n5218 & ~n17822 ) | ( n8813 & ~n17822 ) ;
  assign n40495 = n40494 ^ n5098 ^ 1'b0 ;
  assign n40496 = n40493 & n40495 ;
  assign n40497 = n30463 ^ n12818 ^ n3963 ;
  assign n40498 = n20650 ^ n2831 ^ 1'b0 ;
  assign n40499 = n20366 | n40498 ;
  assign n40500 = n40499 ^ n18592 ^ 1'b0 ;
  assign n40501 = n5824 & ~n10602 ;
  assign n40502 = ( n12578 & n26322 ) | ( n12578 & ~n40501 ) | ( n26322 & ~n40501 ) ;
  assign n40503 = ( n40497 & n40500 ) | ( n40497 & ~n40502 ) | ( n40500 & ~n40502 ) ;
  assign n40504 = ~n11003 & n28492 ;
  assign n40505 = n40504 ^ n18035 ^ 1'b0 ;
  assign n40506 = n40505 ^ n28992 ^ n8892 ;
  assign n40507 = n5075 & n30227 ;
  assign n40508 = n40507 ^ n18627 ^ 1'b0 ;
  assign n40509 = n40508 ^ n36575 ^ 1'b0 ;
  assign n40510 = n11681 ^ n1807 ^ 1'b0 ;
  assign n40511 = n40510 ^ n18911 ^ n17900 ;
  assign n40512 = n514 | n13596 ;
  assign n40513 = n40512 ^ n28795 ^ 1'b0 ;
  assign n40514 = n26720 ^ n26433 ^ n13875 ;
  assign n40515 = ( ~n40511 & n40513 ) | ( ~n40511 & n40514 ) | ( n40513 & n40514 ) ;
  assign n40516 = ~n3458 & n4991 ;
  assign n40518 = n10173 ^ n3809 ^ 1'b0 ;
  assign n40517 = n3832 & n17526 ;
  assign n40519 = n40518 ^ n40517 ^ 1'b0 ;
  assign n40520 = ( n17669 & n24864 ) | ( n17669 & ~n32495 ) | ( n24864 & ~n32495 ) ;
  assign n40521 = n40520 ^ n32372 ^ 1'b0 ;
  assign n40522 = n7832 & ~n40521 ;
  assign n40523 = ( n8826 & n27158 ) | ( n8826 & n40522 ) | ( n27158 & n40522 ) ;
  assign n40527 = n29862 | n31017 ;
  assign n40524 = n22046 & n27449 ;
  assign n40525 = ~n15184 & n15781 ;
  assign n40526 = n40524 & ~n40525 ;
  assign n40528 = n40527 ^ n40526 ^ n998 ;
  assign n40529 = n37138 ^ n27680 ^ 1'b0 ;
  assign n40530 = ( ~n14324 & n17412 ) | ( ~n14324 & n39385 ) | ( n17412 & n39385 ) ;
  assign n40531 = ( n8964 & n10659 ) | ( n8964 & ~n11060 ) | ( n10659 & ~n11060 ) ;
  assign n40532 = ~n15112 & n40531 ;
  assign n40533 = x138 & n32815 ;
  assign n40534 = ~n38979 & n40533 ;
  assign n40535 = n40534 ^ n8003 ^ 1'b0 ;
  assign n40536 = n39125 ^ n32438 ^ n25737 ;
  assign n40537 = n30149 | n40536 ;
  assign n40538 = n12388 | n13399 ;
  assign n40539 = n40538 ^ n3653 ^ 1'b0 ;
  assign n40540 = n4078 ^ n2110 ^ 1'b0 ;
  assign n40541 = n36716 & n40540 ;
  assign n40542 = n40539 & ~n40541 ;
  assign n40543 = n3799 & ~n10027 ;
  assign n40544 = ~n16999 & n40543 ;
  assign n40545 = n399 & n34496 ;
  assign n40546 = n40545 ^ n25423 ^ n11043 ;
  assign n40547 = ~n421 & n13593 ;
  assign n40548 = n40547 ^ x25 ^ 1'b0 ;
  assign n40549 = ( n15378 & n20767 ) | ( n15378 & n40548 ) | ( n20767 & n40548 ) ;
  assign n40550 = ( ~n13543 & n37248 ) | ( ~n13543 & n40549 ) | ( n37248 & n40549 ) ;
  assign n40551 = n14232 ^ n2296 ^ 1'b0 ;
  assign n40552 = n24942 ^ n4619 ^ n2416 ;
  assign n40553 = n17327 ^ n4397 ^ 1'b0 ;
  assign n40554 = n40552 | n40553 ;
  assign n40555 = ( n34504 & n40551 ) | ( n34504 & n40554 ) | ( n40551 & n40554 ) ;
  assign n40556 = ( ~n13097 & n23517 ) | ( ~n13097 & n31314 ) | ( n23517 & n31314 ) ;
  assign n40557 = ( n12841 & n34683 ) | ( n12841 & ~n40556 ) | ( n34683 & ~n40556 ) ;
  assign n40558 = ( n5585 & n5792 ) | ( n5585 & n29844 ) | ( n5792 & n29844 ) ;
  assign n40559 = n15338 ^ n9741 ^ n5728 ;
  assign n40560 = n40559 ^ n21153 ^ n19921 ;
  assign n40561 = n6198 & n6660 ;
  assign n40562 = n5205 | n23192 ;
  assign n40563 = n40561 | n40562 ;
  assign n40564 = ( n37054 & n40560 ) | ( n37054 & n40563 ) | ( n40560 & n40563 ) ;
  assign n40565 = n982 | n40564 ;
  assign n40566 = n24003 & n27222 ;
  assign n40567 = ~n18635 & n39368 ;
  assign n40568 = ~n40566 & n40567 ;
  assign n40569 = ( n11605 & n14279 ) | ( n11605 & ~n20017 ) | ( n14279 & ~n20017 ) ;
  assign n40570 = n40569 ^ n36358 ^ n18191 ;
  assign n40571 = ~n22807 & n40570 ;
  assign n40572 = n40571 ^ n1098 ^ 1'b0 ;
  assign n40573 = n14657 ^ n12143 ^ 1'b0 ;
  assign n40574 = n29227 & n40573 ;
  assign n40575 = ~n10097 & n40574 ;
  assign n40576 = n8791 & n40575 ;
  assign n40577 = n20279 & ~n40576 ;
  assign n40578 = n34985 ^ n27765 ^ n14175 ;
  assign n40579 = n15852 ^ n8423 ^ n3273 ;
  assign n40580 = n10426 & ~n40579 ;
  assign n40581 = ( n15165 & n15456 ) | ( n15165 & ~n24080 ) | ( n15456 & ~n24080 ) ;
  assign n40582 = n23476 & ~n40581 ;
  assign n40583 = n9741 ^ n5446 ^ n459 ;
  assign n40584 = n553 | n40583 ;
  assign n40585 = n40584 ^ n13286 ^ 1'b0 ;
  assign n40586 = ( ~n40580 & n40582 ) | ( ~n40580 & n40585 ) | ( n40582 & n40585 ) ;
  assign n40587 = ( ~n4569 & n11378 ) | ( ~n4569 & n40586 ) | ( n11378 & n40586 ) ;
  assign n40588 = n40587 ^ n27513 ^ 1'b0 ;
  assign n40589 = n39947 ^ n29921 ^ n15676 ;
  assign n40591 = ( ~x164 & n19797 ) | ( ~x164 & n21780 ) | ( n19797 & n21780 ) ;
  assign n40590 = ( ~n18339 & n19518 ) | ( ~n18339 & n33913 ) | ( n19518 & n33913 ) ;
  assign n40592 = n40591 ^ n40590 ^ n4011 ;
  assign n40593 = n37592 ^ n9686 ^ 1'b0 ;
  assign n40594 = ~n21997 & n40593 ;
  assign n40595 = n32609 ^ n17155 ^ n11335 ;
  assign n40596 = n40595 ^ n20840 ^ n7906 ;
  assign n40597 = n5537 & ~n40596 ;
  assign n40598 = n15175 & n16672 ;
  assign n40599 = ( n13455 & n18549 ) | ( n13455 & ~n23742 ) | ( n18549 & ~n23742 ) ;
  assign n40600 = ( n7469 & ~n11269 ) | ( n7469 & n40599 ) | ( ~n11269 & n40599 ) ;
  assign n40601 = ( n7518 & n14870 ) | ( n7518 & ~n16903 ) | ( n14870 & ~n16903 ) ;
  assign n40602 = ( n3026 & n10849 ) | ( n3026 & n24258 ) | ( n10849 & n24258 ) ;
  assign n40603 = n7098 & n17888 ;
  assign n40604 = ~n11259 & n40603 ;
  assign n40605 = n40604 ^ n33707 ^ n5088 ;
  assign n40606 = ( n37986 & n40602 ) | ( n37986 & n40605 ) | ( n40602 & n40605 ) ;
  assign n40607 = ( x192 & n1600 ) | ( x192 & n6077 ) | ( n1600 & n6077 ) ;
  assign n40608 = n40607 ^ n30549 ^ n1511 ;
  assign n40609 = n40608 ^ n26550 ^ n7543 ;
  assign n40610 = n32812 ^ n27833 ^ 1'b0 ;
  assign n40611 = ~n27316 & n40610 ;
  assign n40612 = n15452 | n29951 ;
  assign n40613 = n19966 & ~n40612 ;
  assign n40614 = n16660 ^ n14186 ^ n10240 ;
  assign n40615 = n37027 ^ n15372 ^ 1'b0 ;
  assign n40616 = n40614 | n40615 ;
  assign n40617 = n36350 ^ n6100 ^ 1'b0 ;
  assign n40618 = n5387 & ~n40617 ;
  assign n40619 = n23929 | n25881 ;
  assign n40620 = n23046 & ~n40619 ;
  assign n40621 = n4662 & ~n40620 ;
  assign n40622 = ~n40618 & n40621 ;
  assign n40624 = ( n1171 & n3212 ) | ( n1171 & n6873 ) | ( n3212 & n6873 ) ;
  assign n40623 = ~n7827 & n19190 ;
  assign n40625 = n40624 ^ n40623 ^ n23711 ;
  assign n40626 = n40625 ^ n30175 ^ n15024 ;
  assign n40627 = ( n2229 & n20108 ) | ( n2229 & n40626 ) | ( n20108 & n40626 ) ;
  assign n40629 = ~n1195 & n4063 ;
  assign n40630 = n40629 ^ n3898 ^ 1'b0 ;
  assign n40628 = ( x97 & n10441 ) | ( x97 & ~n24767 ) | ( n10441 & ~n24767 ) ;
  assign n40631 = n40630 ^ n40628 ^ n14507 ;
  assign n40636 = ( n4825 & n6033 ) | ( n4825 & ~n9665 ) | ( n6033 & ~n9665 ) ;
  assign n40637 = n40636 ^ n30133 ^ n29757 ;
  assign n40638 = n18804 & ~n40637 ;
  assign n40632 = ( n2056 & n31355 ) | ( n2056 & n35923 ) | ( n31355 & n35923 ) ;
  assign n40633 = ( ~n13865 & n14150 ) | ( ~n13865 & n40632 ) | ( n14150 & n40632 ) ;
  assign n40634 = n8588 & n40633 ;
  assign n40635 = n40634 ^ n13240 ^ 1'b0 ;
  assign n40639 = n40638 ^ n40635 ^ n30883 ;
  assign n40640 = n4535 ^ n705 ^ 1'b0 ;
  assign n40641 = ~n7887 & n9581 ;
  assign n40642 = ~n25281 & n40641 ;
  assign n40643 = ( n16225 & n40640 ) | ( n16225 & ~n40642 ) | ( n40640 & ~n40642 ) ;
  assign n40644 = n24237 ^ n19933 ^ n9599 ;
  assign n40645 = ( n8336 & ~n23873 ) | ( n8336 & n40644 ) | ( ~n23873 & n40644 ) ;
  assign n40646 = n10722 | n11364 ;
  assign n40647 = n14186 & n40646 ;
  assign n40648 = n40647 ^ n2464 ^ 1'b0 ;
  assign n40649 = ( n12086 & n15225 ) | ( n12086 & n21780 ) | ( n15225 & n21780 ) ;
  assign n40650 = n21388 & n40649 ;
  assign n40651 = ~n25893 & n40650 ;
  assign n40652 = n33757 ^ n33149 ^ n25723 ;
  assign n40653 = n2853 & ~n40652 ;
  assign n40654 = n40653 ^ n25342 ^ 1'b0 ;
  assign n40655 = ~n25282 & n40654 ;
  assign n40656 = ~n35609 & n40655 ;
  assign n40657 = n37167 ^ n12712 ^ n11732 ;
  assign n40658 = ( n3740 & n18752 ) | ( n3740 & n22632 ) | ( n18752 & n22632 ) ;
  assign n40659 = n40658 ^ n9681 ^ n289 ;
  assign n40660 = n40659 ^ n30721 ^ n9018 ;
  assign n40661 = ( n897 & ~n10687 ) | ( n897 & n11901 ) | ( ~n10687 & n11901 ) ;
  assign n40662 = n22449 | n40661 ;
  assign n40665 = ~n2154 & n28242 ;
  assign n40666 = n17555 ^ n7661 ^ n7087 ;
  assign n40667 = ( n20037 & n40665 ) | ( n20037 & ~n40666 ) | ( n40665 & ~n40666 ) ;
  assign n40663 = n4359 & n5998 ;
  assign n40664 = n40663 ^ n25276 ^ 1'b0 ;
  assign n40668 = n40667 ^ n40664 ^ n23594 ;
  assign n40669 = n9365 & n15513 ;
  assign n40670 = n2964 & n40669 ;
  assign n40671 = n3235 | n14325 ;
  assign n40672 = ( n6901 & n40670 ) | ( n6901 & n40671 ) | ( n40670 & n40671 ) ;
  assign n40673 = n16449 | n40672 ;
  assign n40674 = n21276 & n37554 ;
  assign n40675 = n34018 & n40674 ;
  assign n40676 = n6070 & ~n40675 ;
  assign n40677 = n40676 ^ n19413 ^ 1'b0 ;
  assign n40678 = n5700 & n23302 ;
  assign n40679 = n40678 ^ n11973 ^ 1'b0 ;
  assign n40680 = n20984 ^ n11856 ^ n4617 ;
  assign n40681 = n22408 & ~n40680 ;
  assign n40682 = n40681 ^ n27231 ^ 1'b0 ;
  assign n40683 = n39330 & n40682 ;
  assign n40684 = n40683 ^ n34740 ^ 1'b0 ;
  assign n40687 = ~n16972 & n26691 ;
  assign n40688 = ~n11901 & n40687 ;
  assign n40689 = n15098 | n20272 ;
  assign n40690 = n2751 & ~n40689 ;
  assign n40691 = n40690 ^ n5139 ^ 1'b0 ;
  assign n40692 = n40688 | n40691 ;
  assign n40685 = ( x13 & n4688 ) | ( x13 & ~n6815 ) | ( n4688 & ~n6815 ) ;
  assign n40686 = n39435 | n40685 ;
  assign n40693 = n40692 ^ n40686 ^ 1'b0 ;
  assign n40695 = n1727 | n6131 ;
  assign n40694 = n8354 ^ n5881 ^ 1'b0 ;
  assign n40696 = n40695 ^ n40694 ^ n20930 ;
  assign n40697 = n36928 ^ n13366 ^ 1'b0 ;
  assign n40698 = ~n19754 & n40697 ;
  assign n40699 = n22913 ^ n20190 ^ 1'b0 ;
  assign n40700 = n31048 & ~n40699 ;
  assign n40701 = n19394 & n40700 ;
  assign n40702 = n40701 ^ n15694 ^ 1'b0 ;
  assign n40704 = ( n1977 & ~n2002 ) | ( n1977 & n4137 ) | ( ~n2002 & n4137 ) ;
  assign n40705 = n14474 | n40704 ;
  assign n40703 = ~n1864 & n19527 ;
  assign n40706 = n40705 ^ n40703 ^ 1'b0 ;
  assign n40707 = ~n32514 & n40706 ;
  assign n40708 = ~n10197 & n11287 ;
  assign n40709 = n22146 & n40708 ;
  assign n40710 = n40709 ^ n23859 ^ n6564 ;
  assign n40711 = n11680 & ~n22717 ;
  assign n40712 = n40710 & n40711 ;
  assign n40713 = n29077 ^ n23575 ^ n15760 ;
  assign n40714 = n14922 & n26234 ;
  assign n40715 = n40714 ^ n23277 ^ n19725 ;
  assign n40716 = ( n9840 & n40713 ) | ( n9840 & ~n40715 ) | ( n40713 & ~n40715 ) ;
  assign n40717 = n28329 ^ n2271 ^ 1'b0 ;
  assign n40718 = n34146 ^ n14660 ^ x245 ;
  assign n40719 = n17462 | n20948 ;
  assign n40720 = n11635 & ~n40719 ;
  assign n40721 = n1169 | n28370 ;
  assign n40722 = n13893 | n40721 ;
  assign n40723 = n23320 & ~n40722 ;
  assign n40724 = n18708 | n23956 ;
  assign n40725 = n40724 ^ n21899 ^ 1'b0 ;
  assign n40726 = n23120 ^ n19247 ^ 1'b0 ;
  assign n40727 = n40726 ^ n14609 ^ n5502 ;
  assign n40728 = n40727 ^ n5651 ^ n4126 ;
  assign n40729 = n40728 ^ n10207 ^ 1'b0 ;
  assign n40730 = n40729 ^ n37297 ^ n35731 ;
  assign n40731 = ( n15482 & ~n18140 ) | ( n15482 & n24435 ) | ( ~n18140 & n24435 ) ;
  assign n40732 = n40731 ^ n26951 ^ 1'b0 ;
  assign n40733 = n8888 & ~n27950 ;
  assign n40734 = ~n40732 & n40733 ;
  assign n40735 = n40734 ^ n2301 ^ 1'b0 ;
  assign n40736 = n17129 ^ n11273 ^ 1'b0 ;
  assign n40737 = ~n10027 & n10222 ;
  assign n40738 = ~n40736 & n40737 ;
  assign n40739 = n7932 ^ n3228 ^ 1'b0 ;
  assign n40740 = ( n3616 & ~n40738 ) | ( n3616 & n40739 ) | ( ~n40738 & n40739 ) ;
  assign n40741 = ( n4841 & ~n21366 ) | ( n4841 & n30092 ) | ( ~n21366 & n30092 ) ;
  assign n40742 = x31 & ~n12007 ;
  assign n40743 = ( n1297 & ~n8302 ) | ( n1297 & n40742 ) | ( ~n8302 & n40742 ) ;
  assign n40744 = ~n8492 & n40743 ;
  assign n40745 = n11147 ^ n2735 ^ 1'b0 ;
  assign n40746 = ( ~n3760 & n40744 ) | ( ~n3760 & n40745 ) | ( n40744 & n40745 ) ;
  assign n40747 = n40746 ^ n2964 ^ 1'b0 ;
  assign n40748 = ( n36148 & n40741 ) | ( n36148 & ~n40747 ) | ( n40741 & ~n40747 ) ;
  assign n40749 = n40748 ^ n25042 ^ 1'b0 ;
  assign n40750 = ( n1888 & n28695 ) | ( n1888 & n31651 ) | ( n28695 & n31651 ) ;
  assign n40751 = n10990 & ~n40750 ;
  assign n40752 = n37383 ^ n22768 ^ n19818 ;
  assign n40753 = n4195 | n40752 ;
  assign n40754 = n9194 | n12559 ;
  assign n40755 = n29582 & ~n40754 ;
  assign n40756 = ( n11574 & n15035 ) | ( n11574 & ~n25766 ) | ( n15035 & ~n25766 ) ;
  assign n40757 = n40756 ^ n10653 ^ 1'b0 ;
  assign n40758 = n32147 | n34637 ;
  assign n40759 = n26430 ^ n11048 ^ 1'b0 ;
  assign n40760 = n40758 | n40759 ;
  assign n40761 = n40760 ^ n29812 ^ 1'b0 ;
  assign n40762 = n25203 ^ n18706 ^ n6846 ;
  assign n40763 = ( n2466 & n2751 ) | ( n2466 & ~n19045 ) | ( n2751 & ~n19045 ) ;
  assign n40764 = ( n1210 & n2090 ) | ( n1210 & n22286 ) | ( n2090 & n22286 ) ;
  assign n40765 = ~n12779 & n25329 ;
  assign n40766 = ~n40764 & n40765 ;
  assign n40767 = n40766 ^ n3036 ^ 1'b0 ;
  assign n40768 = x169 & n20665 ;
  assign n40769 = n40768 ^ n18409 ^ 1'b0 ;
  assign n40770 = n32273 & n40769 ;
  assign n40772 = n33454 ^ n17086 ^ 1'b0 ;
  assign n40773 = n40772 ^ n22577 ^ n20087 ;
  assign n40771 = ( n6731 & n9892 ) | ( n6731 & n26710 ) | ( n9892 & n26710 ) ;
  assign n40774 = n40773 ^ n40771 ^ n13546 ;
  assign n40775 = n4757 & ~n39469 ;
  assign n40776 = n40775 ^ n26736 ^ 1'b0 ;
  assign n40777 = n24849 | n40776 ;
  assign n40778 = n40774 & ~n40777 ;
  assign n40779 = n18340 | n40778 ;
  assign n40780 = n40393 | n40779 ;
  assign n40781 = n38880 ^ n17567 ^ 1'b0 ;
  assign n40782 = n23746 | n40781 ;
  assign n40783 = n6401 & ~n27237 ;
  assign n40784 = n8282 ^ x88 ^ 1'b0 ;
  assign n40785 = n40784 ^ n15773 ^ n10140 ;
  assign n40786 = n40785 ^ n23403 ^ 1'b0 ;
  assign n40787 = n6923 ^ n2526 ^ 1'b0 ;
  assign n40788 = ( n807 & ~n10215 ) | ( n807 & n40787 ) | ( ~n10215 & n40787 ) ;
  assign n40789 = ~n13848 & n40788 ;
  assign n40791 = ~n16053 & n20739 ;
  assign n40790 = ( x131 & n22091 ) | ( x131 & n22792 ) | ( n22091 & n22792 ) ;
  assign n40792 = n40791 ^ n40790 ^ 1'b0 ;
  assign n40793 = n14250 & ~n40792 ;
  assign n40794 = ~n5345 & n40793 ;
  assign n40795 = n20051 & n40794 ;
  assign n40796 = ~n31480 & n36728 ;
  assign n40797 = ~n6025 & n40796 ;
  assign n40798 = ( n12947 & ~n13899 ) | ( n12947 & n16381 ) | ( ~n13899 & n16381 ) ;
  assign n40799 = n15924 ^ n1351 ^ n318 ;
  assign n40800 = n3476 & n8982 ;
  assign n40801 = ~n40799 & n40800 ;
  assign n40802 = ( n16444 & n40798 ) | ( n16444 & ~n40801 ) | ( n40798 & ~n40801 ) ;
  assign n40803 = ( n1311 & ~n24254 ) | ( n1311 & n39383 ) | ( ~n24254 & n39383 ) ;
  assign n40804 = n3848 & ~n35544 ;
  assign n40805 = ~n13161 & n40804 ;
  assign n40806 = n40805 ^ n17369 ^ n6700 ;
  assign n40807 = n5454 & ~n23193 ;
  assign n40808 = ~n32047 & n40807 ;
  assign n40809 = ( n15323 & n40172 ) | ( n15323 & n40808 ) | ( n40172 & n40808 ) ;
  assign n40810 = n13515 ^ x61 ^ 1'b0 ;
  assign n40811 = n25160 ^ n946 ^ 1'b0 ;
  assign n40812 = n40811 ^ n16188 ^ 1'b0 ;
  assign n40813 = n13404 ^ n9275 ^ 1'b0 ;
  assign n40814 = ~n40812 & n40813 ;
  assign n40815 = n13573 ^ n12198 ^ n6979 ;
  assign n40816 = n5040 | n40815 ;
  assign n40817 = n40816 ^ n32193 ^ 1'b0 ;
  assign n40818 = ( n2199 & ~n3799 ) | ( n2199 & n13712 ) | ( ~n3799 & n13712 ) ;
  assign n40819 = n40817 & n40818 ;
  assign n40820 = n5027 | n40819 ;
  assign n40821 = n29960 ^ n11078 ^ 1'b0 ;
  assign n40822 = n40821 ^ n12656 ^ 1'b0 ;
  assign n40823 = n502 | n40822 ;
  assign n40824 = n9155 | n40823 ;
  assign n40825 = n32829 ^ n10131 ^ n1264 ;
  assign n40826 = ( ~n18040 & n40824 ) | ( ~n18040 & n40825 ) | ( n40824 & n40825 ) ;
  assign n40827 = n27002 ^ n20726 ^ n17425 ;
  assign n40828 = n40111 ^ n24753 ^ n8538 ;
  assign n40829 = ( ~n7634 & n40827 ) | ( ~n7634 & n40828 ) | ( n40827 & n40828 ) ;
  assign n40830 = n29879 ^ n25916 ^ n24032 ;
  assign n40831 = ( ~n34064 & n34793 ) | ( ~n34064 & n35000 ) | ( n34793 & n35000 ) ;
  assign n40832 = n10813 ^ n5353 ^ 1'b0 ;
  assign n40833 = n4244 | n40832 ;
  assign n40834 = n7452 | n40833 ;
  assign n40835 = ( n2716 & n17667 ) | ( n2716 & n40834 ) | ( n17667 & n40834 ) ;
  assign n40836 = n34538 ^ n6570 ^ 1'b0 ;
  assign n40837 = n29831 ^ n16993 ^ 1'b0 ;
  assign n40838 = n2272 | n24543 ;
  assign n40839 = n40837 | n40838 ;
  assign n40840 = n7601 | n13699 ;
  assign n40841 = ( ~n4155 & n8557 ) | ( ~n4155 & n9094 ) | ( n8557 & n9094 ) ;
  assign n40842 = n24147 & ~n40841 ;
  assign n40843 = n40819 & n40842 ;
  assign n40844 = n40843 ^ n34334 ^ n11164 ;
  assign n40845 = n40844 ^ n6237 ^ 1'b0 ;
  assign n40846 = n10636 | n40845 ;
  assign n40847 = n24938 & ~n40846 ;
  assign n40848 = n40847 ^ n36619 ^ 1'b0 ;
  assign n40849 = n3412 | n6187 ;
  assign n40850 = n40849 ^ n14288 ^ 1'b0 ;
  assign n40851 = n40850 ^ n1819 ^ 1'b0 ;
  assign n40852 = ( ~n2177 & n18892 ) | ( ~n2177 & n40851 ) | ( n18892 & n40851 ) ;
  assign n40853 = n26558 ^ n1000 ^ 1'b0 ;
  assign n40854 = ~n7732 & n40853 ;
  assign n40855 = n40854 ^ n14293 ^ n961 ;
  assign n40856 = n4309 | n31494 ;
  assign n40857 = n15802 | n40856 ;
  assign n40858 = n40857 ^ n12775 ^ n7116 ;
  assign n40859 = n30789 ^ n17665 ^ n3814 ;
  assign n40860 = n28160 | n37436 ;
  assign n40861 = x6 & n6871 ;
  assign n40862 = ~n40860 & n40861 ;
  assign n40863 = n40862 ^ n19491 ^ 1'b0 ;
  assign n40864 = n28705 | n36254 ;
  assign n40865 = n21173 ^ n11886 ^ 1'b0 ;
  assign n40866 = ( n3666 & ~n18576 ) | ( n3666 & n20641 ) | ( ~n18576 & n20641 ) ;
  assign n40867 = n6349 | n40866 ;
  assign n40868 = n5427 | n32326 ;
  assign n40869 = ( ~n822 & n7821 ) | ( ~n822 & n40868 ) | ( n7821 & n40868 ) ;
  assign n40870 = n35604 | n35615 ;
  assign n40871 = n40870 ^ n29733 ^ 1'b0 ;
  assign n40872 = ( n17110 & n23059 ) | ( n17110 & n40871 ) | ( n23059 & n40871 ) ;
  assign n40873 = n25131 | n26562 ;
  assign n40874 = n40873 ^ n9050 ^ 1'b0 ;
  assign n40875 = n40874 ^ n10931 ^ n2949 ;
  assign n40876 = n16285 | n31319 ;
  assign n40877 = n40876 ^ n2731 ^ 1'b0 ;
  assign n40878 = ( n9573 & n14844 ) | ( n9573 & n40877 ) | ( n14844 & n40877 ) ;
  assign n40879 = n4603 | n12881 ;
  assign n40880 = n9143 | n40879 ;
  assign n40881 = n40880 ^ n8394 ^ 1'b0 ;
  assign n40882 = n40881 ^ n293 ^ 1'b0 ;
  assign n40883 = n40566 & ~n40882 ;
  assign n40884 = n19730 ^ n11528 ^ 1'b0 ;
  assign n40885 = n40884 ^ n16587 ^ 1'b0 ;
  assign n40886 = n40885 ^ n34272 ^ n16589 ;
  assign n40892 = ~n4673 & n11800 ;
  assign n40893 = n40892 ^ n2337 ^ 1'b0 ;
  assign n40894 = n40893 ^ n17642 ^ 1'b0 ;
  assign n40887 = n5223 & ~n20334 ;
  assign n40888 = n40887 ^ n12831 ^ 1'b0 ;
  assign n40889 = ( n8336 & ~n8922 ) | ( n8336 & n10958 ) | ( ~n8922 & n10958 ) ;
  assign n40890 = n40888 | n40889 ;
  assign n40891 = ( ~n6810 & n28403 ) | ( ~n6810 & n40890 ) | ( n28403 & n40890 ) ;
  assign n40895 = n40894 ^ n40891 ^ n2608 ;
  assign n40896 = n40306 ^ n30478 ^ n7741 ;
  assign n40897 = ( n1482 & n2671 ) | ( n1482 & ~n5353 ) | ( n2671 & ~n5353 ) ;
  assign n40898 = n40897 ^ n34980 ^ n10679 ;
  assign n40899 = n20130 ^ n13092 ^ n7475 ;
  assign n40900 = ~n25594 & n40899 ;
  assign n40901 = n8904 ^ n1133 ^ 1'b0 ;
  assign n40902 = n4464 ^ n1329 ^ n441 ;
  assign n40903 = n40902 ^ n38124 ^ 1'b0 ;
  assign n40904 = n40903 ^ n1189 ^ 1'b0 ;
  assign n40905 = ~n40901 & n40904 ;
  assign n40906 = n11558 & n15959 ;
  assign n40907 = n40906 ^ n36317 ^ 1'b0 ;
  assign n40911 = ~n17140 & n19142 ;
  assign n40912 = n40911 ^ n9059 ^ 1'b0 ;
  assign n40910 = n22864 & n22959 ;
  assign n40908 = n9279 & n16639 ;
  assign n40909 = ( ~n10127 & n40347 ) | ( ~n10127 & n40908 ) | ( n40347 & n40908 ) ;
  assign n40913 = n40912 ^ n40910 ^ n40909 ;
  assign n40914 = n37889 ^ n30290 ^ 1'b0 ;
  assign n40915 = n8984 & ~n40914 ;
  assign n40916 = n11783 & ~n40915 ;
  assign n40917 = n9101 ^ n1705 ^ 1'b0 ;
  assign n40918 = ~n35783 & n40917 ;
  assign n40919 = ~n2671 & n40918 ;
  assign n40920 = n7506 & n40919 ;
  assign n40921 = n6372 | n24822 ;
  assign n40922 = n1786 & ~n40921 ;
  assign n40923 = n1482 & ~n10240 ;
  assign n40924 = n35379 ^ n13484 ^ 1'b0 ;
  assign n40925 = n40923 | n40924 ;
  assign n40926 = n1229 & n9500 ;
  assign n40927 = n30629 ^ n2020 ^ 1'b0 ;
  assign n40928 = n40927 ^ n15443 ^ n8064 ;
  assign n40929 = n7834 ^ n1846 ^ 1'b0 ;
  assign n40930 = n1957 | n10005 ;
  assign n40931 = n40930 ^ n12583 ^ 1'b0 ;
  assign n40932 = n8309 & ~n15338 ;
  assign n40933 = n40932 ^ n26227 ^ 1'b0 ;
  assign n40934 = n928 & ~n11922 ;
  assign n40935 = ~n22735 & n40934 ;
  assign n40936 = n1361 ^ n934 ^ 1'b0 ;
  assign n40937 = n30460 ^ n11756 ^ 1'b0 ;
  assign n40938 = n39310 ^ n34914 ^ n26671 ;
  assign n40939 = ( n16790 & n17973 ) | ( n16790 & ~n36254 ) | ( n17973 & ~n36254 ) ;
  assign n40940 = n952 | n40939 ;
  assign n40941 = n579 & ~n39866 ;
  assign n40942 = n8799 ^ n6004 ^ 1'b0 ;
  assign n40943 = n40942 ^ n11304 ^ 1'b0 ;
  assign n40944 = n40943 ^ n19250 ^ 1'b0 ;
  assign n40945 = n3491 & ~n40944 ;
  assign n40946 = n40945 ^ n10198 ^ n8262 ;
  assign n40947 = ( n3310 & n40941 ) | ( n3310 & ~n40946 ) | ( n40941 & ~n40946 ) ;
  assign n40948 = n13118 & ~n16230 ;
  assign n40949 = n450 & n40948 ;
  assign n40950 = ( ~n13539 & n20522 ) | ( ~n13539 & n31959 ) | ( n20522 & n31959 ) ;
  assign n40951 = ~n40949 & n40950 ;
  assign n40952 = n9869 & ~n9952 ;
  assign n40953 = n40952 ^ n26074 ^ 1'b0 ;
  assign n40954 = n40953 ^ n3123 ^ 1'b0 ;
  assign n40955 = n17193 ^ n10817 ^ 1'b0 ;
  assign n40956 = n10070 & ~n20442 ;
  assign n40957 = ~n19038 & n40956 ;
  assign n40958 = n11775 ^ n7597 ^ x221 ;
  assign n40959 = n13817 & ~n40958 ;
  assign n40960 = n40959 ^ n22234 ^ n9220 ;
  assign n40962 = n5715 ^ x147 ^ 1'b0 ;
  assign n40963 = n7234 & ~n40962 ;
  assign n40964 = n40963 ^ n306 ^ 1'b0 ;
  assign n40965 = n40964 ^ n30334 ^ n14235 ;
  assign n40961 = ~n19608 & n35418 ;
  assign n40966 = n40965 ^ n40961 ^ 1'b0 ;
  assign n40967 = n23570 ^ n8495 ^ 1'b0 ;
  assign n40968 = n25412 & n40967 ;
  assign n40969 = n21422 & n40968 ;
  assign n40970 = n40969 ^ n8033 ^ 1'b0 ;
  assign n40971 = ~n37678 & n40970 ;
  assign n40972 = ( n518 & ~n18087 ) | ( n518 & n22882 ) | ( ~n18087 & n22882 ) ;
  assign n40973 = ~n3846 & n14820 ;
  assign n40974 = ~n40972 & n40973 ;
  assign n40975 = n39083 ^ n31858 ^ n29385 ;
  assign n40976 = ( n14632 & n18592 ) | ( n14632 & n19121 ) | ( n18592 & n19121 ) ;
  assign n40979 = n26070 ^ n23437 ^ n10055 ;
  assign n40977 = n5927 & n18073 ;
  assign n40978 = ~n9235 & n40977 ;
  assign n40980 = n40979 ^ n40978 ^ n12494 ;
  assign n40981 = n40980 ^ n31053 ^ 1'b0 ;
  assign n40982 = n40981 ^ n40745 ^ n29220 ;
  assign n40983 = n23075 | n34440 ;
  assign n40984 = n40983 ^ n19295 ^ 1'b0 ;
  assign n40985 = n5027 & ~n15086 ;
  assign n40986 = n12143 & n40985 ;
  assign n40987 = n11172 ^ n1724 ^ 1'b0 ;
  assign n40988 = n40986 | n40987 ;
  assign n40989 = n1628 | n10765 ;
  assign n40990 = n37004 | n40989 ;
  assign n40991 = ~n4271 & n5495 ;
  assign n40994 = n36684 ^ n7335 ^ 1'b0 ;
  assign n40995 = n768 & n40994 ;
  assign n40992 = n6546 & n8023 ;
  assign n40993 = n40992 ^ n40230 ^ n36614 ;
  assign n40996 = n40995 ^ n40993 ^ n10254 ;
  assign n40997 = n23716 ^ n5863 ^ 1'b0 ;
  assign n40998 = ~n15443 & n40997 ;
  assign n40999 = n21078 | n21456 ;
  assign n41000 = n40999 ^ n34020 ^ 1'b0 ;
  assign n41001 = n33096 & ~n33765 ;
  assign n41002 = ( n20501 & n36614 ) | ( n20501 & n41001 ) | ( n36614 & n41001 ) ;
  assign n41003 = n32796 ^ n19158 ^ n10163 ;
  assign n41004 = ( n4390 & ~n4636 ) | ( n4390 & n28103 ) | ( ~n4636 & n28103 ) ;
  assign n41005 = ( n2986 & n12642 ) | ( n2986 & ~n41004 ) | ( n12642 & ~n41004 ) ;
  assign n41006 = ( ~n5719 & n8349 ) | ( ~n5719 & n31935 ) | ( n8349 & n31935 ) ;
  assign n41007 = n7175 | n41006 ;
  assign n41008 = n18308 & ~n31046 ;
  assign n41009 = n15237 & n41008 ;
  assign n41010 = n4714 & ~n39473 ;
  assign n41011 = n41010 ^ n512 ^ 1'b0 ;
  assign n41012 = n33095 | n41011 ;
  assign n41013 = n37633 ^ n17695 ^ 1'b0 ;
  assign n41014 = n19952 & ~n37038 ;
  assign n41015 = n39613 ^ n32565 ^ n24862 ;
  assign n41016 = n29360 ^ n17141 ^ n13263 ;
  assign n41017 = n22815 ^ n10778 ^ n1603 ;
  assign n41018 = n27618 | n41017 ;
  assign n41019 = n40524 ^ n11363 ^ n4198 ;
  assign n41020 = ~n6097 & n41019 ;
  assign n41021 = ~n17740 & n41020 ;
  assign n41022 = n11883 | n17115 ;
  assign n41023 = n41022 ^ n4173 ^ 1'b0 ;
  assign n41024 = n16064 | n41023 ;
  assign n41025 = n41024 ^ n10187 ^ 1'b0 ;
  assign n41026 = n41025 ^ n37425 ^ n10998 ;
  assign n41027 = n3811 & n19347 ;
  assign n41028 = ( n5153 & n19254 ) | ( n5153 & ~n22121 ) | ( n19254 & ~n22121 ) ;
  assign n41029 = n35642 ^ n7796 ^ 1'b0 ;
  assign n41030 = n41029 ^ n37579 ^ n16795 ;
  assign n41031 = ( n5454 & n20010 ) | ( n5454 & n20991 ) | ( n20010 & n20991 ) ;
  assign n41032 = n5759 & n23526 ;
  assign n41033 = n11200 | n41032 ;
  assign n41034 = n41033 ^ n6257 ^ 1'b0 ;
  assign n41035 = ~n20928 & n29912 ;
  assign n41036 = n41035 ^ n4087 ^ 1'b0 ;
  assign n41037 = ( ~n7255 & n38127 ) | ( ~n7255 & n41036 ) | ( n38127 & n41036 ) ;
  assign n41038 = n20076 ^ n2784 ^ 1'b0 ;
  assign n41039 = n9911 & n41038 ;
  assign n41040 = ~n41037 & n41039 ;
  assign n41041 = n27495 ^ n18571 ^ 1'b0 ;
  assign n41042 = n31817 & ~n41041 ;
  assign n41043 = n5086 | n29151 ;
  assign n41044 = n33427 & ~n41043 ;
  assign n41045 = ( n12373 & n13141 ) | ( n12373 & n31161 ) | ( n13141 & n31161 ) ;
  assign n41046 = ~n29266 & n41045 ;
  assign n41050 = n21252 ^ n13423 ^ 1'b0 ;
  assign n41047 = ( ~n9645 & n11894 ) | ( ~n9645 & n12460 ) | ( n11894 & n12460 ) ;
  assign n41048 = ( n1759 & n17627 ) | ( n1759 & ~n40549 ) | ( n17627 & ~n40549 ) ;
  assign n41049 = n41047 | n41048 ;
  assign n41051 = n41050 ^ n41049 ^ n31710 ;
  assign n41052 = n39960 ^ n16496 ^ n9182 ;
  assign n41053 = n13640 ^ n5782 ^ 1'b0 ;
  assign n41054 = n41053 ^ n11231 ^ 1'b0 ;
  assign n41056 = n16784 ^ n13242 ^ 1'b0 ;
  assign n41057 = n39414 | n41056 ;
  assign n41055 = ~n9045 & n17156 ;
  assign n41058 = n41057 ^ n41055 ^ 1'b0 ;
  assign n41059 = n15468 | n24359 ;
  assign n41060 = n10495 & n22938 ;
  assign n41061 = ~n3010 & n41060 ;
  assign n41062 = n41061 ^ n6259 ^ 1'b0 ;
  assign n41063 = n11099 ^ n1515 ^ n1447 ;
  assign n41064 = ( n5965 & n23772 ) | ( n5965 & ~n41063 ) | ( n23772 & ~n41063 ) ;
  assign n41065 = n20453 & ~n41064 ;
  assign n41066 = n41062 & n41065 ;
  assign n41067 = n31255 ^ n6862 ^ 1'b0 ;
  assign n41068 = ( n8980 & n26517 ) | ( n8980 & n41067 ) | ( n26517 & n41067 ) ;
  assign n41069 = n12487 | n26443 ;
  assign n41070 = ( n425 & ~n3419 ) | ( n425 & n12350 ) | ( ~n3419 & n12350 ) ;
  assign n41071 = n17851 ^ n14807 ^ n5302 ;
  assign n41072 = n14149 & ~n41071 ;
  assign n41073 = n28719 ^ n6234 ^ 1'b0 ;
  assign n41074 = n39934 & n41073 ;
  assign n41075 = n41074 ^ n2205 ^ 1'b0 ;
  assign n41076 = ( n530 & ~n7960 ) | ( n530 & n9482 ) | ( ~n7960 & n9482 ) ;
  assign n41077 = n41076 ^ n664 ^ 1'b0 ;
  assign n41078 = ( n3210 & n24127 ) | ( n3210 & ~n41077 ) | ( n24127 & ~n41077 ) ;
  assign n41079 = n18882 ^ n6432 ^ 1'b0 ;
  assign n41080 = ( ~n9851 & n35581 ) | ( ~n9851 & n41079 ) | ( n35581 & n41079 ) ;
  assign n41081 = n13612 ^ n13161 ^ 1'b0 ;
  assign n41082 = n41081 ^ x181 ^ 1'b0 ;
  assign n41083 = n1648 | n41082 ;
  assign n41084 = n28057 ^ n27599 ^ n6570 ;
  assign n41085 = n33176 ^ n1354 ^ 1'b0 ;
  assign n41086 = n18281 & n41085 ;
  assign n41087 = n20690 ^ n8274 ^ 1'b0 ;
  assign n41088 = n31449 & n41087 ;
  assign n41089 = n753 & n3401 ;
  assign n41090 = ~n3184 & n41089 ;
  assign n41091 = n41090 ^ n9174 ^ 1'b0 ;
  assign n41092 = ~n8480 & n22933 ;
  assign n41093 = n41091 & n41092 ;
  assign n41094 = ~n41088 & n41093 ;
  assign n41095 = ( ~n3314 & n12332 ) | ( ~n3314 & n13351 ) | ( n12332 & n13351 ) ;
  assign n41096 = n41095 ^ n6850 ^ 1'b0 ;
  assign n41097 = n18605 & n41096 ;
  assign n41098 = n12841 ^ n6573 ^ 1'b0 ;
  assign n41099 = n14677 & ~n41098 ;
  assign n41100 = ( ~n1291 & n8824 ) | ( ~n1291 & n41099 ) | ( n8824 & n41099 ) ;
  assign n41103 = ~n2998 & n8231 ;
  assign n41101 = ~n4584 & n26608 ;
  assign n41102 = ~n21574 & n41101 ;
  assign n41104 = n41103 ^ n41102 ^ n29180 ;
  assign n41105 = n24407 ^ n11772 ^ n8907 ;
  assign n41106 = n2832 & n22986 ;
  assign n41107 = n41106 ^ n8695 ^ 1'b0 ;
  assign n41108 = n41107 ^ n24544 ^ n20092 ;
  assign n41109 = n6735 & n36303 ;
  assign n41110 = n41109 ^ n38027 ^ n6892 ;
  assign n41111 = ~n36606 & n36772 ;
  assign n41112 = n41111 ^ n14885 ^ 1'b0 ;
  assign n41114 = n25792 ^ n2298 ^ 1'b0 ;
  assign n41115 = n2002 | n3838 ;
  assign n41116 = n41114 | n41115 ;
  assign n41113 = ( n13209 & n26455 ) | ( n13209 & ~n30989 ) | ( n26455 & ~n30989 ) ;
  assign n41117 = n41116 ^ n41113 ^ 1'b0 ;
  assign n41118 = n7746 | n8201 ;
  assign n41119 = n41118 ^ n13543 ^ 1'b0 ;
  assign n41120 = ~n4414 & n41119 ;
  assign n41121 = ( n25772 & n28040 ) | ( n25772 & n41120 ) | ( n28040 & n41120 ) ;
  assign n41122 = n15400 ^ n11649 ^ 1'b0 ;
  assign n41123 = ( n20840 & ~n41121 ) | ( n20840 & n41122 ) | ( ~n41121 & n41122 ) ;
  assign n41124 = n16274 ^ n5666 ^ 1'b0 ;
  assign n41125 = n41124 ^ n40580 ^ n33030 ;
  assign n41126 = n23250 | n38146 ;
  assign n41127 = n17757 & ~n22157 ;
  assign n41128 = n41127 ^ n30526 ^ 1'b0 ;
  assign n41129 = n34991 ^ n29450 ^ 1'b0 ;
  assign n41130 = n33208 | n41129 ;
  assign n41131 = n6418 | n41130 ;
  assign n41132 = n41131 ^ n2096 ^ 1'b0 ;
  assign n41133 = n3725 | n41132 ;
  assign n41134 = n41133 ^ n13612 ^ 1'b0 ;
  assign n41135 = n6468 & ~n8267 ;
  assign n41136 = n16219 ^ n12802 ^ 1'b0 ;
  assign n41137 = n32856 | n41136 ;
  assign n41138 = n27498 ^ n9727 ^ 1'b0 ;
  assign n41139 = n41138 ^ n900 ^ 1'b0 ;
  assign n41143 = n30803 ^ n16766 ^ 1'b0 ;
  assign n41144 = n5374 & n41143 ;
  assign n41140 = n22373 ^ n13667 ^ 1'b0 ;
  assign n41141 = n22856 & n41140 ;
  assign n41142 = ( n2655 & n22081 ) | ( n2655 & n41141 ) | ( n22081 & n41141 ) ;
  assign n41145 = n41144 ^ n41142 ^ n36434 ;
  assign n41146 = n26269 ^ n11935 ^ 1'b0 ;
  assign n41147 = ~n33472 & n41146 ;
  assign n41148 = ~n5077 & n6037 ;
  assign n41149 = ( n8428 & n41147 ) | ( n8428 & n41148 ) | ( n41147 & n41148 ) ;
  assign n41151 = x183 & ~n38271 ;
  assign n41152 = n41151 ^ n3813 ^ 1'b0 ;
  assign n41150 = n11436 ^ n2828 ^ 1'b0 ;
  assign n41153 = n41152 ^ n41150 ^ n24836 ;
  assign n41154 = n897 & n41153 ;
  assign n41157 = n13661 & n14571 ;
  assign n41158 = n41157 ^ n3638 ^ 1'b0 ;
  assign n41159 = n23074 | n41158 ;
  assign n41160 = n7976 | n41159 ;
  assign n41161 = n12705 ^ n8027 ^ 1'b0 ;
  assign n41162 = ( n6362 & n41160 ) | ( n6362 & ~n41161 ) | ( n41160 & ~n41161 ) ;
  assign n41155 = n8200 & n10474 ;
  assign n41156 = n32281 & n41155 ;
  assign n41163 = n41162 ^ n41156 ^ n14227 ;
  assign n41164 = n20706 ^ n1458 ^ 1'b0 ;
  assign n41165 = n7374 | n22198 ;
  assign n41166 = n41165 ^ n39290 ^ 1'b0 ;
  assign n41167 = n9681 ^ n9602 ^ n4230 ;
  assign n41173 = n16553 ^ n16334 ^ n8924 ;
  assign n41174 = n41173 ^ n5509 ^ 1'b0 ;
  assign n41168 = n16847 ^ n2962 ^ 1'b0 ;
  assign n41169 = n25042 & n41168 ;
  assign n41170 = n41169 ^ n16561 ^ 1'b0 ;
  assign n41171 = n41170 ^ n24149 ^ 1'b0 ;
  assign n41172 = ~n14325 & n41171 ;
  assign n41175 = n41174 ^ n41172 ^ n29842 ;
  assign n41176 = n20535 ^ n6314 ^ 1'b0 ;
  assign n41177 = ( ~n4925 & n6807 ) | ( ~n4925 & n39731 ) | ( n6807 & n39731 ) ;
  assign n41182 = ( n14151 & ~n24349 ) | ( n14151 & n29198 ) | ( ~n24349 & n29198 ) ;
  assign n41178 = n20126 & n21768 ;
  assign n41179 = n1331 & ~n41178 ;
  assign n41180 = n7189 & n41179 ;
  assign n41181 = ( ~n16240 & n16645 ) | ( ~n16240 & n41180 ) | ( n16645 & n41180 ) ;
  assign n41183 = n41182 ^ n41181 ^ 1'b0 ;
  assign n41184 = n10761 & ~n41183 ;
  assign n41185 = n22740 | n27757 ;
  assign n41186 = n41185 ^ n23386 ^ 1'b0 ;
  assign n41187 = ~n1040 & n8299 ;
  assign n41188 = ~n6329 & n41187 ;
  assign n41189 = n38213 ^ n33602 ^ 1'b0 ;
  assign n41190 = n41188 | n41189 ;
  assign n41192 = ( n10463 & n17654 ) | ( n10463 & ~n21136 ) | ( n17654 & ~n21136 ) ;
  assign n41193 = n41192 ^ n3254 ^ 1'b0 ;
  assign n41194 = n9153 | n41193 ;
  assign n41191 = n2819 | n11308 ;
  assign n41195 = n41194 ^ n41191 ^ 1'b0 ;
  assign n41196 = n15033 & ~n38635 ;
  assign n41197 = ( n16929 & n20056 ) | ( n16929 & ~n24663 ) | ( n20056 & ~n24663 ) ;
  assign n41198 = n10990 ^ n2405 ^ 1'b0 ;
  assign n41199 = ~n5949 & n41198 ;
  assign n41200 = ( n7370 & ~n41197 ) | ( n7370 & n41199 ) | ( ~n41197 & n41199 ) ;
  assign n41201 = n18631 ^ n3405 ^ n800 ;
  assign n41202 = ( n7173 & n27231 ) | ( n7173 & ~n41201 ) | ( n27231 & ~n41201 ) ;
  assign n41203 = n36866 ^ n33636 ^ n20143 ;
  assign n41204 = n5391 & n8254 ;
  assign n41205 = n41204 ^ n2661 ^ 1'b0 ;
  assign n41206 = n38485 & ~n41205 ;
  assign n41207 = n41206 ^ n36952 ^ 1'b0 ;
  assign n41208 = ( ~n37375 & n41203 ) | ( ~n37375 & n41207 ) | ( n41203 & n41207 ) ;
  assign n41209 = ( ~n25171 & n25370 ) | ( ~n25171 & n41208 ) | ( n25370 & n41208 ) ;
  assign n41210 = ( n8710 & ~n13612 ) | ( n8710 & n25303 ) | ( ~n13612 & n25303 ) ;
  assign n41211 = n41210 ^ n8409 ^ 1'b0 ;
  assign n41212 = n30496 & n41211 ;
  assign n41213 = n41212 ^ n821 ^ 1'b0 ;
  assign n41214 = n22863 ^ n3877 ^ 1'b0 ;
  assign n41215 = n9011 | n41214 ;
  assign n41216 = n18244 & ~n41215 ;
  assign n41217 = n41216 ^ n18631 ^ 1'b0 ;
  assign n41218 = n30483 ^ n24014 ^ n13335 ;
  assign n41219 = ( n10665 & ~n31033 ) | ( n10665 & n35832 ) | ( ~n31033 & n35832 ) ;
  assign n41220 = n16775 & n41219 ;
  assign n41221 = ~n41218 & n41220 ;
  assign n41222 = n6837 | n41221 ;
  assign n41223 = n32409 & ~n41222 ;
  assign n41224 = n27302 ^ n4592 ^ 1'b0 ;
  assign n41225 = ~n2598 & n11362 ;
  assign n41226 = n41225 ^ n31069 ^ n17213 ;
  assign n41227 = ( n29699 & n33530 ) | ( n29699 & n41226 ) | ( n33530 & n41226 ) ;
  assign n41228 = n32896 ^ n13204 ^ n12902 ;
  assign n41229 = n41228 ^ n28386 ^ n8748 ;
  assign n41234 = ( ~n2091 & n10388 ) | ( ~n2091 & n32371 ) | ( n10388 & n32371 ) ;
  assign n41233 = n5618 | n12962 ;
  assign n41235 = n41234 ^ n41233 ^ 1'b0 ;
  assign n41236 = n20761 & n41235 ;
  assign n41237 = n6124 & n41236 ;
  assign n41230 = n6373 ^ n528 ^ 1'b0 ;
  assign n41231 = n7789 & n41230 ;
  assign n41232 = n41231 ^ n28294 ^ 1'b0 ;
  assign n41238 = n41237 ^ n41232 ^ n20904 ;
  assign n41239 = n41238 ^ n39434 ^ n38643 ;
  assign n41240 = n25536 ^ n7078 ^ 1'b0 ;
  assign n41241 = ( n2811 & ~n7518 ) | ( n2811 & n11659 ) | ( ~n7518 & n11659 ) ;
  assign n41242 = ( n29829 & n41240 ) | ( n29829 & n41241 ) | ( n41240 & n41241 ) ;
  assign n41245 = ~n6665 & n31669 ;
  assign n41246 = n19423 ^ n15623 ^ n14602 ;
  assign n41247 = ~n41245 & n41246 ;
  assign n41248 = ~n15482 & n41247 ;
  assign n41243 = n12590 & n38655 ;
  assign n41244 = n30963 | n41243 ;
  assign n41249 = n41248 ^ n41244 ^ 1'b0 ;
  assign n41250 = ( n6195 & ~n32217 ) | ( n6195 & n38176 ) | ( ~n32217 & n38176 ) ;
  assign n41251 = n10645 & ~n41250 ;
  assign n41252 = n41251 ^ n37920 ^ 1'b0 ;
  assign n41253 = n6452 & ~n41252 ;
  assign n41254 = n41253 ^ n34589 ^ 1'b0 ;
  assign n41255 = n35698 ^ n27206 ^ n893 ;
  assign n41256 = ~n27628 & n41255 ;
  assign n41257 = ~n787 & n41256 ;
  assign n41258 = n7761 ^ n5460 ^ n1228 ;
  assign n41259 = n41258 ^ n6086 ^ n5738 ;
  assign n41260 = ( ~x249 & n3948 ) | ( ~x249 & n40586 ) | ( n3948 & n40586 ) ;
  assign n41261 = n20829 | n21416 ;
  assign n41262 = n41261 ^ n16145 ^ 1'b0 ;
  assign n41263 = ( ~n4044 & n7155 ) | ( ~n4044 & n36457 ) | ( n7155 & n36457 ) ;
  assign n41264 = n21915 & ~n33554 ;
  assign n41265 = n40818 ^ n17479 ^ n9089 ;
  assign n41266 = ~n41264 & n41265 ;
  assign n41267 = n20269 ^ n19646 ^ n5620 ;
  assign n41268 = n11253 ^ n6045 ^ n3666 ;
  assign n41269 = n22536 & n30629 ;
  assign n41270 = n41269 ^ n4217 ^ 1'b0 ;
  assign n41271 = n41268 & ~n41270 ;
  assign n41272 = n41271 ^ n3977 ^ 1'b0 ;
  assign n41273 = ~n41267 & n41272 ;
  assign n41274 = n1647 ^ n751 ^ 1'b0 ;
  assign n41275 = n286 | n26037 ;
  assign n41276 = ( n3028 & n14854 ) | ( n3028 & ~n16830 ) | ( n14854 & ~n16830 ) ;
  assign n41277 = n32144 & ~n41276 ;
  assign n41278 = n18689 & ~n36341 ;
  assign n41279 = n16306 & ~n41278 ;
  assign n41280 = ( n28801 & n41277 ) | ( n28801 & n41279 ) | ( n41277 & n41279 ) ;
  assign n41281 = ( n12796 & n26975 ) | ( n12796 & ~n41280 ) | ( n26975 & ~n41280 ) ;
  assign n41282 = ( n834 & n4848 ) | ( n834 & ~n33547 ) | ( n4848 & ~n33547 ) ;
  assign n41283 = n17594 | n41282 ;
  assign n41285 = n14609 ^ n9732 ^ n796 ;
  assign n41284 = n33643 ^ n25964 ^ n19642 ;
  assign n41286 = n41285 ^ n41284 ^ n10828 ;
  assign n41287 = n37592 ^ n19149 ^ n2615 ;
  assign n41288 = n5176 & ~n9443 ;
  assign n41289 = n18909 ^ n15020 ^ 1'b0 ;
  assign n41290 = n40338 & ~n41289 ;
  assign n41291 = n10785 | n37075 ;
  assign n41292 = n36200 & ~n41291 ;
  assign n41293 = n35189 ^ n30480 ^ n12564 ;
  assign n41294 = n37815 ^ n25867 ^ n19398 ;
  assign n41295 = n41294 ^ n30046 ^ 1'b0 ;
  assign n41296 = n7402 ^ n1722 ^ 1'b0 ;
  assign n41297 = ~n6336 & n41296 ;
  assign n41298 = n41297 ^ n8489 ^ 1'b0 ;
  assign n41299 = ( n41293 & ~n41295 ) | ( n41293 & n41298 ) | ( ~n41295 & n41298 ) ;
  assign n41300 = ~n6824 & n39075 ;
  assign n41301 = n10802 & ~n13811 ;
  assign n41302 = n41301 ^ n24003 ^ 1'b0 ;
  assign n41303 = ( n13720 & n41300 ) | ( n13720 & n41302 ) | ( n41300 & n41302 ) ;
  assign n41304 = n21483 & n34982 ;
  assign n41305 = n14161 & ~n41304 ;
  assign n41306 = n13460 & n41305 ;
  assign n41307 = n31346 ^ n3637 ^ 1'b0 ;
  assign n41308 = n36107 & ~n41307 ;
  assign n41309 = n11965 ^ n8562 ^ 1'b0 ;
  assign n41310 = n18909 & n21631 ;
  assign n41311 = n17051 & n41310 ;
  assign n41312 = ( n674 & ~n14206 ) | ( n674 & n31571 ) | ( ~n14206 & n31571 ) ;
  assign n41313 = ~n2953 & n10198 ;
  assign n41314 = ( n23249 & n31690 ) | ( n23249 & n33506 ) | ( n31690 & n33506 ) ;
  assign n41315 = n11119 & n41314 ;
  assign n41316 = n41315 ^ n34885 ^ 1'b0 ;
  assign n41317 = n9008 & n41316 ;
  assign n41318 = n39580 ^ n22113 ^ n15157 ;
  assign n41329 = n5441 | n19175 ;
  assign n41330 = n14493 | n41329 ;
  assign n41331 = n21053 & n22768 ;
  assign n41332 = ( ~n31491 & n41330 ) | ( ~n31491 & n41331 ) | ( n41330 & n41331 ) ;
  assign n41319 = n15226 & ~n36293 ;
  assign n41320 = n41319 ^ x64 ^ 1'b0 ;
  assign n41321 = n8907 & n24640 ;
  assign n41322 = n41321 ^ n697 ^ 1'b0 ;
  assign n41323 = ( n16160 & n41320 ) | ( n16160 & ~n41322 ) | ( n41320 & ~n41322 ) ;
  assign n41324 = n7605 ^ n7482 ^ n4906 ;
  assign n41325 = ( ~n332 & n11836 ) | ( ~n332 & n41324 ) | ( n11836 & n41324 ) ;
  assign n41326 = ( ~n1981 & n22917 ) | ( ~n1981 & n41325 ) | ( n22917 & n41325 ) ;
  assign n41327 = n36631 ^ n28516 ^ n25136 ;
  assign n41328 = ( ~n41323 & n41326 ) | ( ~n41323 & n41327 ) | ( n41326 & n41327 ) ;
  assign n41333 = n41332 ^ n41328 ^ n27088 ;
  assign n41334 = n1635 | n36381 ;
  assign n41335 = n9176 | n41334 ;
  assign n41336 = n31688 & n41335 ;
  assign n41337 = ~n23528 & n41336 ;
  assign n41338 = ~n9351 & n30913 ;
  assign n41339 = n41257 ^ n25158 ^ 1'b0 ;
  assign n41340 = n12674 | n41339 ;
  assign n41341 = n28021 | n32405 ;
  assign n41342 = n41341 ^ n27502 ^ 1'b0 ;
  assign n41343 = ( n4508 & ~n16573 ) | ( n4508 & n41342 ) | ( ~n16573 & n41342 ) ;
  assign n41344 = n41343 ^ n19811 ^ 1'b0 ;
  assign n41345 = n6219 ^ n4011 ^ 1'b0 ;
  assign n41346 = n1206 | n30234 ;
  assign n41351 = ( ~n2567 & n3843 ) | ( ~n2567 & n13165 ) | ( n3843 & n13165 ) ;
  assign n41350 = ~n4175 & n19952 ;
  assign n41352 = n41351 ^ n41350 ^ n29763 ;
  assign n41347 = ~n1143 & n27185 ;
  assign n41348 = n41347 ^ n6781 ^ 1'b0 ;
  assign n41349 = n33514 & ~n41348 ;
  assign n41353 = n41352 ^ n41349 ^ n25818 ;
  assign n41354 = ( n11324 & ~n13972 ) | ( n11324 & n39151 ) | ( ~n13972 & n39151 ) ;
  assign n41355 = n1124 | n13287 ;
  assign n41356 = n9368 ^ n5101 ^ 1'b0 ;
  assign n41357 = n41356 ^ n30781 ^ 1'b0 ;
  assign n41358 = n41357 ^ n585 ^ 1'b0 ;
  assign n41359 = n6354 & n15357 ;
  assign n41360 = n41359 ^ n9434 ^ 1'b0 ;
  assign n41361 = n41360 ^ n27702 ^ 1'b0 ;
  assign n41362 = n2347 & ~n4327 ;
  assign n41363 = n41362 ^ n13831 ^ 1'b0 ;
  assign n41364 = n41363 ^ n18083 ^ 1'b0 ;
  assign n41365 = n41364 ^ n9883 ^ n4873 ;
  assign n41366 = ~n10218 & n41365 ;
  assign n41367 = n26447 ^ n22641 ^ 1'b0 ;
  assign n41368 = n39289 | n41367 ;
  assign n41369 = n41366 & ~n41368 ;
  assign n41370 = n16500 & ~n32059 ;
  assign n41371 = n41370 ^ n27029 ^ 1'b0 ;
  assign n41372 = n19114 & ~n32892 ;
  assign n41373 = ( n10699 & ~n34768 ) | ( n10699 & n36551 ) | ( ~n34768 & n36551 ) ;
  assign n41374 = n29653 ^ n8260 ^ n5883 ;
  assign n41375 = n41374 ^ n8867 ^ n1002 ;
  assign n41376 = n16400 ^ n1916 ^ 1'b0 ;
  assign n41377 = n41375 | n41376 ;
  assign n41378 = n15338 & ~n17346 ;
  assign n41379 = n41378 ^ n41206 ^ 1'b0 ;
  assign n41380 = ( n27968 & n41377 ) | ( n27968 & ~n41379 ) | ( n41377 & ~n41379 ) ;
  assign n41381 = n41380 ^ n17405 ^ 1'b0 ;
  assign n41382 = n15568 ^ n9876 ^ 1'b0 ;
  assign n41383 = n35647 & n41382 ;
  assign n41384 = n14049 ^ n3462 ^ 1'b0 ;
  assign n41385 = n2691 & ~n41384 ;
  assign n41386 = n15449 ^ n7757 ^ 1'b0 ;
  assign n41387 = ~n41385 & n41386 ;
  assign n41388 = n20832 ^ n19352 ^ 1'b0 ;
  assign n41389 = n22453 & ~n41388 ;
  assign n41390 = n17798 ^ n17776 ^ 1'b0 ;
  assign n41391 = n41389 & n41390 ;
  assign n41392 = n9788 & ~n20203 ;
  assign n41393 = n41392 ^ n4674 ^ 1'b0 ;
  assign n41394 = ~n3632 & n20758 ;
  assign n41395 = n41394 ^ n12303 ^ 1'b0 ;
  assign n41396 = ~n10824 & n40705 ;
  assign n41397 = n41396 ^ n33128 ^ 1'b0 ;
  assign n41398 = n41397 ^ n31629 ^ n384 ;
  assign n41399 = n8882 ^ n8038 ^ n6220 ;
  assign n41400 = ( n12048 & ~n41019 ) | ( n12048 & n41399 ) | ( ~n41019 & n41399 ) ;
  assign n41401 = n23990 ^ n10216 ^ n5020 ;
  assign n41402 = ( n23644 & n27210 ) | ( n23644 & ~n41401 ) | ( n27210 & ~n41401 ) ;
  assign n41407 = ( n4014 & n4632 ) | ( n4014 & ~n9810 ) | ( n4632 & ~n9810 ) ;
  assign n41408 = ( n22326 & ~n22437 ) | ( n22326 & n41407 ) | ( ~n22437 & n41407 ) ;
  assign n41403 = ( n7729 & ~n7747 ) | ( n7729 & n10235 ) | ( ~n7747 & n10235 ) ;
  assign n41404 = n14340 & ~n41403 ;
  assign n41405 = n13000 & ~n41404 ;
  assign n41406 = n41405 ^ n29354 ^ 1'b0 ;
  assign n41409 = n41408 ^ n41406 ^ n17879 ;
  assign n41410 = n37838 ^ n19802 ^ n9331 ;
  assign n41411 = n8327 ^ n5281 ^ 1'b0 ;
  assign n41412 = ~n13900 & n41411 ;
  assign n41413 = n3011 & ~n41412 ;
  assign n41414 = n41413 ^ n2077 ^ 1'b0 ;
  assign n41415 = ~n14189 & n41414 ;
  assign n41418 = n39050 ^ n18776 ^ 1'b0 ;
  assign n41416 = n13277 ^ n7790 ^ n6827 ;
  assign n41417 = ( n13309 & n40569 ) | ( n13309 & n41416 ) | ( n40569 & n41416 ) ;
  assign n41419 = n41418 ^ n41417 ^ n7122 ;
  assign n41420 = n25939 ^ n9466 ^ 1'b0 ;
  assign n41421 = ~n22610 & n41420 ;
  assign n41422 = n4971 & ~n7025 ;
  assign n41423 = ~n41421 & n41422 ;
  assign n41424 = ( n701 & ~n12431 ) | ( n701 & n41423 ) | ( ~n12431 & n41423 ) ;
  assign n41425 = ( n1460 & ~n8064 ) | ( n1460 & n41424 ) | ( ~n8064 & n41424 ) ;
  assign n41426 = ( ~n8049 & n18914 ) | ( ~n8049 & n32409 ) | ( n18914 & n32409 ) ;
  assign n41427 = ( ~n27022 & n29007 ) | ( ~n27022 & n41426 ) | ( n29007 & n41426 ) ;
  assign n41428 = ( n15794 & ~n17532 ) | ( n15794 & n26011 ) | ( ~n17532 & n26011 ) ;
  assign n41429 = n41428 ^ n8000 ^ 1'b0 ;
  assign n41433 = ~n686 & n4769 ;
  assign n41434 = n30951 ^ n3173 ^ 1'b0 ;
  assign n41435 = n41433 & n41434 ;
  assign n41430 = n30814 ^ n21788 ^ n14950 ;
  assign n41431 = n40432 & n41430 ;
  assign n41432 = n36682 & ~n41431 ;
  assign n41436 = n41435 ^ n41432 ^ 1'b0 ;
  assign n41437 = ~n7469 & n16042 ;
  assign n41438 = n32774 ^ n8092 ^ 1'b0 ;
  assign n41439 = n3585 & ~n11006 ;
  assign n41440 = n25192 ^ n5885 ^ 1'b0 ;
  assign n41441 = ( ~n7917 & n19258 ) | ( ~n7917 & n41440 ) | ( n19258 & n41440 ) ;
  assign n41442 = n16803 ^ n15585 ^ n4501 ;
  assign n41443 = n7658 | n41442 ;
  assign n41444 = n41443 ^ n1047 ^ 1'b0 ;
  assign n41445 = n41444 ^ n6360 ^ 1'b0 ;
  assign n41446 = ~n19458 & n41445 ;
  assign n41447 = ~n10261 & n14339 ;
  assign n41448 = ( ~n12912 & n35259 ) | ( ~n12912 & n41447 ) | ( n35259 & n41447 ) ;
  assign n41450 = ( n4586 & n6423 ) | ( n4586 & ~n17249 ) | ( n6423 & ~n17249 ) ;
  assign n41449 = n2537 & ~n13890 ;
  assign n41451 = n41450 ^ n41449 ^ 1'b0 ;
  assign n41452 = n11771 | n41451 ;
  assign n41453 = n36342 & ~n41452 ;
  assign n41454 = ( n13207 & n19854 ) | ( n13207 & n41453 ) | ( n19854 & n41453 ) ;
  assign n41455 = n11567 ^ n8721 ^ 1'b0 ;
  assign n41456 = n41455 ^ n18036 ^ 1'b0 ;
  assign n41457 = n41231 ^ n2438 ^ x232 ;
  assign n41458 = n3139 & ~n30180 ;
  assign n41459 = n41457 & n41458 ;
  assign n41461 = n26979 ^ n23043 ^ n3504 ;
  assign n41460 = n10786 | n32512 ;
  assign n41462 = n41461 ^ n41460 ^ 1'b0 ;
  assign n41463 = n9016 & ~n18732 ;
  assign n41464 = ( n1524 & n16594 ) | ( n1524 & ~n39961 ) | ( n16594 & ~n39961 ) ;
  assign n41465 = ( n4972 & n5267 ) | ( n4972 & ~n35780 ) | ( n5267 & ~n35780 ) ;
  assign n41466 = ( n16664 & ~n34438 ) | ( n16664 & n40747 ) | ( ~n34438 & n40747 ) ;
  assign n41467 = n21157 ^ n12841 ^ n10953 ;
  assign n41468 = ( ~x13 & n22182 ) | ( ~x13 & n31369 ) | ( n22182 & n31369 ) ;
  assign n41469 = ~n842 & n41468 ;
  assign n41470 = ( n1138 & n5581 ) | ( n1138 & n41469 ) | ( n5581 & n41469 ) ;
  assign n41471 = n8501 & ~n41470 ;
  assign n41472 = ~n8260 & n41471 ;
  assign n41473 = n35088 | n41178 ;
  assign n41474 = ( n481 & n7737 ) | ( n481 & n17132 ) | ( n7737 & n17132 ) ;
  assign n41475 = n5690 & ~n41474 ;
  assign n41476 = ~n41473 & n41475 ;
  assign n41477 = ( n9021 & n11402 ) | ( n9021 & ~n22674 ) | ( n11402 & ~n22674 ) ;
  assign n41478 = n27312 ^ n18825 ^ 1'b0 ;
  assign n41479 = ~n41477 & n41478 ;
  assign n41480 = n2106 ^ n1739 ^ 1'b0 ;
  assign n41481 = n41480 ^ n37840 ^ 1'b0 ;
  assign n41485 = n16929 | n28318 ;
  assign n41482 = n10823 ^ n5657 ^ 1'b0 ;
  assign n41483 = n41482 ^ n27192 ^ 1'b0 ;
  assign n41484 = n29389 & n41483 ;
  assign n41486 = n41485 ^ n41484 ^ n4604 ;
  assign n41487 = n14156 ^ n3762 ^ n577 ;
  assign n41488 = n22417 ^ n8871 ^ 1'b0 ;
  assign n41489 = n3300 & ~n41488 ;
  assign n41490 = ( ~n26493 & n38036 ) | ( ~n26493 & n41489 ) | ( n38036 & n41489 ) ;
  assign n41491 = ( n3401 & n4227 ) | ( n3401 & ~n9597 ) | ( n4227 & ~n9597 ) ;
  assign n41492 = n5416 & n41491 ;
  assign n41493 = ~n3116 & n41492 ;
  assign n41494 = n5163 | n30669 ;
  assign n41495 = n17122 ^ n12234 ^ n9234 ;
  assign n41496 = ( n7201 & ~n16099 ) | ( n7201 & n41495 ) | ( ~n16099 & n41495 ) ;
  assign n41497 = n41496 ^ n22624 ^ 1'b0 ;
  assign n41498 = n14322 ^ n6269 ^ n5512 ;
  assign n41499 = ~n2819 & n16708 ;
  assign n41502 = n6789 | n16855 ;
  assign n41500 = n18350 ^ n13269 ^ 1'b0 ;
  assign n41501 = n28233 & n41500 ;
  assign n41503 = n41502 ^ n41501 ^ n24356 ;
  assign n41504 = n10228 & n17523 ;
  assign n41505 = n41504 ^ n31913 ^ n25853 ;
  assign n41506 = n4977 | n41505 ;
  assign n41507 = n34427 & ~n41506 ;
  assign n41508 = n12628 ^ n10974 ^ n2480 ;
  assign n41509 = ~n3997 & n41508 ;
  assign n41510 = n22072 | n41509 ;
  assign n41511 = n23897 & ~n41510 ;
  assign n41512 = n39607 ^ n7653 ^ 1'b0 ;
  assign n41513 = n2515 & ~n31883 ;
  assign n41514 = ( ~n3002 & n22075 ) | ( ~n3002 & n41513 ) | ( n22075 & n41513 ) ;
  assign n41515 = n10491 | n41514 ;
  assign n41516 = n7692 | n24627 ;
  assign n41517 = n41516 ^ n27660 ^ n13786 ;
  assign n41518 = n20799 ^ n6149 ^ 1'b0 ;
  assign n41519 = n4022 & n10739 ;
  assign n41520 = n38602 ^ n33463 ^ 1'b0 ;
  assign n41521 = ~x65 & n41520 ;
  assign n41522 = n11244 ^ n5804 ^ n1523 ;
  assign n41523 = n33721 & n41522 ;
  assign n41524 = ( n13171 & ~n18581 ) | ( n13171 & n41523 ) | ( ~n18581 & n41523 ) ;
  assign n41525 = ( n6255 & n12064 ) | ( n6255 & n29058 ) | ( n12064 & n29058 ) ;
  assign n41526 = n609 | n1682 ;
  assign n41527 = n41525 | n41526 ;
  assign n41528 = n41527 ^ n18827 ^ n4634 ;
  assign n41529 = n17226 ^ n12315 ^ 1'b0 ;
  assign n41530 = ( n924 & ~n9648 ) | ( n924 & n21805 ) | ( ~n9648 & n21805 ) ;
  assign n41531 = n36970 ^ n2377 ^ 1'b0 ;
  assign n41532 = ( n10522 & ~n41530 ) | ( n10522 & n41531 ) | ( ~n41530 & n41531 ) ;
  assign n41536 = ( n3261 & n14941 ) | ( n3261 & ~n24909 ) | ( n14941 & ~n24909 ) ;
  assign n41533 = n22437 & ~n32866 ;
  assign n41534 = ~x56 & n41533 ;
  assign n41535 = n41534 ^ n28344 ^ n11758 ;
  assign n41537 = n41536 ^ n41535 ^ 1'b0 ;
  assign n41538 = ( ~n4310 & n18893 ) | ( ~n4310 & n30607 ) | ( n18893 & n30607 ) ;
  assign n41539 = n11795 & n41538 ;
  assign n41540 = ~n11867 & n41539 ;
  assign n41541 = n32129 ^ n20663 ^ n11562 ;
  assign n41542 = ( n16386 & n23484 ) | ( n16386 & n29946 ) | ( n23484 & n29946 ) ;
  assign n41543 = n21665 ^ n3116 ^ 1'b0 ;
  assign n41544 = n41543 ^ n41237 ^ n3735 ;
  assign n41545 = ( ~n13218 & n25428 ) | ( ~n13218 & n41017 ) | ( n25428 & n41017 ) ;
  assign n41546 = n1995 & n30887 ;
  assign n41548 = ~n3820 & n16351 ;
  assign n41549 = n24961 & n41548 ;
  assign n41550 = n12361 & n37708 ;
  assign n41551 = n41549 & n41550 ;
  assign n41552 = n41551 ^ n16152 ^ 1'b0 ;
  assign n41553 = n5474 & ~n41552 ;
  assign n41547 = n14334 | n38535 ;
  assign n41554 = n41553 ^ n41547 ^ 1'b0 ;
  assign n41555 = n36564 ^ n3984 ^ x173 ;
  assign n41556 = n27389 ^ n25563 ^ 1'b0 ;
  assign n41560 = n8537 ^ n5183 ^ n4060 ;
  assign n41561 = n41560 ^ n25369 ^ 1'b0 ;
  assign n41562 = n22106 & n41561 ;
  assign n41557 = ( n3420 & n4922 ) | ( n3420 & n10372 ) | ( n4922 & n10372 ) ;
  assign n41558 = n3612 & ~n14330 ;
  assign n41559 = n41557 & n41558 ;
  assign n41563 = n41562 ^ n41559 ^ 1'b0 ;
  assign n41564 = ~n6372 & n26377 ;
  assign n41565 = n17058 ^ n3276 ^ 1'b0 ;
  assign n41566 = n41564 & n41565 ;
  assign n41567 = ( n16561 & n17156 ) | ( n16561 & n36781 ) | ( n17156 & n36781 ) ;
  assign n41568 = n40146 ^ n28974 ^ 1'b0 ;
  assign n41569 = ( n23216 & ~n41567 ) | ( n23216 & n41568 ) | ( ~n41567 & n41568 ) ;
  assign n41570 = n27621 & ~n41569 ;
  assign n41571 = n727 & n19908 ;
  assign n41572 = n3601 | n41571 ;
  assign n41573 = n41572 ^ n10458 ^ 1'b0 ;
  assign n41574 = n19144 | n41573 ;
  assign n41575 = n23557 & n41574 ;
  assign n41576 = ~n2885 & n41575 ;
  assign n41580 = n6277 ^ n3627 ^ 1'b0 ;
  assign n41581 = n4936 & n41580 ;
  assign n41582 = n41581 ^ n15377 ^ n3532 ;
  assign n41577 = n3923 & ~n32409 ;
  assign n41578 = n41577 ^ n467 ^ 1'b0 ;
  assign n41579 = ( n6494 & ~n31266 ) | ( n6494 & n41578 ) | ( ~n31266 & n41578 ) ;
  assign n41583 = n41582 ^ n41579 ^ 1'b0 ;
  assign n41584 = n36716 & n41583 ;
  assign n41585 = n27949 ^ n24206 ^ n5159 ;
  assign n41586 = n37384 ^ n21200 ^ 1'b0 ;
  assign n41587 = n41586 ^ n24147 ^ n11122 ;
  assign n41592 = n24519 ^ n9287 ^ n6418 ;
  assign n41593 = n28592 ^ n5676 ^ 1'b0 ;
  assign n41594 = ~n41592 & n41593 ;
  assign n41591 = n16472 ^ n14956 ^ n10480 ;
  assign n41588 = n22025 | n25242 ;
  assign n41589 = n41588 ^ n27564 ^ 1'b0 ;
  assign n41590 = n41589 ^ n32425 ^ n10327 ;
  assign n41595 = n41594 ^ n41591 ^ n41590 ;
  assign n41596 = n2416 & ~n5140 ;
  assign n41597 = n41596 ^ n40743 ^ 1'b0 ;
  assign n41598 = ~n22882 & n25315 ;
  assign n41599 = n29331 & n41067 ;
  assign n41600 = ~n15226 & n41599 ;
  assign n41601 = n15682 & n19095 ;
  assign n41602 = n41601 ^ n12826 ^ 1'b0 ;
  assign n41603 = n19961 | n24669 ;
  assign n41607 = n16871 ^ n12208 ^ 1'b0 ;
  assign n41608 = n22768 & n41607 ;
  assign n41604 = ( ~n533 & n4554 ) | ( ~n533 & n12558 ) | ( n4554 & n12558 ) ;
  assign n41605 = n19235 | n38186 ;
  assign n41606 = n41604 & ~n41605 ;
  assign n41609 = n41608 ^ n41606 ^ n3117 ;
  assign n41610 = n19142 ^ n16307 ^ 1'b0 ;
  assign n41611 = ( n8726 & n19284 ) | ( n8726 & ~n29348 ) | ( n19284 & ~n29348 ) ;
  assign n41612 = n6166 ^ n4678 ^ 1'b0 ;
  assign n41613 = ( n2700 & n6033 ) | ( n2700 & n6190 ) | ( n6033 & n6190 ) ;
  assign n41614 = n41613 ^ n12361 ^ 1'b0 ;
  assign n41615 = ( n21528 & n41612 ) | ( n21528 & n41614 ) | ( n41612 & n41614 ) ;
  assign n41616 = n37779 ^ n36779 ^ 1'b0 ;
  assign n41617 = n12249 & n41616 ;
  assign n41618 = ~n6992 & n13989 ;
  assign n41619 = ( n3883 & ~n16028 ) | ( n3883 & n41618 ) | ( ~n16028 & n41618 ) ;
  assign n41620 = n17421 ^ n11948 ^ 1'b0 ;
  assign n41621 = n4604 & ~n41620 ;
  assign n41622 = n41621 ^ n21805 ^ n18000 ;
  assign n41623 = n20920 & n41622 ;
  assign n41624 = n11044 & n41623 ;
  assign n41625 = n41619 & n41624 ;
  assign n41626 = ~n1746 & n29887 ;
  assign n41627 = n31655 & n41626 ;
  assign n41628 = n34235 ^ n21867 ^ n7291 ;
  assign n41629 = ( ~n23418 & n31624 ) | ( ~n23418 & n32247 ) | ( n31624 & n32247 ) ;
  assign n41632 = ( n8904 & n12820 ) | ( n8904 & ~n14875 ) | ( n12820 & ~n14875 ) ;
  assign n41630 = n10338 & ~n22925 ;
  assign n41631 = ( ~n6581 & n11206 ) | ( ~n6581 & n41630 ) | ( n11206 & n41630 ) ;
  assign n41633 = n41632 ^ n41631 ^ n37009 ;
  assign n41634 = n7103 ^ n5432 ^ 1'b0 ;
  assign n41635 = n16174 & ~n41634 ;
  assign n41636 = ( n17185 & ~n33748 ) | ( n17185 & n41635 ) | ( ~n33748 & n41635 ) ;
  assign n41637 = n41636 ^ n15196 ^ n8926 ;
  assign n41638 = ( n16186 & n22355 ) | ( n16186 & n23729 ) | ( n22355 & n23729 ) ;
  assign n41639 = ( ~n23183 & n30621 ) | ( ~n23183 & n41638 ) | ( n30621 & n41638 ) ;
  assign n41640 = ~n6433 & n22483 ;
  assign n41641 = ~n23598 & n41640 ;
  assign n41642 = n16005 & ~n22627 ;
  assign n41643 = n41641 & n41642 ;
  assign n41644 = n5123 | n39383 ;
  assign n41645 = n41644 ^ n1198 ^ 1'b0 ;
  assign n41646 = n14097 & ~n20226 ;
  assign n41647 = ( n11802 & n21707 ) | ( n11802 & ~n41646 ) | ( n21707 & ~n41646 ) ;
  assign n41648 = ~n13820 & n41647 ;
  assign n41649 = n25346 ^ n582 ^ 1'b0 ;
  assign n41650 = n30968 ^ n16498 ^ n4664 ;
  assign n41651 = n3456 | n5372 ;
  assign n41652 = n10247 | n41651 ;
  assign n41653 = n41652 ^ n27675 ^ n13271 ;
  assign n41654 = n36397 ^ n29287 ^ n547 ;
  assign n41655 = n1834 | n18518 ;
  assign n41656 = n35269 ^ n30964 ^ n28650 ;
  assign n41657 = ( n10327 & n41655 ) | ( n10327 & ~n41656 ) | ( n41655 & ~n41656 ) ;
  assign n41658 = n3228 & n25448 ;
  assign n41659 = n41658 ^ n15101 ^ 1'b0 ;
  assign n41660 = n17696 ^ n1473 ^ n293 ;
  assign n41661 = n41660 ^ n437 ^ 1'b0 ;
  assign n41662 = ~n41659 & n41661 ;
  assign n41663 = ( n994 & n9267 ) | ( n994 & ~n28771 ) | ( n9267 & ~n28771 ) ;
  assign n41664 = n27465 ^ n2256 ^ 1'b0 ;
  assign n41665 = n41664 ^ n37726 ^ n7873 ;
  assign n41666 = n18940 & n41665 ;
  assign n41667 = n41663 & n41666 ;
  assign n41668 = n5912 | n7896 ;
  assign n41669 = n41668 ^ n32391 ^ n18527 ;
  assign n41670 = n14716 & n41669 ;
  assign n41671 = ( n2015 & n12435 ) | ( n2015 & ~n15425 ) | ( n12435 & ~n15425 ) ;
  assign n41672 = ~n7597 & n40580 ;
  assign n41673 = ~n6219 & n41672 ;
  assign n41674 = ( n22878 & ~n41671 ) | ( n22878 & n41673 ) | ( ~n41671 & n41673 ) ;
  assign n41675 = ( ~n1326 & n3590 ) | ( ~n1326 & n41505 ) | ( n3590 & n41505 ) ;
  assign n41676 = n32912 ^ n21703 ^ n4938 ;
  assign n41677 = n40744 ^ n25538 ^ n23416 ;
  assign n41678 = n41677 ^ n18338 ^ 1'b0 ;
  assign n41679 = n13695 & ~n41678 ;
  assign n41680 = ( n20068 & ~n21494 ) | ( n20068 & n25707 ) | ( ~n21494 & n25707 ) ;
  assign n41683 = n28690 ^ n20583 ^ n1482 ;
  assign n41681 = n7270 & ~n11350 ;
  assign n41682 = n13379 & n41681 ;
  assign n41684 = n41683 ^ n41682 ^ n23000 ;
  assign n41685 = n1885 & ~n21388 ;
  assign n41686 = ~n29334 & n41685 ;
  assign n41687 = n41686 ^ n19701 ^ n13802 ;
  assign n41688 = n3475 & n36304 ;
  assign n41689 = n41688 ^ n21122 ^ n12863 ;
  assign n41690 = n41689 ^ n25039 ^ n2642 ;
  assign n41691 = n26494 ^ n9887 ^ 1'b0 ;
  assign n41692 = n8451 | n12460 ;
  assign n41693 = n6519 | n41692 ;
  assign n41694 = n21380 ^ n11653 ^ 1'b0 ;
  assign n41695 = ~n12050 & n41694 ;
  assign n41696 = n41695 ^ n26618 ^ 1'b0 ;
  assign n41697 = n21393 ^ n17031 ^ n4449 ;
  assign n41698 = n41697 ^ n9286 ^ 1'b0 ;
  assign n41699 = ~n7809 & n17968 ;
  assign n41700 = n17216 & ~n41699 ;
  assign n41701 = n17062 | n19225 ;
  assign n41702 = n18599 | n41701 ;
  assign n41703 = n41702 ^ n19152 ^ n1763 ;
  assign n41704 = n41703 ^ n29710 ^ n15973 ;
  assign n41705 = ( n5536 & n13904 ) | ( n5536 & n14299 ) | ( n13904 & n14299 ) ;
  assign n41706 = n33572 ^ n19610 ^ n19235 ;
  assign n41707 = ( ~x193 & n31993 ) | ( ~x193 & n41706 ) | ( n31993 & n41706 ) ;
  assign n41708 = ~n5567 & n39444 ;
  assign n41709 = n23597 ^ n5804 ^ 1'b0 ;
  assign n41710 = n16336 & ~n41709 ;
  assign n41711 = n7521 ^ n873 ^ 1'b0 ;
  assign n41712 = n8171 & ~n12527 ;
  assign n41713 = ( n4456 & n8594 ) | ( n4456 & n41712 ) | ( n8594 & n41712 ) ;
  assign n41714 = n41713 ^ n12945 ^ n4024 ;
  assign n41715 = ( n2596 & n26741 ) | ( n2596 & n41194 ) | ( n26741 & n41194 ) ;
  assign n41716 = n23235 & ~n30051 ;
  assign n41717 = n41716 ^ n6714 ^ 1'b0 ;
  assign n41718 = n19745 ^ n4828 ^ 1'b0 ;
  assign n41719 = n16621 | n41718 ;
  assign n41720 = ( n9973 & ~n37412 ) | ( n9973 & n41719 ) | ( ~n37412 & n41719 ) ;
  assign n41721 = n5725 ^ n4613 ^ n296 ;
  assign n41722 = n8045 & n41721 ;
  assign n41723 = n41722 ^ n14548 ^ 1'b0 ;
  assign n41724 = n22922 & n41723 ;
  assign n41725 = n6892 & n41724 ;
  assign n41726 = n40489 ^ n3011 ^ 1'b0 ;
  assign n41727 = n9877 & n41726 ;
  assign n41728 = ( ~n6481 & n10364 ) | ( ~n6481 & n41727 ) | ( n10364 & n41727 ) ;
  assign n41729 = n24067 ^ n517 ^ x31 ;
  assign n41730 = ( n5459 & n31397 ) | ( n5459 & ~n41729 ) | ( n31397 & ~n41729 ) ;
  assign n41731 = n31937 ^ n1343 ^ 1'b0 ;
  assign n41732 = n23265 ^ n17532 ^ 1'b0 ;
  assign n41733 = n6618 ^ n4458 ^ 1'b0 ;
  assign n41734 = n7731 & ~n41733 ;
  assign n41735 = ~n8247 & n41734 ;
  assign n41736 = ~n41732 & n41735 ;
  assign n41737 = n4095 ^ n2668 ^ 1'b0 ;
  assign n41738 = ~n32580 & n41737 ;
  assign n41739 = n1749 | n18476 ;
  assign n41740 = ( n6592 & ~n34683 ) | ( n6592 & n41739 ) | ( ~n34683 & n41739 ) ;
  assign n41741 = n17681 ^ n7042 ^ 1'b0 ;
  assign n41742 = n22169 & ~n41741 ;
  assign n41743 = ( n10281 & n11446 ) | ( n10281 & ~n41742 ) | ( n11446 & ~n41742 ) ;
  assign n41744 = n10829 | n41743 ;
  assign n41745 = n6448 ^ n2680 ^ 1'b0 ;
  assign n41746 = n24738 & ~n41745 ;
  assign n41747 = n33463 & n41746 ;
  assign n41748 = n41747 ^ n13217 ^ 1'b0 ;
  assign n41750 = ( n689 & n13924 ) | ( n689 & n17966 ) | ( n13924 & n17966 ) ;
  assign n41749 = n34522 ^ n23994 ^ n4868 ;
  assign n41751 = n41750 ^ n41749 ^ n13154 ;
  assign n41752 = n12371 | n16894 ;
  assign n41753 = n41752 ^ n6097 ^ 1'b0 ;
  assign n41754 = ( n35657 & n38255 ) | ( n35657 & n41753 ) | ( n38255 & n41753 ) ;
  assign n41755 = ( n9507 & ~n25484 ) | ( n9507 & n41754 ) | ( ~n25484 & n41754 ) ;
  assign n41756 = n18201 & n25423 ;
  assign n41757 = n4431 & n41756 ;
  assign n41758 = n8355 | n41757 ;
  assign n41759 = ( ~n2330 & n10570 ) | ( ~n2330 & n16911 ) | ( n10570 & n16911 ) ;
  assign n41760 = n41759 ^ n37961 ^ 1'b0 ;
  assign n41761 = n8206 & ~n41760 ;
  assign n41762 = n1073 & ~n41761 ;
  assign n41763 = n5827 & n41762 ;
  assign n41764 = n41763 ^ n7960 ^ 1'b0 ;
  assign n41765 = n19472 ^ n2500 ^ 1'b0 ;
  assign n41766 = n41765 ^ n27999 ^ 1'b0 ;
  assign n41767 = n41141 ^ n38315 ^ 1'b0 ;
  assign n41768 = n18725 & ~n41767 ;
  assign n41769 = n41768 ^ n26893 ^ 1'b0 ;
  assign n41770 = n10061 & n18424 ;
  assign n41771 = n41770 ^ n35601 ^ n21135 ;
  assign n41772 = n1052 & n8472 ;
  assign n41773 = n9184 & n41772 ;
  assign n41774 = n18522 & n26278 ;
  assign n41775 = n41773 & n41774 ;
  assign n41776 = n41775 ^ n35660 ^ 1'b0 ;
  assign n41778 = ( n291 & n1305 ) | ( n291 & n1803 ) | ( n1305 & n1803 ) ;
  assign n41779 = n36991 ^ n14741 ^ 1'b0 ;
  assign n41780 = ~n41778 & n41779 ;
  assign n41777 = ( n1784 & n5454 ) | ( n1784 & ~n28439 ) | ( n5454 & ~n28439 ) ;
  assign n41781 = n41780 ^ n41777 ^ n40772 ;
  assign n41782 = ( n6203 & n9368 ) | ( n6203 & n18823 ) | ( n9368 & n18823 ) ;
  assign n41783 = n41782 ^ n1842 ^ 1'b0 ;
  assign n41784 = n14474 ^ n11809 ^ 1'b0 ;
  assign n41785 = n7329 & ~n41784 ;
  assign n41786 = n41785 ^ n28605 ^ n23586 ;
  assign n41787 = n16359 | n41786 ;
  assign n41788 = ( n7605 & n8835 ) | ( n7605 & ~n38651 ) | ( n8835 & ~n38651 ) ;
  assign n41789 = n12590 | n41788 ;
  assign n41790 = n41789 ^ n27048 ^ 1'b0 ;
  assign n41791 = n16615 ^ n4421 ^ 1'b0 ;
  assign n41792 = n35254 & ~n41791 ;
  assign n41793 = n39068 ^ n26309 ^ n24862 ;
  assign n41794 = n14868 ^ n13563 ^ n11538 ;
  assign n41795 = n3832 | n32900 ;
  assign n41796 = ( n4601 & n15442 ) | ( n4601 & ~n27144 ) | ( n15442 & ~n27144 ) ;
  assign n41797 = n31571 | n34627 ;
  assign n41798 = n41797 ^ x17 ^ 1'b0 ;
  assign n41799 = n28004 | n41798 ;
  assign n41800 = n4820 ^ n957 ^ 1'b0 ;
  assign n41801 = n15976 & ~n41800 ;
  assign n41802 = ( n3750 & n30153 ) | ( n3750 & ~n33013 ) | ( n30153 & ~n33013 ) ;
  assign n41803 = ~n23104 & n41802 ;
  assign n41804 = ( n24676 & ~n41801 ) | ( n24676 & n41803 ) | ( ~n41801 & n41803 ) ;
  assign n41806 = ( ~n29108 & n39436 ) | ( ~n29108 & n39621 ) | ( n39436 & n39621 ) ;
  assign n41805 = n3057 | n3151 ;
  assign n41807 = n41806 ^ n41805 ^ 1'b0 ;
  assign n41808 = n9279 | n39068 ;
  assign n41809 = n35891 & ~n41808 ;
  assign n41810 = n17111 ^ n5218 ^ 1'b0 ;
  assign n41811 = ~n15751 & n41810 ;
  assign n41812 = ( n6778 & n30274 ) | ( n6778 & n41811 ) | ( n30274 & n41811 ) ;
  assign n41813 = n695 & n21036 ;
  assign n41814 = n41813 ^ n7466 ^ 1'b0 ;
  assign n41815 = ~n7523 & n41814 ;
  assign n41816 = ( n805 & ~n3819 ) | ( n805 & n36137 ) | ( ~n3819 & n36137 ) ;
  assign n41817 = n41815 & ~n41816 ;
  assign n41818 = n28507 ^ n23867 ^ n14707 ;
  assign n41820 = n22722 ^ n13817 ^ n12120 ;
  assign n41819 = n3026 & ~n3200 ;
  assign n41821 = n41820 ^ n41819 ^ 1'b0 ;
  assign n41822 = n39305 ^ n9499 ^ n5793 ;
  assign n41823 = n32672 ^ n2898 ^ 1'b0 ;
  assign n41824 = n41822 | n41823 ;
  assign n41825 = n2083 & ~n11460 ;
  assign n41826 = n20473 ^ n5960 ^ n3520 ;
  assign n41827 = n3609 & ~n25004 ;
  assign n41828 = n15184 | n34410 ;
  assign n41829 = n37391 ^ n11594 ^ n8877 ;
  assign n41830 = ( n41827 & ~n41828 ) | ( n41827 & n41829 ) | ( ~n41828 & n41829 ) ;
  assign n41831 = ~n23053 & n37524 ;
  assign n41832 = n22939 & n41831 ;
  assign n41833 = n8665 & n40736 ;
  assign n41834 = n41833 ^ n487 ^ 1'b0 ;
  assign n41835 = ~n6387 & n16469 ;
  assign n41836 = n41835 ^ n1655 ^ 1'b0 ;
  assign n41837 = n12497 | n41836 ;
  assign n41838 = n12854 | n41837 ;
  assign n41839 = ( ~n22712 & n41834 ) | ( ~n22712 & n41838 ) | ( n41834 & n41838 ) ;
  assign n41840 = n25537 ^ n7658 ^ n4553 ;
  assign n41843 = n40685 ^ n2066 ^ 1'b0 ;
  assign n41841 = n9342 | n10761 ;
  assign n41842 = n26820 & ~n41841 ;
  assign n41844 = n41843 ^ n41842 ^ 1'b0 ;
  assign n41845 = n17799 ^ n7825 ^ n5806 ;
  assign n41846 = ( n19905 & n34412 ) | ( n19905 & n41845 ) | ( n34412 & n41845 ) ;
  assign n41847 = n41846 ^ n17695 ^ n12305 ;
  assign n41848 = n41847 ^ n3625 ^ 1'b0 ;
  assign n41849 = ( n9026 & n11810 ) | ( n9026 & n27081 ) | ( n11810 & n27081 ) ;
  assign n41850 = n10742 & ~n12286 ;
  assign n41851 = n41849 & n41850 ;
  assign n41853 = ~n1789 & n16546 ;
  assign n41854 = n41853 ^ n8568 ^ 1'b0 ;
  assign n41852 = n2418 | n39963 ;
  assign n41855 = n41854 ^ n41852 ^ 1'b0 ;
  assign n41856 = ~n18418 & n20305 ;
  assign n41857 = ~n2210 & n41856 ;
  assign n41858 = n23558 ^ n1945 ^ 1'b0 ;
  assign n41859 = ~n41857 & n41858 ;
  assign n41860 = n41859 ^ n30671 ^ n27849 ;
  assign n41861 = n39065 ^ n32859 ^ n18602 ;
  assign n41862 = n41861 ^ n306 ^ 1'b0 ;
  assign n41863 = n38868 ^ n29324 ^ 1'b0 ;
  assign n41864 = ( n8296 & ~n33067 ) | ( n8296 & n39742 ) | ( ~n33067 & n39742 ) ;
  assign n41865 = ~n1524 & n27391 ;
  assign n41866 = ~n8105 & n41865 ;
  assign n41867 = n41866 ^ n22830 ^ n20686 ;
  assign n41868 = n36105 ^ n23719 ^ 1'b0 ;
  assign n41869 = n8835 & n41868 ;
  assign n41870 = n6146 ^ n4587 ^ 1'b0 ;
  assign n41871 = n41870 ^ n4111 ^ n1562 ;
  assign n41872 = n997 | n40614 ;
  assign n41873 = ~n11043 & n20460 ;
  assign n41874 = n41873 ^ n25149 ^ 1'b0 ;
  assign n41875 = ( ~n14052 & n37759 ) | ( ~n14052 & n41874 ) | ( n37759 & n41874 ) ;
  assign n41876 = ( n10009 & ~n29928 ) | ( n10009 & n41875 ) | ( ~n29928 & n41875 ) ;
  assign n41877 = n3188 & n29288 ;
  assign n41878 = ( n5514 & n10521 ) | ( n5514 & ~n41877 ) | ( n10521 & ~n41877 ) ;
  assign n41879 = n41878 ^ n6002 ^ 1'b0 ;
  assign n41880 = n40531 & n41879 ;
  assign n41881 = ( n13612 & n26415 ) | ( n13612 & ~n30175 ) | ( n26415 & ~n30175 ) ;
  assign n41882 = n41881 ^ n14628 ^ 1'b0 ;
  assign n41883 = n41880 & n41882 ;
  assign n41884 = n41883 ^ n18826 ^ n14587 ;
  assign n41885 = n17787 ^ n11479 ^ 1'b0 ;
  assign n41886 = n24980 | n41885 ;
  assign n41887 = n16887 & ~n41886 ;
  assign n41888 = n41887 ^ n38505 ^ n21406 ;
  assign n41889 = ~n2481 & n8134 ;
  assign n41890 = ~n15836 & n41889 ;
  assign n41891 = n41890 ^ n20289 ^ n16512 ;
  assign n41892 = n1885 & n36275 ;
  assign n41893 = n41892 ^ n40936 ^ 1'b0 ;
  assign n41894 = n41891 & ~n41893 ;
  assign n41895 = ( n28163 & n33437 ) | ( n28163 & ~n41894 ) | ( n33437 & ~n41894 ) ;
  assign n41896 = n1264 & n2474 ;
  assign n41897 = n27244 & n41896 ;
  assign n41898 = n19385 & ~n20217 ;
  assign n41899 = n810 & n41898 ;
  assign n41900 = ( n2702 & n9469 ) | ( n2702 & n13595 ) | ( n9469 & n13595 ) ;
  assign n41901 = n30864 & ~n41900 ;
  assign n41902 = n11389 & n17831 ;
  assign n41903 = ( n4965 & ~n15001 ) | ( n4965 & n22744 ) | ( ~n15001 & n22744 ) ;
  assign n41904 = ( n8056 & ~n34312 ) | ( n8056 & n39893 ) | ( ~n34312 & n39893 ) ;
  assign n41905 = n23214 ^ n13074 ^ n4024 ;
  assign n41906 = n41905 ^ n28532 ^ 1'b0 ;
  assign n41907 = ~n5551 & n32436 ;
  assign n41911 = n2143 | n20902 ;
  assign n41912 = n23948 & ~n41911 ;
  assign n41908 = n15603 ^ n5214 ^ n4568 ;
  assign n41909 = ( ~n6853 & n20755 ) | ( ~n6853 & n32516 ) | ( n20755 & n32516 ) ;
  assign n41910 = ( n15277 & n41908 ) | ( n15277 & n41909 ) | ( n41908 & n41909 ) ;
  assign n41913 = n41912 ^ n41910 ^ n30303 ;
  assign n41914 = n36934 ^ n5159 ^ 1'b0 ;
  assign n41915 = n23196 ^ n15153 ^ x196 ;
  assign n41916 = n41915 ^ n31654 ^ n23503 ;
  assign n41917 = ~n31656 & n41019 ;
  assign n41918 = n30785 ^ n16483 ^ 1'b0 ;
  assign n41919 = n41918 ^ n11275 ^ 1'b0 ;
  assign n41920 = n1071 & n41919 ;
  assign n41921 = ( ~n5671 & n15056 ) | ( ~n5671 & n40046 ) | ( n15056 & n40046 ) ;
  assign n41922 = n16580 | n41921 ;
  assign n41923 = n24996 & n35659 ;
  assign n41924 = n41923 ^ n14793 ^ 1'b0 ;
  assign n41925 = ( x45 & n26534 ) | ( x45 & ~n41924 ) | ( n26534 & ~n41924 ) ;
  assign n41926 = n18679 & n41925 ;
  assign n41927 = ~n22312 & n41926 ;
  assign n41928 = ( ~n9374 & n21065 ) | ( ~n9374 & n35770 ) | ( n21065 & n35770 ) ;
  assign n41929 = n30205 ^ n13159 ^ 1'b0 ;
  assign n41930 = n20213 & ~n41929 ;
  assign n41931 = ~n11931 & n41930 ;
  assign n41932 = n19647 ^ n2885 ^ 1'b0 ;
  assign n41933 = n11532 ^ n7735 ^ 1'b0 ;
  assign n41934 = n16042 & n41933 ;
  assign n41935 = n3352 | n10800 ;
  assign n41936 = n41935 ^ n33067 ^ 1'b0 ;
  assign n41937 = ( n23968 & ~n41934 ) | ( n23968 & n41936 ) | ( ~n41934 & n41936 ) ;
  assign n41938 = n25780 & n41937 ;
  assign n41942 = n4079 & ~n7803 ;
  assign n41943 = ~n10205 & n41942 ;
  assign n41941 = n22859 ^ n11760 ^ 1'b0 ;
  assign n41939 = n6399 ^ n3067 ^ 1'b0 ;
  assign n41940 = n41939 ^ n16640 ^ n4265 ;
  assign n41944 = n41943 ^ n41941 ^ n41940 ;
  assign n41945 = n3502 | n5939 ;
  assign n41946 = n5268 | n41945 ;
  assign n41947 = ~n2442 & n7902 ;
  assign n41948 = n41947 ^ n9028 ^ 1'b0 ;
  assign n41949 = ( n10591 & n19692 ) | ( n10591 & ~n34232 ) | ( n19692 & ~n34232 ) ;
  assign n41950 = ( ~n41946 & n41948 ) | ( ~n41946 & n41949 ) | ( n41948 & n41949 ) ;
  assign n41951 = n18735 ^ n12143 ^ n11809 ;
  assign n41952 = n4167 & n28264 ;
  assign n41953 = n12366 & n41952 ;
  assign n41954 = ~n41951 & n41953 ;
  assign n41955 = n28750 ^ n23168 ^ 1'b0 ;
  assign n41956 = n21873 ^ n9259 ^ 1'b0 ;
  assign n41957 = n9731 & n41956 ;
  assign n41958 = n28956 ^ n14789 ^ 1'b0 ;
  assign n41959 = n17981 ^ n14180 ^ n8807 ;
  assign n41960 = ( n388 & ~n5557 ) | ( n388 & n41959 ) | ( ~n5557 & n41959 ) ;
  assign n41961 = n18937 ^ n17520 ^ 1'b0 ;
  assign n41962 = ( n15798 & ~n40510 ) | ( n15798 & n41961 ) | ( ~n40510 & n41961 ) ;
  assign n41963 = ( n15325 & n25853 ) | ( n15325 & ~n41962 ) | ( n25853 & ~n41962 ) ;
  assign n41964 = ( n29344 & ~n39388 ) | ( n29344 & n41963 ) | ( ~n39388 & n41963 ) ;
  assign n41965 = n14571 & ~n16055 ;
  assign n41966 = ~n1288 & n41965 ;
  assign n41967 = n41966 ^ n27182 ^ 1'b0 ;
  assign n41968 = ~n1010 & n41967 ;
  assign n41969 = n1998 | n17155 ;
  assign n41970 = ( n41495 & n41968 ) | ( n41495 & n41969 ) | ( n41968 & n41969 ) ;
  assign n41971 = ( n362 & n11246 ) | ( n362 & ~n26845 ) | ( n11246 & ~n26845 ) ;
  assign n41976 = n4724 & n27872 ;
  assign n41975 = n6765 & ~n32480 ;
  assign n41972 = ~n13247 & n41081 ;
  assign n41973 = ~n9511 & n41972 ;
  assign n41974 = n21272 | n41973 ;
  assign n41977 = n41976 ^ n41975 ^ n41974 ;
  assign n41978 = ~n1294 & n38039 ;
  assign n41979 = n41978 ^ n332 ^ 1'b0 ;
  assign n41980 = ~n8754 & n24898 ;
  assign n41981 = n41980 ^ n30885 ^ 1'b0 ;
  assign n41982 = n27181 ^ n23324 ^ n20611 ;
  assign n41983 = n34992 ^ n17710 ^ n11850 ;
  assign n41984 = ( n550 & n690 ) | ( n550 & ~n41983 ) | ( n690 & ~n41983 ) ;
  assign n41985 = n23615 ^ n20662 ^ n13152 ;
  assign n41986 = n39403 ^ n19158 ^ 1'b0 ;
  assign n41987 = ~n35111 & n41986 ;
  assign n41988 = ( ~n285 & n7796 ) | ( ~n285 & n22150 ) | ( n7796 & n22150 ) ;
  assign n41989 = ( ~n10992 & n24240 ) | ( ~n10992 & n41988 ) | ( n24240 & n41988 ) ;
  assign n41990 = n41989 ^ n13385 ^ 1'b0 ;
  assign n41991 = n41990 ^ n4831 ^ 1'b0 ;
  assign n41992 = n4300 & n41991 ;
  assign n41993 = ( n19799 & n32015 ) | ( n19799 & ~n41992 ) | ( n32015 & ~n41992 ) ;
  assign n41994 = n41987 | n41993 ;
  assign n41995 = n22673 ^ n10138 ^ n983 ;
  assign n41997 = ~n7296 & n17687 ;
  assign n41998 = n27473 & ~n41997 ;
  assign n41999 = ( ~n21805 & n23604 ) | ( ~n21805 & n41998 ) | ( n23604 & n41998 ) ;
  assign n41996 = n12233 & n26033 ;
  assign n42000 = n41999 ^ n41996 ^ 1'b0 ;
  assign n42001 = ~n12725 & n30700 ;
  assign n42002 = n42001 ^ n12740 ^ 1'b0 ;
  assign n42003 = n42002 ^ n12887 ^ 1'b0 ;
  assign n42004 = n6602 & ~n42003 ;
  assign n42005 = n42004 ^ n18015 ^ 1'b0 ;
  assign n42006 = n3854 & ~n16097 ;
  assign n42007 = n12272 & n42006 ;
  assign n42008 = n42007 ^ n35154 ^ n22807 ;
  assign n42009 = ( n6304 & n20792 ) | ( n6304 & ~n22453 ) | ( n20792 & ~n22453 ) ;
  assign n42010 = n35297 ^ n926 ^ 1'b0 ;
  assign n42011 = n23612 ^ n22022 ^ 1'b0 ;
  assign n42012 = ~n3520 & n42011 ;
  assign n42013 = n42012 ^ n13218 ^ 1'b0 ;
  assign n42014 = n12034 | n30663 ;
  assign n42015 = n42014 ^ n9266 ^ n9260 ;
  assign n42016 = n42015 ^ n26493 ^ n15460 ;
  assign n42017 = ( ~n2638 & n18552 ) | ( ~n2638 & n32088 ) | ( n18552 & n32088 ) ;
  assign n42018 = ( ~n22254 & n39007 ) | ( ~n22254 & n42017 ) | ( n39007 & n42017 ) ;
  assign n42019 = ( n1585 & n18355 ) | ( n1585 & ~n42018 ) | ( n18355 & ~n42018 ) ;
  assign n42020 = n26414 ^ n19328 ^ n14500 ;
  assign n42021 = n42020 ^ n32941 ^ 1'b0 ;
  assign n42022 = n25093 & ~n42021 ;
  assign n42023 = n28175 ^ n26647 ^ 1'b0 ;
  assign n42024 = n42023 ^ n38299 ^ 1'b0 ;
  assign n42025 = ~n25918 & n42024 ;
  assign n42026 = n37328 ^ n36849 ^ n25687 ;
  assign n42029 = n22218 ^ n1230 ^ 1'b0 ;
  assign n42030 = ~n4884 & n42029 ;
  assign n42027 = n407 & ~n11541 ;
  assign n42028 = ~n5797 & n42027 ;
  assign n42031 = n42030 ^ n42028 ^ 1'b0 ;
  assign n42032 = ( n5400 & n23265 ) | ( n5400 & n39678 ) | ( n23265 & n39678 ) ;
  assign n42033 = n7295 & ~n19163 ;
  assign n42034 = ( n21399 & n42032 ) | ( n21399 & n42033 ) | ( n42032 & n42033 ) ;
  assign n42035 = n26314 ^ n17513 ^ 1'b0 ;
  assign n42036 = ~n7445 & n15914 ;
  assign n42037 = ~n9916 & n42036 ;
  assign n42038 = ( n6104 & n6204 ) | ( n6104 & ~n39722 ) | ( n6204 & ~n39722 ) ;
  assign n42039 = n30993 ^ n29809 ^ n10939 ;
  assign n42040 = ( ~n34844 & n39388 ) | ( ~n34844 & n42039 ) | ( n39388 & n42039 ) ;
  assign n42041 = ( n17511 & n27208 ) | ( n17511 & ~n42040 ) | ( n27208 & ~n42040 ) ;
  assign n42043 = n12889 | n37104 ;
  assign n42042 = n32736 ^ n17135 ^ n6653 ;
  assign n42044 = n42043 ^ n42042 ^ n27456 ;
  assign n42045 = n42044 ^ n19270 ^ n17430 ;
  assign n42046 = n13048 ^ n4984 ^ n4378 ;
  assign n42047 = n42046 ^ n16878 ^ n14050 ;
  assign n42048 = n42047 ^ n39046 ^ n38232 ;
  assign n42049 = ~n10898 & n11657 ;
  assign n42050 = ~n4033 & n42049 ;
  assign n42051 = n2319 | n19599 ;
  assign n42052 = n42051 ^ n11033 ^ 1'b0 ;
  assign n42053 = ( n24648 & n26534 ) | ( n24648 & n34416 ) | ( n26534 & n34416 ) ;
  assign n42056 = n1312 & ~n4776 ;
  assign n42057 = n42056 ^ n27720 ^ 1'b0 ;
  assign n42054 = ( n1239 & ~n15124 ) | ( n1239 & n37880 ) | ( ~n15124 & n37880 ) ;
  assign n42055 = n42054 ^ n19913 ^ n7702 ;
  assign n42058 = n42057 ^ n42055 ^ n35159 ;
  assign n42059 = n11420 ^ n1516 ^ 1'b0 ;
  assign n42060 = ( n13111 & ~n14379 ) | ( n13111 & n15045 ) | ( ~n14379 & n15045 ) ;
  assign n42061 = n25754 ^ n20047 ^ 1'b0 ;
  assign n42062 = ( n42059 & ~n42060 ) | ( n42059 & n42061 ) | ( ~n42060 & n42061 ) ;
  assign n42063 = n36746 ^ n31835 ^ 1'b0 ;
  assign n42064 = n12307 ^ n7887 ^ 1'b0 ;
  assign n42065 = ~n21780 & n42064 ;
  assign n42066 = n14342 | n28205 ;
  assign n42067 = n42065 & ~n42066 ;
  assign n42068 = ~n6878 & n34731 ;
  assign n42069 = n31890 ^ n14777 ^ n11643 ;
  assign n42070 = n15968 ^ n15879 ^ 1'b0 ;
  assign n42071 = n10269 | n42070 ;
  assign n42072 = n26776 ^ n650 ^ 1'b0 ;
  assign n42073 = n42071 | n42072 ;
  assign n42074 = ( n12099 & ~n24093 ) | ( n12099 & n42073 ) | ( ~n24093 & n42073 ) ;
  assign n42075 = n42074 ^ n39931 ^ n18829 ;
  assign n42079 = ~x194 & n26349 ;
  assign n42078 = n39044 ^ n18200 ^ n16980 ;
  assign n42076 = ( ~n14909 & n15868 ) | ( ~n14909 & n15925 ) | ( n15868 & n15925 ) ;
  assign n42077 = n33507 & n42076 ;
  assign n42080 = n42079 ^ n42078 ^ n42077 ;
  assign n42081 = n20632 & n25334 ;
  assign n42082 = n3320 & n42081 ;
  assign n42083 = n42082 ^ n34338 ^ n33123 ;
  assign n42084 = n19223 ^ n806 ^ 1'b0 ;
  assign n42085 = n3791 & n42084 ;
  assign n42086 = ~n6351 & n11273 ;
  assign n42087 = n42086 ^ n15790 ^ n10025 ;
  assign n42088 = ~n10708 & n12834 ;
  assign n42089 = ~n14023 & n42088 ;
  assign n42090 = n384 & ~n16306 ;
  assign n42091 = n5888 & n31276 ;
  assign n42092 = ( n8889 & ~n32589 ) | ( n8889 & n42091 ) | ( ~n32589 & n42091 ) ;
  assign n42093 = n1227 | n10290 ;
  assign n42094 = n2315 & n42093 ;
  assign n42095 = ~n2964 & n7367 ;
  assign n42096 = n2155 & n42095 ;
  assign n42097 = ( n2155 & n17289 ) | ( n2155 & n42096 ) | ( n17289 & n42096 ) ;
  assign n42098 = n22306 ^ n8689 ^ n4465 ;
  assign n42099 = ( n1108 & ~n2123 ) | ( n1108 & n2671 ) | ( ~n2123 & n2671 ) ;
  assign n42100 = n1416 & n8350 ;
  assign n42101 = n3559 & n42100 ;
  assign n42102 = n22555 & n31485 ;
  assign n42103 = n42102 ^ n8456 ^ 1'b0 ;
  assign n42104 = n9450 & ~n42103 ;
  assign n42105 = n42101 & n42104 ;
  assign n42106 = ( ~x130 & n42099 ) | ( ~x130 & n42105 ) | ( n42099 & n42105 ) ;
  assign n42107 = n23781 ^ n17578 ^ n5645 ;
  assign n42108 = n42107 ^ n40561 ^ n32599 ;
  assign n42109 = n1850 | n42108 ;
  assign n42110 = n9912 & ~n42109 ;
  assign n42111 = n25950 ^ n12350 ^ 1'b0 ;
  assign n42112 = ( n17822 & ~n23732 ) | ( n17822 & n25427 ) | ( ~n23732 & n25427 ) ;
  assign n42113 = n32674 ^ n16204 ^ n8661 ;
  assign n42114 = n18468 ^ n17571 ^ n1233 ;
  assign n42115 = n11801 & n16784 ;
  assign n42116 = n13554 | n32047 ;
  assign n42117 = n42116 ^ n37541 ^ x84 ;
  assign n42118 = ( n30190 & n42115 ) | ( n30190 & ~n42117 ) | ( n42115 & ~n42117 ) ;
  assign n42119 = n7248 | n42118 ;
  assign n42120 = n20803 | n23549 ;
  assign n42121 = n42120 ^ n17081 ^ 1'b0 ;
  assign n42122 = ( ~n19178 & n23683 ) | ( ~n19178 & n42121 ) | ( n23683 & n42121 ) ;
  assign n42123 = n16179 & n28359 ;
  assign n42124 = n42123 ^ n9571 ^ 1'b0 ;
  assign n42125 = n22277 ^ n21741 ^ n3542 ;
  assign n42126 = n42124 | n42125 ;
  assign n42127 = ~n9691 & n31777 ;
  assign n42128 = n42127 ^ n15016 ^ 1'b0 ;
  assign n42129 = n42128 ^ n17706 ^ 1'b0 ;
  assign n42130 = n8015 & n42129 ;
  assign n42131 = ~n14593 & n20024 ;
  assign n42132 = n42131 ^ n23763 ^ 1'b0 ;
  assign n42133 = n1562 & n2392 ;
  assign n42134 = ( n485 & n670 ) | ( n485 & n5001 ) | ( n670 & n5001 ) ;
  assign n42135 = n42134 ^ n20554 ^ 1'b0 ;
  assign n42136 = ( n5786 & n21818 ) | ( n5786 & ~n26066 ) | ( n21818 & ~n26066 ) ;
  assign n42137 = n33675 ^ n2256 ^ 1'b0 ;
  assign n42138 = ( n25027 & ~n30478 ) | ( n25027 & n41522 ) | ( ~n30478 & n41522 ) ;
  assign n42139 = x177 & n8440 ;
  assign n42140 = n42139 ^ n20794 ^ 1'b0 ;
  assign n42141 = ( n4883 & ~n13731 ) | ( n4883 & n27465 ) | ( ~n13731 & n27465 ) ;
  assign n42142 = n42141 ^ n6049 ^ 1'b0 ;
  assign n42143 = n10067 & n42142 ;
  assign n42144 = ( n992 & n7629 ) | ( n992 & n8438 ) | ( n7629 & n8438 ) ;
  assign n42145 = n33010 | n42144 ;
  assign n42146 = n1887 | n42145 ;
  assign n42147 = ( n9317 & n33018 ) | ( n9317 & n42146 ) | ( n33018 & n42146 ) ;
  assign n42148 = ~n10683 & n42147 ;
  assign n42149 = ~n10129 & n42148 ;
  assign n42150 = n3634 & n30520 ;
  assign n42151 = ~n29081 & n42150 ;
  assign n42152 = n42151 ^ n22348 ^ n19973 ;
  assign n42153 = n40310 ^ n29620 ^ n16216 ;
  assign n42154 = n35325 ^ n22746 ^ n20528 ;
  assign n42155 = n42154 ^ n18015 ^ n13165 ;
  assign n42156 = n3569 & ~n38603 ;
  assign n42157 = n37131 ^ n32436 ^ n9572 ;
  assign n42158 = n19407 ^ n14952 ^ 1'b0 ;
  assign n42159 = ~n11353 & n22330 ;
  assign n42160 = ~n6825 & n42159 ;
  assign n42161 = n42160 ^ n12431 ^ 1'b0 ;
  assign n42162 = n6966 & n42161 ;
  assign n42163 = n42162 ^ n33642 ^ 1'b0 ;
  assign n42164 = n8735 | n34239 ;
  assign n42165 = n42163 | n42164 ;
  assign n42166 = n3179 & ~n27190 ;
  assign n42167 = n42166 ^ n9456 ^ 1'b0 ;
  assign n42168 = n8713 & ~n33933 ;
  assign n42169 = n42167 & n42168 ;
  assign n42170 = n32348 ^ n27376 ^ 1'b0 ;
  assign n42171 = n42170 ^ n32040 ^ n15777 ;
  assign n42172 = n9895 & n31472 ;
  assign n42173 = n42172 ^ n20172 ^ 1'b0 ;
  assign n42174 = n42173 ^ n22332 ^ n16951 ;
  assign n42175 = ~n6086 & n18151 ;
  assign n42176 = n42175 ^ n4068 ^ 1'b0 ;
  assign n42177 = n42176 ^ n18138 ^ 1'b0 ;
  assign n42178 = n16715 ^ n5546 ^ 1'b0 ;
  assign n42179 = ( n1737 & n9602 ) | ( n1737 & n42178 ) | ( n9602 & n42178 ) ;
  assign n42180 = n42179 ^ n30545 ^ n24423 ;
  assign n42181 = n9296 | n29846 ;
  assign n42182 = n42181 ^ n3022 ^ 1'b0 ;
  assign n42183 = n38334 ^ n14916 ^ 1'b0 ;
  assign n42184 = ~n16942 & n42183 ;
  assign n42185 = n6024 & n29856 ;
  assign n42186 = ( ~n14207 & n20900 ) | ( ~n14207 & n38442 ) | ( n20900 & n38442 ) ;
  assign n42187 = n42186 ^ n26783 ^ 1'b0 ;
  assign n42188 = ~n9681 & n36495 ;
  assign n42189 = ~n42187 & n42188 ;
  assign n42190 = n40264 ^ n30331 ^ n4604 ;
  assign n42191 = n42190 ^ n40207 ^ n37920 ;
  assign n42192 = n37730 ^ n25440 ^ n22561 ;
  assign n42193 = n14076 & ~n38269 ;
  assign n42194 = n42193 ^ n33524 ^ 1'b0 ;
  assign n42195 = ~n3909 & n26062 ;
  assign n42196 = n42195 ^ n24891 ^ 1'b0 ;
  assign n42197 = ~n1400 & n42196 ;
  assign n42198 = n4084 | n6584 ;
  assign n42202 = n7662 | n25358 ;
  assign n42201 = n22965 ^ n13712 ^ 1'b0 ;
  assign n42199 = n5623 | n33956 ;
  assign n42200 = n26852 & ~n42199 ;
  assign n42203 = n42202 ^ n42201 ^ n42200 ;
  assign n42204 = n20053 ^ n19331 ^ n1299 ;
  assign n42205 = n15821 ^ n12923 ^ 1'b0 ;
  assign n42206 = n3026 & n34938 ;
  assign n42207 = n40170 & n42206 ;
  assign n42208 = n1664 | n42207 ;
  assign n42209 = n36746 | n42208 ;
  assign n42210 = n7663 & ~n15142 ;
  assign n42211 = n3022 & n42210 ;
  assign n42214 = n19523 ^ n12552 ^ n8523 ;
  assign n42212 = ( n2546 & n4449 ) | ( n2546 & n7235 ) | ( n4449 & n7235 ) ;
  assign n42213 = n716 | n42212 ;
  assign n42215 = n42214 ^ n42213 ^ 1'b0 ;
  assign n42216 = n13487 | n42215 ;
  assign n42217 = n42216 ^ n14425 ^ 1'b0 ;
  assign n42218 = n6683 | n11332 ;
  assign n42219 = n12854 & n42218 ;
  assign n42220 = n16011 ^ n12589 ^ 1'b0 ;
  assign n42221 = ( ~n3949 & n22486 ) | ( ~n3949 & n28974 ) | ( n22486 & n28974 ) ;
  assign n42222 = n779 | n42221 ;
  assign n42223 = n18325 | n42222 ;
  assign n42224 = ~n4458 & n12859 ;
  assign n42225 = ~n13132 & n42224 ;
  assign n42226 = ( n5710 & n6077 ) | ( n5710 & n9721 ) | ( n6077 & n9721 ) ;
  assign n42227 = n42226 ^ n10933 ^ n9053 ;
  assign n42228 = n5838 | n42227 ;
  assign n42229 = ~n42225 & n42228 ;
  assign n42230 = ~n42223 & n42229 ;
  assign n42231 = n42230 ^ n20779 ^ n19107 ;
  assign n42232 = n2535 ^ n501 ^ 1'b0 ;
  assign n42233 = ~n19322 & n42232 ;
  assign n42234 = n6740 & ~n7910 ;
  assign n42235 = ~n42233 & n42234 ;
  assign n42236 = n42235 ^ n40316 ^ n37092 ;
  assign n42237 = n27406 ^ n8156 ^ 1'b0 ;
  assign n42238 = n10345 | n10960 ;
  assign n42239 = n42238 ^ n14657 ^ 1'b0 ;
  assign n42240 = ( ~n8906 & n18962 ) | ( ~n8906 & n42239 ) | ( n18962 & n42239 ) ;
  assign n42241 = n18884 & ~n26583 ;
  assign n42242 = ~n29676 & n42241 ;
  assign n42243 = ( n3138 & n21888 ) | ( n3138 & n42242 ) | ( n21888 & n42242 ) ;
  assign n42244 = n8027 & ~n10858 ;
  assign n42245 = n42243 & n42244 ;
  assign n42246 = n42240 & ~n42245 ;
  assign n42247 = n10388 & n42246 ;
  assign n42248 = n26569 & n27169 ;
  assign n42249 = n822 & n31376 ;
  assign n42250 = n42249 ^ n4761 ^ 1'b0 ;
  assign n42251 = n20269 ^ n18030 ^ n9552 ;
  assign n42252 = ( n7671 & n13513 ) | ( n7671 & n42251 ) | ( n13513 & n42251 ) ;
  assign n42253 = ( n13144 & n21072 ) | ( n13144 & n33067 ) | ( n21072 & n33067 ) ;
  assign n42254 = n29526 ^ n12694 ^ n11540 ;
  assign n42255 = n38216 ^ n35846 ^ n5991 ;
  assign n42256 = n35314 ^ n34448 ^ n13351 ;
  assign n42257 = n18306 & n42256 ;
  assign n42258 = ~n4941 & n39797 ;
  assign n42259 = ( n10517 & n19106 ) | ( n10517 & ~n31740 ) | ( n19106 & ~n31740 ) ;
  assign n42260 = n42259 ^ n30497 ^ 1'b0 ;
  assign n42261 = ~n13475 & n42260 ;
  assign n42262 = ~n28232 & n29896 ;
  assign n42263 = n26030 ^ n18747 ^ n17135 ;
  assign n42264 = n33506 ^ n30301 ^ n4967 ;
  assign n42267 = n42154 ^ n3216 ^ 1'b0 ;
  assign n42265 = n2668 & n35156 ;
  assign n42266 = n42265 ^ n14062 ^ 1'b0 ;
  assign n42268 = n42267 ^ n42266 ^ n23064 ;
  assign n42269 = ( x92 & n14169 ) | ( x92 & ~n41298 ) | ( n14169 & ~n41298 ) ;
  assign n42270 = n27345 ^ n19711 ^ n7228 ;
  assign n42271 = n42270 ^ n20019 ^ 1'b0 ;
  assign n42272 = ~n1822 & n16849 ;
  assign n42273 = n17299 & n34426 ;
  assign n42274 = n42272 & n42273 ;
  assign n42275 = n2500 | n9662 ;
  assign n42276 = n42275 ^ n14927 ^ n2569 ;
  assign n42277 = n42276 ^ n13373 ^ 1'b0 ;
  assign n42279 = n4078 ^ n2734 ^ n2722 ;
  assign n42280 = n8296 & n42279 ;
  assign n42281 = n20650 | n42280 ;
  assign n42278 = n12958 & ~n37260 ;
  assign n42282 = n42281 ^ n42278 ^ 1'b0 ;
  assign n42283 = n2179 & ~n9702 ;
  assign n42284 = n42282 & n42283 ;
  assign n42288 = n9784 ^ n7125 ^ 1'b0 ;
  assign n42285 = n24894 ^ n5524 ^ n350 ;
  assign n42286 = ( n2743 & n10372 ) | ( n2743 & n42285 ) | ( n10372 & n42285 ) ;
  assign n42287 = n42286 ^ n30261 ^ 1'b0 ;
  assign n42289 = n42288 ^ n42287 ^ n6558 ;
  assign n42290 = ( n11132 & ~n17636 ) | ( n11132 & n18829 ) | ( ~n17636 & n18829 ) ;
  assign n42291 = ( n11633 & n31228 ) | ( n11633 & n42290 ) | ( n31228 & n42290 ) ;
  assign n42292 = n35608 ^ n35493 ^ n31469 ;
  assign n42293 = n37209 ^ n18403 ^ 1'b0 ;
  assign n42294 = n1185 | n21750 ;
  assign n42295 = n42294 ^ n28106 ^ 1'b0 ;
  assign n42296 = ( ~n13432 & n20129 ) | ( ~n13432 & n42295 ) | ( n20129 & n42295 ) ;
  assign n42297 = n42296 ^ n37399 ^ n31614 ;
  assign n42298 = n40465 ^ n38383 ^ n37711 ;
  assign n42299 = n42298 ^ n1297 ^ 1'b0 ;
  assign n42300 = n41829 | n42299 ;
  assign n42301 = n23551 ^ n14045 ^ 1'b0 ;
  assign n42302 = n42301 ^ n25617 ^ 1'b0 ;
  assign n42303 = n34265 | n42302 ;
  assign n42304 = n31895 | n32070 ;
  assign n42305 = n42304 ^ n14278 ^ 1'b0 ;
  assign n42306 = n30758 & n42305 ;
  assign n42307 = n22416 & n42306 ;
  assign n42308 = n8621 & ~n14232 ;
  assign n42309 = ( n7630 & n38757 ) | ( n7630 & ~n42308 ) | ( n38757 & ~n42308 ) ;
  assign n42310 = n40793 ^ n39938 ^ n896 ;
  assign n42311 = ~n1114 & n12764 ;
  assign n42312 = n4791 & n42311 ;
  assign n42313 = ( n7475 & ~n8672 ) | ( n7475 & n42312 ) | ( ~n8672 & n42312 ) ;
  assign n42314 = ( n20123 & n24953 ) | ( n20123 & n42313 ) | ( n24953 & n42313 ) ;
  assign n42315 = n40618 ^ n28975 ^ 1'b0 ;
  assign n42316 = ( n903 & ~n19738 ) | ( n903 & n33257 ) | ( ~n19738 & n33257 ) ;
  assign n42317 = n42316 ^ n3934 ^ 1'b0 ;
  assign n42318 = n10163 & n42317 ;
  assign n42319 = n30162 ^ n18344 ^ n16508 ;
  assign n42320 = ~n18479 & n22488 ;
  assign n42321 = ( ~n1072 & n42319 ) | ( ~n1072 & n42320 ) | ( n42319 & n42320 ) ;
  assign n42327 = n26450 ^ n21573 ^ n1262 ;
  assign n42328 = n19848 ^ n7288 ^ 1'b0 ;
  assign n42329 = n42327 & ~n42328 ;
  assign n42324 = ( n13241 & ~n20582 ) | ( n13241 & n27035 ) | ( ~n20582 & n27035 ) ;
  assign n42322 = n22873 ^ n5966 ^ n5212 ;
  assign n42323 = n35609 & n42322 ;
  assign n42325 = n42324 ^ n42323 ^ 1'b0 ;
  assign n42326 = n39710 & n42325 ;
  assign n42330 = n42329 ^ n42326 ^ n39677 ;
  assign n42334 = n23758 ^ n6390 ^ n2099 ;
  assign n42331 = n12170 | n19111 ;
  assign n42332 = n42331 ^ n18532 ^ 1'b0 ;
  assign n42333 = ( n2924 & n26207 ) | ( n2924 & n42332 ) | ( n26207 & n42332 ) ;
  assign n42335 = n42334 ^ n42333 ^ n33557 ;
  assign n42336 = ~n2213 & n6716 ;
  assign n42337 = n42336 ^ n9760 ^ 1'b0 ;
  assign n42338 = ( ~n14607 & n17278 ) | ( ~n14607 & n35189 ) | ( n17278 & n35189 ) ;
  assign n42339 = n42337 | n42338 ;
  assign n42340 = ( n9238 & ~n9728 ) | ( n9238 & n34306 ) | ( ~n9728 & n34306 ) ;
  assign n42341 = n4674 ^ n3697 ^ n745 ;
  assign n42342 = ( n15024 & n26699 ) | ( n15024 & ~n42341 ) | ( n26699 & ~n42341 ) ;
  assign n42343 = n13188 | n42342 ;
  assign n42344 = n42343 ^ n37201 ^ 1'b0 ;
  assign n42345 = ~n1713 & n21917 ;
  assign n42346 = n42345 ^ n5146 ^ 1'b0 ;
  assign n42347 = n42346 ^ n2497 ^ 1'b0 ;
  assign n42348 = ( n2895 & n18874 ) | ( n2895 & n21352 ) | ( n18874 & n21352 ) ;
  assign n42349 = ~n12612 & n42348 ;
  assign n42350 = ( n310 & n20063 ) | ( n310 & n42349 ) | ( n20063 & n42349 ) ;
  assign n42351 = n5262 & ~n22656 ;
  assign n42352 = ~n25329 & n42351 ;
  assign n42353 = n8013 | n9148 ;
  assign n42354 = n16438 & ~n42353 ;
  assign n42355 = n42352 | n42354 ;
  assign n42356 = n24040 ^ n19383 ^ n17332 ;
  assign n42357 = n35240 & n40686 ;
  assign n42358 = n42357 ^ n12799 ^ 1'b0 ;
  assign n42359 = n26992 ^ n22996 ^ 1'b0 ;
  assign n42360 = n1331 & ~n42359 ;
  assign n42361 = n42360 ^ n994 ^ 1'b0 ;
  assign n42362 = n17640 & n24640 ;
  assign n42363 = ~n19455 & n42362 ;
  assign n42364 = ( n12424 & ~n24013 ) | ( n12424 & n36790 ) | ( ~n24013 & n36790 ) ;
  assign n42365 = ( n17657 & n42363 ) | ( n17657 & n42364 ) | ( n42363 & n42364 ) ;
  assign n42366 = n19844 ^ n6987 ^ n6367 ;
  assign n42368 = ( n4381 & ~n6855 ) | ( n4381 & n8592 ) | ( ~n6855 & n8592 ) ;
  assign n42367 = n7845 ^ n5946 ^ n3764 ;
  assign n42369 = n42368 ^ n42367 ^ n19584 ;
  assign n42370 = ( n4806 & n20311 ) | ( n4806 & n42369 ) | ( n20311 & n42369 ) ;
  assign n42371 = n21651 & ~n40815 ;
  assign n42372 = n3583 & ~n42371 ;
  assign n42373 = n42372 ^ n36293 ^ 1'b0 ;
  assign n42374 = n29502 & n33246 ;
  assign n42375 = n42373 & n42374 ;
  assign n42376 = n26545 ^ n2900 ^ 1'b0 ;
  assign n42377 = n23078 | n42376 ;
  assign n42378 = n42377 ^ n1572 ^ 1'b0 ;
  assign n42379 = n13700 & ~n26447 ;
  assign n42380 = ~n11392 & n27205 ;
  assign n42381 = n42012 ^ n28390 ^ n683 ;
  assign n42382 = ( n42379 & n42380 ) | ( n42379 & ~n42381 ) | ( n42380 & ~n42381 ) ;
  assign n42383 = n5303 & ~n6711 ;
  assign n42384 = n12636 & ~n14529 ;
  assign n42385 = n42384 ^ n35338 ^ n4575 ;
  assign n42386 = n25073 ^ n12746 ^ 1'b0 ;
  assign n42387 = n42386 ^ n19535 ^ n12128 ;
  assign n42388 = n42387 ^ n31236 ^ n14245 ;
  assign n42389 = ( n15008 & n19189 ) | ( n15008 & n21147 ) | ( n19189 & n21147 ) ;
  assign n42390 = n42388 & ~n42389 ;
  assign n42392 = ( ~n2463 & n11831 ) | ( ~n2463 & n33244 ) | ( n11831 & n33244 ) ;
  assign n42391 = ~n3169 & n3781 ;
  assign n42393 = n42392 ^ n42391 ^ 1'b0 ;
  assign n42394 = ( ~n7758 & n7929 ) | ( ~n7758 & n40011 ) | ( n7929 & n40011 ) ;
  assign n42395 = n42394 ^ n18706 ^ 1'b0 ;
  assign n42396 = n24612 & n42395 ;
  assign n42397 = ( n9226 & n20314 ) | ( n9226 & ~n38414 ) | ( n20314 & ~n38414 ) ;
  assign n42398 = n4118 ^ n2845 ^ n453 ;
  assign n42399 = n30200 ^ n28732 ^ n21820 ;
  assign n42400 = n42399 ^ n33600 ^ n9162 ;
  assign n42401 = n42400 ^ n19585 ^ 1'b0 ;
  assign n42402 = ( ~n12312 & n42398 ) | ( ~n12312 & n42401 ) | ( n42398 & n42401 ) ;
  assign n42403 = ~n14803 & n37543 ;
  assign n42404 = ~n39318 & n42403 ;
  assign n42405 = ( n13160 & ~n16449 ) | ( n13160 & n42404 ) | ( ~n16449 & n42404 ) ;
  assign n42406 = n9074 & n22333 ;
  assign n42407 = n22379 & n42406 ;
  assign n42408 = n17940 ^ n2706 ^ 1'b0 ;
  assign n42409 = n29518 ^ n2327 ^ 1'b0 ;
  assign n42410 = n26957 ^ n15377 ^ 1'b0 ;
  assign n42411 = n42409 & ~n42410 ;
  assign n42412 = n3080 | n4442 ;
  assign n42413 = ( n14279 & ~n14352 ) | ( n14279 & n42412 ) | ( ~n14352 & n42412 ) ;
  assign n42414 = ( ~n17822 & n22506 ) | ( ~n17822 & n40319 ) | ( n22506 & n40319 ) ;
  assign n42415 = n18312 ^ n11952 ^ 1'b0 ;
  assign n42416 = n22722 & n42415 ;
  assign n42417 = n42416 ^ n30516 ^ n12181 ;
  assign n42418 = n22805 ^ n1135 ^ 1'b0 ;
  assign n42419 = ~n8861 & n12001 ;
  assign n42420 = n7423 & n42419 ;
  assign n42421 = n22165 ^ n5050 ^ n838 ;
  assign n42422 = n1821 & ~n4946 ;
  assign n42423 = ~n42421 & n42422 ;
  assign n42428 = n27182 ^ n575 ^ 1'b0 ;
  assign n42429 = n42428 ^ n18525 ^ n1631 ;
  assign n42424 = n2325 ^ x174 ^ 1'b0 ;
  assign n42425 = n42424 ^ n12957 ^ 1'b0 ;
  assign n42426 = n7705 & ~n42425 ;
  assign n42427 = ~n11395 & n42426 ;
  assign n42430 = n42429 ^ n42427 ^ 1'b0 ;
  assign n42431 = n14527 ^ n4520 ^ n1403 ;
  assign n42432 = n15114 & n42431 ;
  assign n42433 = n40881 ^ n10907 ^ n2617 ;
  assign n42434 = n35618 ^ n27725 ^ n1239 ;
  assign n42435 = n1020 & n42434 ;
  assign n42436 = ( n12503 & ~n24304 ) | ( n12503 & n26482 ) | ( ~n24304 & n26482 ) ;
  assign n42437 = ( n10361 & n10800 ) | ( n10361 & ~n26730 ) | ( n10800 & ~n26730 ) ;
  assign n42438 = n4456 & n7110 ;
  assign n42439 = ~n23836 & n42438 ;
  assign n42440 = n15121 & n31286 ;
  assign n42441 = n41057 & n42440 ;
  assign n42442 = n6666 | n18285 ;
  assign n42443 = n42442 ^ n2908 ^ 1'b0 ;
  assign n42444 = n6029 & n42443 ;
  assign n42445 = n42444 ^ n40799 ^ 1'b0 ;
  assign n42446 = n11578 ^ n521 ^ 1'b0 ;
  assign n42447 = n32143 | n42446 ;
  assign n42448 = n8320 & ~n42447 ;
  assign n42450 = ( n1538 & n4831 ) | ( n1538 & ~n33852 ) | ( n4831 & ~n33852 ) ;
  assign n42449 = n7386 & ~n26503 ;
  assign n42451 = n42450 ^ n42449 ^ 1'b0 ;
  assign n42452 = n42451 ^ n40576 ^ n32232 ;
  assign n42453 = n22658 ^ n5783 ^ n696 ;
  assign n42454 = n29178 ^ n22200 ^ n1294 ;
  assign n42455 = n4638 ^ n3545 ^ 1'b0 ;
  assign n42456 = ( n42453 & ~n42454 ) | ( n42453 & n42455 ) | ( ~n42454 & n42455 ) ;
  assign n42457 = n28702 ^ n18046 ^ n7083 ;
  assign n42458 = n32997 & n33629 ;
  assign n42459 = n27751 & ~n40160 ;
  assign n42460 = n26804 | n36162 ;
  assign n42461 = n42460 ^ n21905 ^ 1'b0 ;
  assign n42462 = n29990 ^ n18505 ^ 1'b0 ;
  assign n42463 = ~n27009 & n42462 ;
  assign n42464 = n28398 & n42463 ;
  assign n42465 = n14854 & n16078 ;
  assign n42466 = n23457 & n39367 ;
  assign n42467 = n16414 | n34167 ;
  assign n42468 = n13117 & ~n25479 ;
  assign n42469 = ( ~n1573 & n19892 ) | ( ~n1573 & n42468 ) | ( n19892 & n42468 ) ;
  assign n42470 = n17261 | n19111 ;
  assign n42471 = n42470 ^ n30714 ^ 1'b0 ;
  assign n42472 = n13909 ^ n1419 ^ 1'b0 ;
  assign n42473 = n19446 | n42472 ;
  assign n42474 = n15232 ^ n6285 ^ 1'b0 ;
  assign n42475 = n42473 | n42474 ;
  assign n42476 = ~n14310 & n42116 ;
  assign n42477 = n25534 ^ n18962 ^ n9713 ;
  assign n42478 = n42477 ^ n31132 ^ n25764 ;
  assign n42479 = ( n946 & ~n26143 ) | ( n946 & n27209 ) | ( ~n26143 & n27209 ) ;
  assign n42480 = n42479 ^ n34652 ^ n10377 ;
  assign n42484 = n16310 ^ n12868 ^ n7314 ;
  assign n42485 = ( n5200 & n27515 ) | ( n5200 & ~n42484 ) | ( n27515 & ~n42484 ) ;
  assign n42481 = n17245 ^ n899 ^ 1'b0 ;
  assign n42482 = ( n36287 & n39794 ) | ( n36287 & n41703 ) | ( n39794 & n41703 ) ;
  assign n42483 = ( n18981 & n42481 ) | ( n18981 & n42482 ) | ( n42481 & n42482 ) ;
  assign n42486 = n42485 ^ n42483 ^ 1'b0 ;
  assign n42487 = n12352 ^ n7819 ^ 1'b0 ;
  assign n42489 = n8276 | n11605 ;
  assign n42488 = n7663 & n27381 ;
  assign n42490 = n42489 ^ n42488 ^ n40943 ;
  assign n42491 = ~n11682 & n16856 ;
  assign n42492 = n15405 | n42491 ;
  assign n42493 = n8349 & ~n42492 ;
  assign n42494 = ( ~n30600 & n42490 ) | ( ~n30600 & n42493 ) | ( n42490 & n42493 ) ;
  assign n42495 = n42487 & ~n42494 ;
  assign n42496 = ~n15134 & n42495 ;
  assign n42497 = n34252 ^ x109 ^ 1'b0 ;
  assign n42498 = n9417 & n42497 ;
  assign n42499 = ( n1354 & n24260 ) | ( n1354 & ~n28582 ) | ( n24260 & ~n28582 ) ;
  assign n42500 = ( n805 & n26979 ) | ( n805 & ~n42499 ) | ( n26979 & ~n42499 ) ;
  assign n42501 = x92 & ~n42500 ;
  assign n42502 = n366 & n42501 ;
  assign n42503 = ~n6864 & n16156 ;
  assign n42504 = n42503 ^ n31502 ^ 1'b0 ;
  assign n42505 = n6269 ^ n4336 ^ 1'b0 ;
  assign n42506 = ( ~n6883 & n10948 ) | ( ~n6883 & n16200 ) | ( n10948 & n16200 ) ;
  assign n42510 = ~n6017 & n6027 ;
  assign n42511 = n2444 & n42510 ;
  assign n42512 = ~n17490 & n42511 ;
  assign n42509 = n6320 & ~n21055 ;
  assign n42513 = n42512 ^ n42509 ^ 1'b0 ;
  assign n42507 = n1305 & ~n2788 ;
  assign n42508 = n32709 | n42507 ;
  assign n42514 = n42513 ^ n42508 ^ n41936 ;
  assign n42515 = n15913 | n25610 ;
  assign n42516 = n26389 | n42515 ;
  assign n42517 = n26681 & ~n42516 ;
  assign n42518 = n25358 ^ n2729 ^ n1016 ;
  assign n42519 = n42518 ^ n33019 ^ n30142 ;
  assign n42520 = n41234 ^ n31938 ^ 1'b0 ;
  assign n42521 = ( n704 & ~n17553 ) | ( n704 & n20337 ) | ( ~n17553 & n20337 ) ;
  assign n42522 = n6741 | n10701 ;
  assign n42523 = n5378 | n42522 ;
  assign n42524 = n17665 & ~n42523 ;
  assign n42525 = n6825 & n21817 ;
  assign n42526 = ( ~n21510 & n39205 ) | ( ~n21510 & n42525 ) | ( n39205 & n42525 ) ;
  assign n42528 = n36022 ^ n25698 ^ 1'b0 ;
  assign n42529 = n13077 & ~n42528 ;
  assign n42527 = n6516 & n9347 ;
  assign n42530 = n42529 ^ n42527 ^ n16962 ;
  assign n42532 = n17343 ^ n3529 ^ n1733 ;
  assign n42533 = n42532 ^ n14188 ^ n8475 ;
  assign n42531 = n13647 & ~n26134 ;
  assign n42534 = n42533 ^ n42531 ^ n40381 ;
  assign n42535 = n42534 ^ n580 ^ 1'b0 ;
  assign n42536 = ( n6183 & ~n6304 ) | ( n6183 & n23233 ) | ( ~n6304 & n23233 ) ;
  assign n42537 = ( n3827 & n11992 ) | ( n3827 & n12370 ) | ( n11992 & n12370 ) ;
  assign n42538 = n42537 ^ n26450 ^ n24672 ;
  assign n42539 = ~n23212 & n42538 ;
  assign n42540 = n42539 ^ n19920 ^ n13134 ;
  assign n42541 = n37520 ^ n26638 ^ 1'b0 ;
  assign n42542 = ~n15341 & n42541 ;
  assign n42543 = ~n30916 & n42542 ;
  assign n42544 = n3435 & ~n21650 ;
  assign n42545 = n42544 ^ n28220 ^ 1'b0 ;
  assign n42546 = n23325 & ~n26900 ;
  assign n42547 = ~n21410 & n42546 ;
  assign n42548 = n15597 ^ n8249 ^ n6443 ;
  assign n42549 = n23875 | n42548 ;
  assign n42550 = ~n42547 & n42549 ;
  assign n42551 = n9223 & ~n24785 ;
  assign n42552 = n42551 ^ n18136 ^ 1'b0 ;
  assign n42553 = n4056 & n12737 ;
  assign n42554 = ( n6701 & n35078 ) | ( n6701 & n42553 ) | ( n35078 & n42553 ) ;
  assign n42555 = ( n15454 & n42552 ) | ( n15454 & n42554 ) | ( n42552 & n42554 ) ;
  assign n42556 = ~n10205 & n42555 ;
  assign n42557 = n42556 ^ n23372 ^ n9220 ;
  assign n42558 = n7786 | n9195 ;
  assign n42559 = n42558 ^ n1822 ^ 1'b0 ;
  assign n42560 = ~n21814 & n42559 ;
  assign n42561 = ( n1358 & ~n27147 ) | ( n1358 & n42560 ) | ( ~n27147 & n42560 ) ;
  assign n42562 = n16938 & n17258 ;
  assign n42563 = n42562 ^ n35932 ^ 1'b0 ;
  assign n42564 = n3058 & ~n32952 ;
  assign n42565 = ~n2040 & n19189 ;
  assign n42566 = n41990 & n42565 ;
  assign n42567 = n19932 ^ n14188 ^ n8040 ;
  assign n42568 = n11990 ^ x206 ^ 1'b0 ;
  assign n42569 = ( n7334 & ~n21789 ) | ( n7334 & n42568 ) | ( ~n21789 & n42568 ) ;
  assign n42570 = n42569 ^ n1972 ^ 1'b0 ;
  assign n42571 = n27664 ^ n25353 ^ n21887 ;
  assign n42572 = n13344 ^ n4021 ^ 1'b0 ;
  assign n42573 = n9732 & n42572 ;
  assign n42574 = n22437 ^ n20584 ^ 1'b0 ;
  assign n42575 = ~n19920 & n42574 ;
  assign n42576 = ( n42571 & n42573 ) | ( n42571 & ~n42575 ) | ( n42573 & ~n42575 ) ;
  assign n42577 = ( ~n2310 & n23190 ) | ( ~n2310 & n36128 ) | ( n23190 & n36128 ) ;
  assign n42578 = n14622 ^ n4435 ^ n2244 ;
  assign n42579 = n42578 ^ n12416 ^ 1'b0 ;
  assign n42580 = ( n5810 & ~n18008 ) | ( n5810 & n26534 ) | ( ~n18008 & n26534 ) ;
  assign n42581 = n26689 & n42580 ;
  assign n42582 = n42581 ^ n16353 ^ 1'b0 ;
  assign n42583 = n9790 | n29923 ;
  assign n42584 = n15335 & ~n42583 ;
  assign n42585 = ~n6567 & n8821 ;
  assign n42586 = ~n3856 & n33376 ;
  assign n42587 = n42585 & n42586 ;
  assign n42588 = n16068 ^ n9108 ^ n1064 ;
  assign n42589 = ( n8828 & n15132 ) | ( n8828 & ~n42588 ) | ( n15132 & ~n42588 ) ;
  assign n42590 = n36574 & ~n42589 ;
  assign n42591 = n31402 ^ n2106 ^ 1'b0 ;
  assign n42592 = n38210 ^ n10914 ^ n7155 ;
  assign n42593 = ( ~n2913 & n7768 ) | ( ~n2913 & n18151 ) | ( n7768 & n18151 ) ;
  assign n42594 = ~n16905 & n42593 ;
  assign n42595 = n23966 & ~n24290 ;
  assign n42596 = n15112 | n31843 ;
  assign n42597 = ( n4381 & ~n5570 ) | ( n4381 & n15626 ) | ( ~n5570 & n15626 ) ;
  assign n42598 = n42597 ^ n7549 ^ 1'b0 ;
  assign n42599 = n17843 | n42598 ;
  assign n42600 = n5980 & n17814 ;
  assign n42601 = n42600 ^ n2391 ^ 1'b0 ;
  assign n42602 = n6164 & n23166 ;
  assign n42603 = n42602 ^ n4214 ^ 1'b0 ;
  assign n42604 = ( x80 & n30654 ) | ( x80 & n32326 ) | ( n30654 & n32326 ) ;
  assign n42605 = ~n11381 & n29061 ;
  assign n42606 = n42604 & n42605 ;
  assign n42607 = n42606 ^ n26185 ^ x175 ;
  assign n42608 = n42607 ^ n12484 ^ 1'b0 ;
  assign n42609 = ~n42603 & n42608 ;
  assign n42610 = ( n21199 & n31844 ) | ( n21199 & n42609 ) | ( n31844 & n42609 ) ;
  assign n42611 = n11122 ^ n5140 ^ 1'b0 ;
  assign n42612 = n42611 ^ n18588 ^ 1'b0 ;
  assign n42613 = n42612 ^ n37074 ^ n27181 ;
  assign n42614 = n40288 ^ n26155 ^ n14295 ;
  assign n42615 = n3323 & ~n13398 ;
  assign n42616 = ~n21557 & n42615 ;
  assign n42617 = ( n18644 & ~n29879 ) | ( n18644 & n42616 ) | ( ~n29879 & n42616 ) ;
  assign n42618 = ( n1839 & ~n14159 ) | ( n1839 & n42617 ) | ( ~n14159 & n42617 ) ;
  assign n42619 = n24320 ^ n20326 ^ n8887 ;
  assign n42620 = ( n8621 & n10367 ) | ( n8621 & n42619 ) | ( n10367 & n42619 ) ;
  assign n42621 = ( n12865 & n35688 ) | ( n12865 & ~n42620 ) | ( n35688 & ~n42620 ) ;
  assign n42622 = ( ~n3435 & n8228 ) | ( ~n3435 & n42621 ) | ( n8228 & n42621 ) ;
  assign n42623 = n892 & ~n37432 ;
  assign n42624 = n42623 ^ n41883 ^ 1'b0 ;
  assign n42625 = ( n1138 & n3895 ) | ( n1138 & ~n18715 ) | ( n3895 & ~n18715 ) ;
  assign n42626 = n42625 ^ n13606 ^ 1'b0 ;
  assign n42627 = n19494 & ~n42626 ;
  assign n42628 = n42627 ^ n19352 ^ 1'b0 ;
  assign n42629 = n40097 ^ n21687 ^ n9353 ;
  assign n42630 = n34900 ^ n24342 ^ n10828 ;
  assign n42631 = ~n8738 & n23382 ;
  assign n42632 = ( n2560 & n2749 ) | ( n2560 & ~n4283 ) | ( n2749 & ~n4283 ) ;
  assign n42633 = n42632 ^ n39414 ^ 1'b0 ;
  assign n42634 = n15742 & ~n42633 ;
  assign n42636 = n5501 | n37312 ;
  assign n42637 = n42636 ^ n34410 ^ 1'b0 ;
  assign n42638 = ( ~n20875 & n23392 ) | ( ~n20875 & n42637 ) | ( n23392 & n42637 ) ;
  assign n42635 = ~n2242 & n8501 ;
  assign n42639 = n42638 ^ n42635 ^ 1'b0 ;
  assign n42640 = n24965 | n30082 ;
  assign n42641 = n3011 | n42640 ;
  assign n42642 = ( n11003 & n13502 ) | ( n11003 & n42641 ) | ( n13502 & n42641 ) ;
  assign n42643 = ( n28994 & n40636 ) | ( n28994 & n42642 ) | ( n40636 & n42642 ) ;
  assign n42644 = n31073 ^ n24767 ^ n18101 ;
  assign n42645 = n41715 ^ n40695 ^ n14504 ;
  assign n42646 = ( ~n1257 & n8503 ) | ( ~n1257 & n10657 ) | ( n8503 & n10657 ) ;
  assign n42647 = n29101 ^ n27548 ^ n22842 ;
  assign n42648 = ( n16942 & ~n19191 ) | ( n16942 & n36212 ) | ( ~n19191 & n36212 ) ;
  assign n42649 = n42648 ^ n24766 ^ 1'b0 ;
  assign n42650 = n3223 | n4315 ;
  assign n42651 = n42650 ^ n8303 ^ 1'b0 ;
  assign n42652 = n24283 ^ n22022 ^ n6895 ;
  assign n42653 = ( n26640 & ~n26779 ) | ( n26640 & n42652 ) | ( ~n26779 & n42652 ) ;
  assign n42654 = ( ~x25 & n12141 ) | ( ~x25 & n38447 ) | ( n12141 & n38447 ) ;
  assign n42655 = n37018 ^ n13149 ^ x179 ;
  assign n42656 = ( n7766 & ~n16472 ) | ( n7766 & n42655 ) | ( ~n16472 & n42655 ) ;
  assign n42657 = n15174 | n22404 ;
  assign n42658 = n13257 & ~n34054 ;
  assign n42659 = n42657 & n42658 ;
  assign n42660 = n16808 & ~n35892 ;
  assign n42661 = n42660 ^ n17732 ^ 1'b0 ;
  assign n42662 = n13772 & n42661 ;
  assign n42663 = n42662 ^ n4886 ^ 1'b0 ;
  assign n42664 = n6643 | n36396 ;
  assign n42665 = n19501 | n42664 ;
  assign n42666 = ( ~n2635 & n18678 ) | ( ~n2635 & n31959 ) | ( n18678 & n31959 ) ;
  assign n42667 = ~n8408 & n36368 ;
  assign n42668 = n33795 | n42667 ;
  assign n42669 = n42666 & n42668 ;
  assign n42671 = n32435 ^ n9907 ^ n5325 ;
  assign n42672 = n20476 | n24385 ;
  assign n42673 = n42671 | n42672 ;
  assign n42674 = n42673 ^ n29510 ^ 1'b0 ;
  assign n42670 = n7184 & n36983 ;
  assign n42675 = n42674 ^ n42670 ^ n21693 ;
  assign n42676 = n20200 ^ n12801 ^ 1'b0 ;
  assign n42677 = n2696 & ~n42676 ;
  assign n42678 = ~n34589 & n39653 ;
  assign n42679 = ~n12682 & n42678 ;
  assign n42680 = n17211 & n23301 ;
  assign n42681 = n42680 ^ n20008 ^ 1'b0 ;
  assign n42682 = n42681 ^ n24939 ^ 1'b0 ;
  assign n42683 = ~n42679 & n42682 ;
  assign n42684 = n21561 & ~n36781 ;
  assign n42685 = n14583 & n42684 ;
  assign n42686 = n35406 ^ n23342 ^ n12384 ;
  assign n42687 = n25908 ^ n22135 ^ 1'b0 ;
  assign n42688 = n42687 ^ n5077 ^ n3922 ;
  assign n42689 = n4359 | n7265 ;
  assign n42690 = n17214 & n42689 ;
  assign n42691 = n13594 ^ n693 ^ 1'b0 ;
  assign n42692 = ~n38987 & n42691 ;
  assign n42693 = ~n21848 & n42692 ;
  assign n42694 = n5042 & ~n31436 ;
  assign n42695 = ~n11048 & n42694 ;
  assign n42696 = n13764 ^ n6195 ^ 1'b0 ;
  assign n42697 = ~n42695 & n42696 ;
  assign n42698 = n42697 ^ n26197 ^ 1'b0 ;
  assign n42699 = n416 & n42698 ;
  assign n42700 = n11463 & ~n24544 ;
  assign n42701 = n22853 & n42700 ;
  assign n42702 = ( n13208 & n27547 ) | ( n13208 & n40450 ) | ( n27547 & n40450 ) ;
  assign n42703 = n2801 | n35033 ;
  assign n42706 = n1988 ^ n549 ^ 1'b0 ;
  assign n42704 = ( n14091 & n19565 ) | ( n14091 & n34294 ) | ( n19565 & n34294 ) ;
  assign n42705 = n36030 & n42704 ;
  assign n42707 = n42706 ^ n42705 ^ 1'b0 ;
  assign n42708 = ~n5353 & n32102 ;
  assign n42709 = n38215 & n42708 ;
  assign n42710 = n9044 & ~n42709 ;
  assign n42711 = n7306 & n42710 ;
  assign n42712 = n17036 ^ n10040 ^ 1'b0 ;
  assign n42713 = n42711 | n42712 ;
  assign n42714 = ~n8222 & n16117 ;
  assign n42715 = n19036 ^ n3606 ^ 1'b0 ;
  assign n42716 = n4042 ^ n3143 ^ 1'b0 ;
  assign n42717 = n1164 & n42716 ;
  assign n42718 = n42717 ^ n38712 ^ 1'b0 ;
  assign n42719 = ( n17564 & n19670 ) | ( n17564 & ~n23411 ) | ( n19670 & ~n23411 ) ;
  assign n42720 = ( ~n40161 & n42718 ) | ( ~n40161 & n42719 ) | ( n42718 & n42719 ) ;
  assign n42721 = n13469 | n15774 ;
  assign n42722 = n42721 ^ n16337 ^ 1'b0 ;
  assign n42723 = n10173 & n42722 ;
  assign n42724 = n6190 & ~n19611 ;
  assign n42725 = n42724 ^ n25246 ^ 1'b0 ;
  assign n42726 = n42725 ^ n20008 ^ 1'b0 ;
  assign n42727 = n32635 ^ n26499 ^ n5394 ;
  assign n42728 = n18548 ^ n12037 ^ 1'b0 ;
  assign n42729 = ~n42727 & n42728 ;
  assign n42730 = n23212 ^ n4921 ^ 1'b0 ;
  assign n42731 = ( n16785 & n36218 ) | ( n16785 & ~n42730 ) | ( n36218 & ~n42730 ) ;
  assign n42732 = n40790 ^ n10288 ^ n8724 ;
  assign n42733 = n28136 ^ n20685 ^ n14952 ;
  assign n42734 = n40063 ^ n5417 ^ 1'b0 ;
  assign n42735 = ( n41182 & ~n42733 ) | ( n41182 & n42734 ) | ( ~n42733 & n42734 ) ;
  assign n42736 = n17120 ^ n10653 ^ 1'b0 ;
  assign n42737 = n798 | n42736 ;
  assign n42738 = n36538 ^ n32734 ^ n2711 ;
  assign n42739 = n14552 ^ n8123 ^ 1'b0 ;
  assign n42740 = n20854 | n42739 ;
  assign n42741 = n644 & n25569 ;
  assign n42742 = ~n11814 & n42741 ;
  assign n42743 = n42742 ^ n28614 ^ 1'b0 ;
  assign n42745 = n17117 ^ n11980 ^ 1'b0 ;
  assign n42744 = n12014 | n21945 ;
  assign n42746 = n42745 ^ n42744 ^ 1'b0 ;
  assign n42747 = n11638 ^ n5299 ^ 1'b0 ;
  assign n42748 = ( n15883 & n27394 ) | ( n15883 & n36656 ) | ( n27394 & n36656 ) ;
  assign n42749 = n27471 ^ n14447 ^ 1'b0 ;
  assign n42750 = n42749 ^ n37824 ^ n29023 ;
  assign n42751 = n4906 & ~n10773 ;
  assign n42752 = n42751 ^ n33431 ^ n12808 ;
  assign n42753 = ( n6248 & n28484 ) | ( n6248 & ~n35058 ) | ( n28484 & ~n35058 ) ;
  assign n42754 = ( ~n13712 & n42752 ) | ( ~n13712 & n42753 ) | ( n42752 & n42753 ) ;
  assign n42755 = n1016 & ~n15641 ;
  assign n42756 = n42755 ^ n14276 ^ 1'b0 ;
  assign n42758 = n8508 ^ n8440 ^ 1'b0 ;
  assign n42759 = n11386 & n42758 ;
  assign n42757 = n11195 & ~n29041 ;
  assign n42760 = n42759 ^ n42757 ^ 1'b0 ;
  assign n42761 = n12429 | n31243 ;
  assign n42762 = n16855 | n42761 ;
  assign n42763 = n7504 ^ n4700 ^ 1'b0 ;
  assign n42764 = n42762 & n42763 ;
  assign n42765 = ( n3781 & n6138 ) | ( n3781 & ~n35309 ) | ( n6138 & ~n35309 ) ;
  assign n42766 = ( n15519 & n34589 ) | ( n15519 & n42765 ) | ( n34589 & n42765 ) ;
  assign n42769 = ( n5799 & n14562 ) | ( n5799 & ~n28284 ) | ( n14562 & ~n28284 ) ;
  assign n42770 = n22742 & ~n42769 ;
  assign n42767 = n18000 ^ n9297 ^ n1689 ;
  assign n42768 = ( n744 & n16980 ) | ( n744 & n42767 ) | ( n16980 & n42767 ) ;
  assign n42771 = n42770 ^ n42768 ^ 1'b0 ;
  assign n42772 = n397 & n25933 ;
  assign n42773 = ( ~n11538 & n13988 ) | ( ~n11538 & n26844 ) | ( n13988 & n26844 ) ;
  assign n42774 = n37838 & ~n42773 ;
  assign n42775 = n35922 ^ n13047 ^ n3587 ;
  assign n42776 = n42775 ^ n37476 ^ n35560 ;
  assign n42777 = ( n12504 & n34567 ) | ( n12504 & ~n42776 ) | ( n34567 & ~n42776 ) ;
  assign n42778 = n4456 & ~n6966 ;
  assign n42779 = n32796 ^ n4009 ^ 1'b0 ;
  assign n42780 = n41363 & ~n42779 ;
  assign n42781 = ( n6090 & n19791 ) | ( n6090 & ~n27437 ) | ( n19791 & ~n27437 ) ;
  assign n42782 = n42781 ^ n17468 ^ n536 ;
  assign n42783 = n42782 ^ n2544 ^ 1'b0 ;
  assign n42784 = ( n6033 & ~n18121 ) | ( n6033 & n42783 ) | ( ~n18121 & n42783 ) ;
  assign n42785 = n42780 & ~n42784 ;
  assign n42786 = n42785 ^ n10865 ^ 1'b0 ;
  assign n42788 = n1044 & n9944 ;
  assign n42789 = n16029 & n42788 ;
  assign n42790 = ( n7746 & n20031 ) | ( n7746 & n42789 ) | ( n20031 & n42789 ) ;
  assign n42791 = ( ~n22776 & n34312 ) | ( ~n22776 & n42790 ) | ( n34312 & n42790 ) ;
  assign n42787 = n24289 ^ n19871 ^ n14476 ;
  assign n42792 = n42791 ^ n42787 ^ n16211 ;
  assign n42793 = ( n12962 & ~n28398 ) | ( n12962 & n42792 ) | ( ~n28398 & n42792 ) ;
  assign n42794 = n8110 & n42793 ;
  assign n42795 = n34965 & n42794 ;
  assign n42796 = n39979 ^ n21072 ^ n317 ;
  assign n42804 = ~n344 & n41814 ;
  assign n42799 = ~n922 & n3603 ;
  assign n42800 = n42799 ^ n3600 ^ 1'b0 ;
  assign n42801 = n10463 & ~n42800 ;
  assign n42797 = n29774 ^ n22574 ^ n19280 ;
  assign n42798 = n21798 & n42797 ;
  assign n42802 = n42801 ^ n42798 ^ 1'b0 ;
  assign n42803 = n17672 & n42802 ;
  assign n42805 = n42804 ^ n42803 ^ n32852 ;
  assign n42806 = n27345 ^ n7884 ^ n5276 ;
  assign n42807 = n7970 | n32898 ;
  assign n42808 = n42807 ^ n3123 ^ 1'b0 ;
  assign n42809 = n42808 ^ n2927 ^ 1'b0 ;
  assign n42810 = ~n27040 & n42809 ;
  assign n42811 = n42810 ^ n2265 ^ 1'b0 ;
  assign n42812 = n4173 | n10097 ;
  assign n42813 = n4988 | n42812 ;
  assign n42814 = n42813 ^ n26295 ^ 1'b0 ;
  assign n42815 = ( ~n1351 & n40392 ) | ( ~n1351 & n42814 ) | ( n40392 & n42814 ) ;
  assign n42816 = ~n21650 & n26455 ;
  assign n42817 = n1408 & n42816 ;
  assign n42818 = n13646 | n33883 ;
  assign n42819 = n25522 | n42818 ;
  assign n42820 = n18781 & ~n18813 ;
  assign n42821 = n42820 ^ n30456 ^ 1'b0 ;
  assign n42822 = x252 & ~n22451 ;
  assign n42823 = n42822 ^ n8008 ^ n3123 ;
  assign n42824 = ( ~n13879 & n27762 ) | ( ~n13879 & n42823 ) | ( n27762 & n42823 ) ;
  assign n42825 = n42821 & ~n42824 ;
  assign n42832 = n40372 ^ n3780 ^ n1294 ;
  assign n42831 = ( n652 & n4291 ) | ( n652 & ~n9746 ) | ( n4291 & ~n9746 ) ;
  assign n42826 = n22805 ^ n16647 ^ 1'b0 ;
  assign n42827 = n42826 ^ n8219 ^ n1512 ;
  assign n42828 = n42827 ^ n8428 ^ 1'b0 ;
  assign n42829 = n42828 ^ n34882 ^ n916 ;
  assign n42830 = ( n4129 & n27754 ) | ( n4129 & ~n42829 ) | ( n27754 & ~n42829 ) ;
  assign n42833 = n42832 ^ n42831 ^ n42830 ;
  assign n42834 = n11393 & n19155 ;
  assign n42835 = n42214 ^ n29613 ^ n8212 ;
  assign n42836 = n5832 & ~n10362 ;
  assign n42837 = n42836 ^ n13872 ^ 1'b0 ;
  assign n42838 = n4615 | n26077 ;
  assign n42839 = ~n19328 & n20423 ;
  assign n42840 = ~n42838 & n42839 ;
  assign n42841 = n33589 ^ n20741 ^ 1'b0 ;
  assign n42842 = n29996 | n42841 ;
  assign n42843 = n19644 ^ n8886 ^ x230 ;
  assign n42844 = n42843 ^ n19611 ^ n13194 ;
  assign n42845 = n40461 & n42844 ;
  assign n42846 = n42842 & n42845 ;
  assign n42847 = ~n6887 & n8862 ;
  assign n42848 = ~n8179 & n42847 ;
  assign n42853 = n21298 & ~n34310 ;
  assign n42854 = n42853 ^ n30290 ^ 1'b0 ;
  assign n42855 = n42854 ^ n13747 ^ n11435 ;
  assign n42856 = ( n32501 & ~n38232 ) | ( n32501 & n42855 ) | ( ~n38232 & n42855 ) ;
  assign n42857 = ~n10104 & n42856 ;
  assign n42858 = n14596 & n42857 ;
  assign n42849 = ~n7790 & n33109 ;
  assign n42850 = n42849 ^ n1644 ^ 1'b0 ;
  assign n42851 = n30579 & n42850 ;
  assign n42852 = n42851 ^ n33653 ^ 1'b0 ;
  assign n42859 = n42858 ^ n42852 ^ 1'b0 ;
  assign n42860 = ~n42848 & n42859 ;
  assign n42861 = ( n2350 & n22652 ) | ( n2350 & ~n37353 ) | ( n22652 & ~n37353 ) ;
  assign n42862 = ~n2206 & n7014 ;
  assign n42863 = n32392 & n34193 ;
  assign n42864 = ~x207 & x221 ;
  assign n42865 = n42864 ^ n37100 ^ n10784 ;
  assign n42866 = ( n8063 & ~n23950 ) | ( n8063 & n30545 ) | ( ~n23950 & n30545 ) ;
  assign n42868 = n12243 ^ n8965 ^ n1961 ;
  assign n42867 = n14178 & ~n21890 ;
  assign n42869 = n42868 ^ n42867 ^ 1'b0 ;
  assign n42870 = n42866 & n42869 ;
  assign n42871 = n35988 ^ n5293 ^ 1'b0 ;
  assign n42887 = ( n6242 & n6822 ) | ( n6242 & n7578 ) | ( n6822 & n7578 ) ;
  assign n42888 = ( n18995 & n32878 ) | ( n18995 & ~n42887 ) | ( n32878 & ~n42887 ) ;
  assign n42872 = ( n1511 & ~n2701 ) | ( n1511 & n18380 ) | ( ~n2701 & n18380 ) ;
  assign n42873 = n40704 ^ n24428 ^ n16337 ;
  assign n42874 = n19305 ^ n17843 ^ n5060 ;
  assign n42875 = n13465 & n32475 ;
  assign n42876 = ~n12850 & n42875 ;
  assign n42877 = ( ~n37662 & n42874 ) | ( ~n37662 & n42876 ) | ( n42874 & n42876 ) ;
  assign n42878 = n42877 ^ n5890 ^ 1'b0 ;
  assign n42879 = ~n11732 & n40363 ;
  assign n42880 = n13430 ^ n9452 ^ n7618 ;
  assign n42881 = ( n4120 & ~n13082 ) | ( n4120 & n42880 ) | ( ~n13082 & n42880 ) ;
  assign n42882 = n42881 ^ n4697 ^ 1'b0 ;
  assign n42883 = n42879 | n42882 ;
  assign n42884 = n15426 & ~n42883 ;
  assign n42885 = n42878 & n42884 ;
  assign n42886 = ( ~n42872 & n42873 ) | ( ~n42872 & n42885 ) | ( n42873 & n42885 ) ;
  assign n42889 = n42888 ^ n42886 ^ 1'b0 ;
  assign n42890 = n23598 ^ n12008 ^ n4966 ;
  assign n42891 = n3743 & n4682 ;
  assign n42892 = n42891 ^ n4435 ^ 1'b0 ;
  assign n42893 = n42892 ^ n10367 ^ 1'b0 ;
  assign n42894 = n3107 & ~n36029 ;
  assign n42895 = n42894 ^ n2880 ^ 1'b0 ;
  assign n42896 = ( n5567 & ~n21258 ) | ( n5567 & n36362 ) | ( ~n21258 & n36362 ) ;
  assign n42898 = n17189 ^ n1769 ^ 1'b0 ;
  assign n42899 = n8877 & ~n42898 ;
  assign n42897 = n28173 & ~n30982 ;
  assign n42900 = n42899 ^ n42897 ^ n42312 ;
  assign n42901 = ~n21087 & n22672 ;
  assign n42902 = n16029 & ~n23078 ;
  assign n42903 = n39091 ^ n14868 ^ 1'b0 ;
  assign n42904 = n16578 & ~n42903 ;
  assign n42905 = n42902 & n42904 ;
  assign n42906 = n38039 ^ n10687 ^ 1'b0 ;
  assign n42907 = n30039 ^ n10035 ^ n4783 ;
  assign n42908 = n26262 | n42907 ;
  assign n42909 = n42908 ^ n14067 ^ 1'b0 ;
  assign n42910 = n42909 ^ n20056 ^ 1'b0 ;
  assign n42911 = n24975 | n42910 ;
  assign n42912 = n24251 | n42911 ;
  assign n42913 = n15012 & ~n20824 ;
  assign n42914 = n13164 & n42913 ;
  assign n42915 = n16969 & ~n19622 ;
  assign n42916 = n42914 & n42915 ;
  assign n42917 = n42916 ^ n12010 ^ 1'b0 ;
  assign n42918 = n40821 ^ n16238 ^ 1'b0 ;
  assign n42919 = x71 & n31417 ;
  assign n42920 = n22128 & n42919 ;
  assign n42921 = n42920 ^ n18176 ^ 1'b0 ;
  assign n42922 = n37798 ^ n3499 ^ n1101 ;
  assign n42923 = n19164 ^ n1491 ^ 1'b0 ;
  assign n42924 = n16113 & ~n42923 ;
  assign n42927 = n8526 & ~n18073 ;
  assign n42925 = ( n3525 & n4004 ) | ( n3525 & n23875 ) | ( n4004 & n23875 ) ;
  assign n42926 = n42925 ^ n8549 ^ n6558 ;
  assign n42928 = n42927 ^ n42926 ^ n7660 ;
  assign n42930 = ( n10249 & n14767 ) | ( n10249 & n26264 ) | ( n14767 & n26264 ) ;
  assign n42931 = n15465 | n42930 ;
  assign n42929 = n9264 ^ n8755 ^ 1'b0 ;
  assign n42932 = n42931 ^ n42929 ^ n38515 ;
  assign n42933 = ( n5386 & n21913 ) | ( n5386 & n42932 ) | ( n21913 & n42932 ) ;
  assign n42934 = n20663 & n25542 ;
  assign n42935 = ( n29441 & n32617 ) | ( n29441 & n33621 ) | ( n32617 & n33621 ) ;
  assign n42936 = n2387 & ~n6989 ;
  assign n42937 = n42936 ^ n39342 ^ n21759 ;
  assign n42938 = n12250 | n42937 ;
  assign n42939 = n2655 | n4560 ;
  assign n42940 = n42939 ^ n5305 ^ 1'b0 ;
  assign n42941 = n37399 & ~n42940 ;
  assign n42942 = n16857 ^ n9761 ^ n4478 ;
  assign n42943 = ~n41134 & n42942 ;
  assign n42944 = n19425 & n32939 ;
  assign n42945 = n27610 ^ n23557 ^ n1526 ;
  assign n42946 = n38099 ^ n28993 ^ n17695 ;
  assign n42947 = n3992 | n20507 ;
  assign n42948 = n41652 | n42947 ;
  assign n42949 = ( n12301 & n33210 ) | ( n12301 & n42948 ) | ( n33210 & n42948 ) ;
  assign n42950 = n2426 & n17516 ;
  assign n42951 = n10469 ^ n3021 ^ 1'b0 ;
  assign n42952 = n39936 ^ n36988 ^ n22866 ;
  assign n42953 = n28728 ^ n22632 ^ 1'b0 ;
  assign n42956 = ( ~n3380 & n11275 ) | ( ~n3380 & n15831 ) | ( n11275 & n15831 ) ;
  assign n42954 = n5980 & ~n12717 ;
  assign n42955 = n42954 ^ n9500 ^ 1'b0 ;
  assign n42957 = n42956 ^ n42955 ^ 1'b0 ;
  assign n42959 = n6674 | n12549 ;
  assign n42960 = n42959 ^ n13850 ^ 1'b0 ;
  assign n42961 = n42960 ^ n23946 ^ n1243 ;
  assign n42958 = n37999 & n40046 ;
  assign n42962 = n42961 ^ n42958 ^ 1'b0 ;
  assign n42963 = ~n8398 & n23408 ;
  assign n42964 = n42963 ^ n25492 ^ 1'b0 ;
  assign n42965 = n42964 ^ n1112 ^ 1'b0 ;
  assign n42966 = n29813 & ~n31857 ;
  assign n42967 = ( n2664 & n12277 ) | ( n2664 & n42966 ) | ( n12277 & n42966 ) ;
  assign n42968 = n19463 ^ n2402 ^ 1'b0 ;
  assign n42969 = n9043 & ~n18599 ;
  assign n42970 = n20975 ^ n16790 ^ 1'b0 ;
  assign n42971 = ( n10517 & n26174 ) | ( n10517 & n32498 ) | ( n26174 & n32498 ) ;
  assign n42972 = n36988 ^ n15323 ^ 1'b0 ;
  assign n42973 = ( ~n3633 & n4193 ) | ( ~n3633 & n42972 ) | ( n4193 & n42972 ) ;
  assign n42974 = n42973 ^ n26935 ^ n24578 ;
  assign n42975 = ( n20430 & n21273 ) | ( n20430 & n26227 ) | ( n21273 & n26227 ) ;
  assign n42976 = n35278 ^ n7827 ^ x144 ;
  assign n42977 = ( ~n6230 & n8768 ) | ( ~n6230 & n33176 ) | ( n8768 & n33176 ) ;
  assign n42978 = n42977 ^ n6760 ^ 1'b0 ;
  assign n42979 = n33884 ^ n3544 ^ 1'b0 ;
  assign n42980 = n42979 ^ n19014 ^ n6077 ;
  assign n42981 = ( n19244 & ~n25411 ) | ( n19244 & n36413 ) | ( ~n25411 & n36413 ) ;
  assign n42982 = n42981 ^ n20766 ^ 1'b0 ;
  assign n42990 = ( n8077 & ~n19638 ) | ( n8077 & n26687 ) | ( ~n19638 & n26687 ) ;
  assign n42991 = ( x139 & n30813 ) | ( x139 & n42990 ) | ( n30813 & n42990 ) ;
  assign n42983 = n2490 ^ x106 ^ 1'b0 ;
  assign n42984 = n42983 ^ n15084 ^ n11312 ;
  assign n42985 = n293 | n28477 ;
  assign n42986 = n7929 | n29143 ;
  assign n42987 = n42985 | n42986 ;
  assign n42988 = n42987 ^ n15500 ^ n2107 ;
  assign n42989 = ~n42984 & n42988 ;
  assign n42992 = n42991 ^ n42989 ^ 1'b0 ;
  assign n42993 = ( n4910 & ~n10285 ) | ( n4910 & n37615 ) | ( ~n10285 & n37615 ) ;
  assign n42994 = n7880 & ~n42993 ;
  assign n42995 = n42994 ^ n25496 ^ 1'b0 ;
  assign n42996 = ( n23202 & n30057 ) | ( n23202 & n42995 ) | ( n30057 & n42995 ) ;
  assign n42997 = n13030 & n42996 ;
  assign n42998 = n42997 ^ n22938 ^ 1'b0 ;
  assign n42999 = n1938 & ~n32771 ;
  assign n43000 = n42999 ^ n2869 ^ 1'b0 ;
  assign n43001 = n24929 ^ n10286 ^ 1'b0 ;
  assign n43002 = n43000 & n43001 ;
  assign n43003 = ~n16434 & n43002 ;
  assign n43004 = n42998 & n43003 ;
  assign n43007 = n5452 ^ n4939 ^ 1'b0 ;
  assign n43008 = ( ~n3531 & n34333 ) | ( ~n3531 & n43007 ) | ( n34333 & n43007 ) ;
  assign n43005 = n6941 & n15434 ;
  assign n43006 = n21997 & n43005 ;
  assign n43009 = n43008 ^ n43006 ^ n24018 ;
  assign n43010 = ~n3543 & n43009 ;
  assign n43011 = ( n3953 & ~n19472 ) | ( n3953 & n36910 ) | ( ~n19472 & n36910 ) ;
  assign n43012 = n12763 | n29851 ;
  assign n43013 = ~n43011 & n43012 ;
  assign n43014 = ( ~n4128 & n36311 ) | ( ~n4128 & n43013 ) | ( n36311 & n43013 ) ;
  assign n43015 = n5918 ^ n2014 ^ 1'b0 ;
  assign n43016 = ~n6148 & n39707 ;
  assign n43017 = n2790 | n18763 ;
  assign n43018 = n38552 | n43017 ;
  assign n43019 = ~n732 & n34878 ;
  assign n43020 = ~n29528 & n43019 ;
  assign n43021 = ( ~n2285 & n2609 ) | ( ~n2285 & n33999 ) | ( n2609 & n33999 ) ;
  assign n43022 = n7051 | n43021 ;
  assign n43023 = n11438 & ~n43022 ;
  assign n43024 = n43023 ^ n9374 ^ 1'b0 ;
  assign n43025 = x42 & ~n43024 ;
  assign n43027 = n29942 ^ n23472 ^ n8100 ;
  assign n43026 = ~n15790 & n24642 ;
  assign n43028 = n43027 ^ n43026 ^ 1'b0 ;
  assign n43029 = n32898 ^ n13031 ^ n7672 ;
  assign n43030 = ( n5355 & ~n14767 ) | ( n5355 & n43029 ) | ( ~n14767 & n43029 ) ;
  assign n43031 = ( n13290 & n26920 ) | ( n13290 & n43030 ) | ( n26920 & n43030 ) ;
  assign n43032 = ( ~n5076 & n30356 ) | ( ~n5076 & n43031 ) | ( n30356 & n43031 ) ;
  assign n43033 = ( n3397 & n8828 ) | ( n3397 & n16482 ) | ( n8828 & n16482 ) ;
  assign n43034 = ~n816 & n37155 ;
  assign n43035 = n41589 ^ n41252 ^ n33625 ;
  assign n43043 = n23304 ^ n18456 ^ n1921 ;
  assign n43036 = n13742 ^ n13198 ^ n2528 ;
  assign n43037 = n22769 ^ n12324 ^ n3129 ;
  assign n43038 = ( n13574 & n43036 ) | ( n13574 & n43037 ) | ( n43036 & n43037 ) ;
  assign n43039 = n23967 ^ n16856 ^ n1146 ;
  assign n43040 = ( n17490 & n38622 ) | ( n17490 & n43039 ) | ( n38622 & n43039 ) ;
  assign n43041 = ~n40746 & n43040 ;
  assign n43042 = n43038 & n43041 ;
  assign n43044 = n43043 ^ n43042 ^ n14207 ;
  assign n43045 = ~n13319 & n19765 ;
  assign n43046 = ( n2066 & ~n2987 ) | ( n2066 & n6037 ) | ( ~n2987 & n6037 ) ;
  assign n43047 = ( n9820 & n10998 ) | ( n9820 & ~n43046 ) | ( n10998 & ~n43046 ) ;
  assign n43048 = ( ~n13227 & n34274 ) | ( ~n13227 & n43047 ) | ( n34274 & n43047 ) ;
  assign n43049 = n43045 | n43048 ;
  assign n43050 = n3632 & ~n43049 ;
  assign n43051 = ( n2051 & ~n27187 ) | ( n2051 & n36606 ) | ( ~n27187 & n36606 ) ;
  assign n43052 = n35165 | n43051 ;
  assign n43053 = n31695 | n43052 ;
  assign n43054 = n10004 & ~n18619 ;
  assign n43055 = n14734 & n43054 ;
  assign n43056 = ( n11422 & ~n15284 ) | ( n11422 & n41959 ) | ( ~n15284 & n41959 ) ;
  assign n43057 = n43056 ^ n17357 ^ 1'b0 ;
  assign n43058 = n20392 & ~n43057 ;
  assign n43059 = ( n11046 & n17765 ) | ( n11046 & n43058 ) | ( n17765 & n43058 ) ;
  assign n43060 = ( n824 & n20267 ) | ( n824 & ~n26486 ) | ( n20267 & ~n26486 ) ;
  assign n43061 = n43060 ^ n9848 ^ n433 ;
  assign n43062 = n43061 ^ n32919 ^ n5641 ;
  assign n43063 = n37961 ^ n21736 ^ n18007 ;
  assign n43064 = ~n759 & n43063 ;
  assign n43065 = ( n4199 & n12659 ) | ( n4199 & n17240 ) | ( n12659 & n17240 ) ;
  assign n43066 = ( ~n7471 & n14109 ) | ( ~n7471 & n43065 ) | ( n14109 & n43065 ) ;
  assign n43067 = n43066 ^ n29900 ^ n19888 ;
  assign n43068 = n3124 & ~n5800 ;
  assign n43069 = n42309 ^ x89 ^ 1'b0 ;
  assign n43074 = ~n3241 & n21720 ;
  assign n43075 = n39713 & n43074 ;
  assign n43076 = n4772 & n43075 ;
  assign n43077 = n14320 & ~n43076 ;
  assign n43078 = n18611 & n43077 ;
  assign n43073 = n23545 ^ n22853 ^ 1'b0 ;
  assign n43079 = n43078 ^ n43073 ^ n36385 ;
  assign n43070 = ~n13138 & n13394 ;
  assign n43071 = ( n4068 & n25557 ) | ( n4068 & n43070 ) | ( n25557 & n43070 ) ;
  assign n43072 = n1721 | n43071 ;
  assign n43080 = n43079 ^ n43072 ^ 1'b0 ;
  assign n43081 = n758 & n1171 ;
  assign n43082 = n43081 ^ n8756 ^ 1'b0 ;
  assign n43083 = n17136 & ~n29003 ;
  assign n43084 = ~n43082 & n43083 ;
  assign n43085 = n43084 ^ n27748 ^ 1'b0 ;
  assign n43086 = x144 & ~n43085 ;
  assign n43088 = n10585 | n22366 ;
  assign n43089 = n43088 ^ n14214 ^ n11509 ;
  assign n43087 = n23188 ^ n3927 ^ 1'b0 ;
  assign n43090 = n43089 ^ n43087 ^ n38248 ;
  assign n43091 = n20747 & ~n34744 ;
  assign n43092 = n18376 ^ n13792 ^ 1'b0 ;
  assign n43093 = n43091 | n43092 ;
  assign n43094 = n43093 ^ n35609 ^ n24597 ;
  assign n43095 = n21617 | n41746 ;
  assign n43096 = n25356 ^ n5163 ^ n3950 ;
  assign n43097 = n43096 ^ n14875 ^ 1'b0 ;
  assign n43098 = n5175 | n43097 ;
  assign n43099 = n41250 & ~n43098 ;
  assign n43100 = n20980 ^ n13058 ^ 1'b0 ;
  assign n43101 = n27976 & n43100 ;
  assign n43102 = ( n4931 & n20036 ) | ( n4931 & ~n20368 ) | ( n20036 & ~n20368 ) ;
  assign n43103 = n30370 ^ n2495 ^ 1'b0 ;
  assign n43104 = n43102 & ~n43103 ;
  assign n43105 = ( n380 & n658 ) | ( n380 & ~n6588 ) | ( n658 & ~n6588 ) ;
  assign n43106 = ~n2700 & n40281 ;
  assign n43107 = ( n2174 & ~n6662 ) | ( n2174 & n10078 ) | ( ~n6662 & n10078 ) ;
  assign n43108 = n39295 ^ n6560 ^ 1'b0 ;
  assign n43109 = n43108 ^ n27504 ^ n6948 ;
  assign n43110 = n17056 | n20778 ;
  assign n43111 = n27419 | n43110 ;
  assign n43112 = n23745 ^ n1506 ^ 1'b0 ;
  assign n43113 = n39716 & ~n43112 ;
  assign n43114 = ( ~n12750 & n34920 ) | ( ~n12750 & n43113 ) | ( n34920 & n43113 ) ;
  assign n43115 = ( n4325 & ~n24909 ) | ( n4325 & n25534 ) | ( ~n24909 & n25534 ) ;
  assign n43116 = ( ~n9204 & n16506 ) | ( ~n9204 & n31734 ) | ( n16506 & n31734 ) ;
  assign n43117 = n43116 ^ n19413 ^ n9064 ;
  assign n43118 = n1162 & n35302 ;
  assign n43119 = n43118 ^ n862 ^ 1'b0 ;
  assign n43120 = n6562 & ~n9794 ;
  assign n43121 = n43120 ^ n32683 ^ 1'b0 ;
  assign n43122 = n27676 & n43121 ;
  assign n43128 = n36049 ^ n25253 ^ n6755 ;
  assign n43123 = n12614 | n14758 ;
  assign n43124 = n22370 | n43123 ;
  assign n43125 = n43124 ^ n15407 ^ n3209 ;
  assign n43126 = n43125 ^ n4897 ^ 1'b0 ;
  assign n43127 = n41082 & n43126 ;
  assign n43129 = n43128 ^ n43127 ^ 1'b0 ;
  assign n43130 = n6168 | n26935 ;
  assign n43134 = n700 & n23486 ;
  assign n43131 = n1941 & ~n17482 ;
  assign n43132 = ~x100 & n43131 ;
  assign n43133 = n43132 ^ n30543 ^ n1630 ;
  assign n43135 = n43134 ^ n43133 ^ 1'b0 ;
  assign n43136 = n2811 | n31172 ;
  assign n43137 = n27074 | n38494 ;
  assign n43138 = n43137 ^ n22697 ^ n8531 ;
  assign n43139 = n32952 ^ n18687 ^ n16255 ;
  assign n43140 = n43139 ^ n13009 ^ 1'b0 ;
  assign n43141 = n19992 & ~n41023 ;
  assign n43142 = n29604 ^ n16795 ^ n6092 ;
  assign n43143 = n4750 | n16481 ;
  assign n43144 = n43143 ^ n20262 ^ 1'b0 ;
  assign n43145 = n17102 ^ x110 ^ 1'b0 ;
  assign n43146 = n43144 & n43145 ;
  assign n43147 = n43146 ^ n2070 ^ 1'b0 ;
  assign n43148 = n3959 & ~n43147 ;
  assign n43149 = ~n17497 & n43148 ;
  assign n43150 = ~n4231 & n29103 ;
  assign n43151 = n43150 ^ n12803 ^ 1'b0 ;
  assign n43152 = n40524 ^ n20057 ^ 1'b0 ;
  assign n43153 = n24157 & n43152 ;
  assign n43154 = ( ~n11434 & n25200 ) | ( ~n11434 & n43153 ) | ( n25200 & n43153 ) ;
  assign n43155 = ( ~n5888 & n43151 ) | ( ~n5888 & n43154 ) | ( n43151 & n43154 ) ;
  assign n43156 = n43155 ^ n36638 ^ n16798 ;
  assign n43157 = n16534 & ~n33380 ;
  assign n43158 = n43157 ^ n10222 ^ 1'b0 ;
  assign n43159 = n22237 | n43158 ;
  assign n43160 = n37444 & ~n43159 ;
  assign n43161 = ( n8103 & n18403 ) | ( n8103 & ~n28390 ) | ( n18403 & ~n28390 ) ;
  assign n43162 = n25797 ^ n5828 ^ 1'b0 ;
  assign n43163 = n11216 & ~n43162 ;
  assign n43164 = ( n4017 & n29719 ) | ( n4017 & n41168 ) | ( n29719 & n41168 ) ;
  assign n43165 = n43164 ^ n30837 ^ n4068 ;
  assign n43166 = ( n20873 & n43163 ) | ( n20873 & ~n43165 ) | ( n43163 & ~n43165 ) ;
  assign n43167 = ( n1859 & n10979 ) | ( n1859 & ~n12797 ) | ( n10979 & ~n12797 ) ;
  assign n43168 = n4494 ^ n703 ^ 1'b0 ;
  assign n43169 = ~n3300 & n43168 ;
  assign n43175 = n25479 | n34420 ;
  assign n43176 = n10939 | n43175 ;
  assign n43170 = n41890 ^ n32405 ^ n8330 ;
  assign n43171 = ~n11884 & n38211 ;
  assign n43172 = n43171 ^ n9401 ^ 1'b0 ;
  assign n43173 = n43172 ^ n16373 ^ 1'b0 ;
  assign n43174 = n43170 & ~n43173 ;
  assign n43177 = n43176 ^ n43174 ^ n1107 ;
  assign n43178 = ( n16071 & n19395 ) | ( n16071 & ~n20635 ) | ( n19395 & ~n20635 ) ;
  assign n43179 = n31226 ^ n22424 ^ 1'b0 ;
  assign n43180 = ( n17498 & n43178 ) | ( n17498 & ~n43179 ) | ( n43178 & ~n43179 ) ;
  assign n43181 = ( ~n16422 & n22182 ) | ( ~n16422 & n28344 ) | ( n22182 & n28344 ) ;
  assign n43182 = n23962 ^ n13907 ^ 1'b0 ;
  assign n43183 = ~n2131 & n5254 ;
  assign n43184 = n9081 & n43183 ;
  assign n43185 = n43184 ^ n997 ^ 1'b0 ;
  assign n43186 = n17489 | n28192 ;
  assign n43187 = n28579 | n43186 ;
  assign n43188 = n7604 | n22795 ;
  assign n43189 = n43187 | n43188 ;
  assign n43190 = n8603 ^ n2234 ^ 1'b0 ;
  assign n43191 = n1564 & n43190 ;
  assign n43192 = ~n5209 & n28423 ;
  assign n43193 = n16442 & n43192 ;
  assign n43194 = n17630 | n20925 ;
  assign n43195 = n43194 ^ n5449 ^ 1'b0 ;
  assign n43196 = n21098 ^ n14674 ^ n9996 ;
  assign n43197 = ( n43193 & n43195 ) | ( n43193 & n43196 ) | ( n43195 & n43196 ) ;
  assign n43198 = n5561 & n6504 ;
  assign n43199 = ( n7293 & ~n35821 ) | ( n7293 & n43198 ) | ( ~n35821 & n43198 ) ;
  assign n43202 = n11179 ^ n4015 ^ 1'b0 ;
  assign n43203 = ( n4910 & n16890 ) | ( n4910 & n43202 ) | ( n16890 & n43202 ) ;
  assign n43204 = n43203 ^ n28597 ^ n20847 ;
  assign n43205 = ~n15926 & n20149 ;
  assign n43206 = n43204 & n43205 ;
  assign n43200 = n21481 ^ n12167 ^ 1'b0 ;
  assign n43201 = n8658 & ~n43200 ;
  assign n43207 = n43206 ^ n43201 ^ n5542 ;
  assign n43215 = n39257 ^ n35920 ^ n2095 ;
  assign n43212 = n9257 ^ n6893 ^ n4099 ;
  assign n43213 = ~n7406 & n12243 ;
  assign n43214 = ~n43212 & n43213 ;
  assign n43208 = ~n7618 & n24403 ;
  assign n43209 = n43208 ^ n13166 ^ 1'b0 ;
  assign n43210 = n22025 ^ n1138 ^ 1'b0 ;
  assign n43211 = ( n42312 & n43209 ) | ( n42312 & ~n43210 ) | ( n43209 & ~n43210 ) ;
  assign n43216 = n43215 ^ n43214 ^ n43211 ;
  assign n43217 = n42147 ^ n36276 ^ n10967 ;
  assign n43218 = n14966 & ~n23650 ;
  assign n43219 = n43218 ^ n12631 ^ 1'b0 ;
  assign n43220 = n3107 & ~n43219 ;
  assign n43221 = ( n20663 & n32859 ) | ( n20663 & n37244 ) | ( n32859 & n37244 ) ;
  assign n43223 = ( n3021 & n14125 ) | ( n3021 & n26041 ) | ( n14125 & n26041 ) ;
  assign n43222 = n33960 ^ n2372 ^ 1'b0 ;
  assign n43224 = n43223 ^ n43222 ^ 1'b0 ;
  assign n43225 = ( n3723 & n6211 ) | ( n3723 & ~n19107 ) | ( n6211 & ~n19107 ) ;
  assign n43226 = n34983 ^ n30276 ^ n6692 ;
  assign n43227 = n19558 ^ n13890 ^ n4333 ;
  assign n43228 = n1466 & ~n27595 ;
  assign n43229 = n35281 ^ n15378 ^ 1'b0 ;
  assign n43230 = n43229 ^ n5717 ^ 1'b0 ;
  assign n43231 = n43228 | n43230 ;
  assign n43232 = n12108 & ~n28257 ;
  assign n43233 = n17978 | n25851 ;
  assign n43234 = n19909 | n43233 ;
  assign n43235 = n43234 ^ n14769 ^ x0 ;
  assign n43236 = n43235 ^ x181 ^ 1'b0 ;
  assign n43244 = n7725 & n11474 ;
  assign n43245 = n43244 ^ n15471 ^ n4024 ;
  assign n43242 = n12078 & ~n37345 ;
  assign n43243 = n9564 & n43242 ;
  assign n43240 = n15769 ^ n10088 ^ 1'b0 ;
  assign n43241 = n43240 ^ n5175 ^ 1'b0 ;
  assign n43246 = n43245 ^ n43243 ^ n43241 ;
  assign n43237 = ~n2725 & n14798 ;
  assign n43238 = n43237 ^ n43007 ^ n1538 ;
  assign n43239 = n5129 | n43238 ;
  assign n43247 = n43246 ^ n43239 ^ n17125 ;
  assign n43248 = ( n2911 & n10274 ) | ( n2911 & n13296 ) | ( n10274 & n13296 ) ;
  assign n43249 = n43248 ^ n36551 ^ n12538 ;
  assign n43250 = ( n1796 & ~n20016 ) | ( n1796 & n43249 ) | ( ~n20016 & n43249 ) ;
  assign n43251 = n18865 | n26231 ;
  assign n43252 = n35860 | n43251 ;
  assign n43254 = ( n13338 & n14562 ) | ( n13338 & ~n29272 ) | ( n14562 & ~n29272 ) ;
  assign n43253 = n21961 & n39152 ;
  assign n43255 = n43254 ^ n43253 ^ 1'b0 ;
  assign n43256 = n4804 & n42573 ;
  assign n43257 = n43256 ^ n26896 ^ 1'b0 ;
  assign n43258 = n43257 ^ n9317 ^ 1'b0 ;
  assign n43259 = n31098 & n43258 ;
  assign n43260 = n31834 | n36755 ;
  assign n43261 = ( n15111 & n31833 ) | ( n15111 & ~n43260 ) | ( n31833 & ~n43260 ) ;
  assign n43262 = ( n25286 & ~n35939 ) | ( n25286 & n43240 ) | ( ~n35939 & n43240 ) ;
  assign n43263 = ( n11725 & n23437 ) | ( n11725 & ~n42276 ) | ( n23437 & ~n42276 ) ;
  assign n43264 = n6164 & ~n33547 ;
  assign n43265 = ( n16615 & ~n40005 ) | ( n16615 & n43264 ) | ( ~n40005 & n43264 ) ;
  assign n43266 = ( ~n7681 & n25013 ) | ( ~n7681 & n43265 ) | ( n25013 & n43265 ) ;
  assign n43267 = ~n22451 & n32419 ;
  assign n43268 = n43266 & n43267 ;
  assign n43269 = ( n19873 & n24511 ) | ( n19873 & n43268 ) | ( n24511 & n43268 ) ;
  assign n43270 = n7929 | n22370 ;
  assign n43271 = n33211 ^ n6842 ^ 1'b0 ;
  assign n43272 = n27182 | n43271 ;
  assign n43273 = n18888 & n21885 ;
  assign n43274 = n43273 ^ n2398 ^ 1'b0 ;
  assign n43275 = n36181 ^ n8082 ^ 1'b0 ;
  assign n43276 = n43274 | n43275 ;
  assign n43277 = n13124 | n25351 ;
  assign n43278 = n20599 | n43277 ;
  assign n43279 = n14465 ^ n4833 ^ 1'b0 ;
  assign n43280 = n7291 | n43279 ;
  assign n43281 = ( n3577 & n34859 ) | ( n3577 & ~n43280 ) | ( n34859 & ~n43280 ) ;
  assign n43282 = ( n1352 & ~n8248 ) | ( n1352 & n43281 ) | ( ~n8248 & n43281 ) ;
  assign n43283 = n34442 & n43282 ;
  assign n43284 = n31572 ^ n29704 ^ 1'b0 ;
  assign n43285 = ( n3904 & n8757 ) | ( n3904 & n21001 ) | ( n8757 & n21001 ) ;
  assign n43286 = n43285 ^ n42942 ^ n8276 ;
  assign n43287 = ( n6583 & ~n15594 ) | ( n6583 & n43286 ) | ( ~n15594 & n43286 ) ;
  assign n43288 = n18198 ^ n15639 ^ 1'b0 ;
  assign n43289 = n5108 & ~n43288 ;
  assign n43291 = n10889 | n16866 ;
  assign n43290 = n11915 | n35697 ;
  assign n43292 = n43291 ^ n43290 ^ 1'b0 ;
  assign n43293 = n9941 ^ n1793 ^ 1'b0 ;
  assign n43294 = ( n3067 & n12739 ) | ( n3067 & n18640 ) | ( n12739 & n18640 ) ;
  assign n43295 = n14568 & n20096 ;
  assign n43296 = n20844 | n43295 ;
  assign n43297 = n15817 & ~n43296 ;
  assign n43298 = ( ~n21142 & n43294 ) | ( ~n21142 & n43297 ) | ( n43294 & n43297 ) ;
  assign n43299 = n33790 ^ n33710 ^ 1'b0 ;
  assign n43300 = n41592 ^ n28121 ^ n5397 ;
  assign n43301 = ( n42984 & n43299 ) | ( n42984 & ~n43300 ) | ( n43299 & ~n43300 ) ;
  assign n43302 = n10041 ^ n9931 ^ 1'b0 ;
  assign n43303 = ~n35489 & n43302 ;
  assign n43304 = n3036 & n39647 ;
  assign n43305 = n7859 & n43304 ;
  assign n43306 = ~n8355 & n43305 ;
  assign n43307 = ( n1291 & n43303 ) | ( n1291 & n43306 ) | ( n43303 & n43306 ) ;
  assign n43308 = n14279 ^ n8111 ^ 1'b0 ;
  assign n43309 = n17433 ^ n13461 ^ 1'b0 ;
  assign n43310 = n5809 & n43309 ;
  assign n43311 = n26753 ^ n6642 ^ 1'b0 ;
  assign n43312 = ~n12205 & n43311 ;
  assign n43313 = n1328 & n8555 ;
  assign n43314 = n40012 | n43313 ;
  assign n43315 = n43012 ^ n1934 ^ 1'b0 ;
  assign n43316 = n43315 ^ n28738 ^ 1'b0 ;
  assign n43317 = n37967 ^ n4818 ^ 1'b0 ;
  assign n43318 = n20712 & ~n24092 ;
  assign n43319 = ( n16639 & n20670 ) | ( n16639 & n34436 ) | ( n20670 & n34436 ) ;
  assign n43320 = ( ~n43317 & n43318 ) | ( ~n43317 & n43319 ) | ( n43318 & n43319 ) ;
  assign n43321 = ( n5459 & ~n21337 ) | ( n5459 & n24730 ) | ( ~n21337 & n24730 ) ;
  assign n43326 = ~n2585 & n3984 ;
  assign n43327 = n43326 ^ n2117 ^ 1'b0 ;
  assign n43322 = ~n1294 & n5646 ;
  assign n43323 = n24002 & n43322 ;
  assign n43324 = n43323 ^ n24235 ^ n9075 ;
  assign n43325 = n4969 & n43324 ;
  assign n43328 = n43327 ^ n43325 ^ 1'b0 ;
  assign n43329 = n24366 ^ n8139 ^ 1'b0 ;
  assign n43330 = n8552 ^ n2095 ^ 1'b0 ;
  assign n43331 = n29005 ^ n27842 ^ n8264 ;
  assign n43334 = n5615 | n13064 ;
  assign n43335 = n8033 | n43334 ;
  assign n43336 = n43335 ^ n22461 ^ 1'b0 ;
  assign n43332 = n6702 ^ n1717 ^ 1'b0 ;
  assign n43333 = n12432 & ~n43332 ;
  assign n43337 = n43336 ^ n43333 ^ 1'b0 ;
  assign n43338 = ~n43331 & n43337 ;
  assign n43339 = ( n7421 & n12041 ) | ( n7421 & n35541 ) | ( n12041 & n35541 ) ;
  assign n43340 = n21008 ^ n17073 ^ n8793 ;
  assign n43341 = n43339 & ~n43340 ;
  assign n43342 = ( n13924 & ~n41335 ) | ( n13924 & n43341 ) | ( ~n41335 & n43341 ) ;
  assign n43345 = n5750 | n13203 ;
  assign n43346 = n43345 ^ n7229 ^ 1'b0 ;
  assign n43347 = ( ~n3185 & n42996 ) | ( ~n3185 & n43346 ) | ( n42996 & n43346 ) ;
  assign n43343 = n21917 ^ n19615 ^ n2569 ;
  assign n43344 = ( ~n21071 & n40583 ) | ( ~n21071 & n43343 ) | ( n40583 & n43343 ) ;
  assign n43348 = n43347 ^ n43344 ^ n28307 ;
  assign n43349 = ( n7924 & ~n15799 ) | ( n7924 & n34934 ) | ( ~n15799 & n34934 ) ;
  assign n43350 = ( ~n10710 & n16053 ) | ( ~n10710 & n17021 ) | ( n16053 & n17021 ) ;
  assign n43351 = n32167 ^ n24832 ^ 1'b0 ;
  assign n43352 = n10317 | n11883 ;
  assign n43353 = n43352 ^ n33883 ^ n8281 ;
  assign n43354 = n10482 & n43353 ;
  assign n43356 = n25520 ^ n22010 ^ n15341 ;
  assign n43355 = ~n3611 & n18658 ;
  assign n43357 = n43356 ^ n43355 ^ 1'b0 ;
  assign n43358 = n4963 & n4991 ;
  assign n43359 = n19907 & n26331 ;
  assign n43360 = n43358 & ~n43359 ;
  assign n43361 = n5815 ^ n5093 ^ n3351 ;
  assign n43362 = ( n6176 & n8453 ) | ( n6176 & n43361 ) | ( n8453 & n43361 ) ;
  assign n43363 = n43362 ^ n33387 ^ 1'b0 ;
  assign n43364 = n43363 ^ n23418 ^ n1727 ;
  assign n43365 = ( ~n327 & n12252 ) | ( ~n327 & n43364 ) | ( n12252 & n43364 ) ;
  assign n43366 = n33561 ^ n13049 ^ 1'b0 ;
  assign n43367 = n19646 ^ n13429 ^ 1'b0 ;
  assign n43368 = n9311 & ~n43367 ;
  assign n43369 = ( n5883 & n8276 ) | ( n5883 & ~n19744 ) | ( n8276 & ~n19744 ) ;
  assign n43370 = n43369 ^ n21783 ^ 1'b0 ;
  assign n43371 = ( n880 & n36781 ) | ( n880 & n43370 ) | ( n36781 & n43370 ) ;
  assign n43372 = n43371 ^ n1058 ^ 1'b0 ;
  assign n43373 = ~n35688 & n43372 ;
  assign n43374 = n38135 ^ n32037 ^ 1'b0 ;
  assign n43375 = n41749 ^ n5175 ^ 1'b0 ;
  assign n43376 = n32312 ^ n21318 ^ n16382 ;
  assign n43377 = n43376 ^ n2018 ^ 1'b0 ;
  assign n43378 = n39978 ^ n30057 ^ n10819 ;
  assign n43379 = ( ~x162 & n21023 ) | ( ~x162 & n37897 ) | ( n21023 & n37897 ) ;
  assign n43380 = ( n16063 & n17987 ) | ( n16063 & n43379 ) | ( n17987 & n43379 ) ;
  assign n43381 = n36189 ^ n34389 ^ n25845 ;
  assign n43382 = ( ~n6439 & n8188 ) | ( ~n6439 & n13573 ) | ( n8188 & n13573 ) ;
  assign n43384 = ( n4348 & ~n27201 ) | ( n4348 & n33404 ) | ( ~n27201 & n33404 ) ;
  assign n43385 = n43384 ^ n25805 ^ n6868 ;
  assign n43386 = n43385 ^ n41174 ^ n38990 ;
  assign n43383 = n23964 & n24514 ;
  assign n43387 = n43386 ^ n43383 ^ 1'b0 ;
  assign n43388 = n19112 ^ n13482 ^ 1'b0 ;
  assign n43389 = ~n18637 & n43388 ;
  assign n43390 = n15538 ^ n7070 ^ 1'b0 ;
  assign n43391 = n1317 & ~n43390 ;
  assign n43392 = n43391 ^ n22942 ^ n14320 ;
  assign n43393 = n6096 & ~n17776 ;
  assign n43394 = n11248 ^ n4490 ^ 1'b0 ;
  assign n43395 = n43393 | n43394 ;
  assign n43396 = n26237 ^ n2481 ^ 1'b0 ;
  assign n43397 = n43395 | n43396 ;
  assign n43398 = n43397 ^ n4213 ^ 1'b0 ;
  assign n43399 = n43398 ^ n25122 ^ n13410 ;
  assign n43400 = ~n27895 & n28294 ;
  assign n43402 = n7554 ^ n5086 ^ n2614 ;
  assign n43401 = n24822 ^ n6263 ^ n4256 ;
  assign n43403 = n43402 ^ n43401 ^ n11206 ;
  assign n43404 = n43403 ^ n23796 ^ n19542 ;
  assign n43405 = n28284 ^ n6969 ^ n3116 ;
  assign n43406 = n43405 ^ n24693 ^ 1'b0 ;
  assign n43407 = n8582 | n20217 ;
  assign n43408 = n43406 & ~n43407 ;
  assign n43409 = ( n19453 & ~n30307 ) | ( n19453 & n43408 ) | ( ~n30307 & n43408 ) ;
  assign n43410 = n971 & ~n12799 ;
  assign n43411 = ~n11147 & n43410 ;
  assign n43412 = n10873 | n43411 ;
  assign n43413 = n43412 ^ n20774 ^ 1'b0 ;
  assign n43414 = n43413 ^ n14438 ^ 1'b0 ;
  assign n43415 = n9308 & n43414 ;
  assign n43416 = ~n24089 & n32853 ;
  assign n43417 = n43416 ^ n18144 ^ 1'b0 ;
  assign n43418 = n27040 | n43417 ;
  assign n43419 = n14784 | n43418 ;
  assign n43420 = n21954 ^ n2306 ^ 1'b0 ;
  assign n43421 = n2147 & n43420 ;
  assign n43422 = n43421 ^ n12478 ^ n1937 ;
  assign n43423 = n27738 ^ x21 ^ 1'b0 ;
  assign n43424 = n12739 ^ n3216 ^ 1'b0 ;
  assign n43425 = n4085 & ~n43424 ;
  assign n43426 = n43425 ^ n41926 ^ 1'b0 ;
  assign n43427 = n21742 ^ n7326 ^ x40 ;
  assign n43428 = ( n13502 & ~n23594 ) | ( n13502 & n43427 ) | ( ~n23594 & n43427 ) ;
  assign n43429 = n2824 & n14927 ;
  assign n43431 = ( ~n14657 & n22545 ) | ( ~n14657 & n26283 ) | ( n22545 & n26283 ) ;
  assign n43430 = ( n3013 & ~n31952 ) | ( n3013 & n34949 ) | ( ~n31952 & n34949 ) ;
  assign n43432 = n43431 ^ n43430 ^ 1'b0 ;
  assign n43433 = n963 | n10075 ;
  assign n43434 = n30045 ^ n15015 ^ 1'b0 ;
  assign n43435 = x97 & n43434 ;
  assign n43436 = ~n22370 & n43435 ;
  assign n43437 = ( n1296 & n43433 ) | ( n1296 & ~n43436 ) | ( n43433 & ~n43436 ) ;
  assign n43438 = n3752 ^ n2527 ^ 1'b0 ;
  assign n43439 = ( n21562 & ~n38098 ) | ( n21562 & n43438 ) | ( ~n38098 & n43438 ) ;
  assign n43440 = n23039 & n39645 ;
  assign n43441 = n12368 ^ n701 ^ 1'b0 ;
  assign n43442 = n37456 & n43441 ;
  assign n43443 = n20365 | n43442 ;
  assign n43444 = n11084 & n40539 ;
  assign n43445 = n43444 ^ n18083 ^ 1'b0 ;
  assign n43446 = ( ~n7641 & n15726 ) | ( ~n7641 & n35109 ) | ( n15726 & n35109 ) ;
  assign n43447 = n43446 ^ n42296 ^ n37489 ;
  assign n43448 = n16697 ^ n14923 ^ 1'b0 ;
  assign n43449 = n8388 & ~n43448 ;
  assign n43450 = ( ~n6059 & n17910 ) | ( ~n6059 & n33146 ) | ( n17910 & n33146 ) ;
  assign n43451 = n43449 & n43450 ;
  assign n43452 = n21685 ^ n13971 ^ n11166 ;
  assign n43453 = n11068 ^ n7103 ^ 1'b0 ;
  assign n43454 = ( ~n4179 & n26953 ) | ( ~n4179 & n43453 ) | ( n26953 & n43453 ) ;
  assign n43455 = n39297 ^ n30957 ^ n28724 ;
  assign n43456 = n34001 ^ n27145 ^ 1'b0 ;
  assign n43457 = n37932 & ~n43456 ;
  assign n43458 = ( n2369 & n23009 ) | ( n2369 & ~n43457 ) | ( n23009 & ~n43457 ) ;
  assign n43459 = n13752 ^ n8842 ^ 1'b0 ;
  assign n43460 = ( x185 & ~n439 ) | ( x185 & n4630 ) | ( ~n439 & n4630 ) ;
  assign n43461 = n21386 | n30303 ;
  assign n43462 = n43460 & n43461 ;
  assign n43463 = n43459 & n43462 ;
  assign n43464 = ( n17843 & ~n26642 ) | ( n17843 & n30740 ) | ( ~n26642 & n30740 ) ;
  assign n43465 = ( x218 & n16625 ) | ( x218 & ~n25641 ) | ( n16625 & ~n25641 ) ;
  assign n43466 = ~n7339 & n43465 ;
  assign n43467 = n43464 & n43466 ;
  assign n43468 = n40306 ^ n31361 ^ n9188 ;
  assign n43469 = n15580 ^ n6706 ^ n4310 ;
  assign n43470 = n41265 & ~n43469 ;
  assign n43471 = n28771 ^ n7603 ^ n3729 ;
  assign n43472 = ( n10107 & n12612 ) | ( n10107 & n32912 ) | ( n12612 & n32912 ) ;
  assign n43473 = n33442 & ~n43472 ;
  assign n43474 = n29417 ^ n1949 ^ n1025 ;
  assign n43475 = ( n25501 & n35149 ) | ( n25501 & n43474 ) | ( n35149 & n43474 ) ;
  assign n43476 = ~n18688 & n39030 ;
  assign n43477 = n43476 ^ n8168 ^ 1'b0 ;
  assign n43478 = n19265 ^ n2882 ^ 1'b0 ;
  assign n43479 = n1125 & ~n5325 ;
  assign n43480 = n18690 & n43479 ;
  assign n43484 = n39216 ^ n4975 ^ 1'b0 ;
  assign n43482 = n23620 & n26251 ;
  assign n43483 = n23611 & n43482 ;
  assign n43481 = n6024 | n12207 ;
  assign n43485 = n43484 ^ n43483 ^ n43481 ;
  assign n43486 = n35058 ^ n9544 ^ n5708 ;
  assign n43487 = n43486 ^ n433 ^ 1'b0 ;
  assign n43488 = ~n43485 & n43487 ;
  assign n43489 = ~n11675 & n13555 ;
  assign n43490 = ( ~n3015 & n5768 ) | ( ~n3015 & n42745 ) | ( n5768 & n42745 ) ;
  assign n43491 = n28695 ^ n19159 ^ n1639 ;
  assign n43492 = ( n13296 & n31256 ) | ( n13296 & ~n43491 ) | ( n31256 & ~n43491 ) ;
  assign n43493 = n19560 ^ n16513 ^ n10025 ;
  assign n43494 = ( n470 & n3213 ) | ( n470 & n36033 ) | ( n3213 & n36033 ) ;
  assign n43495 = n11492 & n43494 ;
  assign n43496 = n11261 & n43495 ;
  assign n43497 = ~n4101 & n5217 ;
  assign n43498 = n43497 ^ n21833 ^ 1'b0 ;
  assign n43499 = ( n1408 & n9143 ) | ( n1408 & ~n19486 ) | ( n9143 & ~n19486 ) ;
  assign n43500 = n15845 & n43499 ;
  assign n43501 = n13618 ^ n5910 ^ n2250 ;
  assign n43502 = n10423 ^ n6206 ^ 1'b0 ;
  assign n43503 = n43501 & n43502 ;
  assign n43504 = n27185 ^ n15243 ^ 1'b0 ;
  assign n43505 = n38375 ^ n31846 ^ n1268 ;
  assign n43506 = ( n3329 & n16497 ) | ( n3329 & ~n17476 ) | ( n16497 & ~n17476 ) ;
  assign n43507 = n43506 ^ n8737 ^ 1'b0 ;
  assign n43508 = n29031 ^ n19591 ^ 1'b0 ;
  assign n43509 = ( n10030 & ~n20925 ) | ( n10030 & n43508 ) | ( ~n20925 & n43508 ) ;
  assign n43510 = n25940 ^ n19409 ^ n18518 ;
  assign n43511 = n20873 ^ n11541 ^ n6235 ;
  assign n43512 = n34301 & ~n43511 ;
  assign n43513 = n43512 ^ n19734 ^ 1'b0 ;
  assign n43514 = n9404 ^ n3021 ^ 1'b0 ;
  assign n43515 = n2106 & n43514 ;
  assign n43516 = n2279 | n43515 ;
  assign n43517 = ~n3330 & n43516 ;
  assign n43518 = n43151 ^ n12193 ^ 1'b0 ;
  assign n43519 = n30541 & n38939 ;
  assign n43520 = n43519 ^ n19825 ^ n13087 ;
  assign n43521 = ( n7664 & n7795 ) | ( n7664 & ~n43520 ) | ( n7795 & ~n43520 ) ;
  assign n43522 = n43484 ^ n41014 ^ n11354 ;
  assign n43523 = x210 & ~n43522 ;
  assign n43524 = n2813 & ~n30654 ;
  assign n43525 = n43524 ^ n14770 ^ n12690 ;
  assign n43526 = n43525 ^ n15546 ^ 1'b0 ;
  assign n43527 = n11616 ^ n3261 ^ 1'b0 ;
  assign n43528 = n43527 ^ n13469 ^ n1980 ;
  assign n43529 = n963 & ~n43528 ;
  assign n43530 = n15246 & n22649 ;
  assign n43531 = n36976 ^ n14408 ^ 1'b0 ;
  assign n43532 = n36846 ^ n28007 ^ 1'b0 ;
  assign n43533 = n2604 ^ n2291 ^ 1'b0 ;
  assign n43534 = n8408 | n43533 ;
  assign n43535 = n43534 ^ n24776 ^ 1'b0 ;
  assign n43536 = n43532 & ~n43535 ;
  assign n43537 = n41295 ^ x82 ^ 1'b0 ;
  assign n43538 = n21817 & ~n43537 ;
  assign n43539 = n4502 ^ n3151 ^ 1'b0 ;
  assign n43540 = n31069 ^ n6384 ^ n1839 ;
  assign n43541 = ( n23617 & n40178 ) | ( n23617 & n43540 ) | ( n40178 & n43540 ) ;
  assign n43542 = ( n3314 & n26417 ) | ( n3314 & ~n35237 ) | ( n26417 & ~n35237 ) ;
  assign n43543 = n33584 ^ n17861 ^ 1'b0 ;
  assign n43544 = n15742 ^ n8307 ^ n7664 ;
  assign n43545 = n18217 | n43544 ;
  assign n43546 = n17724 & n30012 ;
  assign n43547 = n18035 & n43546 ;
  assign n43548 = n36882 ^ n26973 ^ 1'b0 ;
  assign n43549 = n31098 & n43548 ;
  assign n43550 = n17221 | n20184 ;
  assign n43551 = n1804 & ~n36426 ;
  assign n43552 = n36072 ^ n15521 ^ n11670 ;
  assign n43553 = ( n3317 & ~n37994 ) | ( n3317 & n43552 ) | ( ~n37994 & n43552 ) ;
  assign n43554 = n12589 & n30847 ;
  assign n43555 = n5069 | n12021 ;
  assign n43556 = ( n13146 & ~n18870 ) | ( n13146 & n37813 ) | ( ~n18870 & n37813 ) ;
  assign n43557 = ( n15932 & n29519 ) | ( n15932 & ~n29689 ) | ( n29519 & ~n29689 ) ;
  assign n43558 = n41482 ^ n33244 ^ 1'b0 ;
  assign n43559 = n9401 & n43558 ;
  assign n43560 = n43559 ^ n8538 ^ 1'b0 ;
  assign n43561 = n22311 | n43244 ;
  assign n43562 = n43561 ^ n23828 ^ 1'b0 ;
  assign n43563 = n8307 | n19663 ;
  assign n43564 = ( ~n24717 & n35720 ) | ( ~n24717 & n43563 ) | ( n35720 & n43563 ) ;
  assign n43565 = n31500 ^ n5584 ^ 1'b0 ;
  assign n43566 = ~n2430 & n26577 ;
  assign n43567 = n43566 ^ n30017 ^ n4930 ;
  assign n43568 = n19382 & ~n41571 ;
  assign n43569 = n21624 & n43568 ;
  assign n43570 = n43569 ^ n36686 ^ n9751 ;
  assign n43571 = n27558 ^ n12028 ^ 1'b0 ;
  assign n43572 = n15090 & n43571 ;
  assign n43573 = ( n11588 & n13036 ) | ( n11588 & ~n37039 ) | ( n13036 & ~n37039 ) ;
  assign n43574 = n43573 ^ n39568 ^ 1'b0 ;
  assign n43575 = n25787 | n43574 ;
  assign n43576 = n9921 ^ n9692 ^ 1'b0 ;
  assign n43577 = n8594 | n43576 ;
  assign n43578 = n11037 ^ n3861 ^ 1'b0 ;
  assign n43579 = n10149 & ~n43578 ;
  assign n43580 = ( n1025 & n22656 ) | ( n1025 & n43579 ) | ( n22656 & n43579 ) ;
  assign n43581 = ~n39352 & n42706 ;
  assign n43582 = n43581 ^ n13586 ^ n4217 ;
  assign n43583 = n25034 ^ x238 ^ 1'b0 ;
  assign n43584 = n36561 ^ n27837 ^ n10766 ;
  assign n43585 = n21363 | n39319 ;
  assign n43586 = ( ~n2350 & n27645 ) | ( ~n2350 & n42847 ) | ( n27645 & n42847 ) ;
  assign n43587 = ( n29466 & n31657 ) | ( n29466 & n43586 ) | ( n31657 & n43586 ) ;
  assign n43588 = n5125 | n5837 ;
  assign n43589 = n41979 | n43588 ;
  assign n43590 = n43587 | n43589 ;
  assign n43591 = n26695 ^ n1980 ^ 1'b0 ;
  assign n43592 = n42892 ^ n38418 ^ 1'b0 ;
  assign n43593 = ~n8398 & n43592 ;
  assign n43594 = n11349 ^ n10886 ^ n10095 ;
  assign n43595 = n7572 | n40297 ;
  assign n43596 = n43595 ^ n27482 ^ 1'b0 ;
  assign n43597 = n43594 & ~n43596 ;
  assign n43598 = n7352 ^ n2126 ^ 1'b0 ;
  assign n43599 = n43598 ^ n17461 ^ n14885 ;
  assign n43600 = ( n427 & n14106 ) | ( n427 & ~n22379 ) | ( n14106 & ~n22379 ) ;
  assign n43601 = n4858 & n16099 ;
  assign n43602 = n43601 ^ n15442 ^ 1'b0 ;
  assign n43603 = n43600 | n43602 ;
  assign n43604 = x87 & n25364 ;
  assign n43605 = n30954 | n43604 ;
  assign n43606 = n43605 ^ n36381 ^ 1'b0 ;
  assign n43607 = n2095 | n4351 ;
  assign n43608 = n13444 | n43607 ;
  assign n43609 = n43608 ^ n12805 ^ 1'b0 ;
  assign n43610 = n43609 ^ n20289 ^ n9176 ;
  assign n43612 = n26013 ^ n24308 ^ n2940 ;
  assign n43611 = n37107 | n39100 ;
  assign n43613 = n43612 ^ n43611 ^ n9709 ;
  assign n43614 = x184 & ~n5975 ;
  assign n43615 = ~n19003 & n43614 ;
  assign n43616 = n43615 ^ n8038 ^ 1'b0 ;
  assign n43617 = ~n26043 & n43616 ;
  assign n43618 = n25131 ^ n24955 ^ n10469 ;
  assign n43619 = n43618 ^ n28113 ^ 1'b0 ;
  assign n43620 = n3274 & ~n43619 ;
  assign n43621 = n32267 ^ n7317 ^ n1137 ;
  assign n43622 = ~n21596 & n43621 ;
  assign n43624 = ( n2165 & n3624 ) | ( n2165 & ~n22839 ) | ( n3624 & ~n22839 ) ;
  assign n43623 = n21840 ^ n20058 ^ n8332 ;
  assign n43625 = n43624 ^ n43623 ^ n13648 ;
  assign n43626 = n6781 & n37961 ;
  assign n43627 = n43626 ^ n1096 ^ 1'b0 ;
  assign n43628 = n17053 | n43627 ;
  assign n43629 = n43628 ^ n41582 ^ n16268 ;
  assign n43634 = ( n27927 & n27995 ) | ( n27927 & ~n39436 ) | ( n27995 & ~n39436 ) ;
  assign n43632 = n8104 & n41416 ;
  assign n43633 = ( n8595 & n25108 ) | ( n8595 & ~n43632 ) | ( n25108 & ~n43632 ) ;
  assign n43630 = n20280 ^ n9693 ^ 1'b0 ;
  assign n43631 = n25095 & n43630 ;
  assign n43635 = n43634 ^ n43633 ^ n43631 ;
  assign n43636 = n4583 | n4931 ;
  assign n43637 = n7474 & ~n26009 ;
  assign n43638 = ( ~n4357 & n27436 ) | ( ~n4357 & n35566 ) | ( n27436 & n35566 ) ;
  assign n43639 = ( ~n43636 & n43637 ) | ( ~n43636 & n43638 ) | ( n43637 & n43638 ) ;
  assign n43640 = n41071 ^ n24848 ^ n2094 ;
  assign n43641 = n32482 ^ n28001 ^ n14783 ;
  assign n43642 = n43641 ^ n315 ^ 1'b0 ;
  assign n43643 = ( n25916 & n43640 ) | ( n25916 & n43642 ) | ( n43640 & n43642 ) ;
  assign n43644 = ~n3958 & n18925 ;
  assign n43645 = n10229 & n18169 ;
  assign n43646 = ( n21287 & n27769 ) | ( n21287 & n30336 ) | ( n27769 & n30336 ) ;
  assign n43647 = n17372 | n43646 ;
  assign n43648 = ( n3353 & ~n11802 ) | ( n3353 & n15225 ) | ( ~n11802 & n15225 ) ;
  assign n43649 = n43648 ^ n16353 ^ 1'b0 ;
  assign n43650 = n1989 | n43649 ;
  assign n43651 = ( n1684 & n17356 ) | ( n1684 & ~n43650 ) | ( n17356 & ~n43650 ) ;
  assign n43652 = n25808 ^ n23355 ^ n12340 ;
  assign n43653 = n31130 ^ n20114 ^ n7702 ;
  assign n43654 = n2538 & n14013 ;
  assign n43655 = ( ~n3309 & n38615 ) | ( ~n3309 & n43654 ) | ( n38615 & n43654 ) ;
  assign n43656 = n25112 ^ n5775 ^ n1003 ;
  assign n43657 = n23418 | n26858 ;
  assign n43658 = n43657 ^ n36896 ^ 1'b0 ;
  assign n43659 = n32299 ^ n6634 ^ n4003 ;
  assign n43660 = n43659 ^ n41418 ^ n34832 ;
  assign n43661 = ~n24597 & n43660 ;
  assign n43662 = n36391 ^ n27749 ^ n14987 ;
  assign n43663 = n31319 ^ n16972 ^ 1'b0 ;
  assign n43664 = n7049 & n35751 ;
  assign n43665 = n35142 ^ n32861 ^ n22275 ;
  assign n43666 = ( n6935 & n23929 ) | ( n6935 & n37229 ) | ( n23929 & n37229 ) ;
  assign n43667 = ( n2029 & n28344 ) | ( n2029 & n43666 ) | ( n28344 & n43666 ) ;
  assign n43668 = ( n6242 & ~n9310 ) | ( n6242 & n22799 ) | ( ~n9310 & n22799 ) ;
  assign n43669 = ~n28163 & n30333 ;
  assign n43670 = n9613 & ~n22458 ;
  assign n43671 = ~n41883 & n43670 ;
  assign n43672 = ~n23437 & n33506 ;
  assign n43673 = n43672 ^ n33983 ^ 1'b0 ;
  assign n43674 = n43673 ^ n23314 ^ n795 ;
  assign n43675 = ( n4772 & ~n15292 ) | ( n4772 & n30318 ) | ( ~n15292 & n30318 ) ;
  assign n43676 = n43675 ^ n39211 ^ 1'b0 ;
  assign n43677 = x198 & n22578 ;
  assign n43678 = n43677 ^ n5022 ^ 1'b0 ;
  assign n43679 = n43678 ^ n30852 ^ 1'b0 ;
  assign n43680 = n11359 ^ n7187 ^ n370 ;
  assign n43681 = n6332 | n15568 ;
  assign n43682 = n17069 & ~n43681 ;
  assign n43683 = n8070 | n33676 ;
  assign n43684 = n43683 ^ n30180 ^ 1'b0 ;
  assign n43685 = n1186 & n7621 ;
  assign n43686 = n2292 & n43685 ;
  assign n43687 = ( n5146 & ~n13768 ) | ( n5146 & n43686 ) | ( ~n13768 & n43686 ) ;
  assign n43688 = ( n3651 & n7127 ) | ( n3651 & n43687 ) | ( n7127 & n43687 ) ;
  assign n43689 = ~n11039 & n43688 ;
  assign n43690 = n43689 ^ n13691 ^ 1'b0 ;
  assign n43691 = n43030 & n43690 ;
  assign n43692 = n5820 | n8360 ;
  assign n43693 = n43692 ^ n7815 ^ 1'b0 ;
  assign n43694 = ( n30931 & n33835 ) | ( n30931 & ~n43693 ) | ( n33835 & ~n43693 ) ;
  assign n43695 = ( n11054 & ~n32022 ) | ( n11054 & n43433 ) | ( ~n32022 & n43433 ) ;
  assign n43696 = n5515 & ~n13866 ;
  assign n43697 = n43696 ^ n24943 ^ 1'b0 ;
  assign n43698 = n22742 ^ n18503 ^ 1'b0 ;
  assign n43699 = ( n10617 & ~n43697 ) | ( n10617 & n43698 ) | ( ~n43697 & n43698 ) ;
  assign n43700 = n31000 ^ n30946 ^ n25979 ;
  assign n43701 = ( n11766 & ~n13273 ) | ( n11766 & n21143 ) | ( ~n13273 & n21143 ) ;
  assign n43702 = n43701 ^ n6100 ^ n1826 ;
  assign n43703 = ( ~n31288 & n43700 ) | ( ~n31288 & n43702 ) | ( n43700 & n43702 ) ;
  assign n43704 = n41618 ^ n2412 ^ 1'b0 ;
  assign n43705 = n43704 ^ n26990 ^ n18460 ;
  assign n43706 = ( ~n23190 & n36649 ) | ( ~n23190 & n36998 ) | ( n36649 & n36998 ) ;
  assign n43707 = n29274 ^ n11742 ^ 1'b0 ;
  assign n43708 = ~n12607 & n41081 ;
  assign n43709 = n43708 ^ n42286 ^ 1'b0 ;
  assign n43710 = ( ~n4198 & n6505 ) | ( ~n4198 & n43709 ) | ( n6505 & n43709 ) ;
  assign n43711 = ( n13921 & n21081 ) | ( n13921 & n29506 ) | ( n21081 & n29506 ) ;
  assign n43712 = n2195 & n34068 ;
  assign n43713 = n43712 ^ x210 ^ 1'b0 ;
  assign n43714 = n43713 ^ n32903 ^ 1'b0 ;
  assign n43715 = ( n25971 & n43711 ) | ( n25971 & n43714 ) | ( n43711 & n43714 ) ;
  assign n43716 = ( ~n25515 & n35689 ) | ( ~n25515 & n43715 ) | ( n35689 & n43715 ) ;
  assign n43717 = n16483 ^ n12934 ^ 1'b0 ;
  assign n43719 = ( ~n1924 & n3278 ) | ( ~n1924 & n10769 ) | ( n3278 & n10769 ) ;
  assign n43720 = ( ~x78 & n24823 ) | ( ~x78 & n43719 ) | ( n24823 & n43719 ) ;
  assign n43718 = n3471 & n11954 ;
  assign n43721 = n43720 ^ n43718 ^ 1'b0 ;
  assign n43722 = ( n15142 & n18562 ) | ( n15142 & n28556 ) | ( n18562 & n28556 ) ;
  assign n43723 = n43722 ^ n22022 ^ 1'b0 ;
  assign n43724 = n9896 & ~n43723 ;
  assign n43725 = ~n26099 & n43724 ;
  assign n43726 = n43725 ^ n27975 ^ 1'b0 ;
  assign n43727 = ( n11364 & ~n27594 ) | ( n11364 & n35066 ) | ( ~n27594 & n35066 ) ;
  assign n43728 = ( n19128 & n38705 ) | ( n19128 & n39684 ) | ( n38705 & n39684 ) ;
  assign n43729 = n18788 & ~n43728 ;
  assign n43730 = n43727 & n43729 ;
  assign n43731 = n25473 ^ n5006 ^ 1'b0 ;
  assign n43732 = n9005 | n43731 ;
  assign n43734 = n28749 ^ n977 ^ 1'b0 ;
  assign n43735 = n20735 & ~n43734 ;
  assign n43733 = n30967 ^ n8722 ^ 1'b0 ;
  assign n43736 = n43735 ^ n43733 ^ n21750 ;
  assign n43737 = x5 & ~n29892 ;
  assign n43738 = ( n11541 & n26157 ) | ( n11541 & n43737 ) | ( n26157 & n43737 ) ;
  assign n43739 = ( n6341 & n18309 ) | ( n6341 & ~n24068 ) | ( n18309 & ~n24068 ) ;
  assign n43740 = n36131 ^ n7956 ^ 1'b0 ;
  assign n43741 = n19309 | n43740 ;
  assign n43742 = n9938 | n43741 ;
  assign n43743 = ~n19296 & n22555 ;
  assign n43744 = n14938 ^ n8561 ^ 1'b0 ;
  assign n43745 = n43744 ^ n25391 ^ n17936 ;
  assign n43746 = n6638 ^ n4946 ^ 1'b0 ;
  assign n43747 = n14311 ^ n1423 ^ 1'b0 ;
  assign n43748 = ~n7597 & n43747 ;
  assign n43749 = n43748 ^ n13829 ^ 1'b0 ;
  assign n43750 = ~n43746 & n43749 ;
  assign n43751 = n3109 & n33555 ;
  assign n43752 = n8594 ^ n440 ^ 1'b0 ;
  assign n43753 = n15482 & ~n43752 ;
  assign n43754 = n43753 ^ n12638 ^ 1'b0 ;
  assign n43755 = n23404 & n38051 ;
  assign n43756 = n43755 ^ n5633 ^ 1'b0 ;
  assign n43757 = n38128 ^ n33433 ^ 1'b0 ;
  assign n43758 = n43756 & ~n43757 ;
  assign n43759 = n20003 ^ n8722 ^ 1'b0 ;
  assign n43760 = n13620 ^ n8215 ^ 1'b0 ;
  assign n43761 = n9685 & n43760 ;
  assign n43762 = n32610 ^ n32066 ^ n4837 ;
  assign n43763 = ( ~n13478 & n36592 ) | ( ~n13478 & n43762 ) | ( n36592 & n43762 ) ;
  assign n43764 = n8416 | n12551 ;
  assign n43765 = ~n8824 & n11958 ;
  assign n43766 = n43765 ^ n513 ^ 1'b0 ;
  assign n43767 = ( ~n1599 & n43764 ) | ( ~n1599 & n43766 ) | ( n43764 & n43766 ) ;
  assign n43768 = n31102 & ~n41653 ;
  assign n43769 = n43768 ^ n28996 ^ 1'b0 ;
  assign n43770 = ~n15111 & n35678 ;
  assign n43771 = n17344 & n43770 ;
  assign n43772 = n26472 ^ n26399 ^ n16491 ;
  assign n43773 = ~n28398 & n43772 ;
  assign n43774 = n26492 ^ n20735 ^ 1'b0 ;
  assign n43775 = n11172 & n43774 ;
  assign n43776 = n43775 ^ n37078 ^ 1'b0 ;
  assign n43777 = n21505 & ~n37906 ;
  assign n43778 = n23185 ^ n17284 ^ 1'b0 ;
  assign n43779 = n32524 ^ n14609 ^ n6723 ;
  assign n43780 = n11318 | n29320 ;
  assign n43781 = ( n11492 & ~n13788 ) | ( n11492 & n43780 ) | ( ~n13788 & n43780 ) ;
  assign n43782 = n9177 | n26834 ;
  assign n43783 = n43782 ^ n33431 ^ 1'b0 ;
  assign n43784 = n13906 | n14443 ;
  assign n43785 = n34294 & n43784 ;
  assign n43786 = n43785 ^ n28842 ^ 1'b0 ;
  assign n43787 = n11265 ^ n3294 ^ 1'b0 ;
  assign n43788 = n43787 ^ n37300 ^ n3500 ;
  assign n43789 = ~n1803 & n2640 ;
  assign n43790 = ~n18593 & n43789 ;
  assign n43791 = n25913 & ~n43790 ;
  assign n43792 = n43791 ^ n14134 ^ 1'b0 ;
  assign n43793 = n43792 ^ n23954 ^ n12131 ;
  assign n43794 = n43793 ^ n13174 ^ 1'b0 ;
  assign n43795 = n43788 & ~n43794 ;
  assign n43796 = n3247 | n20209 ;
  assign n43797 = ( n962 & n10452 ) | ( n962 & ~n11605 ) | ( n10452 & ~n11605 ) ;
  assign n43798 = ( ~n15608 & n18586 ) | ( ~n15608 & n43797 ) | ( n18586 & n43797 ) ;
  assign n43799 = n5227 & n20305 ;
  assign n43800 = ~n12069 & n43799 ;
  assign n43801 = n23202 ^ n3640 ^ 1'b0 ;
  assign n43802 = ~n43800 & n43801 ;
  assign n43803 = ( n31183 & n43798 ) | ( n31183 & n43802 ) | ( n43798 & n43802 ) ;
  assign n43804 = ( ~n21999 & n22398 ) | ( ~n21999 & n32093 ) | ( n22398 & n32093 ) ;
  assign n43805 = ( n6739 & ~n34377 ) | ( n6739 & n43804 ) | ( ~n34377 & n43804 ) ;
  assign n43806 = ( n43796 & ~n43803 ) | ( n43796 & n43805 ) | ( ~n43803 & n43805 ) ;
  assign n43807 = n8276 ^ n1481 ^ 1'b0 ;
  assign n43808 = n43807 ^ n28184 ^ n6059 ;
  assign n43809 = ( n13049 & ~n15360 ) | ( n13049 & n21939 ) | ( ~n15360 & n21939 ) ;
  assign n43810 = ( n27340 & n34922 ) | ( n27340 & ~n43809 ) | ( n34922 & ~n43809 ) ;
  assign n43811 = ( n1670 & ~n41749 ) | ( n1670 & n43810 ) | ( ~n41749 & n43810 ) ;
  assign n43812 = n28930 | n39167 ;
  assign n43813 = ~n1545 & n43182 ;
  assign n43814 = ( n15993 & ~n27354 ) | ( n15993 & n43813 ) | ( ~n27354 & n43813 ) ;
  assign n43815 = n17306 & ~n35550 ;
  assign n43816 = ~n8917 & n43815 ;
  assign n43817 = n21901 & ~n38961 ;
  assign n43818 = n3705 & n43817 ;
  assign n43819 = n15822 ^ n11685 ^ n6224 ;
  assign n43820 = n42392 ^ n28954 ^ n10115 ;
  assign n43821 = ( n7117 & n43819 ) | ( n7117 & n43820 ) | ( n43819 & n43820 ) ;
  assign n43822 = ( n959 & n6066 ) | ( n959 & n43821 ) | ( n6066 & n43821 ) ;
  assign n43823 = ( n988 & n11989 ) | ( n988 & ~n19828 ) | ( n11989 & ~n19828 ) ;
  assign n43824 = n17282 ^ n10556 ^ 1'b0 ;
  assign n43825 = n43823 | n43824 ;
  assign n43826 = n43825 ^ n15887 ^ 1'b0 ;
  assign n43827 = ~n43822 & n43826 ;
  assign n43828 = ~n7461 & n29565 ;
  assign n43829 = n43828 ^ n32008 ^ 1'b0 ;
  assign n43830 = n10917 & n38846 ;
  assign n43831 = n10863 & ~n19957 ;
  assign n43832 = ~n5531 & n43831 ;
  assign n43833 = n43832 ^ n30457 ^ 1'b0 ;
  assign n43834 = n16115 & ~n20621 ;
  assign n43835 = ~n2167 & n43834 ;
  assign n43836 = ( n21046 & ~n29059 ) | ( n21046 & n43835 ) | ( ~n29059 & n43835 ) ;
  assign n43837 = n617 & ~n12764 ;
  assign n43838 = n29602 & ~n43837 ;
  assign n43839 = ( ~n22868 & n35252 ) | ( ~n22868 & n38529 ) | ( n35252 & n38529 ) ;
  assign n43840 = n23728 ^ n16894 ^ n9456 ;
  assign n43841 = n43840 ^ n28556 ^ n20818 ;
  assign n43842 = n8457 ^ n8124 ^ 1'b0 ;
  assign n43843 = ~n19086 & n43842 ;
  assign n43844 = n43843 ^ n20052 ^ n14414 ;
  assign n43845 = n5388 ^ n2707 ^ n1399 ;
  assign n43846 = n43845 ^ n15835 ^ n7871 ;
  assign n43847 = n28519 & ~n32177 ;
  assign n43848 = n43846 & n43847 ;
  assign n43849 = n28800 & ~n42628 ;
  assign n43850 = n43849 ^ n24625 ^ 1'b0 ;
  assign n43851 = n21740 ^ n12401 ^ n1859 ;
  assign n43852 = n32181 & n43851 ;
  assign n43853 = ( n2572 & n14725 ) | ( n2572 & n17017 ) | ( n14725 & n17017 ) ;
  assign n43854 = ( n7600 & n31800 ) | ( n7600 & ~n33598 ) | ( n31800 & ~n33598 ) ;
  assign n43855 = ( n20033 & ~n43853 ) | ( n20033 & n43854 ) | ( ~n43853 & n43854 ) ;
  assign n43856 = n41652 ^ n30091 ^ n2500 ;
  assign n43857 = ( ~n1073 & n2104 ) | ( ~n1073 & n15642 ) | ( n2104 & n15642 ) ;
  assign n43858 = n1832 & ~n2804 ;
  assign n43859 = n19275 | n21320 ;
  assign n43860 = n43859 ^ n42348 ^ n9171 ;
  assign n43861 = n38112 & ~n41657 ;
  assign n43862 = n43861 ^ n6386 ^ 1'b0 ;
  assign n43863 = n14353 ^ n8886 ^ 1'b0 ;
  assign n43864 = n4045 ^ n3263 ^ n1948 ;
  assign n43865 = n15696 ^ n7277 ^ n1278 ;
  assign n43866 = ( n40011 & n43864 ) | ( n40011 & ~n43865 ) | ( n43864 & ~n43865 ) ;
  assign n43867 = n14365 ^ n5135 ^ 1'b0 ;
  assign n43868 = n887 | n43867 ;
  assign n43869 = ( n1340 & ~n2756 ) | ( n1340 & n5986 ) | ( ~n2756 & n5986 ) ;
  assign n43870 = n43869 ^ n35847 ^ n19812 ;
  assign n43871 = n23213 & ~n43870 ;
  assign n43872 = n27058 & n43871 ;
  assign n43873 = n8835 & ~n43872 ;
  assign n43874 = n28395 ^ n11650 ^ n9067 ;
  assign n43875 = n43874 ^ n23372 ^ n518 ;
  assign n43876 = n37994 & ~n43875 ;
  assign n43877 = n43876 ^ n9160 ^ 1'b0 ;
  assign n43878 = n22882 ^ n17564 ^ n7520 ;
  assign n43879 = n7596 & n43878 ;
  assign n43882 = n19027 ^ n18259 ^ n2433 ;
  assign n43880 = ( n7057 & n18154 ) | ( n7057 & ~n34624 ) | ( n18154 & ~n34624 ) ;
  assign n43881 = n43880 ^ n28924 ^ 1'b0 ;
  assign n43883 = n43882 ^ n43881 ^ 1'b0 ;
  assign n43884 = n18148 ^ n13053 ^ n1015 ;
  assign n43885 = ( n6027 & n21379 ) | ( n6027 & ~n43884 ) | ( n21379 & ~n43884 ) ;
  assign n43888 = n30226 ^ n17015 ^ n1052 ;
  assign n43889 = n43888 ^ n33898 ^ n3174 ;
  assign n43886 = n20508 ^ n18358 ^ n2629 ;
  assign n43887 = n43886 ^ n2315 ^ 1'b0 ;
  assign n43890 = n43889 ^ n43887 ^ n37987 ;
  assign n43891 = n11777 & n14800 ;
  assign n43894 = n946 | n35756 ;
  assign n43892 = n2771 | n12377 ;
  assign n43893 = n43892 ^ n6891 ^ 1'b0 ;
  assign n43895 = n43894 ^ n43893 ^ n37602 ;
  assign n43896 = ( n19829 & n21924 ) | ( n19829 & ~n26548 ) | ( n21924 & ~n26548 ) ;
  assign n43897 = n2964 | n28257 ;
  assign n43898 = n43896 & ~n43897 ;
  assign n43899 = n43760 ^ n22031 ^ 1'b0 ;
  assign n43900 = ( n7906 & n29196 ) | ( n7906 & n29814 ) | ( n29196 & n29814 ) ;
  assign n43901 = ( n13219 & n16483 ) | ( n13219 & n28582 ) | ( n16483 & n28582 ) ;
  assign n43902 = n30982 ^ n30707 ^ 1'b0 ;
  assign n43903 = n42364 ^ n32896 ^ n29884 ;
  assign n43904 = ( ~n9072 & n24289 ) | ( ~n9072 & n43501 ) | ( n24289 & n43501 ) ;
  assign n43905 = n37903 ^ n17358 ^ n15560 ;
  assign n43906 = ( n11606 & n31013 ) | ( n11606 & ~n43905 ) | ( n31013 & ~n43905 ) ;
  assign n43907 = n40964 ^ n21656 ^ 1'b0 ;
  assign n43908 = n13351 & n43907 ;
  assign n43911 = n4966 & ~n15332 ;
  assign n43912 = n43911 ^ n22943 ^ 1'b0 ;
  assign n43909 = ~n9046 & n13857 ;
  assign n43910 = n7690 & n43909 ;
  assign n43913 = n43912 ^ n43910 ^ n19096 ;
  assign n43914 = n43146 ^ n20034 ^ n12323 ;
  assign n43915 = n42212 ^ n12162 ^ 1'b0 ;
  assign n43916 = ~n7057 & n43915 ;
  assign n43917 = ( n12574 & n25473 ) | ( n12574 & n31982 ) | ( n25473 & n31982 ) ;
  assign n43918 = n43917 ^ n37667 ^ 1'b0 ;
  assign n43919 = n4613 & ~n18064 ;
  assign n43920 = ~n43918 & n43919 ;
  assign n43921 = n898 | n2393 ;
  assign n43922 = n43921 ^ n28008 ^ 1'b0 ;
  assign n43923 = n43922 ^ n42288 ^ n37637 ;
  assign n43924 = ( n739 & n1995 ) | ( n739 & n17807 ) | ( n1995 & n17807 ) ;
  assign n43925 = ( ~n24422 & n32726 ) | ( ~n24422 & n43924 ) | ( n32726 & n43924 ) ;
  assign n43926 = ~n453 & n23813 ;
  assign n43927 = ( n20272 & n30872 ) | ( n20272 & ~n43926 ) | ( n30872 & ~n43926 ) ;
  assign n43928 = ( n8382 & n21557 ) | ( n8382 & n30711 ) | ( n21557 & n30711 ) ;
  assign n43929 = n10712 ^ n3502 ^ 1'b0 ;
  assign n43930 = n10792 & n43929 ;
  assign n43931 = n19402 ^ n12377 ^ n298 ;
  assign n43932 = ~n8664 & n43931 ;
  assign n43933 = n28397 & ~n43932 ;
  assign n43934 = ( ~n7676 & n8561 ) | ( ~n7676 & n26158 ) | ( n8561 & n26158 ) ;
  assign n43935 = n43581 ^ n17781 ^ n586 ;
  assign n43936 = n40055 ^ n36857 ^ 1'b0 ;
  assign n43937 = n19268 ^ n17430 ^ n7638 ;
  assign n43938 = ( n10314 & n19446 ) | ( n10314 & ~n43937 ) | ( n19446 & ~n43937 ) ;
  assign n43939 = ~n19912 & n23093 ;
  assign n43944 = n23729 ^ n7577 ^ n5712 ;
  assign n43945 = n43944 ^ n32302 ^ n1854 ;
  assign n43942 = n20529 ^ n1818 ^ 1'b0 ;
  assign n43943 = n8331 & n43942 ;
  assign n43940 = n18829 ^ n4727 ^ 1'b0 ;
  assign n43941 = n24371 | n43940 ;
  assign n43946 = n43945 ^ n43943 ^ n43941 ;
  assign n43947 = n29308 ^ n27224 ^ 1'b0 ;
  assign n43948 = n43947 ^ n32276 ^ n25855 ;
  assign n43949 = n34408 ^ n26871 ^ n12680 ;
  assign n43950 = n38580 ^ n23827 ^ n13458 ;
  assign n43951 = ( n7223 & ~n10415 ) | ( n7223 & n15561 ) | ( ~n10415 & n15561 ) ;
  assign n43952 = n3273 & ~n43951 ;
  assign n43953 = n43952 ^ n27552 ^ 1'b0 ;
  assign n43954 = ( ~n14022 & n32227 ) | ( ~n14022 & n43953 ) | ( n32227 & n43953 ) ;
  assign n43955 = n16665 ^ n11559 ^ 1'b0 ;
  assign n43957 = n27475 | n40005 ;
  assign n43958 = n43957 ^ n8104 ^ 1'b0 ;
  assign n43959 = n11154 & ~n43958 ;
  assign n43960 = n43552 & n43959 ;
  assign n43956 = ( n690 & ~n21261 ) | ( n690 & n32891 ) | ( ~n21261 & n32891 ) ;
  assign n43961 = n43960 ^ n43956 ^ 1'b0 ;
  assign n43962 = n30177 & ~n43379 ;
  assign n43963 = ~n7650 & n43962 ;
  assign n43964 = n43963 ^ n39144 ^ 1'b0 ;
  assign n43965 = n37591 ^ n35984 ^ 1'b0 ;
  assign n43966 = ( ~n29605 & n33043 ) | ( ~n29605 & n36346 ) | ( n33043 & n36346 ) ;
  assign n43967 = n30378 ^ n26571 ^ n10150 ;
  assign n43968 = n13414 ^ n3039 ^ 1'b0 ;
  assign n43969 = n43967 & n43968 ;
  assign n43970 = n39169 & ~n43969 ;
  assign n43971 = ( ~x184 & n26412 ) | ( ~x184 & n43970 ) | ( n26412 & n43970 ) ;
  assign n43972 = ( n7703 & n16746 ) | ( n7703 & n17922 ) | ( n16746 & n17922 ) ;
  assign n43973 = ~n10370 & n43972 ;
  assign n43974 = n43973 ^ n31998 ^ 1'b0 ;
  assign n43975 = n43974 ^ n15062 ^ n13694 ;
  assign n43976 = ~n14151 & n21896 ;
  assign n43977 = n3992 | n11897 ;
  assign n43978 = n43977 ^ n14449 ^ 1'b0 ;
  assign n43979 = n39742 ^ n3856 ^ 1'b0 ;
  assign n43980 = n43978 & ~n43979 ;
  assign n43981 = ( n23912 & ~n43976 ) | ( n23912 & n43980 ) | ( ~n43976 & n43980 ) ;
  assign n43982 = n43981 ^ n41325 ^ 1'b0 ;
  assign n43983 = ~n10116 & n43982 ;
  assign n43984 = n15938 ^ n14770 ^ 1'b0 ;
  assign n43985 = ~n40694 & n43984 ;
  assign n43986 = n30447 ^ n22959 ^ 1'b0 ;
  assign n43987 = ~n15245 & n43986 ;
  assign n43988 = n43987 ^ n6058 ^ 1'b0 ;
  assign n43989 = ~n19017 & n43988 ;
  assign n43990 = n43989 ^ n32483 ^ 1'b0 ;
  assign n43991 = n14673 | n43990 ;
  assign n43992 = n12340 ^ n7642 ^ n3637 ;
  assign n43993 = n392 & ~n6196 ;
  assign n43994 = n43992 & n43993 ;
  assign n43995 = ( n947 & n5974 ) | ( n947 & n43994 ) | ( n5974 & n43994 ) ;
  assign n43996 = n9397 & n34952 ;
  assign n43997 = n43996 ^ n43573 ^ n30522 ;
  assign n43998 = n9489 & n36161 ;
  assign n43999 = n43998 ^ n24142 ^ 1'b0 ;
  assign n44000 = n24186 ^ n23353 ^ n10538 ;
  assign n44001 = n16391 | n35513 ;
  assign n44002 = n44001 ^ n35550 ^ 1'b0 ;
  assign n44003 = n3582 & n41891 ;
  assign n44004 = n10169 & n44003 ;
  assign n44005 = n8909 & ~n14740 ;
  assign n44006 = n44005 ^ n13240 ^ n8079 ;
  assign n44007 = n9338 & ~n41836 ;
  assign n44008 = n8008 & n44007 ;
  assign n44009 = n16007 & ~n44008 ;
  assign n44010 = n44009 ^ n18807 ^ n16001 ;
  assign n44011 = n16884 | n44010 ;
  assign n44012 = n44006 & ~n44011 ;
  assign n44013 = n24374 ^ n16341 ^ 1'b0 ;
  assign n44014 = n44013 ^ n34930 ^ n6685 ;
  assign n44015 = ~n19480 & n44014 ;
  assign n44016 = n4032 ^ n2464 ^ 1'b0 ;
  assign n44017 = n22012 & ~n32322 ;
  assign n44018 = ~n15020 & n44017 ;
  assign n44019 = ( n29269 & ~n35946 ) | ( n29269 & n44018 ) | ( ~n35946 & n44018 ) ;
  assign n44020 = n39733 ^ n10602 ^ n8428 ;
  assign n44021 = n18744 & n24845 ;
  assign n44022 = ( n12135 & n36079 ) | ( n12135 & n44021 ) | ( n36079 & n44021 ) ;
  assign n44023 = ( n15494 & n22173 ) | ( n15494 & ~n26793 ) | ( n22173 & ~n26793 ) ;
  assign n44024 = ~n14844 & n41357 ;
  assign n44025 = n15217 & n44024 ;
  assign n44026 = ( n8000 & ~n8095 ) | ( n8000 & n33284 ) | ( ~n8095 & n33284 ) ;
  assign n44027 = n1929 | n44026 ;
  assign n44028 = ( n44023 & n44025 ) | ( n44023 & n44027 ) | ( n44025 & n44027 ) ;
  assign n44029 = ( n3783 & n10480 ) | ( n3783 & n29270 ) | ( n10480 & n29270 ) ;
  assign n44030 = n44029 ^ n28225 ^ n19496 ;
  assign n44031 = n44030 ^ n10739 ^ 1'b0 ;
  assign n44032 = n12108 & ~n39156 ;
  assign n44033 = n44031 & n44032 ;
  assign n44034 = n13606 & n16101 ;
  assign n44035 = ~n31225 & n44034 ;
  assign n44036 = ( n3743 & n15707 ) | ( n3743 & ~n42447 ) | ( n15707 & ~n42447 ) ;
  assign n44037 = ( n6921 & ~n10330 ) | ( n6921 & n39919 ) | ( ~n10330 & n39919 ) ;
  assign n44038 = n9171 & n44037 ;
  assign n44039 = ~n30377 & n44038 ;
  assign n44040 = n44039 ^ n10497 ^ n509 ;
  assign n44041 = n24553 ^ n6018 ^ 1'b0 ;
  assign n44042 = n40140 ^ n25890 ^ 1'b0 ;
  assign n44043 = n44042 ^ n12449 ^ n9264 ;
  assign n44050 = n43880 ^ n30111 ^ n20613 ;
  assign n44051 = n44050 ^ n2597 ^ 1'b0 ;
  assign n44045 = ~n13168 & n42789 ;
  assign n44044 = n19739 ^ n3141 ^ 1'b0 ;
  assign n44046 = n44045 ^ n44044 ^ n29563 ;
  assign n44047 = n37024 ^ n18068 ^ 1'b0 ;
  assign n44048 = n44046 & ~n44047 ;
  assign n44049 = n10019 & n44048 ;
  assign n44052 = n44051 ^ n44049 ^ 1'b0 ;
  assign n44054 = ( n11001 & ~n23896 ) | ( n11001 & n25185 ) | ( ~n23896 & n25185 ) ;
  assign n44053 = n12912 | n43016 ;
  assign n44055 = n44054 ^ n44053 ^ 1'b0 ;
  assign n44056 = ( ~n10755 & n12515 ) | ( ~n10755 & n42387 ) | ( n12515 & n42387 ) ;
  assign n44057 = ( ~n20802 & n29244 ) | ( ~n20802 & n34496 ) | ( n29244 & n34496 ) ;
  assign n44058 = ( n11607 & n19238 ) | ( n11607 & ~n21907 ) | ( n19238 & ~n21907 ) ;
  assign n44059 = n44058 ^ n15886 ^ 1'b0 ;
  assign n44060 = ( n30682 & n42979 ) | ( n30682 & n44059 ) | ( n42979 & n44059 ) ;
  assign n44061 = n29042 ^ n27079 ^ n24213 ;
  assign n44062 = n44061 ^ n20442 ^ n2669 ;
  assign n44063 = ( ~n10651 & n21740 ) | ( ~n10651 & n39234 ) | ( n21740 & n39234 ) ;
  assign n44064 = n21562 & ~n44063 ;
  assign n44065 = ~n20956 & n44064 ;
  assign n44066 = n44065 ^ n30147 ^ n22348 ;
  assign n44067 = n14968 ^ n14074 ^ 1'b0 ;
  assign n44068 = ~n1340 & n44067 ;
  assign n44069 = n1909 & n9017 ;
  assign n44070 = ( ~n1003 & n33480 ) | ( ~n1003 & n44069 ) | ( n33480 & n44069 ) ;
  assign n44071 = ( n25622 & ~n44068 ) | ( n25622 & n44070 ) | ( ~n44068 & n44070 ) ;
  assign n44072 = n27912 & n40512 ;
  assign n44073 = n16521 & ~n27154 ;
  assign n44074 = n44073 ^ n40574 ^ n17369 ;
  assign n44075 = n44074 ^ n16726 ^ 1'b0 ;
  assign n44076 = ~n44072 & n44075 ;
  assign n44077 = n14534 ^ n2908 ^ 1'b0 ;
  assign n44078 = n13399 | n44077 ;
  assign n44079 = n44078 ^ n15501 ^ n14205 ;
  assign n44080 = n44079 ^ n12623 ^ 1'b0 ;
  assign n44081 = n8033 & ~n30463 ;
  assign n44082 = n44081 ^ n1281 ^ 1'b0 ;
  assign n44083 = n32854 | n38247 ;
  assign n44084 = n3687 | n44083 ;
  assign n44085 = n4510 & ~n34914 ;
  assign n44086 = ( n22696 & ~n27201 ) | ( n22696 & n44085 ) | ( ~n27201 & n44085 ) ;
  assign n44087 = n8919 ^ n8576 ^ 1'b0 ;
  assign n44088 = n34535 ^ n9951 ^ n1859 ;
  assign n44089 = ~n16286 & n32111 ;
  assign n44090 = ( ~n17548 & n19314 ) | ( ~n17548 & n40670 ) | ( n19314 & n40670 ) ;
  assign n44091 = n26722 & n44090 ;
  assign n44092 = n44091 ^ n5952 ^ 1'b0 ;
  assign n44094 = ~n8152 & n33096 ;
  assign n44095 = n44094 ^ n13909 ^ n3945 ;
  assign n44096 = n44095 ^ n40881 ^ 1'b0 ;
  assign n44093 = ~n697 & n28854 ;
  assign n44097 = n44096 ^ n44093 ^ 1'b0 ;
  assign n44098 = n9238 ^ n4192 ^ n356 ;
  assign n44099 = n27061 ^ n22439 ^ 1'b0 ;
  assign n44100 = n11322 | n44099 ;
  assign n44101 = ( n28936 & n44098 ) | ( n28936 & ~n44100 ) | ( n44098 & ~n44100 ) ;
  assign n44102 = n43627 ^ n14868 ^ 1'b0 ;
  assign n44103 = n4475 & ~n36194 ;
  assign n44104 = n21800 & n37727 ;
  assign n44105 = n22928 & n44104 ;
  assign n44106 = n38714 ^ n29332 ^ n20141 ;
  assign n44107 = n37938 ^ n18910 ^ 1'b0 ;
  assign n44108 = n31157 & n44107 ;
  assign n44109 = n44108 ^ n33573 ^ n31788 ;
  assign n44110 = n20656 ^ n2857 ^ 1'b0 ;
  assign n44111 = n19038 & n31833 ;
  assign n44112 = ~n2085 & n44111 ;
  assign n44113 = ( n9955 & ~n18375 ) | ( n9955 & n44112 ) | ( ~n18375 & n44112 ) ;
  assign n44114 = n14281 | n14775 ;
  assign n44115 = ~n7565 & n15409 ;
  assign n44116 = n35709 & n39214 ;
  assign n44117 = n44115 & n44116 ;
  assign n44118 = n1896 | n4334 ;
  assign n44119 = n39754 ^ n13543 ^ 1'b0 ;
  assign n44120 = n44119 ^ n22854 ^ n17983 ;
  assign n44121 = n44120 ^ n802 ^ 1'b0 ;
  assign n44122 = n21694 & n44121 ;
  assign n44123 = n22546 ^ n8980 ^ n2199 ;
  assign n44124 = ( ~n11950 & n35855 ) | ( ~n11950 & n44123 ) | ( n35855 & n44123 ) ;
  assign n44125 = ( n2008 & n27224 ) | ( n2008 & n41440 ) | ( n27224 & n41440 ) ;
  assign n44126 = n39983 ^ n1246 ^ 1'b0 ;
  assign n44127 = n44126 ^ n30276 ^ n19804 ;
  assign n44128 = n38851 ^ n19460 ^ 1'b0 ;
  assign n44129 = n21533 | n44128 ;
  assign n44130 = ( n44125 & ~n44127 ) | ( n44125 & n44129 ) | ( ~n44127 & n44129 ) ;
  assign n44131 = ( n11436 & ~n30565 ) | ( n11436 & n36189 ) | ( ~n30565 & n36189 ) ;
  assign n44132 = ( n18105 & ~n43333 ) | ( n18105 & n44131 ) | ( ~n43333 & n44131 ) ;
  assign n44133 = n3355 & n4363 ;
  assign n44134 = n40819 & n44133 ;
  assign n44135 = n44134 ^ n13137 ^ n6767 ;
  assign n44136 = n24875 ^ n3235 ^ n669 ;
  assign n44137 = n5401 & n8268 ;
  assign n44138 = n11601 | n35932 ;
  assign n44139 = n11231 | n44138 ;
  assign n44140 = n44139 ^ n40328 ^ 1'b0 ;
  assign n44141 = n20695 & ~n44140 ;
  assign n44142 = n6930 ^ n305 ^ 1'b0 ;
  assign n44148 = n2968 & ~n9796 ;
  assign n44149 = n44148 ^ n32579 ^ 1'b0 ;
  assign n44144 = n18658 ^ n10508 ^ 1'b0 ;
  assign n44145 = n44144 ^ n4764 ^ 1'b0 ;
  assign n44146 = n7226 | n44145 ;
  assign n44143 = n39310 ^ n16654 ^ n15697 ;
  assign n44147 = n44146 ^ n44143 ^ n1507 ;
  assign n44150 = n44149 ^ n44147 ^ 1'b0 ;
  assign n44151 = n868 & n22208 ;
  assign n44152 = n44151 ^ n36341 ^ 1'b0 ;
  assign n44153 = ( n3495 & ~n8500 ) | ( n3495 & n44152 ) | ( ~n8500 & n44152 ) ;
  assign n44154 = n26695 ^ n23737 ^ 1'b0 ;
  assign n44155 = n10114 | n24107 ;
  assign n44156 = n33957 | n44155 ;
  assign n44157 = ~n37937 & n44156 ;
  assign n44158 = ( n2970 & ~n5333 ) | ( n2970 & n44157 ) | ( ~n5333 & n44157 ) ;
  assign n44159 = ( n5573 & ~n7630 ) | ( n5573 & n7887 ) | ( ~n7630 & n7887 ) ;
  assign n44160 = n44159 ^ n24207 ^ n16548 ;
  assign n44161 = ~n13513 & n44160 ;
  assign n44162 = n2784 | n33519 ;
  assign n44163 = n27727 & ~n44162 ;
  assign n44164 = n14998 | n18779 ;
  assign n44165 = ~n7947 & n10241 ;
  assign n44166 = ( ~n1626 & n6781 ) | ( ~n1626 & n27659 ) | ( n6781 & n27659 ) ;
  assign n44168 = n40607 ^ n3221 ^ n2608 ;
  assign n44167 = ~n4333 & n9643 ;
  assign n44169 = n44168 ^ n44167 ^ n30266 ;
  assign n44170 = n5222 & ~n5670 ;
  assign n44171 = ~n8558 & n44170 ;
  assign n44172 = n44171 ^ n9721 ^ 1'b0 ;
  assign n44173 = n44172 ^ n35840 ^ n10353 ;
  assign n44174 = ( n1545 & n24428 ) | ( n1545 & n44173 ) | ( n24428 & n44173 ) ;
  assign n44175 = ( n3794 & ~n15250 ) | ( n3794 & n26257 ) | ( ~n15250 & n26257 ) ;
  assign n44176 = ( ~n16942 & n27138 ) | ( ~n16942 & n34627 ) | ( n27138 & n34627 ) ;
  assign n44177 = n301 & ~n10781 ;
  assign n44178 = n44176 & n44177 ;
  assign n44179 = n36453 | n40467 ;
  assign n44180 = x7 & ~n781 ;
  assign n44181 = n26074 & n44180 ;
  assign n44182 = n27575 ^ n18586 ^ n11973 ;
  assign n44183 = ~n5931 & n44182 ;
  assign n44184 = n44183 ^ n14967 ^ 1'b0 ;
  assign n44185 = n4043 & ~n28684 ;
  assign n44186 = ~x76 & n44185 ;
  assign n44187 = n14183 & ~n29401 ;
  assign n44188 = n44187 ^ n28002 ^ 1'b0 ;
  assign n44189 = ( n33449 & n44186 ) | ( n33449 & n44188 ) | ( n44186 & n44188 ) ;
  assign n44190 = ( ~n25681 & n31698 ) | ( ~n25681 & n34157 ) | ( n31698 & n34157 ) ;
  assign n44191 = ( ~n6360 & n17767 ) | ( ~n6360 & n37709 ) | ( n17767 & n37709 ) ;
  assign n44193 = n3371 | n7282 ;
  assign n44194 = n44193 ^ n20343 ^ 1'b0 ;
  assign n44195 = n4926 & n44194 ;
  assign n44196 = n44195 ^ n28912 ^ 1'b0 ;
  assign n44192 = n1895 | n9283 ;
  assign n44197 = n44196 ^ n44192 ^ n39861 ;
  assign n44198 = n6021 | n44197 ;
  assign n44199 = ( n25516 & n27353 ) | ( n25516 & n43544 ) | ( n27353 & n43544 ) ;
  assign n44200 = n44199 ^ n19549 ^ 1'b0 ;
  assign n44201 = ~n22884 & n44200 ;
  assign n44202 = n31330 ^ n10896 ^ n9349 ;
  assign n44203 = n44201 & n44202 ;
  assign n44204 = n12466 & ~n37155 ;
  assign n44205 = n14299 | n27872 ;
  assign n44206 = n44205 ^ n4451 ^ 1'b0 ;
  assign n44207 = n44206 ^ n41237 ^ x117 ;
  assign n44208 = ( ~n28189 & n43595 ) | ( ~n28189 & n44207 ) | ( n43595 & n44207 ) ;
  assign n44209 = n41004 ^ n5883 ^ n1909 ;
  assign n44210 = n33534 ^ n14607 ^ 1'b0 ;
  assign n44211 = n1904 & n44210 ;
  assign n44212 = n44211 ^ n35350 ^ n2600 ;
  assign n44213 = n23744 ^ n11240 ^ n7369 ;
  assign n44214 = n44213 ^ n22133 ^ n791 ;
  assign n44215 = n44214 ^ n12494 ^ n917 ;
  assign n44216 = ( n28234 & n31474 ) | ( n28234 & n44215 ) | ( n31474 & n44215 ) ;
  assign n44217 = ( n7019 & n21507 ) | ( n7019 & ~n21957 ) | ( n21507 & ~n21957 ) ;
  assign n44218 = n1854 & ~n35059 ;
  assign n44219 = n44218 ^ n31952 ^ 1'b0 ;
  assign n44220 = n11382 | n12979 ;
  assign n44221 = n11641 | n44220 ;
  assign n44222 = n3371 | n23849 ;
  assign n44223 = n1438 | n2684 ;
  assign n44224 = n44223 ^ n23152 ^ 1'b0 ;
  assign n44225 = n40064 ^ n7792 ^ 1'b0 ;
  assign n44226 = ~n44224 & n44225 ;
  assign n44227 = ~n14757 & n44226 ;
  assign n44228 = n22221 & n44227 ;
  assign n44230 = ( n5355 & n10196 ) | ( n5355 & ~n17256 ) | ( n10196 & ~n17256 ) ;
  assign n44229 = n21805 | n36731 ;
  assign n44231 = n44230 ^ n44229 ^ 1'b0 ;
  assign n44232 = ( n13432 & ~n20212 ) | ( n13432 & n44231 ) | ( ~n20212 & n44231 ) ;
  assign n44233 = n30540 ^ n5542 ^ n3366 ;
  assign n44234 = n25573 & n44233 ;
  assign n44235 = n26185 ^ n24423 ^ 1'b0 ;
  assign n44240 = n8196 & n10368 ;
  assign n44238 = n6078 & n27046 ;
  assign n44239 = n44238 ^ n35491 ^ 1'b0 ;
  assign n44236 = n41192 ^ n14216 ^ 1'b0 ;
  assign n44237 = ( n29647 & ~n42534 ) | ( n29647 & n44236 ) | ( ~n42534 & n44236 ) ;
  assign n44241 = n44240 ^ n44239 ^ n44237 ;
  assign n44242 = n22421 ^ n2110 ^ 1'b0 ;
  assign n44243 = n11429 & n44242 ;
  assign n44244 = n44243 ^ n21312 ^ n540 ;
  assign n44245 = n9338 | n29502 ;
  assign n44246 = ( n11685 & n25318 ) | ( n11685 & ~n44245 ) | ( n25318 & ~n44245 ) ;
  assign n44247 = n33575 ^ n18784 ^ 1'b0 ;
  assign n44248 = n3017 & n38903 ;
  assign n44249 = ~n44247 & n44248 ;
  assign n44250 = n1507 & n19518 ;
  assign n44251 = n19499 ^ n16545 ^ 1'b0 ;
  assign n44252 = n20762 & ~n44251 ;
  assign n44253 = n22310 ^ n4175 ^ 1'b0 ;
  assign n44254 = n20596 & ~n44253 ;
  assign n44255 = n13670 ^ n12244 ^ 1'b0 ;
  assign n44256 = n2440 & n44255 ;
  assign n44257 = n28694 & n44256 ;
  assign n44258 = ( n4395 & ~n6109 ) | ( n4395 & n10391 ) | ( ~n6109 & n10391 ) ;
  assign n44260 = n41777 ^ n5320 ^ 1'b0 ;
  assign n44261 = n11933 | n44260 ;
  assign n44259 = n36880 ^ n24591 ^ n19583 ;
  assign n44262 = n44261 ^ n44259 ^ n1566 ;
  assign n44263 = n7221 | n12729 ;
  assign n44264 = n24913 ^ n15932 ^ 1'b0 ;
  assign n44265 = n28194 & n44264 ;
  assign n44266 = ~n44263 & n44265 ;
  assign n44267 = ~n11153 & n24709 ;
  assign n44268 = n15282 | n31477 ;
  assign n44269 = n6355 & n44268 ;
  assign n44270 = ~n28198 & n44269 ;
  assign n44271 = n28614 ^ n10186 ^ 1'b0 ;
  assign n44272 = n24280 | n44271 ;
  assign n44273 = n4995 | n44272 ;
  assign n44274 = n44273 ^ n43737 ^ 1'b0 ;
  assign n44275 = ( n8190 & ~n13070 ) | ( n8190 & n27322 ) | ( ~n13070 & n27322 ) ;
  assign n44277 = n1747 | n2053 ;
  assign n44278 = n44277 ^ n10918 ^ 1'b0 ;
  assign n44276 = n21169 ^ n20415 ^ 1'b0 ;
  assign n44279 = n44278 ^ n44276 ^ n3636 ;
  assign n44280 = n2318 & ~n26888 ;
  assign n44281 = n2857 & n44280 ;
  assign n44282 = n44281 ^ n38906 ^ n28819 ;
  assign n44283 = n32118 ^ n31161 ^ 1'b0 ;
  assign n44284 = ( n624 & n1481 ) | ( n624 & ~n42940 ) | ( n1481 & ~n42940 ) ;
  assign n44285 = n7465 & n44284 ;
  assign n44286 = ( n3555 & n44283 ) | ( n3555 & ~n44285 ) | ( n44283 & ~n44285 ) ;
  assign n44289 = ( ~n5253 & n29308 ) | ( ~n5253 & n29775 ) | ( n29308 & n29775 ) ;
  assign n44287 = ( n12765 & n24338 ) | ( n12765 & n29247 ) | ( n24338 & n29247 ) ;
  assign n44288 = n40160 & n44287 ;
  assign n44290 = n44289 ^ n44288 ^ 1'b0 ;
  assign n44291 = n27092 ^ n20010 ^ n3130 ;
  assign n44292 = n33095 ^ n14399 ^ 1'b0 ;
  assign n44293 = ~n6714 & n15131 ;
  assign n44294 = ( n5159 & ~n35508 ) | ( n5159 & n44293 ) | ( ~n35508 & n44293 ) ;
  assign n44295 = n5693 | n16970 ;
  assign n44296 = n14587 ^ n13287 ^ n4892 ;
  assign n44297 = n8678 & n15546 ;
  assign n44298 = ~n8130 & n12502 ;
  assign n44299 = n32427 & n44298 ;
  assign n44301 = n10373 ^ n1705 ^ 1'b0 ;
  assign n44302 = n3684 | n44301 ;
  assign n44303 = n14841 & ~n44302 ;
  assign n44300 = n6023 | n24462 ;
  assign n44304 = n44303 ^ n44300 ^ 1'b0 ;
  assign n44305 = n44304 ^ n27371 ^ n13330 ;
  assign n44306 = n789 | n13859 ;
  assign n44307 = n44306 ^ n1154 ^ 1'b0 ;
  assign n44308 = ( ~n18594 & n19379 ) | ( ~n18594 & n44307 ) | ( n19379 & n44307 ) ;
  assign n44309 = n41006 ^ n21507 ^ n10619 ;
  assign n44310 = n44309 ^ n43969 ^ n22633 ;
  assign n44311 = n975 | n11685 ;
  assign n44312 = n44311 ^ n31524 ^ 1'b0 ;
  assign n44313 = n6328 & n43779 ;
  assign n44314 = n4227 & n44313 ;
  assign n44315 = n21952 ^ n19348 ^ 1'b0 ;
  assign n44316 = n5166 & ~n44315 ;
  assign n44317 = n34206 & n44316 ;
  assign n44318 = n44317 ^ n33877 ^ 1'b0 ;
  assign n44319 = n7528 & ~n38872 ;
  assign n44320 = n44319 ^ n4759 ^ 1'b0 ;
  assign n44322 = ~n10036 & n11242 ;
  assign n44323 = n44322 ^ x230 ^ 1'b0 ;
  assign n44321 = n17073 ^ n10235 ^ n3527 ;
  assign n44324 = n44323 ^ n44321 ^ n33272 ;
  assign n44325 = ( n29765 & ~n35768 ) | ( n29765 & n39970 ) | ( ~n35768 & n39970 ) ;
  assign n44326 = ( ~n7019 & n8229 ) | ( ~n7019 & n9192 ) | ( n8229 & n9192 ) ;
  assign n44327 = n5518 & ~n9327 ;
  assign n44328 = n44327 ^ n33809 ^ 1'b0 ;
  assign n44329 = n3873 & n44328 ;
  assign n44330 = ~n28413 & n44329 ;
  assign n44331 = ( ~n7456 & n16055 ) | ( ~n7456 & n28842 ) | ( n16055 & n28842 ) ;
  assign n44332 = n23035 ^ n22914 ^ 1'b0 ;
  assign n44333 = n15255 | n44332 ;
  assign n44334 = n44333 ^ n28315 ^ n22629 ;
  assign n44336 = ( x145 & ~n1015 ) | ( x145 & n12612 ) | ( ~n1015 & n12612 ) ;
  assign n44335 = n9924 & ~n33898 ;
  assign n44337 = n44336 ^ n44335 ^ n24510 ;
  assign n44338 = ~x201 & n13490 ;
  assign n44339 = n17391 ^ n13656 ^ 1'b0 ;
  assign n44340 = ( n2701 & n14838 ) | ( n2701 & n28834 ) | ( n14838 & n28834 ) ;
  assign n44341 = ( n8557 & ~n44339 ) | ( n8557 & n44340 ) | ( ~n44339 & n44340 ) ;
  assign n44342 = ( n547 & n29331 ) | ( n547 & n29740 ) | ( n29331 & n29740 ) ;
  assign n44344 = ( n5909 & n12392 ) | ( n5909 & ~n18653 ) | ( n12392 & ~n18653 ) ;
  assign n44345 = n44344 ^ n26637 ^ n8296 ;
  assign n44346 = n30178 ^ n9622 ^ n2196 ;
  assign n44347 = n44346 ^ n4301 ^ 1'b0 ;
  assign n44348 = ( n350 & n44345 ) | ( n350 & n44347 ) | ( n44345 & n44347 ) ;
  assign n44343 = ~n5653 & n27069 ;
  assign n44349 = n44348 ^ n44343 ^ 1'b0 ;
  assign n44350 = n29143 ^ n17821 ^ 1'b0 ;
  assign n44353 = n39584 ^ n2973 ^ 1'b0 ;
  assign n44354 = ( n30185 & ~n39776 ) | ( n30185 & n44353 ) | ( ~n39776 & n44353 ) ;
  assign n44351 = n6681 | n29119 ;
  assign n44352 = n29146 | n44351 ;
  assign n44355 = n44354 ^ n44352 ^ 1'b0 ;
  assign n44356 = ( x188 & ~n12140 ) | ( x188 & n13573 ) | ( ~n12140 & n13573 ) ;
  assign n44357 = n27310 | n32458 ;
  assign n44358 = n44357 ^ n31310 ^ n20445 ;
  assign n44359 = n44358 ^ n7940 ^ 1'b0 ;
  assign n44360 = n27659 ^ n24040 ^ n3568 ;
  assign n44361 = n44360 ^ n38578 ^ n16043 ;
  assign n44362 = ( ~n24374 & n44359 ) | ( ~n24374 & n44361 ) | ( n44359 & n44361 ) ;
  assign n44363 = ( n21778 & n44356 ) | ( n21778 & n44362 ) | ( n44356 & n44362 ) ;
  assign n44364 = n9558 ^ n436 ^ 1'b0 ;
  assign n44365 = ( n2100 & n15745 ) | ( n2100 & n44364 ) | ( n15745 & n44364 ) ;
  assign n44366 = n7181 & ~n20152 ;
  assign n44368 = n31243 ^ n30951 ^ n25604 ;
  assign n44367 = n25618 | n43076 ;
  assign n44369 = n44368 ^ n44367 ^ 1'b0 ;
  assign n44370 = n34686 & ~n44369 ;
  assign n44371 = n44370 ^ n4697 ^ 1'b0 ;
  assign n44372 = n30173 ^ n5683 ^ 1'b0 ;
  assign n44373 = n39139 ^ n7349 ^ 1'b0 ;
  assign n44374 = ( n2292 & ~n37335 ) | ( n2292 & n44373 ) | ( ~n37335 & n44373 ) ;
  assign n44375 = n28920 ^ n19359 ^ n2080 ;
  assign n44376 = n13011 | n44375 ;
  assign n44377 = n13905 | n27475 ;
  assign n44378 = n44377 ^ n44335 ^ 1'b0 ;
  assign n44379 = x97 & ~n32020 ;
  assign n44380 = n44378 & n44379 ;
  assign n44381 = n22302 | n39991 ;
  assign n44382 = n44381 ^ n39172 ^ 1'b0 ;
  assign n44383 = n3430 & ~n23772 ;
  assign n44384 = n14901 & n44383 ;
  assign n44385 = n44384 ^ n32476 ^ 1'b0 ;
  assign n44386 = ( n6592 & n12620 ) | ( n6592 & n22748 ) | ( n12620 & n22748 ) ;
  assign n44387 = n44386 ^ n32353 ^ n2311 ;
  assign n44388 = ~n1598 & n12441 ;
  assign n44389 = ( n4165 & n23517 ) | ( n4165 & ~n44388 ) | ( n23517 & ~n44388 ) ;
  assign n44390 = n30133 ^ n22479 ^ n13739 ;
  assign n44392 = n4449 & n27224 ;
  assign n44393 = n44392 ^ n30077 ^ 1'b0 ;
  assign n44391 = n22698 ^ n4438 ^ 1'b0 ;
  assign n44394 = n44393 ^ n44391 ^ n22031 ;
  assign n44395 = n19262 ^ n17081 ^ n16503 ;
  assign n44396 = n44395 ^ n29975 ^ 1'b0 ;
  assign n44397 = n21446 & ~n44396 ;
  assign n44398 = n30053 ^ n20517 ^ 1'b0 ;
  assign n44399 = n16925 | n44398 ;
  assign n44400 = n19299 & n44399 ;
  assign n44401 = n24108 ^ n8403 ^ 1'b0 ;
  assign n44402 = n44401 ^ n21238 ^ n15955 ;
  assign n44403 = ( n21415 & n34180 ) | ( n21415 & n44402 ) | ( n34180 & n44402 ) ;
  assign n44404 = n33941 ^ n5388 ^ 1'b0 ;
  assign n44405 = n5505 | n44404 ;
  assign n44406 = n44405 ^ n22933 ^ n21393 ;
  assign n44407 = n33409 ^ n10737 ^ n3942 ;
  assign n44408 = n44407 ^ n28917 ^ n24120 ;
  assign n44410 = n7637 & n11487 ;
  assign n44411 = n27721 & n44410 ;
  assign n44409 = ~n18935 & n26227 ;
  assign n44412 = n44411 ^ n44409 ^ 1'b0 ;
  assign n44413 = n44412 ^ n32671 ^ n20932 ;
  assign n44414 = ( n14499 & ~n18035 ) | ( n14499 & n38594 ) | ( ~n18035 & n38594 ) ;
  assign n44415 = n44414 ^ n588 ^ 1'b0 ;
  assign n44416 = n40026 | n44415 ;
  assign n44417 = n29093 ^ n14159 ^ n4693 ;
  assign n44418 = n44417 ^ n20147 ^ n6505 ;
  assign n44419 = n33511 ^ n29849 ^ 1'b0 ;
  assign n44420 = ~n44418 & n44419 ;
  assign n44421 = n905 | n27029 ;
  assign n44422 = n29234 & ~n44421 ;
  assign n44423 = n37817 ^ n27127 ^ n24107 ;
  assign n44424 = ( n21697 & n32867 ) | ( n21697 & ~n44031 ) | ( n32867 & ~n44031 ) ;
  assign n44430 = ~n1681 & n17864 ;
  assign n44431 = n44430 ^ n17258 ^ 1'b0 ;
  assign n44425 = ( x101 & ~n6392 ) | ( x101 & n8607 ) | ( ~n6392 & n8607 ) ;
  assign n44426 = n5013 | n17710 ;
  assign n44427 = n44426 ^ n15856 ^ 1'b0 ;
  assign n44428 = n44425 | n44427 ;
  assign n44429 = n44428 ^ n5097 ^ 1'b0 ;
  assign n44432 = n44431 ^ n44429 ^ 1'b0 ;
  assign n44433 = n19259 & ~n42062 ;
  assign n44434 = ~n9696 & n44433 ;
  assign n44435 = n4266 ^ x126 ^ 1'b0 ;
  assign n44436 = ~n35804 & n44435 ;
  assign n44437 = ( n11685 & ~n15177 ) | ( n11685 & n23624 ) | ( ~n15177 & n23624 ) ;
  assign n44438 = ( ~n14271 & n20395 ) | ( ~n14271 & n44437 ) | ( n20395 & n44437 ) ;
  assign n44439 = n44438 ^ n23373 ^ 1'b0 ;
  assign n44440 = n7268 & ~n21388 ;
  assign n44441 = n23503 ^ n9156 ^ 1'b0 ;
  assign n44442 = n44441 ^ n1305 ^ 1'b0 ;
  assign n44443 = n44442 ^ n40505 ^ 1'b0 ;
  assign n44444 = n40370 ^ n10517 ^ n8904 ;
  assign n44445 = n7453 ^ n2152 ^ 1'b0 ;
  assign n44446 = n12988 | n44445 ;
  assign n44447 = ( n364 & n14077 ) | ( n364 & ~n44446 ) | ( n14077 & ~n44446 ) ;
  assign n44448 = n44447 ^ n17950 ^ 1'b0 ;
  assign n44449 = n6476 & ~n42827 ;
  assign n44450 = n7612 & n34975 ;
  assign n44451 = n23075 & n44450 ;
  assign n44452 = ( n27989 & n38352 ) | ( n27989 & n44451 ) | ( n38352 & n44451 ) ;
  assign n44453 = n15224 ^ n14168 ^ 1'b0 ;
  assign n44454 = n8155 & ~n44453 ;
  assign n44455 = n29763 ^ n2661 ^ 1'b0 ;
  assign n44456 = n13126 | n44455 ;
  assign n44457 = ( n30745 & ~n35134 ) | ( n30745 & n44456 ) | ( ~n35134 & n44456 ) ;
  assign n44458 = ( ~n40492 & n44454 ) | ( ~n40492 & n44457 ) | ( n44454 & n44457 ) ;
  assign n44459 = n12623 ^ n8888 ^ n8756 ;
  assign n44460 = n44459 ^ n25342 ^ 1'b0 ;
  assign n44461 = n27302 ^ n10088 ^ 1'b0 ;
  assign n44462 = n44460 & ~n44461 ;
  assign n44463 = n44462 ^ n1214 ^ 1'b0 ;
  assign n44464 = n20031 ^ n9310 ^ 1'b0 ;
  assign n44465 = n10907 & n44464 ;
  assign n44466 = n20966 | n24497 ;
  assign n44467 = n1336 & ~n44466 ;
  assign n44468 = n24057 ^ n11514 ^ n280 ;
  assign n44469 = n27835 ^ n19028 ^ n7627 ;
  assign n44470 = ( ~n20726 & n27302 ) | ( ~n20726 & n38931 ) | ( n27302 & n38931 ) ;
  assign n44472 = n350 & ~n9575 ;
  assign n44473 = n4044 & n44472 ;
  assign n44471 = n23029 & ~n25459 ;
  assign n44474 = n44473 ^ n44471 ^ n39584 ;
  assign n44475 = n4771 | n10123 ;
  assign n44476 = n4290 & n44475 ;
  assign n44477 = n44476 ^ n5405 ^ 1'b0 ;
  assign n44478 = n15513 ^ n5742 ^ n3762 ;
  assign n44479 = n44478 ^ n27585 ^ 1'b0 ;
  assign n44480 = n14459 | n44479 ;
  assign n44481 = ( n2243 & n6249 ) | ( n2243 & n8174 ) | ( n6249 & n8174 ) ;
  assign n44482 = n21312 | n44481 ;
  assign n44483 = n12114 ^ n6317 ^ n2315 ;
  assign n44484 = n1431 ^ n1037 ^ 1'b0 ;
  assign n44485 = n44484 ^ n28047 ^ n11245 ;
  assign n44486 = n12222 & n37124 ;
  assign n44487 = ( n1385 & n13131 ) | ( n1385 & ~n23364 ) | ( n13131 & ~n23364 ) ;
  assign n44488 = n44487 ^ n16156 ^ 1'b0 ;
  assign n44489 = n34716 ^ n26812 ^ 1'b0 ;
  assign n44490 = n39959 ^ n15154 ^ n12451 ;
  assign n44491 = ( n2012 & ~n3730 ) | ( n2012 & n8792 ) | ( ~n3730 & n8792 ) ;
  assign n44492 = n44491 ^ n2928 ^ 1'b0 ;
  assign n44493 = n44490 & ~n44492 ;
  assign n44496 = n8438 ^ n943 ^ 1'b0 ;
  assign n44497 = n9869 & n44496 ;
  assign n44494 = ~n8222 & n21698 ;
  assign n44495 = n44494 ^ n31618 ^ 1'b0 ;
  assign n44498 = n44497 ^ n44495 ^ n2094 ;
  assign n44499 = n13059 | n44498 ;
  assign n44500 = n44499 ^ n18621 ^ 1'b0 ;
  assign n44501 = n9076 & ~n44500 ;
  assign n44502 = n39331 ^ n32044 ^ n4169 ;
  assign n44503 = n38652 ^ n35612 ^ n25881 ;
  assign n44504 = ~n2728 & n44503 ;
  assign n44505 = n2922 & ~n30170 ;
  assign n44506 = n44505 ^ n12540 ^ n4848 ;
  assign n44507 = n27658 & ~n34943 ;
  assign n44508 = n9427 & n44507 ;
  assign n44509 = ~n20062 & n34046 ;
  assign n44510 = n24659 & n44509 ;
  assign n44511 = ~n19620 & n44510 ;
  assign n44512 = n8863 | n44511 ;
  assign n44513 = n12229 | n12371 ;
  assign n44514 = n44513 ^ n43956 ^ 1'b0 ;
  assign n44515 = n21079 ^ n2080 ^ 1'b0 ;
  assign n44516 = n1439 & ~n44515 ;
  assign n44517 = n26996 ^ n9691 ^ n6711 ;
  assign n44518 = n32574 ^ n19652 ^ n14645 ;
  assign n44519 = n44176 ^ n21475 ^ n9286 ;
  assign n44520 = n3263 & n28310 ;
  assign n44521 = ~n17101 & n44520 ;
  assign n44522 = n44521 ^ n16715 ^ n2950 ;
  assign n44523 = ( ~n11949 & n12737 ) | ( ~n11949 & n22815 ) | ( n12737 & n22815 ) ;
  assign n44525 = n5056 | n21303 ;
  assign n44524 = n1960 & ~n22601 ;
  assign n44526 = n44525 ^ n44524 ^ 1'b0 ;
  assign n44527 = ( n7627 & n8958 ) | ( n7627 & n13121 ) | ( n8958 & n13121 ) ;
  assign n44528 = n44527 ^ n7609 ^ n3471 ;
  assign n44529 = n13788 | n44528 ;
  assign n44530 = ( n10297 & ~n15615 ) | ( n10297 & n44529 ) | ( ~n15615 & n44529 ) ;
  assign n44531 = ~n37050 & n44530 ;
  assign n44532 = n4743 | n26057 ;
  assign n44534 = n18868 ^ n4553 ^ 1'b0 ;
  assign n44533 = ( ~n6548 & n17155 ) | ( ~n6548 & n34504 ) | ( n17155 & n34504 ) ;
  assign n44535 = n44534 ^ n44533 ^ n9670 ;
  assign n44536 = n44535 ^ n13453 ^ 1'b0 ;
  assign n44537 = n38652 | n44536 ;
  assign n44538 = n28439 ^ n7793 ^ 1'b0 ;
  assign n44539 = ~n28104 & n44538 ;
  assign n44540 = ( ~n388 & n10149 ) | ( ~n388 & n27574 ) | ( n10149 & n27574 ) ;
  assign n44541 = n26990 ^ n12710 ^ n7772 ;
  assign n44542 = n12138 | n21115 ;
  assign n44543 = n44542 ^ n20920 ^ 1'b0 ;
  assign n44544 = n44543 ^ n22049 ^ n11407 ;
  assign n44545 = ( ~n2396 & n6734 ) | ( ~n2396 & n39404 ) | ( n6734 & n39404 ) ;
  assign n44546 = n8575 & ~n34639 ;
  assign n44547 = ( n17031 & ~n23686 ) | ( n17031 & n28191 ) | ( ~n23686 & n28191 ) ;
  assign n44548 = ~n21972 & n44547 ;
  assign n44549 = n44548 ^ n27121 ^ 1'b0 ;
  assign n44550 = ( ~n3814 & n17239 ) | ( ~n3814 & n28368 ) | ( n17239 & n28368 ) ;
  assign n44551 = n44550 ^ n19279 ^ 1'b0 ;
  assign n44552 = n27731 & n41659 ;
  assign n44553 = n44552 ^ n8793 ^ n6159 ;
  assign n44554 = n31294 ^ n28050 ^ 1'b0 ;
  assign n44555 = ( n10833 & n17036 ) | ( n10833 & ~n36279 ) | ( n17036 & ~n36279 ) ;
  assign n44556 = n3655 & ~n9275 ;
  assign n44557 = n20214 ^ n5159 ^ 1'b0 ;
  assign n44558 = n44556 | n44557 ;
  assign n44559 = n13552 & n17081 ;
  assign n44560 = n44559 ^ n14004 ^ 1'b0 ;
  assign n44561 = n19242 & ~n44560 ;
  assign n44562 = ( n3406 & ~n7388 ) | ( n3406 & n17268 ) | ( ~n7388 & n17268 ) ;
  assign n44563 = n15309 & n28447 ;
  assign n44564 = ( n7241 & n15217 ) | ( n7241 & n28979 ) | ( n15217 & n28979 ) ;
  assign n44565 = ( n24893 & ~n28917 ) | ( n24893 & n44564 ) | ( ~n28917 & n44564 ) ;
  assign n44566 = n34538 ^ n3160 ^ 1'b0 ;
  assign n44567 = n35497 ^ n21062 ^ n17905 ;
  assign n44568 = n37326 ^ n32520 ^ n8517 ;
  assign n44569 = n25278 & ~n44568 ;
  assign n44570 = n44569 ^ n17076 ^ 1'b0 ;
  assign n44571 = n35402 ^ n34685 ^ n7389 ;
  assign n44572 = ~n6344 & n44571 ;
  assign n44573 = n44572 ^ n41367 ^ 1'b0 ;
  assign n44574 = ( ~n9487 & n16109 ) | ( ~n9487 & n37141 ) | ( n16109 & n37141 ) ;
  assign n44575 = n44574 ^ n43182 ^ n40664 ;
  assign n44576 = n16504 ^ n9196 ^ 1'b0 ;
  assign n44577 = ~n32758 & n44576 ;
  assign n44578 = ~n6582 & n44577 ;
  assign n44579 = n44578 ^ n10233 ^ 1'b0 ;
  assign n44580 = n7520 & n44579 ;
  assign n44581 = ~n29081 & n44580 ;
  assign n44582 = n44581 ^ n30188 ^ 1'b0 ;
  assign n44583 = n14600 & ~n44582 ;
  assign n44584 = n9328 & ~n9511 ;
  assign n44585 = n36541 ^ n9341 ^ n2428 ;
  assign n44586 = n18130 ^ x19 ^ 1'b0 ;
  assign n44587 = n44585 & n44586 ;
  assign n44588 = n22662 & n26441 ;
  assign n44589 = n44588 ^ n8059 ^ 1'b0 ;
  assign n44590 = ~n10720 & n35971 ;
  assign n44591 = n24512 & n44590 ;
  assign n44592 = n21959 | n37802 ;
  assign n44593 = n44592 ^ n13574 ^ 1'b0 ;
  assign n44594 = n6122 & ~n44593 ;
  assign n44595 = n4680 & ~n23845 ;
  assign n44596 = ~n44577 & n44595 ;
  assign n44597 = ( n19604 & ~n39748 ) | ( n19604 & n44596 ) | ( ~n39748 & n44596 ) ;
  assign n44598 = ( n12324 & n19151 ) | ( n12324 & ~n19655 ) | ( n19151 & ~n19655 ) ;
  assign n44599 = n24565 | n26217 ;
  assign n44600 = n44599 ^ n13272 ^ 1'b0 ;
  assign n44601 = n44600 ^ n40563 ^ 1'b0 ;
  assign n44602 = ~n8479 & n27979 ;
  assign n44603 = n17817 & n44602 ;
  assign n44604 = n40373 ^ n4357 ^ 1'b0 ;
  assign n44605 = n11220 | n44604 ;
  assign n44606 = n43659 ^ n9946 ^ 1'b0 ;
  assign n44607 = n12360 ^ n8364 ^ n1063 ;
  assign n44608 = n35294 ^ n15931 ^ n9971 ;
  assign n44609 = n29736 ^ n17261 ^ 1'b0 ;
  assign n44610 = ( n19473 & ~n44608 ) | ( n19473 & n44609 ) | ( ~n44608 & n44609 ) ;
  assign n44611 = n29866 ^ n9973 ^ n693 ;
  assign n44612 = n18653 ^ n1108 ^ 1'b0 ;
  assign n44613 = n44612 ^ n27117 ^ n20554 ;
  assign n44614 = n7776 ^ n1427 ^ 1'b0 ;
  assign n44615 = ( ~x25 & n24005 ) | ( ~x25 & n28031 ) | ( n24005 & n28031 ) ;
  assign n44616 = n44615 ^ n4564 ^ 1'b0 ;
  assign n44617 = n44614 & n44616 ;
  assign n44618 = n30604 ^ n19065 ^ n9584 ;
  assign n44619 = n19278 & n36947 ;
  assign n44620 = ~n29681 & n44619 ;
  assign n44621 = n15729 | n21065 ;
  assign n44622 = n44621 ^ n11767 ^ 1'b0 ;
  assign n44623 = n38085 ^ n16053 ^ 1'b0 ;
  assign n44624 = ~n21642 & n44623 ;
  assign n44625 = ( n627 & ~n4840 ) | ( n627 & n17058 ) | ( ~n4840 & n17058 ) ;
  assign n44626 = ( n6907 & n9381 ) | ( n6907 & ~n16113 ) | ( n9381 & ~n16113 ) ;
  assign n44627 = n44626 ^ n37008 ^ n8085 ;
  assign n44628 = ( n10522 & n12498 ) | ( n10522 & n26166 ) | ( n12498 & n26166 ) ;
  assign n44629 = ( n2607 & ~n2760 ) | ( n2607 & n7406 ) | ( ~n2760 & n7406 ) ;
  assign n44630 = n44629 ^ n38412 ^ n8647 ;
  assign n44631 = n44630 ^ n17439 ^ 1'b0 ;
  assign n44632 = ~n8796 & n24898 ;
  assign n44633 = ~n3146 & n44632 ;
  assign n44634 = ( ~n2132 & n27795 ) | ( ~n2132 & n35015 ) | ( n27795 & n35015 ) ;
  assign n44635 = n44634 ^ n42341 ^ n25030 ;
  assign n44636 = n2637 & ~n44635 ;
  assign n44637 = n44636 ^ n19214 ^ 1'b0 ;
  assign n44638 = n3303 | n11332 ;
  assign n44639 = n44637 | n44638 ;
  assign n44640 = n14103 ^ n5317 ^ n2930 ;
  assign n44641 = n4326 ^ n2174 ^ 1'b0 ;
  assign n44642 = n44640 & n44641 ;
  assign n44643 = n42376 ^ n36191 ^ n4691 ;
  assign n44644 = n273 | n24801 ;
  assign n44645 = n44644 ^ n9911 ^ 1'b0 ;
  assign n44646 = n24531 ^ n16244 ^ n15601 ;
  assign n44647 = ( n6677 & n22829 ) | ( n6677 & n44646 ) | ( n22829 & n44646 ) ;
  assign n44648 = ( n2034 & ~n44645 ) | ( n2034 & n44647 ) | ( ~n44645 & n44647 ) ;
  assign n44649 = ( ~n1888 & n28948 ) | ( ~n1888 & n44648 ) | ( n28948 & n44648 ) ;
  assign n44650 = ( ~n9301 & n24521 ) | ( ~n9301 & n39406 ) | ( n24521 & n39406 ) ;
  assign n44651 = ( ~n9930 & n27275 ) | ( ~n9930 & n31343 ) | ( n27275 & n31343 ) ;
  assign n44652 = n10829 | n15457 ;
  assign n44653 = n16580 & ~n44652 ;
  assign n44654 = n44653 ^ n39662 ^ n16448 ;
  assign n44655 = ( ~n2394 & n7259 ) | ( ~n2394 & n29472 ) | ( n7259 & n29472 ) ;
  assign n44656 = n40786 & n44655 ;
  assign n44657 = n44656 ^ n36183 ^ 1'b0 ;
  assign n44658 = n44384 ^ n22799 ^ 1'b0 ;
  assign n44659 = n7606 | n44658 ;
  assign n44660 = ~n4356 & n8928 ;
  assign n44661 = ~n11040 & n44660 ;
  assign n44662 = n44661 ^ n14040 ^ 1'b0 ;
  assign n44663 = n39685 ^ n27503 ^ 1'b0 ;
  assign n44664 = n40092 ^ n15479 ^ 1'b0 ;
  assign n44665 = ~n17110 & n44664 ;
  assign n44666 = n44665 ^ n31105 ^ 1'b0 ;
  assign n44667 = n30477 ^ n25684 ^ 1'b0 ;
  assign n44668 = n2857 | n7423 ;
  assign n44669 = n44668 ^ n7849 ^ 1'b0 ;
  assign n44670 = n44669 ^ n27174 ^ n23193 ;
  assign n44671 = n6488 | n9530 ;
  assign n44672 = n8234 ^ n6341 ^ 1'b0 ;
  assign n44673 = n44672 ^ n17708 ^ 1'b0 ;
  assign n44674 = n30607 & n44673 ;
  assign n44675 = n37808 ^ n24402 ^ 1'b0 ;
  assign n44676 = x63 & n44675 ;
  assign n44677 = n6560 ^ n3992 ^ 1'b0 ;
  assign n44678 = ~n16119 & n44677 ;
  assign n44679 = n44678 ^ n14837 ^ 1'b0 ;
  assign n44680 = n20314 | n39357 ;
  assign n44681 = n44680 ^ n6867 ^ 1'b0 ;
  assign n44682 = ( n14870 & n37348 ) | ( n14870 & n44681 ) | ( n37348 & n44681 ) ;
  assign n44684 = ( ~n3305 & n11584 ) | ( ~n3305 & n14356 ) | ( n11584 & n14356 ) ;
  assign n44683 = n2493 & n4153 ;
  assign n44685 = n44684 ^ n44683 ^ n34813 ;
  assign n44686 = n44685 ^ n28416 ^ n14868 ;
  assign n44687 = ~n304 & n12499 ;
  assign n44688 = n44687 ^ n29182 ^ n13796 ;
  assign n44689 = n33973 ^ n21410 ^ n6615 ;
  assign n44690 = n24290 ^ n848 ^ 1'b0 ;
  assign n44691 = n20161 & n44690 ;
  assign n44692 = ~n29502 & n44691 ;
  assign n44693 = n43333 ^ n35454 ^ 1'b0 ;
  assign n44694 = n2069 | n44693 ;
  assign n44695 = n28259 ^ n9298 ^ 1'b0 ;
  assign n44696 = n587 & n44695 ;
  assign n44697 = n42612 ^ n12690 ^ 1'b0 ;
  assign n44698 = n8059 | n44697 ;
  assign n44699 = n6121 & n8137 ;
  assign n44700 = n44699 ^ n4000 ^ 1'b0 ;
  assign n44701 = ~n36501 & n44700 ;
  assign n44702 = n27376 ^ n13373 ^ n2598 ;
  assign n44703 = n11473 | n44702 ;
  assign n44704 = n6072 ^ n1722 ^ 1'b0 ;
  assign n44705 = n5155 & ~n44704 ;
  assign n44706 = n44705 ^ n9405 ^ n1611 ;
  assign n44707 = n7085 ^ n4466 ^ n1328 ;
  assign n44708 = n44707 ^ n26842 ^ n2816 ;
  assign n44709 = n36370 ^ n25165 ^ n2215 ;
  assign n44710 = n36362 ^ n15142 ^ 1'b0 ;
  assign n44711 = n36658 | n44710 ;
  assign n44712 = ( n17816 & ~n29068 ) | ( n17816 & n33608 ) | ( ~n29068 & n33608 ) ;
  assign n44718 = n37383 ^ n11287 ^ n6889 ;
  assign n44713 = n43036 ^ n22154 ^ n313 ;
  assign n44714 = n43210 ^ n973 ^ 1'b0 ;
  assign n44715 = ~n34029 & n44714 ;
  assign n44716 = ~n40877 & n44715 ;
  assign n44717 = n44713 & n44716 ;
  assign n44719 = n44718 ^ n44717 ^ n12558 ;
  assign n44720 = ( n35030 & n37192 ) | ( n35030 & ~n38365 ) | ( n37192 & ~n38365 ) ;
  assign n44721 = ( ~n20175 & n39124 ) | ( ~n20175 & n44720 ) | ( n39124 & n44720 ) ;
  assign n44723 = n10432 ^ n1706 ^ 1'b0 ;
  assign n44722 = ~n20932 & n43972 ;
  assign n44724 = n44723 ^ n44722 ^ n10949 ;
  assign n44725 = n44724 ^ n18294 ^ n7429 ;
  assign n44726 = ( n10649 & n44721 ) | ( n10649 & ~n44725 ) | ( n44721 & ~n44725 ) ;
  assign n44727 = ( ~n9077 & n14219 ) | ( ~n9077 & n33698 ) | ( n14219 & n33698 ) ;
  assign n44728 = ( ~n9197 & n11918 ) | ( ~n9197 & n14571 ) | ( n11918 & n14571 ) ;
  assign n44729 = n40626 ^ n21986 ^ 1'b0 ;
  assign n44730 = n4329 & n44729 ;
  assign n44731 = n38294 & ~n38652 ;
  assign n44732 = n8320 & n17839 ;
  assign n44733 = ~n5760 & n44732 ;
  assign n44734 = n24110 | n42482 ;
  assign n44735 = n44734 ^ n4601 ^ 1'b0 ;
  assign n44736 = n21399 ^ n7419 ^ n1789 ;
  assign n44737 = n17940 & n44736 ;
  assign n44738 = n10545 | n44737 ;
  assign n44739 = n44738 ^ n41081 ^ 1'b0 ;
  assign n44740 = n44739 ^ n10904 ^ 1'b0 ;
  assign n44741 = n9477 ^ n7709 ^ n3810 ;
  assign n44743 = n23811 ^ n2606 ^ 1'b0 ;
  assign n44742 = n13707 & ~n31256 ;
  assign n44744 = n44743 ^ n44742 ^ 1'b0 ;
  assign n44745 = n21833 ^ n11673 ^ 1'b0 ;
  assign n44746 = n27576 & ~n44745 ;
  assign n44747 = ( n10372 & n20471 ) | ( n10372 & n44746 ) | ( n20471 & n44746 ) ;
  assign n44748 = ( ~n26827 & n44744 ) | ( ~n26827 & n44747 ) | ( n44744 & n44747 ) ;
  assign n44749 = n24482 ^ n5833 ^ n4501 ;
  assign n44750 = ( n38571 & n44685 ) | ( n38571 & ~n44749 ) | ( n44685 & ~n44749 ) ;
  assign n44751 = ( x122 & ~n7009 ) | ( x122 & n14695 ) | ( ~n7009 & n14695 ) ;
  assign n44752 = n37856 ^ n6308 ^ n2301 ;
  assign n44753 = n44752 ^ n16600 ^ 1'b0 ;
  assign n44754 = ~n44751 & n44753 ;
  assign n44760 = ( n3861 & ~n23925 ) | ( n3861 & n39341 ) | ( ~n23925 & n39341 ) ;
  assign n44755 = n8156 & ~n25024 ;
  assign n44756 = n44755 ^ n19044 ^ 1'b0 ;
  assign n44757 = n31430 ^ n14091 ^ 1'b0 ;
  assign n44758 = n31516 & n44757 ;
  assign n44759 = n44756 & n44758 ;
  assign n44761 = n44760 ^ n44759 ^ 1'b0 ;
  assign n44762 = n37276 ^ n12661 ^ 1'b0 ;
  assign n44763 = ( n1970 & n7086 ) | ( n1970 & ~n43624 ) | ( n7086 & ~n43624 ) ;
  assign n44764 = n44763 ^ n31432 ^ n3887 ;
  assign n44765 = n12879 & ~n38368 ;
  assign n44766 = n44765 ^ n33482 ^ 1'b0 ;
  assign n44767 = n2190 ^ n1414 ^ n606 ;
  assign n44768 = n5183 & n44767 ;
  assign n44769 = n4253 & n9502 ;
  assign n44770 = n44768 & n44769 ;
  assign n44771 = n13510 & ~n44770 ;
  assign n44772 = n42672 & n44771 ;
  assign n44773 = n6281 | n26167 ;
  assign n44774 = n40841 & ~n44773 ;
  assign n44775 = n19480 & ~n44774 ;
  assign n44776 = n1494 & ~n13499 ;
  assign n44777 = ~n1995 & n44776 ;
  assign n44778 = n44777 ^ n44429 ^ 1'b0 ;
  assign n44779 = n10521 & ~n44778 ;
  assign n44780 = n21438 & n44779 ;
  assign n44781 = ~n44775 & n44780 ;
  assign n44782 = n15849 ^ n9573 ^ 1'b0 ;
  assign n44783 = n665 | n27604 ;
  assign n44784 = ( n18105 & n25371 ) | ( n18105 & n38834 ) | ( n25371 & n38834 ) ;
  assign n44785 = ( n5311 & n10778 ) | ( n5311 & ~n15880 ) | ( n10778 & ~n15880 ) ;
  assign n44786 = ( n322 & n23012 ) | ( n322 & n35294 ) | ( n23012 & n35294 ) ;
  assign n44787 = n44786 ^ n43648 ^ n31895 ;
  assign n44788 = ( n42290 & n44785 ) | ( n42290 & n44787 ) | ( n44785 & n44787 ) ;
  assign n44789 = n13099 ^ n6115 ^ 1'b0 ;
  assign n44790 = n41734 ^ n6118 ^ 1'b0 ;
  assign n44791 = n44789 & n44790 ;
  assign n44792 = ~n897 & n18377 ;
  assign n44793 = ~n24288 & n44792 ;
  assign n44794 = n21218 & n30473 ;
  assign n44795 = ~n8262 & n44794 ;
  assign n44796 = n18551 & n35836 ;
  assign n44797 = n3240 & n44796 ;
  assign n44798 = n44797 ^ n25588 ^ n13794 ;
  assign n44799 = n38027 ^ n20409 ^ n6365 ;
  assign n44801 = n14088 ^ n5798 ^ 1'b0 ;
  assign n44802 = n30328 & ~n44801 ;
  assign n44800 = n16820 | n19949 ;
  assign n44803 = n44802 ^ n44800 ^ 1'b0 ;
  assign n44804 = n654 | n7956 ;
  assign n44805 = ( n1236 & ~n19522 ) | ( n1236 & n44804 ) | ( ~n19522 & n44804 ) ;
  assign n44806 = n20742 ^ n10769 ^ 1'b0 ;
  assign n44807 = n40029 | n44806 ;
  assign n44808 = ( ~n18607 & n44805 ) | ( ~n18607 & n44807 ) | ( n44805 & n44807 ) ;
  assign n44809 = n44808 ^ n41025 ^ n9360 ;
  assign n44810 = n28431 ^ n25883 ^ 1'b0 ;
  assign n44811 = ~n25262 & n44810 ;
  assign n44812 = n44811 ^ n20848 ^ 1'b0 ;
  assign n44813 = n23375 | n31485 ;
  assign n44814 = n44813 ^ n34944 ^ 1'b0 ;
  assign n44815 = n38652 ^ n25142 ^ 1'b0 ;
  assign n44816 = n22015 & n44815 ;
  assign n44817 = n7213 & n10533 ;
  assign n44818 = ~n14740 & n44817 ;
  assign n44819 = n6511 & ~n44818 ;
  assign n44820 = n39584 ^ n23442 ^ n6872 ;
  assign n44821 = n44820 ^ n10536 ^ n1439 ;
  assign n44823 = n9928 ^ n6594 ^ n593 ;
  assign n44822 = ( n31992 & n36101 ) | ( n31992 & n39871 ) | ( n36101 & n39871 ) ;
  assign n44824 = n44823 ^ n44822 ^ 1'b0 ;
  assign n44825 = n8890 & n44824 ;
  assign n44826 = n44825 ^ n35894 ^ n5375 ;
  assign n44827 = n8126 & ~n40174 ;
  assign n44828 = n44827 ^ n35052 ^ n9872 ;
  assign n44829 = ( n3474 & ~n13235 ) | ( n3474 & n27872 ) | ( ~n13235 & n27872 ) ;
  assign n44830 = n20495 & n26486 ;
  assign n44831 = n31563 ^ n23346 ^ n4814 ;
  assign n44832 = n12418 & n44831 ;
  assign n44833 = ~n6275 & n44832 ;
  assign n44834 = ~n27781 & n44350 ;
  assign n44835 = n44834 ^ n19713 ^ 1'b0 ;
  assign n44836 = ( n1393 & ~n13061 ) | ( n1393 & n21222 ) | ( ~n13061 & n21222 ) ;
  assign n44837 = n7626 | n44836 ;
  assign n44838 = n44837 ^ n9483 ^ 1'b0 ;
  assign n44839 = n37013 ^ n36227 ^ 1'b0 ;
  assign n44840 = ~n2813 & n44839 ;
  assign n44841 = n29776 | n44840 ;
  assign n44844 = ~n3902 & n25534 ;
  assign n44845 = n5873 & n44844 ;
  assign n44842 = n35751 & n40881 ;
  assign n44843 = ~n3410 & n44842 ;
  assign n44846 = n44845 ^ n44843 ^ 1'b0 ;
  assign n44847 = n16163 ^ n13816 ^ n13558 ;
  assign n44848 = ( ~n9248 & n34611 ) | ( ~n9248 & n44847 ) | ( n34611 & n44847 ) ;
  assign n44849 = n44848 ^ n30384 ^ 1'b0 ;
  assign n44850 = n9147 | n16163 ;
  assign n44851 = n44850 ^ n9233 ^ 1'b0 ;
  assign n44852 = ( ~n13347 & n38782 ) | ( ~n13347 & n44851 ) | ( n38782 & n44851 ) ;
  assign n44853 = n38229 ^ n6979 ^ 1'b0 ;
  assign n44854 = n8419 & ~n44853 ;
  assign n44855 = n3342 & n21444 ;
  assign n44856 = n16634 & n44855 ;
  assign n44857 = ( n18308 & n21218 ) | ( n18308 & n32104 ) | ( n21218 & n32104 ) ;
  assign n44860 = n34237 ^ n29582 ^ n13906 ;
  assign n44858 = ~n3526 & n4023 ;
  assign n44859 = n44858 ^ n30835 ^ 1'b0 ;
  assign n44861 = n44860 ^ n44859 ^ n35351 ;
  assign n44863 = n14206 ^ n3307 ^ 1'b0 ;
  assign n44864 = ~n16284 & n44863 ;
  assign n44862 = n19746 ^ n7578 ^ n3910 ;
  assign n44865 = n44864 ^ n44862 ^ n6865 ;
  assign n44866 = ( n2986 & ~n20535 ) | ( n2986 & n28512 ) | ( ~n20535 & n28512 ) ;
  assign n44867 = n23294 ^ n7120 ^ 1'b0 ;
  assign n44868 = n4804 & ~n44867 ;
  assign n44869 = ( ~n478 & n10113 ) | ( ~n478 & n44868 ) | ( n10113 & n44868 ) ;
  assign n44870 = n44869 ^ n14772 ^ n6516 ;
  assign n44871 = n7551 | n20508 ;
  assign n44872 = n23668 | n44871 ;
  assign n44873 = ( n7175 & n28322 ) | ( n7175 & n44872 ) | ( n28322 & n44872 ) ;
  assign n44874 = ~n10420 & n39584 ;
  assign n44875 = n28819 & n44874 ;
  assign n44876 = n8970 & ~n31737 ;
  assign n44877 = n44876 ^ n24746 ^ 1'b0 ;
  assign n44878 = ~n8506 & n18330 ;
  assign n44879 = ~n44877 & n44878 ;
  assign n44881 = ~n5595 & n11429 ;
  assign n44880 = n15413 & ~n41367 ;
  assign n44882 = n44881 ^ n44880 ^ 1'b0 ;
  assign n44883 = ( n1339 & n30179 ) | ( n1339 & n44882 ) | ( n30179 & n44882 ) ;
  assign n44884 = ( n1036 & ~n12985 ) | ( n1036 & n35121 ) | ( ~n12985 & n35121 ) ;
  assign n44885 = ( ~n19315 & n35656 ) | ( ~n19315 & n44884 ) | ( n35656 & n44884 ) ;
  assign n44888 = n11467 & n12557 ;
  assign n44889 = n44888 ^ n6927 ^ 1'b0 ;
  assign n44886 = n2042 | n24869 ;
  assign n44887 = ( n17855 & ~n30001 ) | ( n17855 & n44886 ) | ( ~n30001 & n44886 ) ;
  assign n44890 = n44889 ^ n44887 ^ 1'b0 ;
  assign n44891 = n11800 & ~n44890 ;
  assign n44892 = ( ~n11357 & n15142 ) | ( ~n11357 & n26975 ) | ( n15142 & n26975 ) ;
  assign n44893 = ( ~n21259 & n44891 ) | ( ~n21259 & n44892 ) | ( n44891 & n44892 ) ;
  assign n44894 = n10452 ^ n3847 ^ 1'b0 ;
  assign n44895 = n5704 | n6048 ;
  assign n44896 = n44894 & ~n44895 ;
  assign n44897 = ( n1901 & n14185 ) | ( n1901 & n18043 ) | ( n14185 & n18043 ) ;
  assign n44898 = n3117 | n44897 ;
  assign n44899 = n5889 & ~n44898 ;
  assign n44900 = n2785 & n36918 ;
  assign n44901 = n44899 & n44900 ;
  assign n44902 = ~n11613 & n12882 ;
  assign n44903 = n31660 ^ n520 ^ 1'b0 ;
  assign n44904 = ( n2574 & ~n24290 ) | ( n2574 & n44243 ) | ( ~n24290 & n44243 ) ;
  assign n44905 = n44904 ^ n41150 ^ n9469 ;
  assign n44909 = n10926 ^ n2353 ^ n1612 ;
  assign n44906 = n17047 ^ n1592 ^ 1'b0 ;
  assign n44907 = n10974 & n16323 ;
  assign n44908 = ~n44906 & n44907 ;
  assign n44910 = n44909 ^ n44908 ^ n42961 ;
  assign n44911 = n13218 | n20026 ;
  assign n44912 = n9736 & n40595 ;
  assign n44913 = n12261 & n44912 ;
  assign n44914 = ~n20378 & n44913 ;
  assign n44915 = n40292 ^ n32362 ^ n6364 ;
  assign n44916 = n42287 ^ n39080 ^ 1'b0 ;
  assign n44917 = n15427 & n44916 ;
  assign n44918 = n9670 | n36953 ;
  assign n44919 = n386 | n18875 ;
  assign n44920 = ~n25732 & n33122 ;
  assign n44921 = ( n7485 & n33932 ) | ( n7485 & ~n44920 ) | ( n33932 & ~n44920 ) ;
  assign n44922 = n43869 ^ n3154 ^ 1'b0 ;
  assign n44923 = n35488 ^ n34820 ^ 1'b0 ;
  assign n44924 = n24279 | n34489 ;
  assign n44925 = n44924 ^ n5835 ^ 1'b0 ;
  assign n44926 = n12089 & ~n24441 ;
  assign n44927 = ( n26154 & ~n44925 ) | ( n26154 & n44926 ) | ( ~n44925 & n44926 ) ;
  assign n44928 = ( ~n443 & n10048 ) | ( ~n443 & n12247 ) | ( n10048 & n12247 ) ;
  assign n44929 = ~n5865 & n44928 ;
  assign n44930 = n25004 & n44929 ;
  assign n44931 = n11384 & ~n44930 ;
  assign n44932 = n3196 & n44931 ;
  assign n44933 = ~n938 & n11118 ;
  assign n44934 = n44933 ^ n9456 ^ 1'b0 ;
  assign n44935 = ( n1630 & n15941 ) | ( n1630 & ~n36045 ) | ( n15941 & ~n36045 ) ;
  assign n44936 = ( n12205 & n15456 ) | ( n12205 & n17807 ) | ( n15456 & n17807 ) ;
  assign n44937 = n7880 & n34616 ;
  assign n44938 = n44937 ^ n25605 ^ 1'b0 ;
  assign n44939 = ( n20679 & n44936 ) | ( n20679 & n44938 ) | ( n44936 & n44938 ) ;
  assign n44940 = n40766 ^ n15383 ^ n2775 ;
  assign n44941 = ( n1500 & ~n5618 ) | ( n1500 & n31033 ) | ( ~n5618 & n31033 ) ;
  assign n44942 = n11099 & ~n36078 ;
  assign n44943 = n9930 | n38719 ;
  assign n44944 = n34798 & ~n44943 ;
  assign n44945 = ( n547 & n22096 ) | ( n547 & n24553 ) | ( n22096 & n24553 ) ;
  assign n44946 = n44945 ^ n28503 ^ n3160 ;
  assign n44947 = n36128 | n41990 ;
  assign n44948 = n44946 | n44947 ;
  assign n44949 = ~n22202 & n37592 ;
  assign n44950 = n11644 & n16341 ;
  assign n44951 = n44950 ^ n7977 ^ 1'b0 ;
  assign n44952 = ( n21428 & n39970 ) | ( n21428 & ~n44951 ) | ( n39970 & ~n44951 ) ;
  assign n44953 = n37927 ^ n34579 ^ 1'b0 ;
  assign n44954 = n39877 ^ n8836 ^ n8453 ;
  assign n44955 = n2394 & ~n35968 ;
  assign n44956 = ~n20213 & n43631 ;
  assign n44957 = n6868 & n27679 ;
  assign n44958 = n16149 ^ n841 ^ 1'b0 ;
  assign n44959 = x58 & ~n30356 ;
  assign n44960 = n44959 ^ n37903 ^ 1'b0 ;
  assign n44961 = n3352 ^ n1333 ^ 1'b0 ;
  assign n44962 = ( ~n4239 & n18644 ) | ( ~n4239 & n22170 ) | ( n18644 & n22170 ) ;
  assign n44963 = n39551 ^ n21178 ^ 1'b0 ;
  assign n44964 = n44962 | n44963 ;
  assign n44965 = ( n4642 & n22776 ) | ( n4642 & ~n44964 ) | ( n22776 & ~n44964 ) ;
  assign n44966 = n44961 & n44965 ;
  assign n44967 = n19824 ^ n11058 ^ n1690 ;
  assign n44968 = n15124 & n44967 ;
  assign n44969 = ( n23746 & ~n24927 ) | ( n23746 & n44968 ) | ( ~n24927 & n44968 ) ;
  assign n44970 = n20102 ^ n8104 ^ 1'b0 ;
  assign n44971 = n2428 & n44970 ;
  assign n44972 = n44971 ^ n14859 ^ 1'b0 ;
  assign n44973 = n29035 ^ n21840 ^ n15799 ;
  assign n44974 = n1819 | n21957 ;
  assign n44975 = n44973 & ~n44974 ;
  assign n44976 = n6539 & n17152 ;
  assign n44977 = n44976 ^ n14836 ^ 1'b0 ;
  assign n44978 = ( ~n1645 & n15962 ) | ( ~n1645 & n25281 ) | ( n15962 & n25281 ) ;
  assign n44979 = n22621 ^ n8512 ^ n7359 ;
  assign n44980 = ( n1229 & ~n38112 ) | ( n1229 & n44979 ) | ( ~n38112 & n44979 ) ;
  assign n44981 = ( n22455 & n42491 ) | ( n22455 & n44980 ) | ( n42491 & n44980 ) ;
  assign n44982 = ~n23348 & n28087 ;
  assign n44983 = n1924 & ~n16556 ;
  assign n44984 = n5013 | n6947 ;
  assign n44985 = n44984 ^ n32619 ^ n22717 ;
  assign n44986 = n7365 & n13202 ;
  assign n44987 = n44986 ^ n7456 ^ 1'b0 ;
  assign n44988 = n23552 ^ n23286 ^ 1'b0 ;
  assign n44989 = n6036 | n44988 ;
  assign n44990 = n44989 ^ n2926 ^ 1'b0 ;
  assign n44991 = n17600 & ~n25722 ;
  assign n44992 = ~n38713 & n44991 ;
  assign n44993 = n38681 ^ n30151 ^ 1'b0 ;
  assign n44994 = ( n3370 & n12932 ) | ( n3370 & ~n22382 ) | ( n12932 & ~n22382 ) ;
  assign n44997 = ( x75 & n4846 ) | ( x75 & ~n5846 ) | ( n4846 & ~n5846 ) ;
  assign n44995 = n28301 ^ n25749 ^ n17882 ;
  assign n44996 = n44995 ^ n34125 ^ n18511 ;
  assign n44998 = n44997 ^ n44996 ^ n2329 ;
  assign n44999 = n10693 | n13070 ;
  assign n45000 = n11472 & ~n44999 ;
  assign n45001 = ( n4508 & ~n36666 ) | ( n4508 & n45000 ) | ( ~n36666 & n45000 ) ;
  assign n45002 = n22307 & ~n25242 ;
  assign n45003 = n8019 & ~n36986 ;
  assign n45004 = n45003 ^ n14744 ^ 1'b0 ;
  assign n45005 = n30235 ^ n8686 ^ n5197 ;
  assign n45006 = ~n10019 & n45005 ;
  assign n45007 = n35922 ^ n29059 ^ n16158 ;
  assign n45008 = n13990 & ~n29691 ;
  assign n45009 = n45008 ^ n11858 ^ 1'b0 ;
  assign n45010 = n45009 ^ n14905 ^ n9031 ;
  assign n45011 = n17480 ^ n10594 ^ 1'b0 ;
  assign n45012 = n13387 & ~n45011 ;
  assign n45013 = ( n7391 & n14485 ) | ( n7391 & ~n30076 ) | ( n14485 & ~n30076 ) ;
  assign n45014 = ( n6213 & ~n26155 ) | ( n6213 & n43264 ) | ( ~n26155 & n43264 ) ;
  assign n45015 = n35046 ^ n14010 ^ x234 ;
  assign n45016 = ( n45013 & n45014 ) | ( n45013 & n45015 ) | ( n45014 & n45015 ) ;
  assign n45017 = n24551 ^ n19983 ^ 1'b0 ;
  assign n45018 = n10103 | n18695 ;
  assign n45019 = n22234 & ~n45018 ;
  assign n45020 = n23029 | n35346 ;
  assign n45021 = n5574 | n45020 ;
  assign n45022 = ~n31789 & n45021 ;
  assign n45024 = n27576 ^ n8827 ^ 1'b0 ;
  assign n45025 = n34856 & ~n45024 ;
  assign n45023 = n22662 ^ n13667 ^ n4659 ;
  assign n45026 = n45025 ^ n45023 ^ 1'b0 ;
  assign n45027 = n10040 & ~n42713 ;
  assign n45028 = ( n11820 & n31755 ) | ( n11820 & n45027 ) | ( n31755 & n45027 ) ;
  assign n45029 = n22156 ^ n16136 ^ 1'b0 ;
  assign n45030 = n24133 | n32505 ;
  assign n45031 = ( n22974 & n28694 ) | ( n22974 & ~n45030 ) | ( n28694 & ~n45030 ) ;
  assign n45032 = ( n36897 & n45029 ) | ( n36897 & ~n45031 ) | ( n45029 & ~n45031 ) ;
  assign n45033 = n2291 & n5005 ;
  assign n45034 = ( ~n17156 & n25628 ) | ( ~n17156 & n28836 ) | ( n25628 & n28836 ) ;
  assign n45035 = n23961 ^ n16237 ^ 1'b0 ;
  assign n45036 = n2224 & n12380 ;
  assign n45037 = ( n1440 & n4117 ) | ( n1440 & ~n45036 ) | ( n4117 & ~n45036 ) ;
  assign n45038 = n28252 ^ n27334 ^ 1'b0 ;
  assign n45039 = n3182 & n45038 ;
  assign n45040 = ( n35071 & n35916 ) | ( n35071 & n45039 ) | ( n35916 & n45039 ) ;
  assign n45041 = n45040 ^ n13224 ^ n3212 ;
  assign n45042 = ( n9005 & ~n9584 ) | ( n9005 & n20484 ) | ( ~n9584 & n20484 ) ;
  assign n45043 = n11819 & n44435 ;
  assign n45044 = n24156 ^ n10179 ^ 1'b0 ;
  assign n45045 = n30008 | n45044 ;
  assign n45046 = n21168 & ~n31978 ;
  assign n45047 = n15593 | n17564 ;
  assign n45048 = n5584 & ~n45047 ;
  assign n45049 = n34887 ^ n21525 ^ n6149 ;
  assign n45050 = n43280 ^ n5339 ^ n632 ;
  assign n45051 = n45050 ^ n43469 ^ n12751 ;
  assign n45052 = ~n15457 & n45051 ;
  assign n45053 = ~n45049 & n45052 ;
  assign n45054 = n31872 ^ n6390 ^ 1'b0 ;
  assign n45055 = ( n2455 & ~n12244 ) | ( n2455 & n15226 ) | ( ~n12244 & n15226 ) ;
  assign n45056 = n15142 | n20263 ;
  assign n45057 = n45056 ^ n44913 ^ 1'b0 ;
  assign n45058 = n3939 | n4498 ;
  assign n45059 = ( ~n7480 & n38205 ) | ( ~n7480 & n45058 ) | ( n38205 & n45058 ) ;
  assign n45060 = ( n14622 & n20797 ) | ( n14622 & n45059 ) | ( n20797 & n45059 ) ;
  assign n45061 = n9473 | n19525 ;
  assign n45062 = n45061 ^ n1724 ^ 1'b0 ;
  assign n45063 = ( n12683 & n14883 ) | ( n12683 & n45062 ) | ( n14883 & n45062 ) ;
  assign n45064 = ( ~n29436 & n45060 ) | ( ~n29436 & n45063 ) | ( n45060 & n45063 ) ;
  assign n45065 = n1637 & n29598 ;
  assign n45066 = n45065 ^ n41410 ^ n28920 ;
  assign n45068 = ( ~n6510 & n12411 ) | ( ~n6510 & n26639 ) | ( n12411 & n26639 ) ;
  assign n45067 = n14942 & n30700 ;
  assign n45069 = n45068 ^ n45067 ^ 1'b0 ;
  assign n45070 = n29689 ^ n12360 ^ 1'b0 ;
  assign n45071 = n6033 | n45070 ;
  assign n45072 = ( ~n960 & n8354 ) | ( ~n960 & n36457 ) | ( n8354 & n36457 ) ;
  assign n45075 = n8646 ^ n3756 ^ 1'b0 ;
  assign n45076 = n15494 & n45075 ;
  assign n45073 = n7671 & n26353 ;
  assign n45074 = n45073 ^ n17700 ^ 1'b0 ;
  assign n45077 = n45076 ^ n45074 ^ n18385 ;
  assign n45078 = n39030 ^ n26020 ^ n6001 ;
  assign n45079 = n5504 & ~n20995 ;
  assign n45080 = n34894 ^ n28752 ^ 1'b0 ;
  assign n45081 = n45080 ^ n34243 ^ n28720 ;
  assign n45082 = n32520 ^ n21799 ^ n19161 ;
  assign n45083 = x160 & ~n45082 ;
  assign n45084 = ~n25438 & n45083 ;
  assign n45085 = n15796 & ~n45084 ;
  assign n45086 = n14381 & n45085 ;
  assign n45087 = n14723 ^ n13019 ^ 1'b0 ;
  assign n45088 = n11863 & n45087 ;
  assign n45089 = n31976 | n45088 ;
  assign n45090 = n29025 & ~n45089 ;
  assign n45091 = n45090 ^ n3221 ^ 1'b0 ;
  assign n45092 = n8128 & ~n22410 ;
  assign n45093 = n39228 ^ n32852 ^ n23015 ;
  assign n45094 = n45093 ^ n5446 ^ 1'b0 ;
  assign n45095 = n9602 ^ n3313 ^ 1'b0 ;
  assign n45096 = ( ~n4519 & n37434 ) | ( ~n4519 & n45095 ) | ( n37434 & n45095 ) ;
  assign n45097 = ( ~n10790 & n29690 ) | ( ~n10790 & n33790 ) | ( n29690 & n33790 ) ;
  assign n45098 = ( ~n40057 & n45096 ) | ( ~n40057 & n45097 ) | ( n45096 & n45097 ) ;
  assign n45099 = n20247 ^ n16023 ^ n2705 ;
  assign n45100 = ~n14762 & n34481 ;
  assign n45101 = n30406 ^ n22012 ^ n21303 ;
  assign n45102 = n1786 & n45101 ;
  assign n45103 = ( n10898 & n27192 ) | ( n10898 & ~n27949 ) | ( n27192 & ~n27949 ) ;
  assign n45104 = n7019 ^ n2166 ^ 1'b0 ;
  assign n45106 = n37673 ^ n14960 ^ n1826 ;
  assign n45105 = n23625 & ~n34087 ;
  assign n45107 = n45106 ^ n45105 ^ 1'b0 ;
  assign n45110 = n23221 ^ n22439 ^ 1'b0 ;
  assign n45111 = n45110 ^ n32775 ^ n4759 ;
  assign n45112 = n45111 ^ n28932 ^ n21458 ;
  assign n45108 = n16864 ^ n14585 ^ x253 ;
  assign n45109 = ~n23985 & n45108 ;
  assign n45113 = n45112 ^ n45109 ^ 1'b0 ;
  assign n45114 = n13217 | n17643 ;
  assign n45115 = n45114 ^ n29373 ^ 1'b0 ;
  assign n45116 = n9263 & n17814 ;
  assign n45117 = n10292 & n45116 ;
  assign n45118 = ( n2831 & n11567 ) | ( n2831 & ~n45117 ) | ( n11567 & ~n45117 ) ;
  assign n45119 = n20135 ^ n16202 ^ n8543 ;
  assign n45120 = n6832 & ~n15491 ;
  assign n45121 = n45120 ^ n14381 ^ 1'b0 ;
  assign n45122 = ~n27673 & n45121 ;
  assign n45123 = ~n17753 & n45122 ;
  assign n45124 = ~n35461 & n45123 ;
  assign n45125 = ( n6723 & n45119 ) | ( n6723 & ~n45124 ) | ( n45119 & ~n45124 ) ;
  assign n45126 = n25567 & ~n42245 ;
  assign n45127 = n13852 & ~n17378 ;
  assign n45128 = n11980 & n19254 ;
  assign n45129 = n45128 ^ n16979 ^ 1'b0 ;
  assign n45130 = n45129 ^ n36350 ^ n10584 ;
  assign n45131 = ( n19663 & n45127 ) | ( n19663 & ~n45130 ) | ( n45127 & ~n45130 ) ;
  assign n45132 = n29332 ^ n20509 ^ n13929 ;
  assign n45133 = n45132 ^ n36818 ^ n3339 ;
  assign n45134 = n43254 ^ n22947 ^ 1'b0 ;
  assign n45135 = ~n23300 & n45134 ;
  assign n45136 = n33045 ^ n12014 ^ n11244 ;
  assign n45137 = n45136 ^ n37041 ^ n25392 ;
  assign n45138 = ~n11378 & n20663 ;
  assign n45139 = ~n4938 & n45138 ;
  assign n45140 = n12221 & ~n40760 ;
  assign n45141 = n45140 ^ n15373 ^ 1'b0 ;
  assign n45142 = n45139 | n45141 ;
  assign n45143 = n45137 & ~n45142 ;
  assign n45144 = n15971 | n30384 ;
  assign n45145 = ~n25588 & n30776 ;
  assign n45146 = ( n13004 & n14941 ) | ( n13004 & n21687 ) | ( n14941 & n21687 ) ;
  assign n45149 = n16754 ^ n2691 ^ 1'b0 ;
  assign n45150 = n24338 & n45149 ;
  assign n45147 = ( ~n1653 & n1814 ) | ( ~n1653 & n11614 ) | ( n1814 & n11614 ) ;
  assign n45148 = n7133 & n45147 ;
  assign n45151 = n45150 ^ n45148 ^ n29251 ;
  assign n45152 = n6887 & n15390 ;
  assign n45153 = ( ~n10824 & n14300 ) | ( ~n10824 & n45152 ) | ( n14300 & n45152 ) ;
  assign n45154 = n31651 ^ n11368 ^ 1'b0 ;
  assign n45155 = ( n33417 & n45153 ) | ( n33417 & n45154 ) | ( n45153 & n45154 ) ;
  assign n45156 = n34383 ^ n16565 ^ n5524 ;
  assign n45157 = n45152 ^ n27202 ^ n2922 ;
  assign n45158 = ( n9402 & n20399 ) | ( n9402 & ~n29324 ) | ( n20399 & ~n29324 ) ;
  assign n45159 = n45157 & n45158 ;
  assign n45160 = n1886 & ~n21241 ;
  assign n45161 = n45160 ^ n5688 ^ 1'b0 ;
  assign n45162 = ~n10565 & n35711 ;
  assign n45163 = n45162 ^ n18780 ^ n11629 ;
  assign n45164 = n10010 & n45163 ;
  assign n45165 = n4789 | n45164 ;
  assign n45166 = n14105 & ~n45165 ;
  assign n45167 = ~n2000 & n25132 ;
  assign n45168 = ~n1146 & n45167 ;
  assign n45169 = n25098 ^ n16904 ^ n15505 ;
  assign n45170 = n18241 ^ n12321 ^ n7122 ;
  assign n45171 = n25605 & ~n32069 ;
  assign n45172 = n4892 & n45171 ;
  assign n45173 = n45172 ^ n27158 ^ n17764 ;
  assign n45174 = n11794 & n19643 ;
  assign n45175 = n41090 | n45174 ;
  assign n45176 = ( n45170 & n45173 ) | ( n45170 & ~n45175 ) | ( n45173 & ~n45175 ) ;
  assign n45177 = n18935 ^ n12768 ^ n1288 ;
  assign n45178 = n37620 ^ n27600 ^ x141 ;
  assign n45179 = n17571 ^ n4332 ^ 1'b0 ;
  assign n45180 = n13499 ^ n9974 ^ n9577 ;
  assign n45181 = n18329 ^ n1763 ^ 1'b0 ;
  assign n45182 = n45180 & n45181 ;
  assign n45183 = n30478 ^ n19176 ^ 1'b0 ;
  assign n45184 = n37784 & ~n45183 ;
  assign n45185 = n17750 & ~n20051 ;
  assign n45186 = n7660 & n45185 ;
  assign n45187 = ( n2677 & ~n17135 ) | ( n2677 & n42907 ) | ( ~n17135 & n42907 ) ;
  assign n45188 = n45187 ^ n25595 ^ 1'b0 ;
  assign n45189 = n22406 | n45188 ;
  assign n45190 = n1098 | n45189 ;
  assign n45191 = n42553 & ~n45190 ;
  assign n45192 = n25887 ^ n2293 ^ 1'b0 ;
  assign n45193 = n3398 | n45192 ;
  assign n45194 = ~n1648 & n6837 ;
  assign n45195 = n45194 ^ n30287 ^ 1'b0 ;
  assign n45196 = ( ~n1400 & n4528 ) | ( ~n1400 & n15340 ) | ( n4528 & n15340 ) ;
  assign n45197 = ( n11751 & n45195 ) | ( n11751 & n45196 ) | ( n45195 & n45196 ) ;
  assign n45198 = ( n10494 & n19709 ) | ( n10494 & n20237 ) | ( n19709 & n20237 ) ;
  assign n45199 = n45198 ^ n2594 ^ 1'b0 ;
  assign n45200 = ( n3897 & n8523 ) | ( n3897 & n45199 ) | ( n8523 & n45199 ) ;
  assign n45201 = n27359 ^ n9684 ^ 1'b0 ;
  assign n45202 = n15821 & ~n32581 ;
  assign n45203 = n7677 & ~n15492 ;
  assign n45204 = n2585 & n8919 ;
  assign n45205 = ( n15811 & ~n45203 ) | ( n15811 & n45204 ) | ( ~n45203 & n45204 ) ;
  assign n45206 = ( n42632 & ~n45202 ) | ( n42632 & n45205 ) | ( ~n45202 & n45205 ) ;
  assign n45207 = n11998 | n38304 ;
  assign n45208 = n20487 ^ n10792 ^ n7157 ;
  assign n45209 = n45208 ^ n31589 ^ n18655 ;
  assign n45214 = ~n7874 & n36906 ;
  assign n45215 = n45214 ^ n7471 ^ 1'b0 ;
  assign n45210 = n602 & ~n7739 ;
  assign n45211 = ~n14194 & n45210 ;
  assign n45212 = n2770 & ~n16364 ;
  assign n45213 = ( n2107 & n45211 ) | ( n2107 & n45212 ) | ( n45211 & n45212 ) ;
  assign n45216 = n45215 ^ n45213 ^ n9952 ;
  assign n45217 = n27924 & n45216 ;
  assign n45218 = n5671 | n18695 ;
  assign n45219 = n41104 ^ n22213 ^ n13954 ;
  assign n45220 = ( ~n7018 & n18542 ) | ( ~n7018 & n28588 ) | ( n18542 & n28588 ) ;
  assign n45221 = n6704 | n23856 ;
  assign n45222 = n45221 ^ n26415 ^ n19271 ;
  assign n45223 = n10200 ^ n5978 ^ 1'b0 ;
  assign n45224 = n45222 & ~n45223 ;
  assign n45225 = ( n13450 & ~n18558 ) | ( n13450 & n45224 ) | ( ~n18558 & n45224 ) ;
  assign n45226 = n24299 | n32076 ;
  assign n45227 = n12431 & ~n45226 ;
  assign n45228 = n21050 ^ n16350 ^ 1'b0 ;
  assign n45229 = n31861 ^ n10302 ^ n7010 ;
  assign n45230 = ( ~n8366 & n18570 ) | ( ~n8366 & n45229 ) | ( n18570 & n45229 ) ;
  assign n45231 = n45230 ^ n12026 ^ n9883 ;
  assign n45232 = n42147 ^ n8984 ^ n5176 ;
  assign n45233 = ~n17139 & n41351 ;
  assign n45234 = n7056 & n45233 ;
  assign n45235 = n45234 ^ n7440 ^ 1'b0 ;
  assign n45236 = n45235 ^ n27048 ^ n14047 ;
  assign n45237 = n6787 | n7726 ;
  assign n45238 = n29270 & ~n45237 ;
  assign n45239 = n45238 ^ n10274 ^ n6969 ;
  assign n45240 = n30034 ^ n28080 ^ 1'b0 ;
  assign n45241 = n45240 ^ n25198 ^ n17018 ;
  assign n45242 = n21292 | n45241 ;
  assign n45250 = ( n10180 & n11204 ) | ( n10180 & ~n24719 ) | ( n11204 & ~n24719 ) ;
  assign n45243 = ( ~n8911 & n10777 ) | ( ~n8911 & n11859 ) | ( n10777 & n11859 ) ;
  assign n45244 = n45243 ^ n15527 ^ 1'b0 ;
  assign n45245 = n10570 & ~n45244 ;
  assign n45246 = n45245 ^ n5314 ^ 1'b0 ;
  assign n45247 = ~n488 & n45246 ;
  assign n45248 = n45247 ^ n21793 ^ 1'b0 ;
  assign n45249 = n36996 & ~n45248 ;
  assign n45251 = n45250 ^ n45249 ^ 1'b0 ;
  assign n45252 = ( n12486 & ~n23337 ) | ( n12486 & n35326 ) | ( ~n23337 & n35326 ) ;
  assign n45253 = n10263 & n45252 ;
  assign n45254 = n27738 & n45253 ;
  assign n45255 = n27257 ^ n3659 ^ n1089 ;
  assign n45256 = n11297 & n21096 ;
  assign n45257 = n45256 ^ n15214 ^ n12323 ;
  assign n45258 = n11788 ^ n11584 ^ n5576 ;
  assign n45259 = ( ~n5309 & n12363 ) | ( ~n5309 & n45258 ) | ( n12363 & n45258 ) ;
  assign n45260 = n22970 ^ n20034 ^ 1'b0 ;
  assign n45261 = n13025 | n45260 ;
  assign n45263 = ( ~n8558 & n11752 ) | ( ~n8558 & n12059 ) | ( n11752 & n12059 ) ;
  assign n45264 = ~n16953 & n45263 ;
  assign n45265 = n45264 ^ n6161 ^ 1'b0 ;
  assign n45262 = n37603 ^ n32704 ^ n5126 ;
  assign n45266 = n45265 ^ n45262 ^ n28541 ;
  assign n45267 = ( n15506 & n31206 ) | ( n15506 & ~n43945 ) | ( n31206 & ~n43945 ) ;
  assign n45268 = n45267 ^ n33604 ^ n19214 ;
  assign n45270 = ( n1543 & ~n8468 ) | ( n1543 & n12186 ) | ( ~n8468 & n12186 ) ;
  assign n45269 = ( n8049 & n19581 ) | ( n8049 & n24723 ) | ( n19581 & n24723 ) ;
  assign n45271 = n45270 ^ n45269 ^ 1'b0 ;
  assign n45272 = ( n1195 & ~n6158 ) | ( n1195 & n19411 ) | ( ~n6158 & n19411 ) ;
  assign n45273 = n45272 ^ n19638 ^ n8740 ;
  assign n45274 = ( n12128 & n43720 ) | ( n12128 & n45273 ) | ( n43720 & n45273 ) ;
  assign n45275 = n42079 ^ n5042 ^ 1'b0 ;
  assign n45276 = n24340 ^ n8334 ^ 1'b0 ;
  assign n45277 = n8756 | n45276 ;
  assign n45278 = ~n6838 & n35396 ;
  assign n45279 = n45278 ^ n18631 ^ 1'b0 ;
  assign n45280 = n12071 ^ n1183 ^ 1'b0 ;
  assign n45281 = ~n634 & n45280 ;
  assign n45282 = ( n13271 & ~n45279 ) | ( n13271 & n45281 ) | ( ~n45279 & n45281 ) ;
  assign n45283 = n26121 ^ n6038 ^ 1'b0 ;
  assign n45284 = n45283 ^ n37927 ^ 1'b0 ;
  assign n45285 = n45282 & ~n45284 ;
  assign n45286 = n44090 ^ n27827 ^ n19706 ;
  assign n45287 = ( n29841 & n31417 ) | ( n29841 & ~n45286 ) | ( n31417 & ~n45286 ) ;
  assign n45288 = ( n2350 & n10187 ) | ( n2350 & n38662 ) | ( n10187 & n38662 ) ;
  assign n45289 = ( ~n16117 & n20288 ) | ( ~n16117 & n35662 ) | ( n20288 & n35662 ) ;
  assign n45290 = n45139 ^ n43158 ^ 1'b0 ;
  assign n45291 = n7795 ^ n4780 ^ n2617 ;
  assign n45292 = n332 & n45291 ;
  assign n45293 = n45292 ^ n2349 ^ 1'b0 ;
  assign n45294 = n36391 | n45293 ;
  assign n45295 = n1587 | n45294 ;
  assign n45296 = n33771 | n34302 ;
  assign n45297 = n8688 & ~n9100 ;
  assign n45298 = n45297 ^ n3829 ^ 1'b0 ;
  assign n45299 = n28451 ^ n17831 ^ n10774 ;
  assign n45300 = n45299 ^ n36673 ^ n28144 ;
  assign n45301 = n40291 ^ n17245 ^ 1'b0 ;
  assign n45302 = n37464 & ~n45301 ;
  assign n45303 = n21326 ^ n20156 ^ n8979 ;
  assign n45304 = n16530 ^ n12675 ^ 1'b0 ;
  assign n45305 = n7398 & n45304 ;
  assign n45306 = ~n18964 & n45305 ;
  assign n45307 = n45306 ^ n34306 ^ 1'b0 ;
  assign n45308 = n19038 & ~n44442 ;
  assign n45309 = n3408 & n8644 ;
  assign n45310 = ~n45308 & n45309 ;
  assign n45311 = n12721 | n16385 ;
  assign n45312 = n40768 | n45311 ;
  assign n45313 = n2301 & n4428 ;
  assign n45314 = n3577 & n45313 ;
  assign n45315 = n36734 | n43045 ;
  assign n45316 = n45315 ^ n721 ^ 1'b0 ;
  assign n45317 = ( ~n19972 & n45314 ) | ( ~n19972 & n45316 ) | ( n45314 & n45316 ) ;
  assign n45318 = n20258 ^ n15519 ^ 1'b0 ;
  assign n45319 = n19944 ^ n19521 ^ n5956 ;
  assign n45320 = ( n5002 & n33013 ) | ( n5002 & ~n34891 ) | ( n33013 & ~n34891 ) ;
  assign n45321 = ( n22382 & n41573 ) | ( n22382 & ~n45320 ) | ( n41573 & ~n45320 ) ;
  assign n45322 = n37632 ^ n16737 ^ n10261 ;
  assign n45323 = n45322 ^ n27825 ^ 1'b0 ;
  assign n45324 = n5517 & n45323 ;
  assign n45325 = n35106 ^ n19367 ^ n19348 ;
  assign n45326 = ( n33854 & n45324 ) | ( n33854 & n45325 ) | ( n45324 & n45325 ) ;
  assign n45327 = n22234 ^ n18367 ^ n8536 ;
  assign n45328 = ( n8062 & ~n26908 ) | ( n8062 & n45327 ) | ( ~n26908 & n45327 ) ;
  assign n45329 = n17222 & ~n24743 ;
  assign n45330 = n45329 ^ n27063 ^ 1'b0 ;
  assign n45331 = n14613 | n44970 ;
  assign n45332 = n19629 | n20799 ;
  assign n45333 = n22577 ^ n17105 ^ n10667 ;
  assign n45334 = n30649 ^ n21661 ^ n12422 ;
  assign n45335 = n45334 ^ n18069 ^ n822 ;
  assign n45336 = n45335 ^ n18778 ^ n11022 ;
  assign n45337 = ( ~n11046 & n45333 ) | ( ~n11046 & n45336 ) | ( n45333 & n45336 ) ;
  assign n45338 = n2320 & ~n31729 ;
  assign n45339 = n45338 ^ n11534 ^ 1'b0 ;
  assign n45340 = n45339 ^ n1410 ^ 1'b0 ;
  assign n45341 = n30320 ^ n24364 ^ n1667 ;
  assign n45342 = n26314 ^ n9963 ^ 1'b0 ;
  assign n45343 = n45341 & n45342 ;
  assign n45344 = n40418 ^ n39209 ^ n7862 ;
  assign n45345 = n1932 & n26880 ;
  assign n45346 = n18630 & n45345 ;
  assign n45347 = n34481 & ~n37910 ;
  assign n45348 = n45347 ^ n20027 ^ 1'b0 ;
  assign n45349 = n1087 ^ x136 ^ 1'b0 ;
  assign n45350 = n20076 ^ n17826 ^ n3420 ;
  assign n45351 = n11379 ^ n10054 ^ 1'b0 ;
  assign n45352 = n45350 | n45351 ;
  assign n45353 = n45352 ^ n15364 ^ 1'b0 ;
  assign n45354 = n21533 ^ n20777 ^ 1'b0 ;
  assign n45355 = n17928 | n45354 ;
  assign n45356 = ( ~n16905 & n45198 ) | ( ~n16905 & n45355 ) | ( n45198 & n45355 ) ;
  assign n45357 = n7079 & ~n9633 ;
  assign n45358 = n45357 ^ n3653 ^ 1'b0 ;
  assign n45359 = ( n21552 & n29566 ) | ( n21552 & n45358 ) | ( n29566 & n45358 ) ;
  assign n45360 = n18249 ^ n14973 ^ n9277 ;
  assign n45361 = n45360 ^ n3592 ^ 1'b0 ;
  assign n45362 = n24687 ^ n13907 ^ n2535 ;
  assign n45363 = ~n31779 & n45362 ;
  assign n45364 = n1235 & n37559 ;
  assign n45365 = ( n2475 & n45363 ) | ( n2475 & ~n45364 ) | ( n45363 & ~n45364 ) ;
  assign n45366 = n7579 ^ n3674 ^ 1'b0 ;
  assign n45367 = n9329 & ~n45366 ;
  assign n45368 = n39582 ^ n27587 ^ 1'b0 ;
  assign n45369 = n28289 | n45368 ;
  assign n45370 = n16467 & n45369 ;
  assign n45371 = n8434 ^ n3997 ^ n1297 ;
  assign n45372 = n45371 ^ n8892 ^ 1'b0 ;
  assign n45373 = n5730 & ~n42128 ;
  assign n45374 = ~n15897 & n45373 ;
  assign n45375 = n45374 ^ n25567 ^ n10680 ;
  assign n45376 = n18143 & n30810 ;
  assign n45377 = n40640 ^ n6938 ^ n2131 ;
  assign n45378 = ( n21441 & n26724 ) | ( n21441 & n45377 ) | ( n26724 & n45377 ) ;
  assign n45379 = n29970 ^ n15154 ^ n6139 ;
  assign n45380 = ( n7024 & ~n37171 ) | ( n7024 & n45379 ) | ( ~n37171 & n45379 ) ;
  assign n45381 = n17497 ^ n7065 ^ 1'b0 ;
  assign n45382 = n23559 | n44965 ;
  assign n45383 = n45382 ^ n38001 ^ 1'b0 ;
  assign n45384 = n1793 & ~n29666 ;
  assign n45385 = n29678 & n45384 ;
  assign n45386 = n14912 ^ n1593 ^ 1'b0 ;
  assign n45387 = ~n3905 & n10173 ;
  assign n45388 = n45387 ^ n5486 ^ 1'b0 ;
  assign n45389 = n45388 ^ n31660 ^ 1'b0 ;
  assign n45390 = ( ~n37814 & n40422 ) | ( ~n37814 & n45389 ) | ( n40422 & n45389 ) ;
  assign n45391 = n30754 ^ n9708 ^ 1'b0 ;
  assign n45392 = n41509 | n43662 ;
  assign n45393 = n45392 ^ n16714 ^ 1'b0 ;
  assign n45395 = n20669 ^ n12158 ^ 1'b0 ;
  assign n45396 = n12653 | n45395 ;
  assign n45394 = ~n6287 & n10163 ;
  assign n45397 = n45396 ^ n45394 ^ n15035 ;
  assign n45398 = ~n28915 & n36604 ;
  assign n45399 = n31013 & n45398 ;
  assign n45400 = ( n6450 & n40454 ) | ( n6450 & ~n45399 ) | ( n40454 & ~n45399 ) ;
  assign n45402 = n34053 ^ n25070 ^ n19010 ;
  assign n45401 = ~n1682 & n8830 ;
  assign n45403 = n45402 ^ n45401 ^ 1'b0 ;
  assign n45404 = n871 | n45403 ;
  assign n45405 = n14123 ^ n6983 ^ 1'b0 ;
  assign n45406 = n13241 ^ n3874 ^ n732 ;
  assign n45407 = n13720 ^ n8927 ^ 1'b0 ;
  assign n45408 = ~n45406 & n45407 ;
  assign n45409 = ( n29180 & ~n33117 ) | ( n29180 & n45408 ) | ( ~n33117 & n45408 ) ;
  assign n45410 = n45058 ^ n33413 ^ n25273 ;
  assign n45411 = n6304 & n26724 ;
  assign n45412 = n45410 & n45411 ;
  assign n45413 = n39610 ^ n15774 ^ 1'b0 ;
  assign n45414 = ~n6984 & n45413 ;
  assign n45415 = ( n20881 & n25176 ) | ( n20881 & ~n35292 ) | ( n25176 & ~n35292 ) ;
  assign n45416 = ~n11366 & n45362 ;
  assign n45417 = n23710 & ~n45416 ;
  assign n45418 = n45415 & n45417 ;
  assign n45419 = n19303 | n22512 ;
  assign n45420 = n35532 ^ n16086 ^ 1'b0 ;
  assign n45421 = ~n3050 & n45420 ;
  assign n45422 = ( ~n44401 & n45419 ) | ( ~n44401 & n45421 ) | ( n45419 & n45421 ) ;
  assign n45429 = ( n7913 & ~n13315 ) | ( n7913 & n18564 ) | ( ~n13315 & n18564 ) ;
  assign n45430 = n21662 ^ n17855 ^ n11218 ;
  assign n45431 = ~n45429 & n45430 ;
  assign n45425 = n1754 | n4500 ;
  assign n45426 = n45425 ^ n25940 ^ n11678 ;
  assign n45427 = n39490 & ~n45426 ;
  assign n45428 = n45427 ^ n27851 ^ 1'b0 ;
  assign n45423 = n31824 ^ n5212 ^ 1'b0 ;
  assign n45424 = n42789 | n45423 ;
  assign n45432 = n45431 ^ n45428 ^ n45424 ;
  assign n45434 = n12768 ^ n10191 ^ n3767 ;
  assign n45433 = ( n1157 & n12089 ) | ( n1157 & ~n18887 ) | ( n12089 & ~n18887 ) ;
  assign n45435 = n45434 ^ n45433 ^ n37596 ;
  assign n45436 = n18008 ^ n9238 ^ 1'b0 ;
  assign n45437 = ( ~n24767 & n28478 ) | ( ~n24767 & n45436 ) | ( n28478 & n45436 ) ;
  assign n45438 = ( n30166 & n45435 ) | ( n30166 & ~n45437 ) | ( n45435 & ~n45437 ) ;
  assign n45439 = ( n14904 & ~n17540 ) | ( n14904 & n19855 ) | ( ~n17540 & n19855 ) ;
  assign n45440 = n45439 ^ n7003 ^ 1'b0 ;
  assign n45441 = n13674 ^ n10303 ^ n4095 ;
  assign n45442 = n11971 ^ n3290 ^ 1'b0 ;
  assign n45443 = n12008 ^ n9260 ^ 1'b0 ;
  assign n45444 = n18013 & n45443 ;
  assign n45445 = n11892 & ~n19053 ;
  assign n45449 = n36746 ^ n28503 ^ n13193 ;
  assign n45446 = n21139 ^ n8594 ^ 1'b0 ;
  assign n45447 = ~n25375 & n45446 ;
  assign n45448 = n1042 & n45447 ;
  assign n45450 = n45449 ^ n45448 ^ 1'b0 ;
  assign n45451 = n12213 ^ n10103 ^ n7955 ;
  assign n45452 = n7457 & ~n15500 ;
  assign n45453 = ~n30569 & n45452 ;
  assign n45454 = ( ~n13926 & n23254 ) | ( ~n13926 & n40041 ) | ( n23254 & n40041 ) ;
  assign n45455 = ( n16900 & ~n17077 ) | ( n16900 & n27335 ) | ( ~n17077 & n27335 ) ;
  assign n45456 = n9340 & n45455 ;
  assign n45457 = n26257 | n43358 ;
  assign n45458 = ~n31261 & n35082 ;
  assign n45459 = n3468 & ~n3832 ;
  assign n45460 = ( n10266 & n27705 ) | ( n10266 & n45459 ) | ( n27705 & n45459 ) ;
  assign n45461 = n11107 & n16595 ;
  assign n45462 = n43040 & n45461 ;
  assign n45463 = n45460 & n45462 ;
  assign n45464 = n17720 ^ n15014 ^ n9311 ;
  assign n45465 = n45464 ^ n16045 ^ 1'b0 ;
  assign n45466 = n5952 & n45465 ;
  assign n45467 = n45466 ^ n10244 ^ n8965 ;
  assign n45469 = n11062 ^ n3983 ^ 1'b0 ;
  assign n45470 = ~n7810 & n45469 ;
  assign n45468 = n26266 & n26909 ;
  assign n45471 = n45470 ^ n45468 ^ 1'b0 ;
  assign n45472 = n45471 ^ n22662 ^ 1'b0 ;
  assign n45473 = n40297 ^ n12200 ^ 1'b0 ;
  assign n45474 = ( n15546 & n29276 ) | ( n15546 & ~n34298 ) | ( n29276 & ~n34298 ) ;
  assign n45475 = n30745 ^ n16547 ^ n3923 ;
  assign n45476 = n15410 & n45475 ;
  assign n45477 = n3121 & ~n12481 ;
  assign n45478 = n45477 ^ n6209 ^ 1'b0 ;
  assign n45479 = ~n25246 & n45478 ;
  assign n45480 = n36063 ^ n18235 ^ 1'b0 ;
  assign n45481 = ~n22237 & n45480 ;
  assign n45482 = ( ~n45476 & n45479 ) | ( ~n45476 & n45481 ) | ( n45479 & n45481 ) ;
  assign n45483 = n25567 & n43336 ;
  assign n45484 = n11598 | n21837 ;
  assign n45485 = n45484 ^ n39138 ^ 1'b0 ;
  assign n45486 = n37637 & n45485 ;
  assign n45487 = n36372 ^ n27751 ^ n27628 ;
  assign n45488 = n1810 & ~n5402 ;
  assign n45489 = ~n3064 & n45488 ;
  assign n45490 = ( n10423 & n23976 ) | ( n10423 & n28430 ) | ( n23976 & n28430 ) ;
  assign n45491 = ( n615 & ~n17019 ) | ( n615 & n45490 ) | ( ~n17019 & n45490 ) ;
  assign n45492 = n23756 | n30665 ;
  assign n45495 = n21112 ^ n13979 ^ 1'b0 ;
  assign n45493 = n11092 ^ n896 ^ 1'b0 ;
  assign n45494 = n4498 & ~n45493 ;
  assign n45496 = n45495 ^ n45494 ^ n18013 ;
  assign n45497 = n38916 ^ n6761 ^ 1'b0 ;
  assign n45498 = ( n9087 & n16296 ) | ( n9087 & n19667 ) | ( n16296 & n19667 ) ;
  assign n45499 = n45498 ^ n23075 ^ 1'b0 ;
  assign n45500 = n15114 & n20501 ;
  assign n45501 = n45500 ^ n36561 ^ 1'b0 ;
  assign n45502 = n24883 ^ n21722 ^ 1'b0 ;
  assign n45503 = n17554 & n45502 ;
  assign n45504 = ( n11366 & n40014 ) | ( n11366 & ~n45503 ) | ( n40014 & ~n45503 ) ;
  assign n45505 = ( n14054 & ~n22693 ) | ( n14054 & n24018 ) | ( ~n22693 & n24018 ) ;
  assign n45507 = n24756 ^ n12196 ^ n1839 ;
  assign n45506 = n15474 & n34553 ;
  assign n45508 = n45507 ^ n45506 ^ 1'b0 ;
  assign n45509 = ~n11404 & n25584 ;
  assign n45510 = ~n45508 & n45509 ;
  assign n45511 = n12701 & n45510 ;
  assign n45512 = n3689 & ~n4946 ;
  assign n45513 = ~n3689 & n45512 ;
  assign n45514 = n45513 ^ n2146 ^ 1'b0 ;
  assign n45515 = n7729 & n45514 ;
  assign n45516 = n12089 & n16894 ;
  assign n45517 = n45516 ^ n12331 ^ 1'b0 ;
  assign n45518 = n11434 ^ n11329 ^ 1'b0 ;
  assign n45519 = ~n10887 & n45518 ;
  assign n45520 = n32963 ^ n26439 ^ n8302 ;
  assign n45521 = n30633 | n45520 ;
  assign n45522 = n6721 & ~n24382 ;
  assign n45523 = n45522 ^ n13724 ^ 1'b0 ;
  assign n45524 = n45523 ^ n40103 ^ n14097 ;
  assign n45525 = n44357 ^ n9329 ^ n8900 ;
  assign n45526 = n43076 ^ n11257 ^ n10716 ;
  assign n45528 = ( n13857 & ~n28186 ) | ( n13857 & n39139 ) | ( ~n28186 & n39139 ) ;
  assign n45529 = n45528 ^ n22423 ^ n12447 ;
  assign n45527 = n15256 ^ n3400 ^ 1'b0 ;
  assign n45530 = n45529 ^ n45527 ^ n7822 ;
  assign n45531 = n44459 ^ n14461 ^ 1'b0 ;
  assign n45532 = ( ~n477 & n11406 ) | ( ~n477 & n20778 ) | ( n11406 & n20778 ) ;
  assign n45533 = n41048 ^ n14745 ^ 1'b0 ;
  assign n45534 = n45532 | n45533 ;
  assign n45535 = ~n14902 & n33400 ;
  assign n45536 = n17191 & n45535 ;
  assign n45537 = n27360 ^ n16159 ^ n3164 ;
  assign n45538 = ( n8984 & n15769 ) | ( n8984 & n45537 ) | ( n15769 & n45537 ) ;
  assign n45539 = ~n27196 & n43889 ;
  assign n45540 = n45539 ^ n14244 ^ 1'b0 ;
  assign n45541 = n45540 ^ n39234 ^ n5533 ;
  assign n45544 = ( n1442 & n20068 ) | ( n1442 & ~n22062 ) | ( n20068 & ~n22062 ) ;
  assign n45542 = ~n14244 & n26464 ;
  assign n45543 = n45542 ^ n18133 ^ 1'b0 ;
  assign n45545 = n45544 ^ n45543 ^ n5182 ;
  assign n45546 = ( ~n6704 & n11021 ) | ( ~n6704 & n29844 ) | ( n11021 & n29844 ) ;
  assign n45547 = ( n19842 & n20621 ) | ( n19842 & n45546 ) | ( n20621 & n45546 ) ;
  assign n45548 = n23220 & ~n24965 ;
  assign n45551 = n16298 & ~n36303 ;
  assign n45552 = ( ~n13336 & n28954 ) | ( ~n13336 & n45551 ) | ( n28954 & n45551 ) ;
  assign n45553 = n19751 & n22101 ;
  assign n45554 = ( ~n34675 & n45552 ) | ( ~n34675 & n45553 ) | ( n45552 & n45553 ) ;
  assign n45549 = n23612 ^ n9429 ^ 1'b0 ;
  assign n45550 = n27912 | n45549 ;
  assign n45555 = n45554 ^ n45550 ^ n3864 ;
  assign n45556 = ( ~n18192 & n45548 ) | ( ~n18192 & n45555 ) | ( n45548 & n45555 ) ;
  assign n45557 = ( ~n5515 & n37823 ) | ( ~n5515 & n45556 ) | ( n37823 & n45556 ) ;
  assign n45558 = n13680 ^ n10604 ^ 1'b0 ;
  assign n45559 = ( ~n4858 & n28860 ) | ( ~n4858 & n45558 ) | ( n28860 & n45558 ) ;
  assign n45560 = ( n17198 & ~n30894 ) | ( n17198 & n45559 ) | ( ~n30894 & n45559 ) ;
  assign n45561 = n45560 ^ n20222 ^ 1'b0 ;
  assign n45562 = ~n15311 & n45561 ;
  assign n45563 = ( n711 & n2329 ) | ( n711 & n4960 ) | ( n2329 & n4960 ) ;
  assign n45564 = n28651 & n45563 ;
  assign n45565 = n12688 & n33946 ;
  assign n45566 = n20802 | n35456 ;
  assign n45567 = n45565 | n45566 ;
  assign n45568 = n10336 & n20086 ;
  assign n45569 = ( n1447 & ~n17637 ) | ( n1447 & n20019 ) | ( ~n17637 & n20019 ) ;
  assign n45570 = n10563 ^ n10454 ^ 1'b0 ;
  assign n45571 = n36717 & n45570 ;
  assign n45572 = n20135 ^ n1756 ^ n592 ;
  assign n45573 = n478 & n3221 ;
  assign n45574 = n45573 ^ n7904 ^ 1'b0 ;
  assign n45575 = ( ~n14258 & n15092 ) | ( ~n14258 & n45574 ) | ( n15092 & n45574 ) ;
  assign n45576 = ~n12341 & n17917 ;
  assign n45577 = n45576 ^ n7310 ^ 1'b0 ;
  assign n45578 = n3697 & n33094 ;
  assign n45579 = n9390 & n45578 ;
  assign n45580 = n18477 & ~n22237 ;
  assign n45581 = n11995 & n45580 ;
  assign n45582 = ~n7396 & n20091 ;
  assign n45583 = n45582 ^ n12370 ^ 1'b0 ;
  assign n45584 = n4841 & ~n45583 ;
  assign n45585 = n45584 ^ n10139 ^ 1'b0 ;
  assign n45586 = ~n2315 & n21034 ;
  assign n45587 = ( n2317 & n4084 ) | ( n2317 & ~n29433 ) | ( n4084 & ~n29433 ) ;
  assign n45588 = n11583 & n12821 ;
  assign n45589 = n45588 ^ n31116 ^ 1'b0 ;
  assign n45590 = n45589 ^ n36787 ^ n26202 ;
  assign n45591 = n45248 ^ n28870 ^ n15852 ;
  assign n45592 = n38034 ^ n662 ^ 1'b0 ;
  assign n45593 = n31669 ^ n31185 ^ n10192 ;
  assign n45596 = n9134 & ~n32283 ;
  assign n45597 = ( n27475 & n42437 ) | ( n27475 & ~n45596 ) | ( n42437 & ~n45596 ) ;
  assign n45594 = n16451 ^ n14550 ^ x129 ;
  assign n45595 = n2501 & ~n45594 ;
  assign n45598 = n45597 ^ n45595 ^ 1'b0 ;
  assign n45600 = ( n2639 & n27892 ) | ( n2639 & ~n28060 ) | ( n27892 & ~n28060 ) ;
  assign n45599 = n4981 | n21190 ;
  assign n45601 = n45600 ^ n45599 ^ 1'b0 ;
  assign n45602 = n10326 & ~n45601 ;
  assign n45603 = n45602 ^ n45503 ^ 1'b0 ;
  assign n45604 = n44192 ^ n31488 ^ n14767 ;
  assign n45605 = n3927 & ~n34387 ;
  assign n45606 = n45605 ^ n40103 ^ 1'b0 ;
  assign n45607 = ( n9509 & n17753 ) | ( n9509 & ~n45606 ) | ( n17753 & ~n45606 ) ;
  assign n45608 = n25948 ^ n11881 ^ 1'b0 ;
  assign n45609 = n27658 & ~n34284 ;
  assign n45610 = ~n27495 & n45609 ;
  assign n45612 = n26162 ^ n13014 ^ n1297 ;
  assign n45611 = n13148 | n34435 ;
  assign n45613 = n45612 ^ n45611 ^ 1'b0 ;
  assign n45614 = n7217 | n10372 ;
  assign n45615 = n45614 ^ n7821 ^ 1'b0 ;
  assign n45616 = n5871 & ~n45615 ;
  assign n45617 = n18889 & n45616 ;
  assign n45618 = ~n7295 & n45617 ;
  assign n45619 = n11129 & n36542 ;
  assign n45620 = n42983 & n45619 ;
  assign n45621 = n24680 & ~n41014 ;
  assign n45622 = n38518 ^ n2279 ^ 1'b0 ;
  assign n45623 = n45622 ^ n28936 ^ n11166 ;
  assign n45624 = n41277 ^ n37879 ^ n25548 ;
  assign n45625 = n32274 ^ n27940 ^ 1'b0 ;
  assign n45626 = ( n24890 & ~n26702 ) | ( n24890 & n30022 ) | ( ~n26702 & n30022 ) ;
  assign n45627 = n35472 ^ n12141 ^ 1'b0 ;
  assign n45628 = n20639 | n45627 ;
  assign n45629 = ~n5642 & n11244 ;
  assign n45630 = ~n15917 & n45629 ;
  assign n45631 = n22370 ^ n11290 ^ 1'b0 ;
  assign n45632 = ~n34605 & n45631 ;
  assign n45633 = ~n3083 & n45632 ;
  assign n45634 = n45633 ^ n30714 ^ 1'b0 ;
  assign n45635 = n16501 & n21204 ;
  assign n45636 = n20317 & n45635 ;
  assign n45637 = n36868 | n45636 ;
  assign n45638 = ( n3324 & n9167 ) | ( n3324 & n14789 ) | ( n9167 & n14789 ) ;
  assign n45639 = n45638 ^ n42709 ^ n12007 ;
  assign n45640 = n17696 ^ n5917 ^ 1'b0 ;
  assign n45641 = n28537 ^ n12915 ^ 1'b0 ;
  assign n45642 = ~n45640 & n45641 ;
  assign n45643 = n45642 ^ n21378 ^ 1'b0 ;
  assign n45644 = n1604 | n2873 ;
  assign n45645 = n45644 ^ n27763 ^ n8553 ;
  assign n45646 = ( n14995 & ~n24181 ) | ( n14995 & n32749 ) | ( ~n24181 & n32749 ) ;
  assign n45647 = n45646 ^ n22339 ^ n10926 ;
  assign n45648 = ( n14150 & n24674 ) | ( n14150 & n43800 ) | ( n24674 & n43800 ) ;
  assign n45649 = ( n3436 & ~n16923 ) | ( n3436 & n42868 ) | ( ~n16923 & n42868 ) ;
  assign n45650 = n2511 | n45649 ;
  assign n45651 = n17440 & ~n45650 ;
  assign n45652 = n18491 | n45651 ;
  assign n45653 = n42984 ^ n13486 ^ 1'b0 ;
  assign n45654 = n34299 | n45653 ;
  assign n45655 = n31225 | n45654 ;
  assign n45656 = ~n36486 & n42409 ;
  assign n45657 = n45656 ^ n14260 ^ n3616 ;
  assign n45658 = ~n13085 & n16073 ;
  assign n45659 = n45657 & n45658 ;
  assign n45660 = n6166 | n32438 ;
  assign n45661 = n16839 | n45660 ;
  assign n45662 = n8386 & n17452 ;
  assign n45663 = n45662 ^ n22801 ^ 1'b0 ;
  assign n45664 = ( ~n21533 & n23072 ) | ( ~n21533 & n45663 ) | ( n23072 & n45663 ) ;
  assign n45670 = n12394 ^ n11619 ^ 1'b0 ;
  assign n45671 = n8084 & n45670 ;
  assign n45672 = n45671 ^ n27384 ^ n5018 ;
  assign n45668 = n12759 & ~n32704 ;
  assign n45669 = n7618 & n45668 ;
  assign n45665 = n3671 & ~n13803 ;
  assign n45666 = n28899 & n45665 ;
  assign n45667 = ( n16920 & ~n19157 ) | ( n16920 & n45666 ) | ( ~n19157 & n45666 ) ;
  assign n45673 = n45672 ^ n45669 ^ n45667 ;
  assign n45674 = ( ~n4839 & n23680 ) | ( ~n4839 & n41894 ) | ( n23680 & n41894 ) ;
  assign n45676 = n3562 ^ n1694 ^ 1'b0 ;
  assign n45677 = n1815 | n45676 ;
  assign n45675 = n36680 ^ n29525 ^ n25058 ;
  assign n45678 = n45677 ^ n45675 ^ n26202 ;
  assign n45679 = n1949 | n14978 ;
  assign n45680 = n8980 | n21470 ;
  assign n45681 = n10809 ^ n4745 ^ 1'b0 ;
  assign n45682 = ( n403 & n3752 ) | ( n403 & ~n6439 ) | ( n3752 & ~n6439 ) ;
  assign n45683 = n29823 & ~n31180 ;
  assign n45684 = n25645 ^ n17343 ^ 1'b0 ;
  assign n45685 = n45684 ^ n15234 ^ 1'b0 ;
  assign n45686 = n40844 ^ n38918 ^ 1'b0 ;
  assign n45687 = n5224 & ~n45686 ;
  assign n45688 = n8723 ^ n7633 ^ n6621 ;
  assign n45689 = ( n37883 & n45687 ) | ( n37883 & n45688 ) | ( n45687 & n45688 ) ;
  assign n45690 = n33284 ^ n20590 ^ 1'b0 ;
  assign n45691 = n45690 ^ n38987 ^ n37761 ;
  assign n45692 = ~n4892 & n13847 ;
  assign n45693 = n45692 ^ n7019 ^ 1'b0 ;
  assign n45694 = ~n9917 & n45693 ;
  assign n45695 = n45691 & n45694 ;
  assign n45696 = ( ~n1139 & n1157 ) | ( ~n1139 & n10013 ) | ( n1157 & n10013 ) ;
  assign n45697 = n45696 ^ n22237 ^ n10338 ;
  assign n45698 = n14890 & ~n30578 ;
  assign n45699 = ~n30537 & n45698 ;
  assign n45700 = n35234 | n45699 ;
  assign n45701 = n45697 & ~n45700 ;
  assign n45702 = n2124 & ~n5205 ;
  assign n45703 = n5205 & n45702 ;
  assign n45704 = n40862 | n45703 ;
  assign n45705 = n45704 ^ n22350 ^ 1'b0 ;
  assign n45710 = ( ~n1104 & n2544 ) | ( ~n1104 & n38349 ) | ( n2544 & n38349 ) ;
  assign n45709 = n20135 ^ n3644 ^ n2123 ;
  assign n45706 = ( n3148 & ~n5730 ) | ( n3148 & n36868 ) | ( ~n5730 & n36868 ) ;
  assign n45707 = n38985 ^ n18207 ^ n15810 ;
  assign n45708 = ( n11861 & n45706 ) | ( n11861 & n45707 ) | ( n45706 & n45707 ) ;
  assign n45711 = n45710 ^ n45709 ^ n45708 ;
  assign n45712 = n23709 | n43042 ;
  assign n45713 = ( n21149 & n37730 ) | ( n21149 & ~n45712 ) | ( n37730 & ~n45712 ) ;
  assign n45714 = n44127 ^ n31457 ^ n11422 ;
  assign n45715 = n25192 & ~n37868 ;
  assign n45716 = n45714 & n45715 ;
  assign n45717 = ( n14842 & n38612 ) | ( n14842 & ~n45716 ) | ( n38612 & ~n45716 ) ;
  assign n45718 = n37613 ^ n22757 ^ 1'b0 ;
  assign n45719 = n45718 ^ n39662 ^ n24438 ;
  assign n45720 = n29592 | n31524 ;
  assign n45721 = n19933 | n45720 ;
  assign n45722 = ~n21627 & n38396 ;
  assign n45723 = ( ~n8414 & n14548 ) | ( ~n8414 & n21017 ) | ( n14548 & n21017 ) ;
  assign n45724 = ( n737 & ~n20304 ) | ( n737 & n45723 ) | ( ~n20304 & n45723 ) ;
  assign n45725 = n3455 | n8056 ;
  assign n45726 = ~n559 & n45725 ;
  assign n45727 = n20310 & ~n28065 ;
  assign n45728 = n18640 ^ n8880 ^ 1'b0 ;
  assign n45729 = n45727 & n45728 ;
  assign n45730 = n45729 ^ n12216 ^ n7679 ;
  assign n45731 = n25524 ^ n11990 ^ 1'b0 ;
  assign n45732 = n17174 ^ n4203 ^ 1'b0 ;
  assign n45733 = n22200 ^ n8415 ^ n1162 ;
  assign n45734 = n3426 & n24734 ;
  assign n45735 = ~n45733 & n45734 ;
  assign n45736 = n16739 & ~n43306 ;
  assign n45737 = n45736 ^ n11650 ^ 1'b0 ;
  assign n45738 = ~n26331 & n43333 ;
  assign n45739 = n45738 ^ n514 ^ 1'b0 ;
  assign n45740 = n20272 ^ x171 ^ 1'b0 ;
  assign n45741 = ( n16918 & n31449 ) | ( n16918 & ~n45740 ) | ( n31449 & ~n45740 ) ;
  assign n45742 = ( ~n18342 & n25176 ) | ( ~n18342 & n43433 ) | ( n25176 & n43433 ) ;
  assign n45743 = n40592 ^ n26237 ^ n24004 ;
  assign n45744 = ~n1010 & n27587 ;
  assign n45745 = n2230 & ~n45744 ;
  assign n45746 = ( n7746 & n7754 ) | ( n7746 & ~n36768 ) | ( n7754 & ~n36768 ) ;
  assign n45747 = n14629 & n24698 ;
  assign n45748 = ( n1953 & ~n6589 ) | ( n1953 & n9865 ) | ( ~n6589 & n9865 ) ;
  assign n45749 = n45748 ^ n29127 ^ 1'b0 ;
  assign n45750 = n6888 | n16519 ;
  assign n45751 = n45750 ^ n40103 ^ 1'b0 ;
  assign n45752 = n28384 ^ n27637 ^ n4053 ;
  assign n45753 = n6811 | n9475 ;
  assign n45754 = n45753 ^ n2832 ^ 1'b0 ;
  assign n45755 = n45084 ^ n30255 ^ n7693 ;
  assign n45756 = ( n45752 & n45754 ) | ( n45752 & n45755 ) | ( n45754 & n45755 ) ;
  assign n45757 = n19642 ^ n18778 ^ n1156 ;
  assign n45758 = ( n3229 & ~n16357 ) | ( n3229 & n42718 ) | ( ~n16357 & n42718 ) ;
  assign n45759 = ( n3906 & n3994 ) | ( n3906 & ~n4271 ) | ( n3994 & ~n4271 ) ;
  assign n45760 = ~n12794 & n45759 ;
  assign n45761 = n19982 ^ n14185 ^ n10710 ;
  assign n45762 = ( n17391 & ~n32985 ) | ( n17391 & n45761 ) | ( ~n32985 & n45761 ) ;
  assign n45763 = ( ~n5171 & n6266 ) | ( ~n5171 & n24705 ) | ( n6266 & n24705 ) ;
  assign n45764 = ( ~n2669 & n43238 ) | ( ~n2669 & n45763 ) | ( n43238 & n45763 ) ;
  assign n45765 = n10462 ^ n8777 ^ 1'b0 ;
  assign n45766 = ~n29584 & n45765 ;
  assign n45767 = n18795 ^ n17234 ^ 1'b0 ;
  assign n45768 = n32665 | n45767 ;
  assign n45769 = ~n2080 & n36836 ;
  assign n45770 = n45769 ^ n42897 ^ n31923 ;
  assign n45771 = n45770 ^ n2624 ^ 1'b0 ;
  assign n45772 = ( n10831 & n31069 ) | ( n10831 & ~n36317 ) | ( n31069 & ~n36317 ) ;
  assign n45773 = n45772 ^ n23064 ^ 1'b0 ;
  assign n45774 = ~n45771 & n45773 ;
  assign n45775 = n34419 ^ n18312 ^ 1'b0 ;
  assign n45776 = ~n13022 & n45775 ;
  assign n45777 = ~n36502 & n45776 ;
  assign n45778 = n27806 & n45777 ;
  assign n45779 = n19443 ^ n18789 ^ 1'b0 ;
  assign n45780 = ~n45778 & n45779 ;
  assign n45781 = ( n5889 & n9390 ) | ( n5889 & ~n13836 ) | ( n9390 & ~n13836 ) ;
  assign n45782 = n17854 & ~n25974 ;
  assign n45783 = n45782 ^ n18167 ^ 1'b0 ;
  assign n45784 = ( n20677 & ~n45781 ) | ( n20677 & n45783 ) | ( ~n45781 & n45783 ) ;
  assign n45785 = n10163 ^ n7633 ^ n6819 ;
  assign n45786 = ( n14232 & n17129 ) | ( n14232 & ~n45785 ) | ( n17129 & ~n45785 ) ;
  assign n45787 = n43063 & n45786 ;
  assign n45788 = ( n2787 & n12970 ) | ( n2787 & n16964 ) | ( n12970 & n16964 ) ;
  assign n45789 = n10032 & ~n45788 ;
  assign n45790 = n32624 ^ n5153 ^ n1282 ;
  assign n45791 = n24894 & ~n45790 ;
  assign n45794 = n12201 | n44078 ;
  assign n45792 = ( ~n12175 & n20747 ) | ( ~n12175 & n21672 ) | ( n20747 & n21672 ) ;
  assign n45793 = ~n33772 & n45792 ;
  assign n45795 = n45794 ^ n45793 ^ 1'b0 ;
  assign n45796 = n5717 | n6897 ;
  assign n45797 = n28597 & ~n45796 ;
  assign n45798 = ( n3090 & n36016 ) | ( n3090 & ~n45797 ) | ( n36016 & ~n45797 ) ;
  assign n45799 = n35011 ^ n27326 ^ 1'b0 ;
  assign n45800 = n17872 | n45799 ;
  assign n45801 = ~n2662 & n17976 ;
  assign n45802 = n7675 | n15642 ;
  assign n45803 = n40442 ^ n16695 ^ 1'b0 ;
  assign n45804 = ~n45802 & n45803 ;
  assign n45805 = n33013 ^ n3290 ^ 1'b0 ;
  assign n45806 = n17593 | n45805 ;
  assign n45807 = n45168 ^ n6476 ^ 1'b0 ;
  assign n45808 = n1403 & ~n45807 ;
  assign n45809 = n32611 ^ n19154 ^ n6080 ;
  assign n45810 = n5786 & n11838 ;
  assign n45811 = n17853 & ~n18832 ;
  assign n45812 = n45811 ^ n42955 ^ n2440 ;
  assign n45813 = n20546 ^ n18436 ^ 1'b0 ;
  assign n45814 = n10863 & n45813 ;
  assign n45815 = n1544 & ~n45814 ;
  assign n45818 = n30126 ^ n13512 ^ 1'b0 ;
  assign n45819 = ~n29183 & n45818 ;
  assign n45816 = ( ~n18853 & n19187 ) | ( ~n18853 & n40120 ) | ( n19187 & n40120 ) ;
  assign n45817 = n2378 & ~n45816 ;
  assign n45820 = n45819 ^ n45817 ^ 1'b0 ;
  assign n45821 = n17935 ^ n14134 ^ 1'b0 ;
  assign n45822 = n17496 & ~n45821 ;
  assign n45823 = n37265 | n40415 ;
  assign n45824 = n973 & ~n45823 ;
  assign n45825 = ~n18929 & n27279 ;
  assign n45830 = ( n13645 & ~n16143 ) | ( n13645 & n25079 ) | ( ~n16143 & n25079 ) ;
  assign n45826 = n4222 ^ n2997 ^ 1'b0 ;
  assign n45827 = n725 & ~n45826 ;
  assign n45828 = n45827 ^ n5901 ^ 1'b0 ;
  assign n45829 = ~n17130 & n45828 ;
  assign n45831 = n45830 ^ n45829 ^ 1'b0 ;
  assign n45832 = ( ~n9680 & n36824 ) | ( ~n9680 & n45831 ) | ( n36824 & n45831 ) ;
  assign n45834 = n8581 ^ n7588 ^ n4902 ;
  assign n45833 = n21781 ^ n21766 ^ n9976 ;
  assign n45835 = n45834 ^ n45833 ^ n17681 ;
  assign n45836 = n41174 ^ n29027 ^ n1796 ;
  assign n45837 = n6673 ^ n3385 ^ n1198 ;
  assign n45838 = ( ~n32093 & n36691 ) | ( ~n32093 & n45837 ) | ( n36691 & n45837 ) ;
  assign n45839 = n6076 | n45838 ;
  assign n45840 = n45839 ^ n10045 ^ 1'b0 ;
  assign n45841 = n45840 ^ n30651 ^ n6888 ;
  assign n45842 = ( n10915 & ~n17449 ) | ( n10915 & n33797 ) | ( ~n17449 & n33797 ) ;
  assign n45843 = ( n12572 & ~n19648 ) | ( n12572 & n45842 ) | ( ~n19648 & n45842 ) ;
  assign n45844 = n25174 & ~n41153 ;
  assign n45845 = n45844 ^ n6482 ^ 1'b0 ;
  assign n45846 = n40626 ^ n25475 ^ 1'b0 ;
  assign n45847 = ~n39567 & n45846 ;
  assign n45848 = n7881 & ~n20581 ;
  assign n45849 = n31675 ^ n30814 ^ n2096 ;
  assign n45850 = ( n18132 & n23452 ) | ( n18132 & n25310 ) | ( n23452 & n25310 ) ;
  assign n45851 = n29049 ^ n2824 ^ n2313 ;
  assign n45852 = n16288 & ~n45851 ;
  assign n45853 = n26276 ^ n12472 ^ n803 ;
  assign n45854 = ( x117 & n23039 ) | ( x117 & ~n45853 ) | ( n23039 & ~n45853 ) ;
  assign n45855 = ~n4676 & n33554 ;
  assign n45856 = n45855 ^ n18058 ^ 1'b0 ;
  assign n45857 = n41063 ^ n6281 ^ 1'b0 ;
  assign n45858 = n19916 ^ n9286 ^ 1'b0 ;
  assign n45859 = n45857 | n45858 ;
  assign n45860 = n5132 ^ n721 ^ 1'b0 ;
  assign n45861 = ~n6333 & n45860 ;
  assign n45862 = ( n8644 & n16051 ) | ( n8644 & n45861 ) | ( n16051 & n45861 ) ;
  assign n45863 = n24913 ^ n15422 ^ x247 ;
  assign n45864 = ( n29858 & n44909 ) | ( n29858 & ~n45863 ) | ( n44909 & ~n45863 ) ;
  assign n45865 = n14262 & ~n19583 ;
  assign n45866 = n45865 ^ n5278 ^ 1'b0 ;
  assign n45867 = n45866 ^ n8466 ^ 1'b0 ;
  assign n45868 = n44303 ^ n36433 ^ n26573 ;
  assign n45869 = n45868 ^ n21034 ^ n18795 ;
  assign n45873 = ~n13877 & n22815 ;
  assign n45874 = n45873 ^ n16125 ^ 1'b0 ;
  assign n45870 = n40995 ^ n6136 ^ 1'b0 ;
  assign n45871 = n7697 & n37738 ;
  assign n45872 = ~n45870 & n45871 ;
  assign n45875 = n45874 ^ n45872 ^ n31170 ;
  assign n45876 = n788 & ~n27196 ;
  assign n45877 = n6657 ^ n1709 ^ n866 ;
  assign n45878 = n17780 & n45877 ;
  assign n45879 = n41806 & n45878 ;
  assign n45880 = n23118 & n28363 ;
  assign n45881 = n14033 & n45880 ;
  assign n45883 = n12000 ^ n959 ^ 1'b0 ;
  assign n45884 = n45883 ^ n35870 ^ n15496 ;
  assign n45885 = n45884 ^ n14883 ^ n1162 ;
  assign n45886 = ( n8076 & n37040 ) | ( n8076 & ~n45885 ) | ( n37040 & ~n45885 ) ;
  assign n45887 = ( n17979 & n22660 ) | ( n17979 & n25893 ) | ( n22660 & n25893 ) ;
  assign n45888 = n27751 & n45887 ;
  assign n45889 = ~n45886 & n45888 ;
  assign n45882 = n15745 & n33361 ;
  assign n45890 = n45889 ^ n45882 ^ n1545 ;
  assign n45891 = n18800 ^ n14916 ^ 1'b0 ;
  assign n45892 = n45891 ^ n29280 ^ n29040 ;
  assign n45893 = n44108 ^ n15993 ^ n9328 ;
  assign n45894 = n24472 & ~n43722 ;
  assign n45895 = n35046 ^ n5108 ^ 1'b0 ;
  assign n45896 = n34308 & n45895 ;
  assign n45897 = n2492 | n8978 ;
  assign n45898 = n9781 | n45897 ;
  assign n45899 = ~n22011 & n45898 ;
  assign n45900 = n45899 ^ n26285 ^ 1'b0 ;
  assign n45901 = n27554 ^ n22458 ^ 1'b0 ;
  assign n45902 = n24229 & n45901 ;
  assign n45903 = ( n1969 & n22928 ) | ( n1969 & n45062 ) | ( n22928 & n45062 ) ;
  assign n45904 = n30615 ^ n18776 ^ n1495 ;
  assign n45905 = n33847 ^ n11974 ^ n6376 ;
  assign n45906 = ( n45903 & ~n45904 ) | ( n45903 & n45905 ) | ( ~n45904 & n45905 ) ;
  assign n45907 = ( ~n5076 & n19443 ) | ( ~n5076 & n35062 ) | ( n19443 & n35062 ) ;
  assign n45908 = n20866 ^ n8148 ^ n2290 ;
  assign n45909 = n45908 ^ n33993 ^ n15144 ;
  assign n45910 = n15109 | n23169 ;
  assign n45911 = n45910 ^ n29972 ^ 1'b0 ;
  assign n45912 = n28865 & n31064 ;
  assign n45913 = ~n2627 & n45912 ;
  assign n45914 = ( n16969 & n37528 ) | ( n16969 & n45913 ) | ( n37528 & n45913 ) ;
  assign n45915 = n26043 | n45914 ;
  assign n45916 = n45915 ^ n17809 ^ 1'b0 ;
  assign n45917 = n39195 & ~n43135 ;
  assign n45918 = ~n18375 & n45917 ;
  assign n45919 = ( ~n8810 & n24966 ) | ( ~n8810 & n28605 ) | ( n24966 & n28605 ) ;
  assign n45920 = n45919 ^ n22430 ^ 1'b0 ;
  assign n45921 = n31795 ^ n17076 ^ 1'b0 ;
  assign n45922 = n14339 ^ n4117 ^ 1'b0 ;
  assign n45923 = n45921 | n45922 ;
  assign n45924 = n35712 ^ n17775 ^ n15282 ;
  assign n45925 = ( ~n15229 & n16873 ) | ( ~n15229 & n45924 ) | ( n16873 & n45924 ) ;
  assign n45926 = n21421 & n28225 ;
  assign n45927 = n2493 & ~n11308 ;
  assign n45928 = ( ~n27302 & n28051 ) | ( ~n27302 & n45927 ) | ( n28051 & n45927 ) ;
  assign n45929 = n44357 ^ n31619 ^ 1'b0 ;
  assign n45930 = n11585 & ~n13698 ;
  assign n45931 = n18025 & n45930 ;
  assign n45932 = n45931 ^ n25273 ^ 1'b0 ;
  assign n45933 = ( n9031 & n28648 ) | ( n9031 & ~n45932 ) | ( n28648 & ~n45932 ) ;
  assign n45934 = n12647 | n28976 ;
  assign n45935 = n45934 ^ n14021 ^ 1'b0 ;
  assign n45936 = n18876 & n24447 ;
  assign n45937 = n45710 & n45936 ;
  assign n45938 = n21683 ^ n6946 ^ 1'b0 ;
  assign n45939 = n44144 & ~n45938 ;
  assign n45940 = ( n10451 & ~n14630 ) | ( n10451 & n17503 ) | ( ~n14630 & n17503 ) ;
  assign n45941 = n45940 ^ n1004 ^ 1'b0 ;
  assign n45942 = n5958 & ~n30788 ;
  assign n45943 = n45942 ^ n1867 ^ 1'b0 ;
  assign n45944 = n45943 ^ n21578 ^ n19472 ;
  assign n45945 = ~n11821 & n45283 ;
  assign n45946 = n7007 | n7101 ;
  assign n45947 = n20748 | n45946 ;
  assign n45948 = ( n15560 & ~n45213 ) | ( n15560 & n45947 ) | ( ~n45213 & n45947 ) ;
  assign n45949 = n20493 ^ n12399 ^ n12097 ;
  assign n45950 = n45949 ^ n37138 ^ 1'b0 ;
  assign n45951 = n43978 & ~n45950 ;
  assign n45952 = n8817 & ~n30703 ;
  assign n45953 = n45952 ^ n43640 ^ 1'b0 ;
  assign n45954 = n29381 ^ n10295 ^ 1'b0 ;
  assign n45955 = n13648 & n45954 ;
  assign n45956 = n45955 ^ n12658 ^ 1'b0 ;
  assign n45957 = ~n29833 & n30963 ;
  assign n45958 = n1400 & n12616 ;
  assign n45959 = n30537 ^ n24480 ^ n18436 ;
  assign n45960 = n10628 ^ n2908 ^ 1'b0 ;
  assign n45961 = n11196 ^ n7817 ^ 1'b0 ;
  assign n45962 = n3612 & n45961 ;
  assign n45963 = n21718 | n45962 ;
  assign n45964 = n15971 ^ n9786 ^ 1'b0 ;
  assign n45965 = ( ~n16781 & n17221 ) | ( ~n16781 & n31613 ) | ( n17221 & n31613 ) ;
  assign n45966 = n20100 & ~n25483 ;
  assign n45967 = ~n45965 & n45966 ;
  assign n45968 = n6312 | n6342 ;
  assign n45969 = n4136 | n45968 ;
  assign n45973 = n4729 | n6709 ;
  assign n45974 = n14418 & ~n45973 ;
  assign n45970 = n22391 ^ n6399 ^ 1'b0 ;
  assign n45971 = n32320 & n45970 ;
  assign n45972 = n11756 & ~n45971 ;
  assign n45975 = n45974 ^ n45972 ^ n9261 ;
  assign n45976 = n15495 ^ n11962 ^ n2877 ;
  assign n45977 = n45976 ^ n18306 ^ 1'b0 ;
  assign n45978 = ( n10443 & n11038 ) | ( n10443 & ~n15296 ) | ( n11038 & ~n15296 ) ;
  assign n45979 = ( n11189 & n43588 ) | ( n11189 & n45978 ) | ( n43588 & n45978 ) ;
  assign n45982 = n18157 & n26716 ;
  assign n45983 = n45982 ^ n18542 ^ 1'b0 ;
  assign n45980 = ~n1111 & n4816 ;
  assign n45981 = n45980 ^ n21791 ^ 1'b0 ;
  assign n45984 = n45983 ^ n45981 ^ 1'b0 ;
  assign n45985 = ( n7531 & n25795 ) | ( n7531 & ~n45749 ) | ( n25795 & ~n45749 ) ;
  assign n45986 = n20119 ^ n18144 ^ n5779 ;
  assign n45987 = n3472 & n3814 ;
  assign n45988 = n9349 & n22426 ;
  assign n45989 = n45988 ^ n20879 ^ 1'b0 ;
  assign n45990 = ~n11263 & n34448 ;
  assign n45991 = n32807 ^ n4213 ^ 1'b0 ;
  assign n45992 = ~n9096 & n10641 ;
  assign n45993 = n45992 ^ n22145 ^ 1'b0 ;
  assign n45994 = n45993 ^ n8374 ^ n5028 ;
  assign n45995 = n45994 ^ n34071 ^ 1'b0 ;
  assign n45996 = n10849 | n45529 ;
  assign n45997 = n29587 ^ n10667 ^ n6037 ;
  assign n45999 = n31564 ^ n21652 ^ n18940 ;
  assign n45998 = ~n6705 & n22382 ;
  assign n46000 = n45999 ^ n45998 ^ 1'b0 ;
  assign n46001 = n8475 ^ n6450 ^ n1249 ;
  assign n46002 = n46001 ^ n13722 ^ n11643 ;
  assign n46003 = ~n314 & n46002 ;
  assign n46004 = n46003 ^ n30486 ^ 1'b0 ;
  assign n46005 = n34820 ^ n29274 ^ n5316 ;
  assign n46006 = n46005 ^ n23312 ^ 1'b0 ;
  assign n46007 = ~n40659 & n46006 ;
  assign n46008 = ~n30096 & n30406 ;
  assign n46009 = ~n3775 & n17477 ;
  assign n46010 = ( ~n2707 & n16789 ) | ( ~n2707 & n21235 ) | ( n16789 & n21235 ) ;
  assign n46014 = n25174 ^ n22931 ^ n15264 ;
  assign n46013 = n18384 & n19757 ;
  assign n46015 = n46014 ^ n46013 ^ 1'b0 ;
  assign n46011 = n33874 ^ n31922 ^ n29215 ;
  assign n46012 = n46011 ^ n1328 ^ 1'b0 ;
  assign n46016 = n46015 ^ n46012 ^ n1722 ;
  assign n46017 = n26036 & ~n30647 ;
  assign n46018 = n39037 ^ n11649 ^ n4772 ;
  assign n46019 = n27121 ^ n6124 ^ x48 ;
  assign n46020 = n9760 ^ n805 ^ 1'b0 ;
  assign n46021 = ~n2515 & n46020 ;
  assign n46022 = n46021 ^ n1861 ^ 1'b0 ;
  assign n46023 = ( n8011 & ~n35291 ) | ( n8011 & n44281 ) | ( ~n35291 & n44281 ) ;
  assign n46024 = ( n1135 & n2384 ) | ( n1135 & n38311 ) | ( n2384 & n38311 ) ;
  assign n46025 = n46024 ^ n43469 ^ n4723 ;
  assign n46026 = n1472 | n25027 ;
  assign n46027 = n16311 & ~n46026 ;
  assign n46028 = n46027 ^ n23680 ^ n1375 ;
  assign n46029 = ( n13224 & n18388 ) | ( n13224 & n40148 ) | ( n18388 & n40148 ) ;
  assign n46030 = n42827 ^ n29364 ^ n22129 ;
  assign n46031 = n46030 ^ n18710 ^ n12621 ;
  assign n46032 = ( n8960 & n32782 ) | ( n8960 & n34122 ) | ( n32782 & n34122 ) ;
  assign n46033 = n25940 ^ n1631 ^ 1'b0 ;
  assign n46034 = n10773 & n46033 ;
  assign n46035 = n24005 ^ n3317 ^ n512 ;
  assign n46036 = ( ~n19133 & n30476 ) | ( ~n19133 & n46035 ) | ( n30476 & n46035 ) ;
  assign n46037 = ~n37141 & n46036 ;
  assign n46038 = n34832 & n46037 ;
  assign n46039 = n1325 & ~n46038 ;
  assign n46040 = n25908 & n46039 ;
  assign n46041 = n5337 & ~n46040 ;
  assign n46042 = n40950 & n46041 ;
  assign n46043 = n22629 ^ n4004 ^ 1'b0 ;
  assign n46044 = n46043 ^ n14967 ^ 1'b0 ;
  assign n46045 = ( n14379 & ~n18710 ) | ( n14379 & n19602 ) | ( ~n18710 & n19602 ) ;
  assign n46046 = ~n40604 & n43810 ;
  assign n46050 = ( n6414 & n8239 ) | ( n6414 & ~n24860 ) | ( n8239 & ~n24860 ) ;
  assign n46051 = n46050 ^ n6462 ^ 1'b0 ;
  assign n46052 = n20724 & ~n46051 ;
  assign n46053 = ~n6307 & n46052 ;
  assign n46048 = n6468 & n34172 ;
  assign n46049 = n46048 ^ n12179 ^ 1'b0 ;
  assign n46047 = n43327 ^ n40427 ^ n26124 ;
  assign n46054 = n46053 ^ n46049 ^ n46047 ;
  assign n46055 = n30755 ^ n18125 ^ 1'b0 ;
  assign n46056 = n15201 ^ n8511 ^ 1'b0 ;
  assign n46057 = n30183 | n46056 ;
  assign n46059 = n16648 ^ n8208 ^ n7335 ;
  assign n46060 = ( n12001 & ~n16113 ) | ( n12001 & n46059 ) | ( ~n16113 & n46059 ) ;
  assign n46058 = n18765 ^ n14684 ^ 1'b0 ;
  assign n46061 = n46060 ^ n46058 ^ 1'b0 ;
  assign n46062 = n46057 | n46061 ;
  assign n46063 = n16333 ^ n10675 ^ n7139 ;
  assign n46064 = n17507 ^ n11101 ^ n3193 ;
  assign n46065 = n28989 ^ n16585 ^ n6009 ;
  assign n46066 = n46065 ^ n15898 ^ 1'b0 ;
  assign n46067 = n19494 & n40257 ;
  assign n46068 = n46067 ^ n34668 ^ n12970 ;
  assign n46069 = n45426 ^ n25431 ^ 1'b0 ;
  assign n46070 = ~n16555 & n21914 ;
  assign n46071 = n46070 ^ n39674 ^ 1'b0 ;
  assign n46072 = n22061 ^ n7683 ^ 1'b0 ;
  assign n46073 = n33550 & ~n46072 ;
  assign n46074 = n10690 ^ n5165 ^ 1'b0 ;
  assign n46075 = n4825 & n46074 ;
  assign n46076 = n19438 ^ n5695 ^ 1'b0 ;
  assign n46077 = n46075 & n46076 ;
  assign n46078 = n46077 ^ n41900 ^ 1'b0 ;
  assign n46079 = ~n28480 & n46078 ;
  assign n46080 = n5952 & n46079 ;
  assign n46081 = n40499 & n46080 ;
  assign n46082 = n9237 ^ n5338 ^ 1'b0 ;
  assign n46083 = ~n7633 & n46082 ;
  assign n46084 = n46083 ^ n24148 ^ 1'b0 ;
  assign n46085 = n10720 | n46084 ;
  assign n46086 = n6678 & ~n34929 ;
  assign n46087 = n15000 & n46086 ;
  assign n46088 = ~n12722 & n22266 ;
  assign n46089 = n46088 ^ n3111 ^ 1'b0 ;
  assign n46090 = n16334 ^ n15170 ^ n1099 ;
  assign n46091 = ( n16063 & ~n46089 ) | ( n16063 & n46090 ) | ( ~n46089 & n46090 ) ;
  assign n46092 = n30334 ^ n11090 ^ n11077 ;
  assign n46093 = n46092 ^ n17377 ^ n275 ;
  assign n46094 = n18458 ^ n10185 ^ n4038 ;
  assign n46096 = n14875 ^ n8087 ^ 1'b0 ;
  assign n46097 = n5521 & n46096 ;
  assign n46095 = n36340 ^ n6424 ^ 1'b0 ;
  assign n46098 = n46097 ^ n46095 ^ n15070 ;
  assign n46100 = n21607 ^ n8601 ^ n4011 ;
  assign n46099 = ~n16236 & n16795 ;
  assign n46101 = n46100 ^ n46099 ^ 1'b0 ;
  assign n46102 = n46101 ^ n42487 ^ n7899 ;
  assign n46103 = ( n10888 & ~n13557 ) | ( n10888 & n33913 ) | ( ~n13557 & n33913 ) ;
  assign n46104 = n20139 ^ n13610 ^ 1'b0 ;
  assign n46105 = n35331 | n46104 ;
  assign n46106 = n32150 ^ n5660 ^ 1'b0 ;
  assign n46107 = n14892 | n46106 ;
  assign n46108 = n43449 ^ n18468 ^ n4753 ;
  assign n46109 = ( ~n16307 & n21637 ) | ( ~n16307 & n46108 ) | ( n21637 & n46108 ) ;
  assign n46110 = ~n9980 & n13384 ;
  assign n46111 = ~n20161 & n46110 ;
  assign n46112 = n12158 | n46111 ;
  assign n46113 = n46112 ^ n39942 ^ n12638 ;
  assign n46114 = n41655 ^ n33053 ^ 1'b0 ;
  assign n46115 = n20412 ^ n12046 ^ 1'b0 ;
  assign n46116 = n15445 | n46115 ;
  assign n46117 = ( n42639 & n46114 ) | ( n42639 & ~n46116 ) | ( n46114 & ~n46116 ) ;
  assign n46118 = n748 & n6920 ;
  assign n46119 = n2188 & n46118 ;
  assign n46120 = n4404 | n46119 ;
  assign n46121 = ( n8847 & n33876 ) | ( n8847 & ~n34969 ) | ( n33876 & ~n34969 ) ;
  assign n46122 = ( n5581 & ~n17947 ) | ( n5581 & n40945 ) | ( ~n17947 & n40945 ) ;
  assign n46123 = n9353 ^ n1219 ^ 1'b0 ;
  assign n46124 = ~n21227 & n46123 ;
  assign n46125 = n10806 ^ n10426 ^ 1'b0 ;
  assign n46126 = n33826 & ~n46125 ;
  assign n46127 = ( ~n7138 & n8848 ) | ( ~n7138 & n9242 ) | ( n8848 & n9242 ) ;
  assign n46128 = n46127 ^ n33356 ^ n32743 ;
  assign n46129 = ( n23767 & n30304 ) | ( n23767 & ~n35781 ) | ( n30304 & ~n35781 ) ;
  assign n46130 = ( ~n11984 & n43846 ) | ( ~n11984 & n45970 ) | ( n43846 & n45970 ) ;
  assign n46131 = n41811 & ~n46130 ;
  assign n46132 = n46131 ^ n31017 ^ 1'b0 ;
  assign n46133 = ( n2917 & n46129 ) | ( n2917 & ~n46132 ) | ( n46129 & ~n46132 ) ;
  assign n46134 = n41557 ^ n19620 ^ 1'b0 ;
  assign n46135 = n7312 | n8257 ;
  assign n46136 = n46135 ^ n6138 ^ 1'b0 ;
  assign n46137 = n3025 & n24442 ;
  assign n46138 = n46137 ^ n26009 ^ 1'b0 ;
  assign n46143 = n6778 ^ n5999 ^ 1'b0 ;
  assign n46144 = n19524 & n46143 ;
  assign n46145 = n46144 ^ n29530 ^ 1'b0 ;
  assign n46141 = n10755 & ~n21001 ;
  assign n46142 = n46141 ^ n10990 ^ 1'b0 ;
  assign n46146 = n46145 ^ n46142 ^ n9835 ;
  assign n46139 = ( n2690 & ~n8678 ) | ( n2690 & n24802 ) | ( ~n8678 & n24802 ) ;
  assign n46140 = n46139 ^ n2968 ^ 1'b0 ;
  assign n46147 = n46146 ^ n46140 ^ n33279 ;
  assign n46148 = n45744 & n45947 ;
  assign n46149 = ~n18601 & n46148 ;
  assign n46150 = n46149 ^ n45015 ^ n4196 ;
  assign n46153 = ~n397 & n498 ;
  assign n46151 = n7608 | n15825 ;
  assign n46152 = n17669 | n46151 ;
  assign n46154 = n46153 ^ n46152 ^ n41335 ;
  assign n46158 = n12825 & ~n29853 ;
  assign n46159 = n46158 ^ n16890 ^ n12138 ;
  assign n46155 = n26471 ^ n23402 ^ 1'b0 ;
  assign n46156 = n40021 & n46155 ;
  assign n46157 = n46156 ^ n12962 ^ n9842 ;
  assign n46160 = n46159 ^ n46157 ^ n20537 ;
  assign n46161 = n46160 ^ n6601 ^ 1'b0 ;
  assign n46162 = n4884 | n6546 ;
  assign n46163 = n46162 ^ n29956 ^ n16586 ;
  assign n46164 = ( n2401 & n8224 ) | ( n2401 & n40690 ) | ( n8224 & n40690 ) ;
  assign n46168 = ( n21273 & n24836 ) | ( n21273 & ~n38850 ) | ( n24836 & ~n38850 ) ;
  assign n46165 = ( n1030 & n13862 ) | ( n1030 & n35324 ) | ( n13862 & n35324 ) ;
  assign n46166 = ( ~n24745 & n37900 ) | ( ~n24745 & n46165 ) | ( n37900 & n46165 ) ;
  assign n46167 = ~n10452 & n46166 ;
  assign n46169 = n46168 ^ n46167 ^ 1'b0 ;
  assign n46170 = n22701 & ~n40088 ;
  assign n46171 = n5257 & ~n19077 ;
  assign n46172 = ~n11663 & n46171 ;
  assign n46173 = n29983 ^ n19187 ^ 1'b0 ;
  assign n46174 = n2166 & n46173 ;
  assign n46175 = ~n1642 & n46174 ;
  assign n46176 = ~n32273 & n46175 ;
  assign n46177 = ( n8444 & n23145 ) | ( n8444 & n46176 ) | ( n23145 & n46176 ) ;
  assign n46178 = n36049 ^ n26758 ^ n12464 ;
  assign n46179 = n37602 & ~n46178 ;
  assign n46180 = n6399 & n6521 ;
  assign n46181 = n2574 & n46180 ;
  assign n46182 = ( ~n14682 & n42709 ) | ( ~n14682 & n46181 ) | ( n42709 & n46181 ) ;
  assign n46183 = n34417 ^ n20318 ^ n9632 ;
  assign n46184 = n23009 | n42930 ;
  assign n46185 = n46183 & ~n46184 ;
  assign n46186 = n46185 ^ n42580 ^ n27520 ;
  assign n46187 = n26190 ^ n518 ^ 1'b0 ;
  assign n46188 = ( n20448 & n23166 ) | ( n20448 & n30378 ) | ( n23166 & n30378 ) ;
  assign n46189 = n46188 ^ n39502 ^ 1'b0 ;
  assign n46190 = n40672 | n41474 ;
  assign n46191 = n46190 ^ n4094 ^ 1'b0 ;
  assign n46192 = n21207 & ~n46191 ;
  assign n46194 = n5111 | n6241 ;
  assign n46195 = n46194 ^ n33093 ^ 1'b0 ;
  assign n46193 = n6459 | n37805 ;
  assign n46196 = n46195 ^ n46193 ^ n38753 ;
  assign n46197 = ( n17262 & n23540 ) | ( n17262 & ~n24630 ) | ( n23540 & ~n24630 ) ;
  assign n46198 = n33958 ^ n25542 ^ 1'b0 ;
  assign n46199 = n19763 & ~n23680 ;
  assign n46200 = n46199 ^ n18311 ^ n11888 ;
  assign n46201 = n33985 ^ n25058 ^ n11757 ;
  assign n46202 = ( n43926 & n46200 ) | ( n43926 & n46201 ) | ( n46200 & n46201 ) ;
  assign n46203 = ( ~n805 & n19404 ) | ( ~n805 & n44751 ) | ( n19404 & n44751 ) ;
  assign n46204 = n20491 | n46203 ;
  assign n46205 = n46204 ^ n46176 ^ n26474 ;
  assign n46206 = n16193 & n40259 ;
  assign n46207 = n20748 & ~n37720 ;
  assign n46208 = ~n6519 & n46207 ;
  assign n46209 = n10230 | n19157 ;
  assign n46210 = n46209 ^ n4972 ^ 1'b0 ;
  assign n46212 = ( ~n3590 & n7554 ) | ( ~n3590 & n21215 ) | ( n7554 & n21215 ) ;
  assign n46211 = n835 | n35926 ;
  assign n46213 = n46212 ^ n46211 ^ n2456 ;
  assign n46214 = n46213 ^ n38955 ^ n28921 ;
  assign n46215 = n500 & ~n46214 ;
  assign n46216 = n15111 | n46092 ;
  assign n46217 = n24181 ^ n9064 ^ 1'b0 ;
  assign n46218 = ~n7076 & n46217 ;
  assign n46219 = ( n11985 & n31357 ) | ( n11985 & n46218 ) | ( n31357 & n46218 ) ;
  assign n46220 = ( n8149 & ~n17612 ) | ( n8149 & n45510 ) | ( ~n17612 & n45510 ) ;
  assign n46221 = n33270 ^ n32020 ^ n4336 ;
  assign n46222 = n4044 | n15609 ;
  assign n46223 = n41451 & ~n46222 ;
  assign n46224 = n34844 ^ n21053 ^ n5428 ;
  assign n46225 = ~n16962 & n46224 ;
  assign n46226 = n17854 & n35823 ;
  assign n46227 = n46226 ^ n10495 ^ 1'b0 ;
  assign n46228 = n15930 ^ n3054 ^ 1'b0 ;
  assign n46229 = n30522 ^ n29350 ^ n11040 ;
  assign n46230 = n18138 & n32907 ;
  assign n46231 = n31659 ^ n26430 ^ 1'b0 ;
  assign n46232 = n8784 & ~n22403 ;
  assign n46233 = n46232 ^ n43303 ^ 1'b0 ;
  assign n46234 = n14029 ^ n8672 ^ x135 ;
  assign n46235 = n29383 & n46234 ;
  assign n46236 = n46235 ^ n41197 ^ 1'b0 ;
  assign n46237 = n28363 ^ n11320 ^ n7834 ;
  assign n46238 = ~n7104 & n46237 ;
  assign n46239 = n46238 ^ n34318 ^ 1'b0 ;
  assign n46240 = n10590 & ~n18829 ;
  assign n46245 = n44884 ^ n35868 ^ n13039 ;
  assign n46241 = n35280 ^ n11110 ^ n10551 ;
  assign n46242 = n5767 & n46241 ;
  assign n46243 = n46242 ^ n27754 ^ 1'b0 ;
  assign n46244 = n46243 ^ n42028 ^ n10939 ;
  assign n46246 = n46245 ^ n46244 ^ n34322 ;
  assign n46247 = n27991 ^ n12457 ^ 1'b0 ;
  assign n46248 = n8344 & ~n24967 ;
  assign n46249 = n39284 ^ n14326 ^ 1'b0 ;
  assign n46250 = ( ~n9489 & n46248 ) | ( ~n9489 & n46249 ) | ( n46248 & n46249 ) ;
  assign n46251 = n29626 ^ n9271 ^ 1'b0 ;
  assign n46252 = n26916 ^ n9528 ^ 1'b0 ;
  assign n46253 = n3654 & n46252 ;
  assign n46254 = n46253 ^ n17985 ^ 1'b0 ;
  assign n46255 = n34659 ^ n15621 ^ 1'b0 ;
  assign n46256 = n10205 & n46255 ;
  assign n46257 = n38773 ^ n5046 ^ 1'b0 ;
  assign n46258 = n3047 & n46257 ;
  assign n46259 = n43831 & n46258 ;
  assign n46260 = n46259 ^ n33851 ^ 1'b0 ;
  assign n46261 = ( n2640 & n20135 ) | ( n2640 & ~n26563 ) | ( n20135 & ~n26563 ) ;
  assign n46262 = n8491 ^ n7796 ^ 1'b0 ;
  assign n46263 = n4316 & ~n31705 ;
  assign n46264 = n34644 ^ n3586 ^ 1'b0 ;
  assign n46265 = ( n8757 & n18006 ) | ( n8757 & ~n46264 ) | ( n18006 & ~n46264 ) ;
  assign n46266 = ( ~n12694 & n12775 ) | ( ~n12694 & n29617 ) | ( n12775 & n29617 ) ;
  assign n46267 = n6039 ^ x12 ^ 1'b0 ;
  assign n46268 = n5337 & n46267 ;
  assign n46269 = n22042 ^ n400 ^ 1'b0 ;
  assign n46270 = n37035 & n46269 ;
  assign n46271 = ( n3152 & n19398 ) | ( n3152 & n33992 ) | ( n19398 & n33992 ) ;
  assign n46272 = n3516 | n10278 ;
  assign n46273 = n6944 & ~n46272 ;
  assign n46274 = n46273 ^ n35686 ^ n4734 ;
  assign n46275 = ( ~n43698 & n46271 ) | ( ~n43698 & n46274 ) | ( n46271 & n46274 ) ;
  assign n46276 = n34074 & ~n38183 ;
  assign n46277 = ( n23449 & n33487 ) | ( n23449 & ~n37572 ) | ( n33487 & ~n37572 ) ;
  assign n46278 = n32226 ^ n7677 ^ n5818 ;
  assign n46279 = n32291 & ~n41636 ;
  assign n46280 = n31461 ^ n28749 ^ n3690 ;
  assign n46281 = n2163 | n46280 ;
  assign n46282 = ~n5414 & n12692 ;
  assign n46283 = ~n6825 & n46282 ;
  assign n46284 = n46283 ^ n27888 ^ n25634 ;
  assign n46285 = ~n18107 & n46284 ;
  assign n46286 = n46285 ^ n30772 ^ 1'b0 ;
  assign n46287 = ~n14828 & n21316 ;
  assign n46288 = n46287 ^ n38750 ^ 1'b0 ;
  assign n46289 = n33149 & n46288 ;
  assign n46290 = n22514 ^ n7644 ^ 1'b0 ;
  assign n46291 = ( n26044 & n28651 ) | ( n26044 & n46290 ) | ( n28651 & n46290 ) ;
  assign n46293 = n23535 ^ n10708 ^ n4119 ;
  assign n46292 = n45642 ^ n45544 ^ n32878 ;
  assign n46294 = n46293 ^ n46292 ^ 1'b0 ;
  assign n46295 = n46294 ^ n18348 ^ n9286 ;
  assign n46296 = n21537 ^ n10814 ^ 1'b0 ;
  assign n46297 = ( n6781 & n14477 ) | ( n6781 & n15714 ) | ( n14477 & n15714 ) ;
  assign n46298 = n1864 & n4930 ;
  assign n46299 = ~n46297 & n46298 ;
  assign n46300 = n5758 & n23242 ;
  assign n46301 = n10069 & ~n16779 ;
  assign n46302 = ~n46300 & n46301 ;
  assign n46303 = n8095 & n8209 ;
  assign n46304 = ( n3499 & ~n11008 ) | ( n3499 & n23041 ) | ( ~n11008 & n23041 ) ;
  assign n46305 = n26187 ^ n807 ^ 1'b0 ;
  assign n46306 = n46305 ^ n40548 ^ 1'b0 ;
  assign n46307 = ( ~n28284 & n34639 ) | ( ~n28284 & n46306 ) | ( n34639 & n46306 ) ;
  assign n46308 = ( n31062 & n37062 ) | ( n31062 & n42042 ) | ( n37062 & n42042 ) ;
  assign n46309 = n34382 ^ n943 ^ 1'b0 ;
  assign n46310 = n17840 ^ n1799 ^ 1'b0 ;
  assign n46311 = ~n16066 & n46310 ;
  assign n46312 = ( ~n11593 & n18025 ) | ( ~n11593 & n35297 ) | ( n18025 & n35297 ) ;
  assign n46313 = ( n3707 & n9821 ) | ( n3707 & n46312 ) | ( n9821 & n46312 ) ;
  assign n46314 = n32507 ^ n26534 ^ n14741 ;
  assign n46315 = ~n36007 & n36677 ;
  assign n46316 = n46315 ^ n42611 ^ 1'b0 ;
  assign n46317 = n17914 & n30044 ;
  assign n46318 = n46317 ^ n3084 ^ 1'b0 ;
  assign n46319 = n46318 ^ n25162 ^ n9997 ;
  assign n46320 = ( n31572 & n39216 ) | ( n31572 & n39939 ) | ( n39216 & n39939 ) ;
  assign n46322 = n29608 ^ n29147 ^ 1'b0 ;
  assign n46323 = n46322 ^ n41081 ^ n5660 ;
  assign n46321 = n6406 | n28153 ;
  assign n46324 = n46323 ^ n46321 ^ 1'b0 ;
  assign n46325 = n4483 & n10854 ;
  assign n46326 = n38904 ^ n34578 ^ 1'b0 ;
  assign n46327 = n30415 ^ n19427 ^ 1'b0 ;
  assign n46328 = n23858 ^ n998 ^ 1'b0 ;
  assign n46329 = n17554 ^ n13859 ^ 1'b0 ;
  assign n46330 = n46329 ^ n6714 ^ n3073 ;
  assign n46331 = n36575 ^ n17327 ^ n17322 ;
  assign n46332 = n46331 ^ n271 ^ 1'b0 ;
  assign n46333 = ~n9469 & n46332 ;
  assign n46334 = n3460 ^ n2311 ^ 1'b0 ;
  assign n46335 = n24189 | n46334 ;
  assign n46336 = ( x54 & n1352 ) | ( x54 & ~n41750 ) | ( n1352 & ~n41750 ) ;
  assign n46337 = n8138 ^ n4920 ^ 1'b0 ;
  assign n46338 = ~n29664 & n46337 ;
  assign n46339 = ~n947 & n46338 ;
  assign n46340 = n46336 & n46339 ;
  assign n46341 = n1429 | n6621 ;
  assign n46342 = n46341 ^ n22930 ^ 1'b0 ;
  assign n46343 = n40033 & n46342 ;
  assign n46344 = n971 & n11818 ;
  assign n46345 = n46344 ^ n5015 ^ 1'b0 ;
  assign n46346 = n46345 ^ n3618 ^ n2180 ;
  assign n46347 = n38335 ^ n6647 ^ 1'b0 ;
  assign n46348 = n46347 ^ n18968 ^ n1502 ;
  assign n46349 = n23600 ^ n13972 ^ n7042 ;
  assign n46350 = n46349 ^ n23254 ^ 1'b0 ;
  assign n46351 = n20206 ^ n13271 ^ 1'b0 ;
  assign n46352 = n16093 ^ n10911 ^ 1'b0 ;
  assign n46353 = n35039 ^ n18625 ^ 1'b0 ;
  assign n46354 = n42305 & n46353 ;
  assign n46355 = ~n9568 & n20773 ;
  assign n46356 = n46355 ^ n681 ^ 1'b0 ;
  assign n46357 = n19254 & ~n36350 ;
  assign n46358 = n46357 ^ n8276 ^ 1'b0 ;
  assign n46359 = n5815 ^ n3427 ^ 1'b0 ;
  assign n46360 = ( n28512 & ~n46358 ) | ( n28512 & n46359 ) | ( ~n46358 & n46359 ) ;
  assign n46361 = n25218 ^ n21853 ^ 1'b0 ;
  assign n46362 = n15930 ^ n11083 ^ n6642 ;
  assign n46363 = ~n10484 & n13603 ;
  assign n46364 = ( ~n12263 & n16684 ) | ( ~n12263 & n39198 ) | ( n16684 & n39198 ) ;
  assign n46368 = ( n2933 & n6042 ) | ( n2933 & n10736 ) | ( n6042 & n10736 ) ;
  assign n46369 = n30229 ^ n8770 ^ 1'b0 ;
  assign n46370 = n46368 & n46369 ;
  assign n46365 = n29656 ^ n26603 ^ n11680 ;
  assign n46366 = n41591 & ~n46365 ;
  assign n46367 = n46366 ^ n4161 ^ 1'b0 ;
  assign n46371 = n46370 ^ n46367 ^ n42996 ;
  assign n46372 = n37416 ^ n22878 ^ 1'b0 ;
  assign n46373 = n20060 ^ n8414 ^ 1'b0 ;
  assign n46374 = n16327 & ~n46373 ;
  assign n46375 = n11185 & n46374 ;
  assign n46376 = n25516 ^ n5370 ^ 1'b0 ;
  assign n46377 = ( n19904 & n37947 ) | ( n19904 & ~n46376 ) | ( n37947 & ~n46376 ) ;
  assign n46378 = n17159 ^ n7641 ^ n3324 ;
  assign n46381 = ( ~x107 & n4847 ) | ( ~x107 & n30268 ) | ( n4847 & n30268 ) ;
  assign n46379 = n1912 ^ n268 ^ 1'b0 ;
  assign n46380 = n46379 ^ n13481 ^ n5536 ;
  assign n46382 = n46381 ^ n46380 ^ 1'b0 ;
  assign n46383 = ( n43780 & n46378 ) | ( n43780 & n46382 ) | ( n46378 & n46382 ) ;
  assign n46384 = ~n2720 & n46383 ;
  assign n46385 = ~n20554 & n20880 ;
  assign n46386 = n46385 ^ n24627 ^ 1'b0 ;
  assign n46388 = ~n633 & n18730 ;
  assign n46389 = n46388 ^ n26412 ^ 1'b0 ;
  assign n46387 = n298 & n11817 ;
  assign n46390 = n46389 ^ n46387 ^ 1'b0 ;
  assign n46391 = n768 & n7454 ;
  assign n46392 = ( n14741 & n20752 ) | ( n14741 & ~n46391 ) | ( n20752 & ~n46391 ) ;
  assign n46393 = ( n882 & n13994 ) | ( n882 & ~n36303 ) | ( n13994 & ~n36303 ) ;
  assign n46394 = n46393 ^ n11735 ^ n10266 ;
  assign n46398 = ( n13173 & ~n21076 ) | ( n13173 & n33515 ) | ( ~n21076 & n33515 ) ;
  assign n46395 = n1722 | n17393 ;
  assign n46396 = ~n9404 & n19576 ;
  assign n46397 = n46395 & n46396 ;
  assign n46399 = n46398 ^ n46397 ^ n39428 ;
  assign n46400 = n4599 & ~n11099 ;
  assign n46401 = ( ~n4523 & n19670 ) | ( ~n4523 & n20533 ) | ( n19670 & n20533 ) ;
  assign n46402 = n46401 ^ n17503 ^ 1'b0 ;
  assign n46403 = ~n10578 & n21258 ;
  assign n46404 = n32943 & n46403 ;
  assign n46405 = n46404 ^ n38139 ^ 1'b0 ;
  assign n46407 = n17179 ^ n7421 ^ n2629 ;
  assign n46408 = n20507 | n46407 ;
  assign n46409 = n46408 ^ n12371 ^ n9037 ;
  assign n46406 = n3994 & n41957 ;
  assign n46410 = n46409 ^ n46406 ^ 1'b0 ;
  assign n46411 = n15698 & ~n33746 ;
  assign n46412 = n31440 & ~n46411 ;
  assign n46413 = ~n12213 & n19512 ;
  assign n46414 = ~n33480 & n46413 ;
  assign n46415 = n15181 ^ n9698 ^ n7980 ;
  assign n46416 = n46415 ^ n3529 ^ 1'b0 ;
  assign n46417 = n1536 | n27228 ;
  assign n46418 = n46416 | n46417 ;
  assign n46419 = n16846 | n25189 ;
  assign n46421 = ( ~n16129 & n16188 ) | ( ~n16129 & n23538 ) | ( n16188 & n23538 ) ;
  assign n46422 = ( ~n20431 & n34035 ) | ( ~n20431 & n46421 ) | ( n34035 & n46421 ) ;
  assign n46420 = n21234 | n28002 ;
  assign n46423 = n46422 ^ n46420 ^ 1'b0 ;
  assign n46424 = n46423 ^ n9996 ^ n1728 ;
  assign n46426 = ( n2933 & n9195 ) | ( n2933 & n13005 ) | ( n9195 & n13005 ) ;
  assign n46425 = n25514 ^ n19154 ^ n18623 ;
  assign n46427 = n46426 ^ n46425 ^ 1'b0 ;
  assign n46428 = n37534 & ~n39994 ;
  assign n46429 = n848 & n46428 ;
  assign n46430 = ( n35598 & n41780 ) | ( n35598 & ~n46429 ) | ( n41780 & ~n46429 ) ;
  assign n46431 = n30361 ^ n20210 ^ n7867 ;
  assign n46432 = n46431 ^ n39041 ^ n8789 ;
  assign n46433 = ~n15636 & n22690 ;
  assign n46434 = ~n9454 & n46433 ;
  assign n46435 = n46434 ^ n42028 ^ n2723 ;
  assign n46436 = n12485 & ~n37967 ;
  assign n46437 = n22201 | n22725 ;
  assign n46438 = n32567 | n46437 ;
  assign n46439 = n31791 & n46438 ;
  assign n46440 = n46439 ^ n2984 ^ 1'b0 ;
  assign n46441 = ( ~n4075 & n6103 ) | ( ~n4075 & n30261 ) | ( n6103 & n30261 ) ;
  assign n46442 = n46441 ^ n22514 ^ 1'b0 ;
  assign n46443 = n10944 ^ n2696 ^ 1'b0 ;
  assign n46444 = n46442 | n46443 ;
  assign n46445 = ~n5761 & n9623 ;
  assign n46446 = n46445 ^ n7114 ^ 1'b0 ;
  assign n46447 = n46446 ^ n35187 ^ n9067 ;
  assign n46450 = n15674 ^ n9565 ^ 1'b0 ;
  assign n46449 = ( n8245 & n16878 ) | ( n8245 & n46050 ) | ( n16878 & n46050 ) ;
  assign n46451 = n46450 ^ n46449 ^ n15655 ;
  assign n46448 = n31377 ^ n30460 ^ n11335 ;
  assign n46452 = n46451 ^ n46448 ^ n26095 ;
  assign n46453 = n37961 ^ n21517 ^ n19740 ;
  assign n46454 = n46453 ^ n28227 ^ 1'b0 ;
  assign n46455 = n46258 ^ n19798 ^ 1'b0 ;
  assign n46456 = n35147 & n43987 ;
  assign n46457 = ~n16675 & n46456 ;
  assign n46458 = ~n8416 & n20371 ;
  assign n46459 = ~n11700 & n46458 ;
  assign n46460 = n46459 ^ n33985 ^ n4566 ;
  assign n46461 = ( ~n2895 & n14905 ) | ( ~n2895 & n22280 ) | ( n14905 & n22280 ) ;
  assign n46462 = ( n1685 & n21139 ) | ( n1685 & ~n39238 ) | ( n21139 & ~n39238 ) ;
  assign n46463 = ~n3983 & n23007 ;
  assign n46464 = n46463 ^ n5403 ^ 1'b0 ;
  assign n46465 = n46464 ^ n36029 ^ n16754 ;
  assign n46466 = n4121 & n20827 ;
  assign n46467 = ( n24001 & n29381 ) | ( n24001 & ~n46466 ) | ( n29381 & ~n46466 ) ;
  assign n46468 = n20457 ^ n11373 ^ 1'b0 ;
  assign n46469 = n25613 | n46468 ;
  assign n46470 = n46469 ^ n23446 ^ n14595 ;
  assign n46471 = n12614 ^ n3963 ^ 1'b0 ;
  assign n46472 = n46470 | n46471 ;
  assign n46474 = ( n3696 & ~n8229 ) | ( n3696 & n36319 ) | ( ~n8229 & n36319 ) ;
  assign n46473 = n5249 ^ n4913 ^ n1646 ;
  assign n46475 = n46474 ^ n46473 ^ 1'b0 ;
  assign n46476 = ( ~n11908 & n25230 ) | ( ~n11908 & n29899 ) | ( n25230 & n29899 ) ;
  assign n46477 = n31449 ^ n5732 ^ 1'b0 ;
  assign n46478 = n36511 ^ n29380 ^ 1'b0 ;
  assign n46479 = n16434 | n46478 ;
  assign n46480 = n15377 | n30355 ;
  assign n46481 = n46480 ^ n5654 ^ 1'b0 ;
  assign n46482 = ~n13634 & n26377 ;
  assign n46483 = n39408 ^ n16775 ^ 1'b0 ;
  assign n46484 = n46482 | n46483 ;
  assign n46485 = n10470 | n46484 ;
  assign n46486 = n20865 & ~n31962 ;
  assign n46487 = n5992 & ~n23995 ;
  assign n46488 = n32372 ^ n17839 ^ 1'b0 ;
  assign n46489 = ~n46487 & n46488 ;
  assign n46490 = ( ~n6628 & n27765 ) | ( ~n6628 & n46305 ) | ( n27765 & n46305 ) ;
  assign n46491 = ( n8858 & ~n20263 ) | ( n8858 & n33254 ) | ( ~n20263 & n33254 ) ;
  assign n46492 = ~n22629 & n27954 ;
  assign n46493 = n12659 & ~n16136 ;
  assign n46494 = ~n2080 & n46493 ;
  assign n46495 = n27497 ^ n20235 ^ 1'b0 ;
  assign n46496 = ( n21358 & ~n46494 ) | ( n21358 & n46495 ) | ( ~n46494 & n46495 ) ;
  assign n46497 = ( ~n11328 & n46492 ) | ( ~n11328 & n46496 ) | ( n46492 & n46496 ) ;
  assign n46498 = n9285 | n42679 ;
  assign n46499 = n31598 ^ n30570 ^ n1598 ;
  assign n46501 = n46404 ^ n35613 ^ n30328 ;
  assign n46500 = n3604 & ~n18681 ;
  assign n46502 = n46501 ^ n46500 ^ 1'b0 ;
  assign n46504 = n6951 ^ n4924 ^ n426 ;
  assign n46503 = n23195 & ~n46320 ;
  assign n46505 = n46504 ^ n46503 ^ 1'b0 ;
  assign n46506 = n2775 | n20222 ;
  assign n46507 = n36094 & ~n46506 ;
  assign n46508 = n2027 | n46507 ;
  assign n46509 = n46508 ^ n34038 ^ 1'b0 ;
  assign n46510 = n8082 | n34383 ;
  assign n46511 = n16281 ^ n6765 ^ 1'b0 ;
  assign n46512 = n46510 & n46511 ;
  assign n46513 = ( n41551 & n42826 ) | ( n41551 & n46512 ) | ( n42826 & n46512 ) ;
  assign n46518 = n14165 ^ n8784 ^ 1'b0 ;
  assign n46514 = n15323 & n45666 ;
  assign n46515 = n20340 ^ n16064 ^ n5937 ;
  assign n46516 = ~n46514 & n46515 ;
  assign n46517 = n35253 & n46516 ;
  assign n46519 = n46518 ^ n46517 ^ 1'b0 ;
  assign n46520 = n17755 ^ n14553 ^ 1'b0 ;
  assign n46521 = n32094 ^ n8713 ^ 1'b0 ;
  assign n46522 = n20108 & ~n21221 ;
  assign n46523 = n46521 & n46522 ;
  assign n46524 = ( n8785 & ~n22313 ) | ( n8785 & n46523 ) | ( ~n22313 & n46523 ) ;
  assign n46525 = ( ~n24461 & n34595 ) | ( ~n24461 & n45870 ) | ( n34595 & n45870 ) ;
  assign n46528 = n42844 ^ n33537 ^ n12148 ;
  assign n46526 = n9557 & ~n14106 ;
  assign n46527 = n11296 | n46526 ;
  assign n46529 = n46528 ^ n46527 ^ 1'b0 ;
  assign n46530 = n9288 | n12461 ;
  assign n46531 = n29639 ^ n27691 ^ n5914 ;
  assign n46532 = n16836 ^ n13543 ^ n2381 ;
  assign n46533 = ~n13537 & n46532 ;
  assign n46534 = ( n13506 & ~n18237 ) | ( n13506 & n27299 ) | ( ~n18237 & n27299 ) ;
  assign n46535 = n41053 ^ n21512 ^ n17449 ;
  assign n46536 = ~n19970 & n46535 ;
  assign n46537 = n30796 & n46536 ;
  assign n46538 = ( n6747 & n23261 ) | ( n6747 & n46537 ) | ( n23261 & n46537 ) ;
  assign n46539 = n1945 | n5779 ;
  assign n46540 = n46539 ^ n40736 ^ n32072 ;
  assign n46541 = ( n13163 & n22939 ) | ( n13163 & n44889 ) | ( n22939 & n44889 ) ;
  assign n46542 = n17496 & n46541 ;
  assign n46543 = n29983 | n33876 ;
  assign n46544 = n24697 | n46543 ;
  assign n46545 = n46544 ^ n25645 ^ 1'b0 ;
  assign n46546 = n15930 ^ n6750 ^ 1'b0 ;
  assign n46547 = n30955 | n46546 ;
  assign n46548 = n29457 ^ n9424 ^ 1'b0 ;
  assign n46549 = n46548 ^ n34984 ^ n6885 ;
  assign n46550 = n10553 & n24391 ;
  assign n46551 = n46550 ^ n3854 ^ 1'b0 ;
  assign n46552 = n46549 | n46551 ;
  assign n46553 = n24465 | n36759 ;
  assign n46554 = n7874 & ~n46553 ;
  assign n46555 = n8906 & n22930 ;
  assign n46556 = ( n22788 & n46554 ) | ( n22788 & ~n46555 ) | ( n46554 & ~n46555 ) ;
  assign n46557 = ( n2900 & n10507 ) | ( n2900 & n21422 ) | ( n10507 & n21422 ) ;
  assign n46558 = n10139 ^ n6723 ^ 1'b0 ;
  assign n46559 = n46558 ^ n26880 ^ n19129 ;
  assign n46560 = ~n43146 & n46559 ;
  assign n46561 = n38067 ^ n24049 ^ n19786 ;
  assign n46563 = ( n3720 & ~n4570 ) | ( n3720 & n7873 ) | ( ~n4570 & n7873 ) ;
  assign n46562 = n35326 ^ n32560 ^ n25379 ;
  assign n46564 = n46563 ^ n46562 ^ n44582 ;
  assign n46565 = n10991 & n17122 ;
  assign n46566 = n46565 ^ n8581 ^ 1'b0 ;
  assign n46567 = ( n1411 & ~n26686 ) | ( n1411 & n35771 ) | ( ~n26686 & n35771 ) ;
  assign n46568 = n3821 & ~n46567 ;
  assign n46569 = ( n21158 & n31313 ) | ( n21158 & n38255 ) | ( n31313 & n38255 ) ;
  assign n46570 = n15594 & n41522 ;
  assign n46571 = n46570 ^ n32322 ^ 1'b0 ;
  assign n46572 = n23155 ^ n5238 ^ 1'b0 ;
  assign n46573 = n34895 & ~n46572 ;
  assign n46574 = ~n46571 & n46573 ;
  assign n46575 = n46574 ^ n10011 ^ 1'b0 ;
  assign n46576 = n46569 & n46575 ;
  assign n46577 = ~n1563 & n17155 ;
  assign n46578 = n35112 & n46577 ;
  assign n46579 = n28482 & ~n46578 ;
  assign n46580 = n33566 & n46579 ;
  assign n46581 = n11155 ^ n4214 ^ 1'b0 ;
  assign n46582 = n19823 | n46581 ;
  assign n46583 = n20329 | n46582 ;
  assign n46584 = n10943 | n19848 ;
  assign n46585 = n15165 | n46584 ;
  assign n46586 = ( n6921 & n8414 ) | ( n6921 & ~n10108 ) | ( n8414 & ~n10108 ) ;
  assign n46587 = n43264 ^ n20396 ^ 1'b0 ;
  assign n46588 = n46586 | n46587 ;
  assign n46589 = n37899 & ~n46588 ;
  assign n46590 = n41389 ^ n23022 ^ n17949 ;
  assign n46593 = n7186 ^ n5914 ^ 1'b0 ;
  assign n46592 = n12583 & ~n17943 ;
  assign n46594 = n46593 ^ n46592 ^ 1'b0 ;
  assign n46595 = n46594 ^ n27328 ^ n8574 ;
  assign n46591 = ~n1984 & n10526 ;
  assign n46596 = n46595 ^ n46591 ^ 1'b0 ;
  assign n46597 = n46596 ^ n28502 ^ n11298 ;
  assign n46598 = n2638 | n34709 ;
  assign n46599 = n4546 & n30076 ;
  assign n46600 = ( ~n39138 & n46598 ) | ( ~n39138 & n46599 ) | ( n46598 & n46599 ) ;
  assign n46601 = ( n12659 & n14093 ) | ( n12659 & n16149 ) | ( n14093 & n16149 ) ;
  assign n46602 = n46601 ^ n43713 ^ n1547 ;
  assign n46603 = ( ~n8917 & n34874 ) | ( ~n8917 & n46602 ) | ( n34874 & n46602 ) ;
  assign n46604 = n31570 ^ n20851 ^ 1'b0 ;
  assign n46605 = n14887 ^ n4064 ^ 1'b0 ;
  assign n46606 = n6554 | n46605 ;
  assign n46607 = n46606 ^ n22350 ^ 1'b0 ;
  assign n46608 = ~n17180 & n33985 ;
  assign n46609 = n4490 & n46608 ;
  assign n46610 = n46609 ^ n12144 ^ 1'b0 ;
  assign n46611 = n31739 ^ n16752 ^ 1'b0 ;
  assign n46612 = n46610 & n46611 ;
  assign n46613 = n45802 ^ n2733 ^ 1'b0 ;
  assign n46614 = n46612 & ~n46613 ;
  assign n46615 = n18322 ^ n13506 ^ 1'b0 ;
  assign n46616 = n46615 ^ n37092 ^ n4490 ;
  assign n46617 = n4674 | n12681 ;
  assign n46618 = n46616 | n46617 ;
  assign n46619 = ( ~n360 & n16280 ) | ( ~n360 & n18537 ) | ( n16280 & n18537 ) ;
  assign n46620 = n46619 ^ n4629 ^ n1125 ;
  assign n46621 = ( n15111 & n20123 ) | ( n15111 & ~n28591 ) | ( n20123 & ~n28591 ) ;
  assign n46622 = n20503 ^ n17094 ^ n10804 ;
  assign n46623 = n15431 ^ n10574 ^ n8828 ;
  assign n46624 = ( n3633 & n5561 ) | ( n3633 & n30577 ) | ( n5561 & n30577 ) ;
  assign n46625 = n46624 ^ n30749 ^ n25746 ;
  assign n46626 = ( n2544 & n6973 ) | ( n2544 & ~n22983 ) | ( n6973 & ~n22983 ) ;
  assign n46629 = ~n13327 & n34349 ;
  assign n46630 = n11720 & n46629 ;
  assign n46627 = n10676 & ~n42312 ;
  assign n46628 = ~n37434 & n46627 ;
  assign n46631 = n46630 ^ n46628 ^ 1'b0 ;
  assign n46632 = n46626 | n46631 ;
  assign n46633 = n16295 ^ n12096 ^ 1'b0 ;
  assign n46634 = n16023 ^ n14986 ^ 1'b0 ;
  assign n46635 = n46633 & ~n46634 ;
  assign n46636 = n38020 ^ n37507 ^ n8103 ;
  assign n46637 = ~n5112 & n46636 ;
  assign n46638 = n46637 ^ n21238 ^ 1'b0 ;
  assign n46639 = n35351 ^ n5020 ^ 1'b0 ;
  assign n46640 = ~n15938 & n26032 ;
  assign n46641 = ~n23678 & n46640 ;
  assign n46642 = ( n5363 & n25319 ) | ( n5363 & n46641 ) | ( n25319 & n46641 ) ;
  assign n46643 = ( n1474 & ~n30055 ) | ( n1474 & n46642 ) | ( ~n30055 & n46642 ) ;
  assign n46644 = n3258 & n46643 ;
  assign n46645 = n46644 ^ n17283 ^ 1'b0 ;
  assign n46646 = n39993 ^ n39422 ^ n14951 ;
  assign n46647 = ~n33585 & n37503 ;
  assign n46649 = n23968 & n44860 ;
  assign n46650 = n46649 ^ n18970 ^ 1'b0 ;
  assign n46648 = n22694 & n40497 ;
  assign n46651 = n46650 ^ n46648 ^ 1'b0 ;
  assign n46652 = ( ~n2779 & n17204 ) | ( ~n2779 & n46651 ) | ( n17204 & n46651 ) ;
  assign n46653 = ( ~n37749 & n44145 ) | ( ~n37749 & n46652 ) | ( n44145 & n46652 ) ;
  assign n46654 = n23106 & ~n26704 ;
  assign n46655 = n46654 ^ n10430 ^ 1'b0 ;
  assign n46656 = n23113 ^ n5583 ^ 1'b0 ;
  assign n46657 = n36141 & ~n46656 ;
  assign n46658 = n39582 ^ n10584 ^ 1'b0 ;
  assign n46659 = n46657 & n46658 ;
  assign n46660 = ( n1382 & ~n5343 ) | ( n1382 & n12100 ) | ( ~n5343 & n12100 ) ;
  assign n46661 = n23332 ^ n19368 ^ 1'b0 ;
  assign n46662 = ( n20272 & n46660 ) | ( n20272 & ~n46661 ) | ( n46660 & ~n46661 ) ;
  assign n46663 = ( ~n1296 & n1573 ) | ( ~n1296 & n32530 ) | ( n1573 & n32530 ) ;
  assign n46664 = n33227 ^ n1670 ^ x29 ;
  assign n46665 = n2110 & ~n46664 ;
  assign n46666 = n22404 ^ n14859 ^ 1'b0 ;
  assign n46667 = n46666 ^ n28909 ^ n28272 ;
  assign n46668 = n46667 ^ n19743 ^ 1'b0 ;
  assign n46669 = n4711 & ~n19189 ;
  assign n46670 = n13031 ^ n12047 ^ 1'b0 ;
  assign n46671 = n28021 ^ n15626 ^ 1'b0 ;
  assign n46672 = n46670 & n46671 ;
  assign n46675 = n3927 & ~n26699 ;
  assign n46676 = n3408 & n46675 ;
  assign n46673 = ~n29792 & n39231 ;
  assign n46674 = n18519 | n46673 ;
  assign n46677 = n46676 ^ n46674 ^ 1'b0 ;
  assign n46678 = ~n7856 & n34891 ;
  assign n46679 = n46677 & n46678 ;
  assign n46680 = n41340 ^ n13645 ^ 1'b0 ;
  assign n46681 = n10289 ^ n1510 ^ 1'b0 ;
  assign n46682 = n25712 & n46681 ;
  assign n46683 = n37770 ^ n13117 ^ x205 ;
  assign n46684 = ~n4674 & n8177 ;
  assign n46685 = n26548 ^ n5787 ^ 1'b0 ;
  assign n46686 = n12371 ^ n2430 ^ 1'b0 ;
  assign n46687 = n1506 & ~n28640 ;
  assign n46688 = ( n5053 & n46686 ) | ( n5053 & ~n46687 ) | ( n46686 & ~n46687 ) ;
  assign n46689 = n11387 ^ n325 ^ 1'b0 ;
  assign n46690 = ~n12148 & n46689 ;
  assign n46691 = ( n13004 & n22511 ) | ( n13004 & ~n46690 ) | ( n22511 & ~n46690 ) ;
  assign n46692 = n16136 | n37137 ;
  assign n46693 = n34969 | n46692 ;
  assign n46694 = ( n19347 & n41120 ) | ( n19347 & ~n46693 ) | ( n41120 & ~n46693 ) ;
  assign n46695 = n34516 | n46694 ;
  assign n46696 = n46695 ^ n32646 ^ 1'b0 ;
  assign n46697 = n12818 & ~n45263 ;
  assign n46698 = n38677 ^ n1697 ^ 1'b0 ;
  assign n46699 = ~n20690 & n46698 ;
  assign n46700 = n20827 ^ n11649 ^ 1'b0 ;
  assign n46701 = n6476 & n46700 ;
  assign n46702 = ~n32535 & n46701 ;
  assign n46703 = ( ~n3806 & n17434 ) | ( ~n3806 & n38528 ) | ( n17434 & n38528 ) ;
  assign n46704 = ( n20450 & n22821 ) | ( n20450 & n25735 ) | ( n22821 & n25735 ) ;
  assign n46705 = ( n1965 & n15698 ) | ( n1965 & n27294 ) | ( n15698 & n27294 ) ;
  assign n46706 = n26208 ^ n12917 ^ 1'b0 ;
  assign n46707 = ( ~n10869 & n11978 ) | ( ~n10869 & n26716 ) | ( n11978 & n26716 ) ;
  assign n46708 = ( n30800 & n46706 ) | ( n30800 & ~n46707 ) | ( n46706 & ~n46707 ) ;
  assign n46709 = n13235 | n41102 ;
  assign n46710 = n43061 & ~n46709 ;
  assign n46711 = n6833 & ~n46205 ;
  assign n46712 = n28288 & n46711 ;
  assign n46713 = n7447 ^ n2377 ^ 1'b0 ;
  assign n46714 = n13114 ^ n9633 ^ n1257 ;
  assign n46715 = n46714 ^ n19588 ^ n18156 ;
  assign n46716 = ( n34694 & n42571 ) | ( n34694 & ~n46715 ) | ( n42571 & ~n46715 ) ;
  assign n46717 = n3658 & n46716 ;
  assign n46718 = ( n10534 & ~n46713 ) | ( n10534 & n46717 ) | ( ~n46713 & n46717 ) ;
  assign n46719 = n15924 ^ n7468 ^ 1'b0 ;
  assign n46720 = n3241 | n46719 ;
  assign n46721 = ( ~n2928 & n23882 ) | ( ~n2928 & n46720 ) | ( n23882 & n46720 ) ;
  assign n46722 = n20158 ^ n13147 ^ 1'b0 ;
  assign n46723 = n13413 | n17001 ;
  assign n46724 = n46723 ^ n21228 ^ 1'b0 ;
  assign n46725 = n4217 & ~n37493 ;
  assign n46726 = ( ~n46722 & n46724 ) | ( ~n46722 & n46725 ) | ( n46724 & n46725 ) ;
  assign n46727 = ( n5071 & n27462 ) | ( n5071 & ~n30890 ) | ( n27462 & ~n30890 ) ;
  assign n46729 = n24926 & ~n46425 ;
  assign n46728 = n17346 ^ n11810 ^ n355 ;
  assign n46730 = n46729 ^ n46728 ^ n20994 ;
  assign n46731 = n22096 ^ n4808 ^ 1'b0 ;
  assign n46732 = n5769 & ~n18704 ;
  assign n46733 = n46732 ^ n2095 ^ 1'b0 ;
  assign n46734 = n13558 | n15136 ;
  assign n46735 = n46734 ^ n19568 ^ 1'b0 ;
  assign n46736 = ~n21211 & n24243 ;
  assign n46737 = ~n40082 & n46736 ;
  assign n46738 = n1614 | n15700 ;
  assign n46739 = n46738 ^ n33232 ^ 1'b0 ;
  assign n46740 = n34420 ^ n26268 ^ 1'b0 ;
  assign n46741 = n36789 ^ n8095 ^ n1659 ;
  assign n46742 = ( n13298 & ~n46280 ) | ( n13298 & n46741 ) | ( ~n46280 & n46741 ) ;
  assign n46743 = n28442 ^ n11065 ^ x59 ;
  assign n46744 = n33960 ^ n12040 ^ n9571 ;
  assign n46745 = n8173 & n46744 ;
  assign n46746 = n35544 ^ n15766 ^ n13305 ;
  assign n46747 = n46746 ^ n12841 ^ n12373 ;
  assign n46748 = n9852 & n37359 ;
  assign n46749 = n40477 & n46748 ;
  assign n46750 = n28386 & n37734 ;
  assign n46751 = n46750 ^ n1401 ^ 1'b0 ;
  assign n46752 = ~n4958 & n16616 ;
  assign n46753 = n46752 ^ n45402 ^ 1'b0 ;
  assign n46754 = n21156 & ~n37695 ;
  assign n46755 = n45484 ^ n9560 ^ 1'b0 ;
  assign n46756 = n24492 ^ n9420 ^ 1'b0 ;
  assign n46757 = n42342 | n46756 ;
  assign n46758 = n11762 ^ n8638 ^ 1'b0 ;
  assign n46759 = ( n744 & n10579 ) | ( n744 & ~n30354 ) | ( n10579 & ~n30354 ) ;
  assign n46760 = n46759 ^ n28192 ^ n27529 ;
  assign n46761 = n18488 & ~n21041 ;
  assign n46762 = n20593 ^ n17994 ^ 1'b0 ;
  assign n46763 = ~n46761 & n46762 ;
  assign n46764 = n19179 ^ n15813 ^ 1'b0 ;
  assign n46765 = n21526 & n46764 ;
  assign n46766 = n28185 ^ n11697 ^ n9850 ;
  assign n46767 = n8597 | n14542 ;
  assign n46768 = n6232 & ~n46767 ;
  assign n46769 = n21172 | n46768 ;
  assign n46770 = n46769 ^ n21135 ^ n17725 ;
  assign n46771 = n46770 ^ n8693 ^ x13 ;
  assign n46773 = ~n2329 & n16222 ;
  assign n46774 = n5275 & n46773 ;
  assign n46772 = n19614 ^ n17769 ^ 1'b0 ;
  assign n46775 = n46774 ^ n46772 ^ n18728 ;
  assign n46779 = n31654 ^ n14432 ^ 1'b0 ;
  assign n46778 = ~n18255 & n26454 ;
  assign n46776 = ( ~n3445 & n3748 ) | ( ~n3445 & n16046 ) | ( n3748 & n16046 ) ;
  assign n46777 = n46776 ^ n37662 ^ n18884 ;
  assign n46780 = n46779 ^ n46778 ^ n46777 ;
  assign n46781 = n38164 ^ n34233 ^ n27671 ;
  assign n46782 = n19843 ^ n9647 ^ 1'b0 ;
  assign n46783 = n46781 & n46782 ;
  assign n46784 = n13047 & n24967 ;
  assign n46785 = n40431 & n46784 ;
  assign n46786 = ( ~n3878 & n3955 ) | ( ~n3878 & n46785 ) | ( n3955 & n46785 ) ;
  assign n46787 = n46786 ^ n33324 ^ 1'b0 ;
  assign n46788 = ( ~n29188 & n46783 ) | ( ~n29188 & n46787 ) | ( n46783 & n46787 ) ;
  assign n46790 = ( ~n3138 & n3677 ) | ( ~n3138 & n16176 ) | ( n3677 & n16176 ) ;
  assign n46791 = n32802 & ~n34417 ;
  assign n46792 = n46790 & n46791 ;
  assign n46793 = n46792 ^ n3220 ^ 1'b0 ;
  assign n46789 = n46395 ^ n9320 ^ 1'b0 ;
  assign n46794 = n46793 ^ n46789 ^ n10450 ;
  assign n46795 = n9834 & n34720 ;
  assign n46796 = ( n19667 & n36262 ) | ( n19667 & ~n37638 ) | ( n36262 & ~n37638 ) ;
  assign n46797 = n43779 & ~n46796 ;
  assign n46798 = n46797 ^ n12906 ^ 1'b0 ;
  assign n46799 = n32630 ^ n9115 ^ n2045 ;
  assign n46800 = ( n23763 & n35321 ) | ( n23763 & ~n45478 ) | ( n35321 & ~n45478 ) ;
  assign n46801 = ( ~n19604 & n46799 ) | ( ~n19604 & n46800 ) | ( n46799 & n46800 ) ;
  assign n46802 = n44369 ^ n20382 ^ n1076 ;
  assign n46803 = n44568 ^ n11101 ^ n4435 ;
  assign n46804 = n31731 ^ n20141 ^ n13581 ;
  assign n46805 = n45360 ^ n10565 ^ n7013 ;
  assign n46806 = n46804 & ~n46805 ;
  assign n46807 = n34713 ^ n17443 ^ n10030 ;
  assign n46808 = n24442 ^ n15810 ^ n1797 ;
  assign n46809 = n40551 ^ n34571 ^ n8703 ;
  assign n46810 = n15431 & ~n46809 ;
  assign n46811 = ~n46808 & n46810 ;
  assign n46812 = n16655 | n46811 ;
  assign n46813 = n9744 | n36637 ;
  assign n46814 = n28498 ^ n7458 ^ 1'b0 ;
  assign n46815 = ( n25351 & n32924 ) | ( n25351 & ~n40860 ) | ( n32924 & ~n40860 ) ;
  assign n46816 = n46815 ^ n1262 ^ x243 ;
  assign n46817 = ~n9656 & n14669 ;
  assign n46818 = n21518 & n46817 ;
  assign n46819 = n46818 ^ n46808 ^ n26202 ;
  assign n46820 = n1462 & ~n7886 ;
  assign n46821 = ~n8600 & n46820 ;
  assign n46822 = ( ~n3988 & n41734 ) | ( ~n3988 & n46821 ) | ( n41734 & n46821 ) ;
  assign n46823 = n15681 & ~n31115 ;
  assign n46824 = n14770 & n46823 ;
  assign n46825 = n46824 ^ n24044 ^ 1'b0 ;
  assign n46826 = n44044 ^ n2907 ^ 1'b0 ;
  assign n46827 = ( n11060 & n12485 ) | ( n11060 & ~n25452 ) | ( n12485 & ~n25452 ) ;
  assign n46828 = n7289 | n36397 ;
  assign n46829 = ( n6973 & n46827 ) | ( n6973 & n46828 ) | ( n46827 & n46828 ) ;
  assign n46830 = n13461 | n24184 ;
  assign n46831 = n46829 & ~n46830 ;
  assign n46832 = ~n12737 & n13786 ;
  assign n46833 = ~n17617 & n46832 ;
  assign n46834 = n5756 | n46833 ;
  assign n46835 = n7763 | n46834 ;
  assign n46836 = n45699 ^ n2778 ^ 1'b0 ;
  assign n46837 = n18242 ^ n16871 ^ 1'b0 ;
  assign n46838 = n5521 & n46837 ;
  assign n46839 = n26789 & n46838 ;
  assign n46840 = ( ~n3986 & n5249 ) | ( ~n3986 & n22143 ) | ( n5249 & n22143 ) ;
  assign n46841 = n23503 | n32823 ;
  assign n46842 = ~n4673 & n20808 ;
  assign n46843 = n37161 & n46842 ;
  assign n46844 = n46843 ^ n14344 ^ 1'b0 ;
  assign n46845 = n43313 ^ n22229 ^ n15744 ;
  assign n46846 = ~n45725 & n46845 ;
  assign n46847 = ( ~n520 & n14437 ) | ( ~n520 & n46846 ) | ( n14437 & n46846 ) ;
  assign n46848 = n46847 ^ n42320 ^ n16268 ;
  assign n46849 = n34402 ^ n31069 ^ n31058 ;
  assign n46850 = ~n7073 & n29963 ;
  assign n46851 = n46850 ^ n46759 ^ n4282 ;
  assign n46852 = ( ~n7449 & n30008 ) | ( ~n7449 & n33609 ) | ( n30008 & n33609 ) ;
  assign n46853 = n15322 | n46852 ;
  assign n46854 = n1905 | n46853 ;
  assign n46855 = n16834 ^ n8063 ^ 1'b0 ;
  assign n46856 = n2657 & ~n13024 ;
  assign n46857 = n46856 ^ n42593 ^ 1'b0 ;
  assign n46858 = n12727 | n29392 ;
  assign n46859 = n46858 ^ n42534 ^ n7049 ;
  assign n46860 = n23276 ^ n9614 ^ n4409 ;
  assign n46862 = n35418 ^ n24549 ^ 1'b0 ;
  assign n46861 = n1433 | n3948 ;
  assign n46863 = n46862 ^ n46861 ^ n13985 ;
  assign n46864 = n46863 ^ n40790 ^ n19730 ;
  assign n46865 = ~n15614 & n17930 ;
  assign n46866 = n46865 ^ n36095 ^ 1'b0 ;
  assign n46867 = n16259 & n22066 ;
  assign n46868 = ~n12667 & n46867 ;
  assign n46869 = n46868 ^ n30930 ^ 1'b0 ;
  assign n46870 = ~n39990 & n46869 ;
  assign n46871 = ( n4579 & n4931 ) | ( n4579 & ~n5352 ) | ( n4931 & ~n5352 ) ;
  assign n46872 = n13115 ^ n7259 ^ 1'b0 ;
  assign n46873 = n46871 | n46872 ;
  assign n46874 = n1985 & ~n15318 ;
  assign n46875 = n46874 ^ n20222 ^ n7692 ;
  assign n46876 = n34827 & ~n46875 ;
  assign n46877 = n18619 ^ n14406 ^ n4976 ;
  assign n46878 = n46877 ^ n33043 ^ n23274 ;
  assign n46879 = ( n1071 & n19533 ) | ( n1071 & ~n46878 ) | ( n19533 & ~n46878 ) ;
  assign n46880 = n8748 | n46879 ;
  assign n46881 = n5601 ^ n3979 ^ n588 ;
  assign n46882 = n31811 ^ n937 ^ 1'b0 ;
  assign n46883 = ( n4729 & n9954 ) | ( n4729 & ~n37054 ) | ( n9954 & ~n37054 ) ;
  assign n46884 = ~n20047 & n46883 ;
  assign n46885 = n46884 ^ n3466 ^ 1'b0 ;
  assign n46886 = n46885 ^ n6324 ^ n1064 ;
  assign n46887 = n42718 ^ n26113 ^ n14667 ;
  assign n46888 = n23090 ^ n17296 ^ 1'b0 ;
  assign n46889 = n18755 | n46888 ;
  assign n46890 = n2166 & ~n3416 ;
  assign n46891 = n46890 ^ n35731 ^ n5036 ;
  assign n46892 = ( n16136 & ~n46889 ) | ( n16136 & n46891 ) | ( ~n46889 & n46891 ) ;
  assign n46893 = n9166 & n19670 ;
  assign n46894 = ~n43178 & n46893 ;
  assign n46895 = n18154 & ~n31342 ;
  assign n46896 = n9048 & n46895 ;
  assign n46897 = ( ~n3864 & n27209 ) | ( ~n3864 & n44904 ) | ( n27209 & n44904 ) ;
  assign n46898 = ( ~n8349 & n12426 ) | ( ~n8349 & n13217 ) | ( n12426 & n13217 ) ;
  assign n46899 = ( n17262 & n17480 ) | ( n17262 & ~n46898 ) | ( n17480 & ~n46898 ) ;
  assign n46900 = n8400 & n38326 ;
  assign n46901 = n46900 ^ n14868 ^ n8221 ;
  assign n46902 = n5431 & ~n23737 ;
  assign n46904 = n4284 & ~n18239 ;
  assign n46905 = n46904 ^ n2572 ^ 1'b0 ;
  assign n46906 = ( ~n17613 & n31603 ) | ( ~n17613 & n46905 ) | ( n31603 & n46905 ) ;
  assign n46903 = ~n43051 & n44840 ;
  assign n46907 = n46906 ^ n46903 ^ 1'b0 ;
  assign n46908 = n28225 ^ n17556 ^ n8291 ;
  assign n46909 = n46908 ^ n7535 ^ 1'b0 ;
  assign n46910 = n17079 & n46909 ;
  assign n46911 = n30731 & ~n38381 ;
  assign n46912 = ( n20405 & n45495 ) | ( n20405 & n46911 ) | ( n45495 & n46911 ) ;
  assign n46913 = ( ~n2115 & n22320 ) | ( ~n2115 & n35045 ) | ( n22320 & n35045 ) ;
  assign n46914 = n4636 & ~n5984 ;
  assign n46915 = ~n33511 & n46914 ;
  assign n46916 = ( n31420 & ~n42671 ) | ( n31420 & n46915 ) | ( ~n42671 & n46915 ) ;
  assign n46919 = ~n19879 & n33537 ;
  assign n46920 = n46919 ^ n3486 ^ 1'b0 ;
  assign n46921 = n46920 ^ n37824 ^ n25249 ;
  assign n46917 = n2228 | n22200 ;
  assign n46918 = n46917 ^ n10604 ^ 1'b0 ;
  assign n46922 = n46921 ^ n46918 ^ n9028 ;
  assign n46923 = n43229 ^ n5128 ^ 1'b0 ;
  assign n46924 = ~n34932 & n46923 ;
  assign n46925 = ( n30103 & ~n46922 ) | ( n30103 & n46924 ) | ( ~n46922 & n46924 ) ;
  assign n46926 = n20017 ^ n10151 ^ 1'b0 ;
  assign n46927 = n4033 & n46926 ;
  assign n46928 = n15036 & n46927 ;
  assign n46929 = ~n43460 & n46928 ;
  assign n46930 = n19898 & ~n37223 ;
  assign n46931 = n46929 & n46930 ;
  assign n46932 = n20014 ^ n2483 ^ 1'b0 ;
  assign n46933 = ( ~n2200 & n3834 ) | ( ~n2200 & n6074 ) | ( n3834 & n6074 ) ;
  assign n46934 = n46932 & n46933 ;
  assign n46936 = ( n7887 & n11460 ) | ( n7887 & n33823 ) | ( n11460 & n33823 ) ;
  assign n46937 = ( ~n3880 & n42842 ) | ( ~n3880 & n46936 ) | ( n42842 & n46936 ) ;
  assign n46935 = n12594 | n28652 ;
  assign n46938 = n46937 ^ n46935 ^ 1'b0 ;
  assign n46939 = ( n5076 & ~n38381 ) | ( n5076 & n45495 ) | ( ~n38381 & n45495 ) ;
  assign n46940 = n16146 & n16423 ;
  assign n46941 = ~n36141 & n46940 ;
  assign n46942 = n46941 ^ n14073 ^ 1'b0 ;
  assign n46943 = ( ~n3075 & n3922 ) | ( ~n3075 & n20321 ) | ( n3922 & n20321 ) ;
  assign n46944 = ( n12144 & ~n26195 ) | ( n12144 & n37917 ) | ( ~n26195 & n37917 ) ;
  assign n46945 = n24867 | n38159 ;
  assign n46946 = n13506 | n46945 ;
  assign n46947 = n31659 ^ n8761 ^ 1'b0 ;
  assign n46948 = ~n41036 & n46947 ;
  assign n46949 = n20440 & n40698 ;
  assign n46950 = n46949 ^ n34875 ^ 1'b0 ;
  assign n46951 = n2679 ^ n426 ^ 1'b0 ;
  assign n46952 = n24776 ^ n10599 ^ 1'b0 ;
  assign n46953 = n18841 & ~n41482 ;
  assign n46954 = ~n9447 & n46953 ;
  assign n46956 = n21698 ^ n7890 ^ 1'b0 ;
  assign n46957 = ~n3046 & n46956 ;
  assign n46955 = ( n1765 & n26009 ) | ( n1765 & n45763 ) | ( n26009 & n45763 ) ;
  assign n46958 = n46957 ^ n46955 ^ n7509 ;
  assign n46959 = ( n3343 & n20167 ) | ( n3343 & n46958 ) | ( n20167 & n46958 ) ;
  assign n46960 = n46959 ^ n32312 ^ n22813 ;
  assign n46961 = ( n33687 & ~n46954 ) | ( n33687 & n46960 ) | ( ~n46954 & n46960 ) ;
  assign n46962 = n738 ^ n286 ^ 1'b0 ;
  assign n46963 = n14973 & ~n17311 ;
  assign n46964 = ( n8978 & n15945 ) | ( n8978 & ~n46963 ) | ( n15945 & ~n46963 ) ;
  assign n46965 = ( ~n9507 & n46962 ) | ( ~n9507 & n46964 ) | ( n46962 & n46964 ) ;
  assign n46966 = n2832 | n20953 ;
  assign n46967 = ( ~n14966 & n21952 ) | ( ~n14966 & n30032 ) | ( n21952 & n30032 ) ;
  assign n46968 = ( n8969 & n10241 ) | ( n8969 & ~n46967 ) | ( n10241 & ~n46967 ) ;
  assign n46969 = n26107 ^ n2592 ^ n2171 ;
  assign n46970 = n13176 ^ n5363 ^ n1073 ;
  assign n46971 = ~n20461 & n46970 ;
  assign n46972 = n46971 ^ n20867 ^ 1'b0 ;
  assign n46973 = n16138 & n18083 ;
  assign n46974 = n46973 ^ n14757 ^ 1'b0 ;
  assign n46975 = ~n30350 & n44744 ;
  assign n46976 = n25794 & n46975 ;
  assign n46977 = n14772 | n33694 ;
  assign n46978 = n8612 | n46977 ;
  assign n46979 = n46978 ^ n24785 ^ 1'b0 ;
  assign n46980 = ( x225 & ~n570 ) | ( x225 & n3405 ) | ( ~n570 & n3405 ) ;
  assign n46981 = n46980 ^ n28639 ^ 1'b0 ;
  assign n46982 = ~n46979 & n46981 ;
  assign n46984 = n15641 | n21101 ;
  assign n46985 = n46984 ^ n18191 ^ 1'b0 ;
  assign n46983 = n26797 ^ n24341 ^ 1'b0 ;
  assign n46986 = n46985 ^ n46983 ^ n22401 ;
  assign n46987 = n46986 ^ n3889 ^ 1'b0 ;
  assign n46988 = n16309 ^ n11937 ^ 1'b0 ;
  assign n46989 = ( ~n39684 & n42525 ) | ( ~n39684 & n46988 ) | ( n42525 & n46988 ) ;
  assign n46990 = n2448 & ~n6791 ;
  assign n46991 = ~n20398 & n46990 ;
  assign n46992 = n46991 ^ n42223 ^ n14202 ;
  assign n46993 = n44240 ^ n31750 ^ n8496 ;
  assign n46994 = ~n14272 & n46993 ;
  assign n46995 = ( n6031 & n26939 ) | ( n6031 & n35679 ) | ( n26939 & n35679 ) ;
  assign n47005 = n35566 ^ n15180 ^ n9369 ;
  assign n47006 = ~n14579 & n20696 ;
  assign n47007 = n47005 | n47006 ;
  assign n47008 = n47007 ^ n24672 ^ 1'b0 ;
  assign n47009 = ( n1138 & ~n13406 ) | ( n1138 & n47008 ) | ( ~n13406 & n47008 ) ;
  assign n46996 = ~n7290 & n9337 ;
  assign n46997 = n19215 & n46996 ;
  assign n46998 = n20524 & ~n46997 ;
  assign n46999 = n25947 & n46998 ;
  assign n47000 = n46999 ^ n18708 ^ n4271 ;
  assign n47001 = n33699 ^ n2784 ^ 1'b0 ;
  assign n47002 = n1416 & n47001 ;
  assign n47003 = n47002 ^ n7094 ^ 1'b0 ;
  assign n47004 = n47000 | n47003 ;
  assign n47010 = n47009 ^ n47004 ^ n9357 ;
  assign n47011 = n47010 ^ n46157 ^ n28694 ;
  assign n47012 = n14311 ^ n14093 ^ 1'b0 ;
  assign n47013 = n2096 | n36991 ;
  assign n47014 = n47012 | n47013 ;
  assign n47015 = n47014 ^ n3069 ^ 1'b0 ;
  assign n47016 = ~n3841 & n47015 ;
  assign n47017 = n47016 ^ n11888 ^ n1007 ;
  assign n47018 = n47017 ^ n13648 ^ n4123 ;
  assign n47019 = n7579 | n43898 ;
  assign n47020 = n47018 & ~n47019 ;
  assign n47021 = n42979 ^ n9724 ^ 1'b0 ;
  assign n47022 = n26230 | n47021 ;
  assign n47030 = n30025 ^ n24489 ^ 1'b0 ;
  assign n47031 = n15943 & n47030 ;
  assign n47023 = ~n6446 & n16464 ;
  assign n47024 = ( n1884 & n5850 ) | ( n1884 & ~n47023 ) | ( n5850 & ~n47023 ) ;
  assign n47025 = n12199 & n22096 ;
  assign n47026 = ( ~n3271 & n47024 ) | ( ~n3271 & n47025 ) | ( n47024 & n47025 ) ;
  assign n47027 = n16712 | n47026 ;
  assign n47028 = n47027 ^ x0 ^ 1'b0 ;
  assign n47029 = n7047 & n47028 ;
  assign n47032 = n47031 ^ n47029 ^ 1'b0 ;
  assign n47033 = n19831 & ~n30931 ;
  assign n47034 = ( n3261 & n24388 ) | ( n3261 & ~n28225 ) | ( n24388 & ~n28225 ) ;
  assign n47035 = n31234 ^ n21833 ^ n11831 ;
  assign n47036 = n47035 ^ n43612 ^ n43534 ;
  assign n47037 = ( n8691 & n12280 ) | ( n8691 & n12874 ) | ( n12280 & n12874 ) ;
  assign n47038 = n42781 | n47037 ;
  assign n47040 = ( n9564 & n37823 ) | ( n9564 & ~n45940 ) | ( n37823 & ~n45940 ) ;
  assign n47039 = n8854 | n31344 ;
  assign n47041 = n47040 ^ n47039 ^ 1'b0 ;
  assign n47042 = n35484 & ~n47041 ;
  assign n47043 = n47042 ^ n37389 ^ n19061 ;
  assign n47044 = ~n15245 & n36036 ;
  assign n47045 = n32432 ^ n19786 ^ n17543 ;
  assign n47046 = n47045 ^ n7496 ^ 1'b0 ;
  assign n47047 = n23104 | n47046 ;
  assign n47048 = n42920 ^ n20848 ^ 1'b0 ;
  assign n47049 = ~n12082 & n47048 ;
  assign n47050 = n9801 & n40116 ;
  assign n47051 = ( ~n18335 & n19558 ) | ( ~n18335 & n25596 ) | ( n19558 & n25596 ) ;
  assign n47052 = n47051 ^ n35234 ^ n21190 ;
  assign n47053 = n34930 | n43996 ;
  assign n47054 = ( n7330 & n19799 ) | ( n7330 & n47053 ) | ( n19799 & n47053 ) ;
  assign n47055 = ( n10640 & n28743 ) | ( n10640 & n31482 ) | ( n28743 & n31482 ) ;
  assign n47056 = ( n6720 & ~n18215 ) | ( n6720 & n38670 ) | ( ~n18215 & n38670 ) ;
  assign n47057 = n18284 ^ n1367 ^ 1'b0 ;
  assign n47058 = n19238 & n47057 ;
  assign n47059 = ( n4272 & ~n40116 ) | ( n4272 & n47058 ) | ( ~n40116 & n47058 ) ;
  assign n47063 = n36512 ^ n14946 ^ 1'b0 ;
  assign n47060 = n25199 ^ n2977 ^ 1'b0 ;
  assign n47061 = n9166 & n47060 ;
  assign n47062 = ~n9530 & n47061 ;
  assign n47064 = n47063 ^ n47062 ^ 1'b0 ;
  assign n47065 = n2333 & ~n17201 ;
  assign n47066 = n47065 ^ n14142 ^ 1'b0 ;
  assign n47067 = n18370 & n18562 ;
  assign n47068 = ~n9132 & n47067 ;
  assign n47069 = ( n566 & n2409 ) | ( n566 & ~n17169 ) | ( n2409 & ~n17169 ) ;
  assign n47070 = ( ~n737 & n13519 ) | ( ~n737 & n16452 ) | ( n13519 & n16452 ) ;
  assign n47071 = ( n8222 & n16448 ) | ( n8222 & ~n47070 ) | ( n16448 & ~n47070 ) ;
  assign n47072 = ( n4613 & ~n47069 ) | ( n4613 & n47071 ) | ( ~n47069 & n47071 ) ;
  assign n47075 = ( n8260 & ~n33146 ) | ( n8260 & n43951 ) | ( ~n33146 & n43951 ) ;
  assign n47073 = n16052 ^ n3052 ^ 1'b0 ;
  assign n47074 = n17787 | n47073 ;
  assign n47076 = n47075 ^ n47074 ^ 1'b0 ;
  assign n47077 = n44967 ^ n25053 ^ n1206 ;
  assign n47078 = ~n11043 & n21054 ;
  assign n47079 = n47078 ^ n10201 ^ 1'b0 ;
  assign n47080 = n47079 ^ n21221 ^ n16677 ;
  assign n47081 = ( n2084 & ~n3993 ) | ( n2084 & n4568 ) | ( ~n3993 & n4568 ) ;
  assign n47082 = n47081 ^ n4630 ^ 1'b0 ;
  assign n47083 = n47080 | n47082 ;
  assign n47084 = ( n34592 & n39378 ) | ( n34592 & n45316 ) | ( n39378 & n45316 ) ;
  assign n47089 = n35719 ^ n32599 ^ n29493 ;
  assign n47085 = n1264 & n8509 ;
  assign n47086 = n17205 & n47085 ;
  assign n47087 = n47086 ^ n672 ^ 1'b0 ;
  assign n47088 = ( n8494 & ~n14595 ) | ( n8494 & n47087 ) | ( ~n14595 & n47087 ) ;
  assign n47090 = n47089 ^ n47088 ^ n21230 ;
  assign n47091 = n24083 | n39656 ;
  assign n47092 = n43460 | n47091 ;
  assign n47093 = n28021 ^ n681 ^ 1'b0 ;
  assign n47094 = ~n14934 & n47093 ;
  assign n47095 = ( ~n1628 & n15170 ) | ( ~n1628 & n25570 ) | ( n15170 & n25570 ) ;
  assign n47096 = n47095 ^ n27537 ^ 1'b0 ;
  assign n47097 = n13112 & ~n14130 ;
  assign n47098 = ( ~n23890 & n27138 ) | ( ~n23890 & n29094 ) | ( n27138 & n29094 ) ;
  assign n47099 = n14728 ^ n14090 ^ n9096 ;
  assign n47100 = ( ~n729 & n15726 ) | ( ~n729 & n47099 ) | ( n15726 & n47099 ) ;
  assign n47101 = n32640 & n35739 ;
  assign n47102 = n47101 ^ n22313 ^ 1'b0 ;
  assign n47103 = n47102 ^ n22251 ^ 1'b0 ;
  assign n47104 = n47103 ^ n7922 ^ 1'b0 ;
  assign n47105 = n24522 & n47104 ;
  assign n47106 = n31317 & ~n34580 ;
  assign n47107 = n47106 ^ n15795 ^ 1'b0 ;
  assign n47108 = ~n9087 & n16913 ;
  assign n47109 = n18977 | n47108 ;
  assign n47110 = n47109 ^ n46449 ^ 1'b0 ;
  assign n47111 = ~n29274 & n30478 ;
  assign n47112 = n8646 & n47111 ;
  assign n47114 = n8127 | n23963 ;
  assign n47115 = n47114 ^ n33509 ^ 1'b0 ;
  assign n47113 = n29357 & n32613 ;
  assign n47116 = n47115 ^ n47113 ^ 1'b0 ;
  assign n47117 = ~n7653 & n13438 ;
  assign n47118 = n47117 ^ n17640 ^ 1'b0 ;
  assign n47119 = ~n45246 & n47118 ;
  assign n47120 = n32029 ^ n6879 ^ n6184 ;
  assign n47121 = n25491 ^ n22248 ^ n15624 ;
  assign n47122 = n30354 ^ n30019 ^ n25288 ;
  assign n47123 = ~n437 & n3761 ;
  assign n47124 = n47123 ^ n27180 ^ 1'b0 ;
  assign n47125 = ( n1289 & n13047 ) | ( n1289 & ~n47124 ) | ( n13047 & ~n47124 ) ;
  assign n47126 = ( n9266 & n21298 ) | ( n9266 & n21835 ) | ( n21298 & n21835 ) ;
  assign n47127 = ( n21172 & ~n23926 ) | ( n21172 & n24581 ) | ( ~n23926 & n24581 ) ;
  assign n47128 = n47127 ^ n19438 ^ n6255 ;
  assign n47129 = ( n45168 & ~n47126 ) | ( n45168 & n47128 ) | ( ~n47126 & n47128 ) ;
  assign n47130 = n8922 & ~n47129 ;
  assign n47131 = n47125 & n47130 ;
  assign n47132 = n47131 ^ n29101 ^ n18139 ;
  assign n47133 = n34353 ^ n13438 ^ n6421 ;
  assign n47134 = n7502 | n13733 ;
  assign n47135 = n4974 & ~n47134 ;
  assign n47136 = n6670 & n9011 ;
  assign n47137 = ~n14115 & n47136 ;
  assign n47138 = n29813 ^ n12537 ^ 1'b0 ;
  assign n47139 = n24033 ^ n20295 ^ n6046 ;
  assign n47140 = n19541 ^ n15028 ^ 1'b0 ;
  assign n47141 = n1916 | n8132 ;
  assign n47142 = n47141 ^ n32567 ^ n11625 ;
  assign n47143 = n47142 ^ n18487 ^ n6458 ;
  assign n47144 = ~n24058 & n29317 ;
  assign n47145 = n47144 ^ n22138 ^ 1'b0 ;
  assign n47146 = n27672 | n47145 ;
  assign n47147 = n40031 | n47146 ;
  assign n47148 = n2797 & ~n18611 ;
  assign n47149 = n47148 ^ n43428 ^ 1'b0 ;
  assign n47150 = ~n21945 & n47149 ;
  assign n47151 = n38651 ^ n8546 ^ n1733 ;
  assign n47152 = n47151 ^ n26117 ^ n2060 ;
  assign n47153 = n47152 ^ n35326 ^ n35099 ;
  assign n47154 = ( n2113 & n12860 ) | ( n2113 & n36100 ) | ( n12860 & n36100 ) ;
  assign n47155 = n5907 & ~n19122 ;
  assign n47156 = n47155 ^ n18382 ^ 1'b0 ;
  assign n47157 = n22427 ^ n12682 ^ 1'b0 ;
  assign n47158 = ( n5054 & n5881 ) | ( n5054 & ~n27697 ) | ( n5881 & ~n27697 ) ;
  assign n47159 = ( ~n47156 & n47157 ) | ( ~n47156 & n47158 ) | ( n47157 & n47158 ) ;
  assign n47160 = ( n5657 & n9279 ) | ( n5657 & n16526 ) | ( n9279 & n16526 ) ;
  assign n47161 = n20202 ^ n5551 ^ 1'b0 ;
  assign n47162 = ~n33928 & n47161 ;
  assign n47163 = n47162 ^ n29886 ^ n8935 ;
  assign n47164 = n44864 ^ n32507 ^ 1'b0 ;
  assign n47165 = ~n6851 & n42868 ;
  assign n47166 = n44333 & n47165 ;
  assign n47167 = n31183 ^ n22162 ^ n5781 ;
  assign n47169 = n17475 ^ n14716 ^ n1826 ;
  assign n47168 = ~n290 & n13312 ;
  assign n47170 = n47169 ^ n47168 ^ 1'b0 ;
  assign n47171 = n47167 & n47170 ;
  assign n47172 = n14287 & n47171 ;
  assign n47173 = n18148 & ~n47172 ;
  assign n47175 = n33543 ^ n23156 ^ 1'b0 ;
  assign n47176 = n47175 ^ n20218 ^ 1'b0 ;
  assign n47177 = ~n26126 & n47176 ;
  assign n47174 = ~n23196 & n43154 ;
  assign n47178 = n47177 ^ n47174 ^ n4539 ;
  assign n47179 = n35984 ^ n28927 ^ n10083 ;
  assign n47180 = n19656 ^ n4572 ^ 1'b0 ;
  assign n47181 = n5266 | n47180 ;
  assign n47182 = n47181 ^ n14393 ^ 1'b0 ;
  assign n47183 = ( n40093 & n47179 ) | ( n40093 & n47182 ) | ( n47179 & n47182 ) ;
  assign n47184 = n18697 ^ n18072 ^ n12585 ;
  assign n47185 = n14255 | n20791 ;
  assign n47186 = n15018 | n47185 ;
  assign n47187 = n47186 ^ n24724 ^ n13729 ;
  assign n47188 = ( ~n1988 & n16369 ) | ( ~n1988 & n18688 ) | ( n16369 & n18688 ) ;
  assign n47190 = ~n6351 & n34196 ;
  assign n47189 = n11270 & ~n14972 ;
  assign n47191 = n47190 ^ n47189 ^ 1'b0 ;
  assign n47192 = n6522 & n46770 ;
  assign n47193 = ~n33741 & n47192 ;
  assign n47194 = n775 & n38706 ;
  assign n47195 = n9288 & n47194 ;
  assign n47196 = n39551 ^ n11122 ^ n1908 ;
  assign n47197 = n47196 ^ n29423 ^ 1'b0 ;
  assign n47198 = ( ~n24213 & n34859 ) | ( ~n24213 & n39121 ) | ( n34859 & n39121 ) ;
  assign n47199 = n47198 ^ n44860 ^ 1'b0 ;
  assign n47200 = n16108 ^ n14456 ^ n7509 ;
  assign n47201 = ( ~x112 & n40415 ) | ( ~x112 & n43286 ) | ( n40415 & n43286 ) ;
  assign n47202 = n7370 & n13483 ;
  assign n47203 = n47202 ^ n10396 ^ 1'b0 ;
  assign n47204 = n47203 ^ n34659 ^ n18388 ;
  assign n47206 = ( n6789 & n7289 ) | ( n6789 & n13870 ) | ( n7289 & n13870 ) ;
  assign n47207 = ~n5800 & n47206 ;
  assign n47205 = n24519 ^ n20385 ^ 1'b0 ;
  assign n47208 = n47207 ^ n47205 ^ n14819 ;
  assign n47209 = n12812 | n22403 ;
  assign n47210 = n4629 & n7446 ;
  assign n47211 = n36619 ^ n13499 ^ 1'b0 ;
  assign n47212 = n12479 | n47211 ;
  assign n47213 = n38139 ^ n31980 ^ n13000 ;
  assign n47214 = ( n47210 & ~n47212 ) | ( n47210 & n47213 ) | ( ~n47212 & n47213 ) ;
  assign n47215 = n47214 ^ n9043 ^ 1'b0 ;
  assign n47216 = n10445 ^ n4902 ^ 1'b0 ;
  assign n47217 = ~n3136 & n16378 ;
  assign n47218 = n47217 ^ n6107 ^ 1'b0 ;
  assign n47220 = ( n18409 & n18628 ) | ( n18409 & n20123 ) | ( n18628 & n20123 ) ;
  assign n47219 = n18428 & ~n35340 ;
  assign n47221 = n47220 ^ n47219 ^ 1'b0 ;
  assign n47222 = ( n3111 & n8639 ) | ( n3111 & ~n37060 ) | ( n8639 & ~n37060 ) ;
  assign n47223 = ~n23223 & n24692 ;
  assign n47224 = n33790 ^ n27206 ^ n13279 ;
  assign n47225 = ( n8634 & n28272 ) | ( n8634 & n47224 ) | ( n28272 & n47224 ) ;
  assign n47226 = n33765 ^ n19404 ^ n15688 ;
  assign n47227 = n11381 ^ n3046 ^ 1'b0 ;
  assign n47228 = n423 & n47227 ;
  assign n47229 = n47228 ^ n10111 ^ 1'b0 ;
  assign n47230 = n15467 & ~n47229 ;
  assign n47231 = n30933 ^ n23074 ^ n3085 ;
  assign n47232 = n24851 ^ n17067 ^ n12838 ;
  assign n47233 = ( n15258 & n47231 ) | ( n15258 & n47232 ) | ( n47231 & n47232 ) ;
  assign n47234 = n40402 ^ n13149 ^ n824 ;
  assign n47235 = n19820 ^ n3761 ^ n1961 ;
  assign n47236 = n17065 & ~n31698 ;
  assign n47237 = n14113 ^ n306 ^ 1'b0 ;
  assign n47238 = n1284 | n47237 ;
  assign n47239 = n34780 & ~n47238 ;
  assign n47240 = n47239 ^ n32845 ^ 1'b0 ;
  assign n47241 = n13716 | n47240 ;
  assign n47242 = ~n7993 & n25772 ;
  assign n47243 = n47242 ^ n26080 ^ 1'b0 ;
  assign n47244 = n25396 ^ n2359 ^ 1'b0 ;
  assign n47245 = ~n38275 & n47244 ;
  assign n47246 = ~n17321 & n47245 ;
  assign n47247 = n14031 | n42512 ;
  assign n47248 = n910 | n47247 ;
  assign n47249 = n37704 ^ n35253 ^ n29957 ;
  assign n47250 = n22097 & ~n30401 ;
  assign n47251 = n26803 | n47250 ;
  assign n47252 = n12837 ^ n2539 ^ 1'b0 ;
  assign n47253 = ( n26991 & n46677 ) | ( n26991 & ~n47252 ) | ( n46677 & ~n47252 ) ;
  assign n47254 = n12916 ^ n8177 ^ n7308 ;
  assign n47255 = n47254 ^ n14991 ^ n6550 ;
  assign n47256 = ( n17998 & ~n26500 ) | ( n17998 & n42337 ) | ( ~n26500 & n42337 ) ;
  assign n47257 = ( ~n38876 & n40585 ) | ( ~n38876 & n47256 ) | ( n40585 & n47256 ) ;
  assign n47258 = ( n4313 & n14433 ) | ( n4313 & ~n19328 ) | ( n14433 & ~n19328 ) ;
  assign n47259 = n42114 ^ n16184 ^ 1'b0 ;
  assign n47260 = ~n33664 & n47259 ;
  assign n47261 = n14318 ^ n391 ^ 1'b0 ;
  assign n47262 = n20601 & n47261 ;
  assign n47263 = n47262 ^ n24104 ^ 1'b0 ;
  assign n47264 = ( n4124 & n16684 ) | ( n4124 & ~n18842 ) | ( n16684 & ~n18842 ) ;
  assign n47265 = n32570 | n47264 ;
  assign n47266 = n33694 | n47265 ;
  assign n47267 = n36170 | n45252 ;
  assign n47268 = n40293 ^ n28002 ^ n24251 ;
  assign n47269 = n38673 ^ n18436 ^ n10169 ;
  assign n47270 = ( ~n6282 & n22047 ) | ( ~n6282 & n47269 ) | ( n22047 & n47269 ) ;
  assign n47271 = ( n4912 & n8901 ) | ( n4912 & n47270 ) | ( n8901 & n47270 ) ;
  assign n47272 = n12767 & ~n39812 ;
  assign n47275 = n41704 ^ n30984 ^ 1'b0 ;
  assign n47273 = ( n1282 & ~n4791 ) | ( n1282 & n28291 ) | ( ~n4791 & n28291 ) ;
  assign n47274 = ( n22891 & n23251 ) | ( n22891 & ~n47273 ) | ( n23251 & ~n47273 ) ;
  assign n47276 = n47275 ^ n47274 ^ n1832 ;
  assign n47277 = n27441 ^ n26095 ^ n2582 ;
  assign n47278 = ( n1772 & n5637 ) | ( n1772 & n6908 ) | ( n5637 & n6908 ) ;
  assign n47279 = ~n3627 & n47278 ;
  assign n47280 = n42697 & n47279 ;
  assign n47281 = n35938 ^ n25565 ^ n22091 ;
  assign n47282 = n47281 ^ n30047 ^ n29666 ;
  assign n47283 = n47282 ^ n41891 ^ 1'b0 ;
  assign n47285 = ~n4642 & n18286 ;
  assign n47286 = n47285 ^ n2885 ^ 1'b0 ;
  assign n47284 = n42138 | n42207 ;
  assign n47287 = n47286 ^ n47284 ^ 1'b0 ;
  assign n47288 = n14609 ^ n9427 ^ 1'b0 ;
  assign n47289 = n3342 & n26776 ;
  assign n47290 = n6984 & n47289 ;
  assign n47291 = ~n9786 & n37485 ;
  assign n47292 = n47291 ^ n33284 ^ 1'b0 ;
  assign n47293 = n45816 ^ n37066 ^ 1'b0 ;
  assign n47294 = ~n2873 & n22405 ;
  assign n47295 = n3398 & n13464 ;
  assign n47296 = n37906 ^ n33598 ^ n5890 ;
  assign n47297 = n44648 ^ n41335 ^ n10029 ;
  assign n47298 = n41223 ^ n31961 ^ 1'b0 ;
  assign n47299 = n15912 & ~n47298 ;
  assign n47300 = n47299 ^ n23635 ^ 1'b0 ;
  assign n47301 = ~n14456 & n47300 ;
  assign n47302 = n44477 ^ n21366 ^ 1'b0 ;
  assign n47303 = n32790 & n47302 ;
  assign n47304 = ~n5002 & n12224 ;
  assign n47305 = n12576 & ~n31983 ;
  assign n47306 = n24130 & n47305 ;
  assign n47307 = n47306 ^ n20882 ^ n8857 ;
  assign n47308 = ( n16723 & n20581 ) | ( n16723 & n38535 ) | ( n20581 & n38535 ) ;
  assign n47309 = n19844 ^ n7286 ^ 1'b0 ;
  assign n47310 = ( n6528 & n15225 ) | ( n6528 & n47309 ) | ( n15225 & n47309 ) ;
  assign n47311 = n3750 & n5559 ;
  assign n47312 = ~n47124 & n47311 ;
  assign n47313 = n47312 ^ n24864 ^ n567 ;
  assign n47314 = ( n3632 & n8329 ) | ( n3632 & n14690 ) | ( n8329 & n14690 ) ;
  assign n47315 = n47314 ^ n20131 ^ 1'b0 ;
  assign n47316 = n35917 & ~n47315 ;
  assign n47317 = n7659 & ~n10361 ;
  assign n47318 = ~n31516 & n47317 ;
  assign n47319 = n22770 & n30947 ;
  assign n47320 = n38096 ^ n9102 ^ n6673 ;
  assign n47321 = n16169 | n29829 ;
  assign n47322 = ( n18187 & n21342 ) | ( n18187 & n47321 ) | ( n21342 & n47321 ) ;
  assign n47323 = ( n3487 & n25882 ) | ( n3487 & ~n44120 ) | ( n25882 & ~n44120 ) ;
  assign n47324 = n14515 ^ n12887 ^ 1'b0 ;
  assign n47325 = n317 & ~n47324 ;
  assign n47326 = n40116 ^ n37320 ^ n24887 ;
  assign n47327 = ( n16000 & n47325 ) | ( n16000 & n47326 ) | ( n47325 & n47326 ) ;
  assign n47328 = ( n1725 & n3575 ) | ( n1725 & n23605 ) | ( n3575 & n23605 ) ;
  assign n47329 = n41877 ^ x218 ^ 1'b0 ;
  assign n47330 = n35444 | n47329 ;
  assign n47331 = ( n9312 & n25081 ) | ( n9312 & n47330 ) | ( n25081 & n47330 ) ;
  assign n47332 = n47331 ^ n6444 ^ n2999 ;
  assign n47333 = ( n2464 & ~n22570 ) | ( n2464 & n26414 ) | ( ~n22570 & n26414 ) ;
  assign n47334 = n47333 ^ n13685 ^ 1'b0 ;
  assign n47335 = ~n22652 & n47334 ;
  assign n47336 = n47335 ^ n33782 ^ 1'b0 ;
  assign n47337 = n15667 & n47336 ;
  assign n47338 = n35531 ^ n7863 ^ 1'b0 ;
  assign n47339 = n35711 ^ n35085 ^ n12833 ;
  assign n47340 = n26195 ^ n5722 ^ 1'b0 ;
  assign n47341 = ~n47339 & n47340 ;
  assign n47342 = n9770 & n26315 ;
  assign n47343 = n40297 ^ n6762 ^ 1'b0 ;
  assign n47344 = ( n18784 & ~n20044 ) | ( n18784 & n23295 ) | ( ~n20044 & n23295 ) ;
  assign n47345 = n47344 ^ n39893 ^ n25988 ;
  assign n47346 = n43967 ^ n19907 ^ 1'b0 ;
  assign n47347 = ( ~n7692 & n33152 ) | ( ~n7692 & n45488 ) | ( n33152 & n45488 ) ;
  assign n47348 = ( n12252 & n16376 ) | ( n12252 & n47347 ) | ( n16376 & n47347 ) ;
  assign n47349 = ( ~n1227 & n38876 ) | ( ~n1227 & n43588 ) | ( n38876 & n43588 ) ;
  assign n47350 = n47349 ^ n9375 ^ n9142 ;
  assign n47351 = n47350 ^ n38670 ^ n15078 ;
  assign n47352 = n23465 ^ n23382 ^ 1'b0 ;
  assign n47353 = n4300 & ~n47352 ;
  assign n47354 = n47353 ^ n37846 ^ 1'b0 ;
  assign n47355 = ~n6569 & n12606 ;
  assign n47356 = ~n47354 & n47355 ;
  assign n47357 = n1193 | n29314 ;
  assign n47358 = n43030 ^ n30681 ^ 1'b0 ;
  assign n47359 = ~n47357 & n47358 ;
  assign n47360 = n15707 | n41158 ;
  assign n47361 = n34758 & ~n47360 ;
  assign n47362 = ( n6237 & ~n20968 ) | ( n6237 & n37298 ) | ( ~n20968 & n37298 ) ;
  assign n47365 = n15449 ^ n9941 ^ 1'b0 ;
  assign n47366 = n1450 & n47365 ;
  assign n47363 = ~n1664 & n6293 ;
  assign n47364 = ~n7587 & n47363 ;
  assign n47367 = n47366 ^ n47364 ^ n13400 ;
  assign n47368 = ( n8034 & ~n19238 ) | ( n8034 & n30248 ) | ( ~n19238 & n30248 ) ;
  assign n47369 = ( n7393 & n22621 ) | ( n7393 & n27556 ) | ( n22621 & n27556 ) ;
  assign n47370 = n30757 & n46983 ;
  assign n47371 = ( ~n10004 & n47369 ) | ( ~n10004 & n47370 ) | ( n47369 & n47370 ) ;
  assign n47372 = n3099 & n35187 ;
  assign n47373 = ( n6149 & ~n13806 ) | ( n6149 & n18046 ) | ( ~n13806 & n18046 ) ;
  assign n47374 = n32671 & ~n47373 ;
  assign n47375 = n9285 ^ n2076 ^ 1'b0 ;
  assign n47376 = n2463 & ~n3093 ;
  assign n47377 = n47375 & n47376 ;
  assign n47378 = n29159 | n47377 ;
  assign n47379 = ( n16663 & n21748 ) | ( n16663 & n46650 ) | ( n21748 & n46650 ) ;
  assign n47380 = n25991 ^ n9069 ^ n1193 ;
  assign n47381 = ( ~x235 & n17156 ) | ( ~x235 & n23064 ) | ( n17156 & n23064 ) ;
  assign n47382 = n47381 ^ n16155 ^ 1'b0 ;
  assign n47383 = ( n15880 & n22849 ) | ( n15880 & ~n24434 ) | ( n22849 & ~n24434 ) ;
  assign n47384 = ~n9794 & n13207 ;
  assign n47385 = n17179 & n47384 ;
  assign n47386 = ( n8732 & n27128 ) | ( n8732 & n47385 ) | ( n27128 & n47385 ) ;
  assign n47388 = n3626 ^ n2903 ^ x102 ;
  assign n47389 = ( n17609 & n42873 ) | ( n17609 & n47388 ) | ( n42873 & n47388 ) ;
  assign n47387 = n20759 & n40893 ;
  assign n47390 = n47389 ^ n47387 ^ 1'b0 ;
  assign n47391 = n12244 & n47390 ;
  assign n47392 = n37050 ^ n7922 ^ 1'b0 ;
  assign n47393 = n37386 & n47392 ;
  assign n47394 = n8761 & ~n24092 ;
  assign n47395 = n32291 & ~n47394 ;
  assign n47396 = ~n34619 & n47395 ;
  assign n47397 = n5388 | n11371 ;
  assign n47398 = n47397 ^ n2595 ^ 1'b0 ;
  assign n47399 = ( ~n5387 & n21750 ) | ( ~n5387 & n23906 ) | ( n21750 & n23906 ) ;
  assign n47400 = ( ~x165 & n1279 ) | ( ~x165 & n14439 ) | ( n1279 & n14439 ) ;
  assign n47401 = ( ~n16507 & n47399 ) | ( ~n16507 & n47400 ) | ( n47399 & n47400 ) ;
  assign n47402 = n37878 ^ n28794 ^ n6975 ;
  assign n47403 = n39473 ^ n21944 ^ 1'b0 ;
  assign n47404 = n11113 ^ n9064 ^ 1'b0 ;
  assign n47405 = n13781 & n47404 ;
  assign n47406 = ( n25322 & n47403 ) | ( n25322 & n47405 ) | ( n47403 & n47405 ) ;
  assign n47407 = n37203 ^ n16943 ^ 1'b0 ;
  assign n47408 = n47407 ^ n21867 ^ n10497 ;
  assign n47409 = n15910 & ~n36503 ;
  assign n47410 = n47409 ^ n38152 ^ 1'b0 ;
  assign n47411 = n11740 | n15296 ;
  assign n47412 = n21093 ^ n5725 ^ 1'b0 ;
  assign n47413 = n47411 & ~n47412 ;
  assign n47414 = n2257 & ~n17151 ;
  assign n47415 = n23013 & n47414 ;
  assign n47416 = n28301 ^ n26584 ^ 1'b0 ;
  assign n47417 = n37124 & ~n47416 ;
  assign n47418 = n6336 ^ n2365 ^ 1'b0 ;
  assign n47419 = n23446 & ~n47418 ;
  assign n47420 = n47419 ^ n5989 ^ x5 ;
  assign n47421 = ( n7042 & n47417 ) | ( n7042 & ~n47420 ) | ( n47417 & ~n47420 ) ;
  assign n47422 = n24533 ^ n5817 ^ 1'b0 ;
  assign n47423 = n24590 & ~n27727 ;
  assign n47424 = ~n339 & n47423 ;
  assign n47425 = ( n5717 & ~n17963 ) | ( n5717 & n47424 ) | ( ~n17963 & n47424 ) ;
  assign n47426 = n17854 & ~n22637 ;
  assign n47427 = n47426 ^ n22840 ^ 1'b0 ;
  assign n47428 = n47427 ^ n45914 ^ n18527 ;
  assign n47429 = ( ~n3040 & n6195 ) | ( ~n3040 & n16216 ) | ( n6195 & n16216 ) ;
  assign n47430 = n47429 ^ n33292 ^ n17795 ;
  assign n47431 = ( n4373 & ~n5617 ) | ( n4373 & n29757 ) | ( ~n5617 & n29757 ) ;
  assign n47432 = n13989 ^ n6356 ^ n3845 ;
  assign n47433 = ~n5633 & n47432 ;
  assign n47434 = n26599 & n47433 ;
  assign n47435 = n47434 ^ n36955 ^ n35719 ;
  assign n47436 = n36753 ^ n32864 ^ 1'b0 ;
  assign n47437 = n26884 & ~n47436 ;
  assign n47438 = ~n47435 & n47437 ;
  assign n47439 = n5797 & ~n42950 ;
  assign n47440 = n47439 ^ n36385 ^ 1'b0 ;
  assign n47441 = n7657 | n31172 ;
  assign n47442 = ( n15378 & n23575 ) | ( n15378 & ~n27200 ) | ( n23575 & ~n27200 ) ;
  assign n47443 = n31393 | n47442 ;
  assign n47444 = n47441 | n47443 ;
  assign n47445 = ( ~n10717 & n15378 ) | ( ~n10717 & n35945 ) | ( n15378 & n35945 ) ;
  assign n47446 = ( n3840 & ~n6354 ) | ( n3840 & n11277 ) | ( ~n6354 & n11277 ) ;
  assign n47447 = n21298 & ~n27363 ;
  assign n47448 = n3331 & n27489 ;
  assign n47449 = ( n12538 & n31918 ) | ( n12538 & ~n40489 ) | ( n31918 & ~n40489 ) ;
  assign n47450 = n4995 | n39292 ;
  assign n47451 = n47450 ^ n40154 ^ 1'b0 ;
  assign n47453 = n36368 ^ n7042 ^ 1'b0 ;
  assign n47454 = ~n652 & n47453 ;
  assign n47452 = n2495 | n14057 ;
  assign n47455 = n47454 ^ n47452 ^ 1'b0 ;
  assign n47456 = ~n10758 & n14050 ;
  assign n47457 = n34519 & n47456 ;
  assign n47458 = n47457 ^ n13469 ^ 1'b0 ;
  assign n47459 = n5655 | n47458 ;
  assign n47460 = n16168 ^ n9909 ^ 1'b0 ;
  assign n47461 = n11314 & ~n47460 ;
  assign n47462 = n47461 ^ n14319 ^ n13020 ;
  assign n47463 = n47462 ^ n7356 ^ 1'b0 ;
  assign n47464 = n13885 & ~n47463 ;
  assign n47465 = ( n1905 & ~n23274 ) | ( n1905 & n47464 ) | ( ~n23274 & n47464 ) ;
  assign n47466 = ( n9730 & n26461 ) | ( n9730 & n44828 ) | ( n26461 & n44828 ) ;
  assign n47469 = n11696 | n22778 ;
  assign n47470 = n47469 ^ n9742 ^ 1'b0 ;
  assign n47467 = n911 | n20807 ;
  assign n47468 = n1894 | n47467 ;
  assign n47471 = n47470 ^ n47468 ^ n36666 ;
  assign n47472 = ( ~n2137 & n13360 ) | ( ~n2137 & n47471 ) | ( n13360 & n47471 ) ;
  assign n47473 = ( n12756 & n28766 ) | ( n12756 & n37348 ) | ( n28766 & n37348 ) ;
  assign n47475 = n39025 ^ n25581 ^ n18359 ;
  assign n47476 = n8438 & n47475 ;
  assign n47474 = ( n14543 & ~n22311 ) | ( n14543 & n41282 ) | ( ~n22311 & n41282 ) ;
  assign n47477 = n47476 ^ n47474 ^ n18828 ;
  assign n47478 = ~n14768 & n35228 ;
  assign n47479 = n47478 ^ n7146 ^ 1'b0 ;
  assign n47480 = ~n5467 & n8894 ;
  assign n47481 = n11777 ^ n10835 ^ n5197 ;
  assign n47482 = ( ~n14674 & n15278 ) | ( ~n14674 & n27171 ) | ( n15278 & n27171 ) ;
  assign n47483 = ~n22041 & n47344 ;
  assign n47484 = n35550 ^ n15504 ^ 1'b0 ;
  assign n47485 = n7912 ^ n5409 ^ 1'b0 ;
  assign n47487 = ( n4171 & n4337 ) | ( n4171 & ~n9028 ) | ( n4337 & ~n9028 ) ;
  assign n47488 = n7587 & n47487 ;
  assign n47489 = ~n6934 & n47488 ;
  assign n47486 = n15122 | n42711 ;
  assign n47490 = n47489 ^ n47486 ^ 1'b0 ;
  assign n47491 = ( n533 & n10533 ) | ( n533 & n22755 ) | ( n10533 & n22755 ) ;
  assign n47492 = x88 & n5160 ;
  assign n47493 = ( n23212 & n47491 ) | ( n23212 & ~n47492 ) | ( n47491 & ~n47492 ) ;
  assign n47494 = ( n14909 & n17263 ) | ( n14909 & ~n20649 ) | ( n17263 & ~n20649 ) ;
  assign n47495 = n47494 ^ n27473 ^ 1'b0 ;
  assign n47496 = n19033 ^ n1152 ^ x29 ;
  assign n47497 = n5305 | n32427 ;
  assign n47498 = n47497 ^ n31071 ^ 1'b0 ;
  assign n47499 = n34562 ^ n21238 ^ n5440 ;
  assign n47500 = n23797 ^ n20739 ^ 1'b0 ;
  assign n47501 = n6859 & ~n19027 ;
  assign n47502 = ~n47500 & n47501 ;
  assign n47503 = n12683 & ~n47502 ;
  assign n47504 = n27825 & n47503 ;
  assign n47505 = n47504 ^ n27790 ^ n1095 ;
  assign n47506 = n695 & ~n16936 ;
  assign n47507 = n12344 & n47506 ;
  assign n47508 = ( ~n1011 & n12931 ) | ( ~n1011 & n23492 ) | ( n12931 & n23492 ) ;
  assign n47509 = ~n8130 & n47508 ;
  assign n47510 = n47509 ^ n6986 ^ 1'b0 ;
  assign n47511 = n47507 | n47510 ;
  assign n47512 = n39555 | n41014 ;
  assign n47513 = n25548 ^ n17707 ^ n7832 ;
  assign n47514 = n12899 | n13372 ;
  assign n47515 = n6357 | n20302 ;
  assign n47516 = n8723 | n47515 ;
  assign n47517 = n8010 & n47516 ;
  assign n47521 = n4806 | n9732 ;
  assign n47518 = n22296 ^ n8643 ^ n8403 ;
  assign n47519 = n19568 | n47518 ;
  assign n47520 = n28308 | n47519 ;
  assign n47522 = n47521 ^ n47520 ^ x179 ;
  assign n47523 = n42823 ^ n18306 ^ n17330 ;
  assign n47524 = n47523 ^ n18961 ^ n12574 ;
  assign n47525 = ( n9380 & ~n37100 ) | ( n9380 & n47524 ) | ( ~n37100 & n47524 ) ;
  assign n47526 = ( n3005 & n28584 ) | ( n3005 & ~n43928 ) | ( n28584 & ~n43928 ) ;
  assign n47527 = ~n8987 & n20970 ;
  assign n47528 = n15535 & ~n25182 ;
  assign n47529 = n47528 ^ n24578 ^ 1'b0 ;
  assign n47530 = ~n13828 & n17949 ;
  assign n47531 = n18613 & n47530 ;
  assign n47532 = n47531 ^ n38664 ^ 1'b0 ;
  assign n47533 = n1014 & ~n3174 ;
  assign n47534 = n47533 ^ n30885 ^ 1'b0 ;
  assign n47535 = n12113 & ~n47534 ;
  assign n47536 = n5388 ^ n5227 ^ x214 ;
  assign n47537 = n47536 ^ n45121 ^ n40596 ;
  assign n47538 = ( n33287 & ~n42824 ) | ( n33287 & n47537 ) | ( ~n42824 & n47537 ) ;
  assign n47539 = n28716 ^ n25899 ^ 1'b0 ;
  assign n47540 = n5043 | n47539 ;
  assign n47541 = ( ~n11641 & n43248 ) | ( ~n11641 & n47540 ) | ( n43248 & n47540 ) ;
  assign n47542 = n4933 & ~n22276 ;
  assign n47543 = n47542 ^ n6582 ^ n1030 ;
  assign n47544 = n25027 ^ n13741 ^ 1'b0 ;
  assign n47545 = n16321 | n47544 ;
  assign n47552 = x133 & n4393 ;
  assign n47553 = n47552 ^ n14624 ^ 1'b0 ;
  assign n47554 = n47553 ^ n24734 ^ 1'b0 ;
  assign n47547 = n39787 ^ n23967 ^ 1'b0 ;
  assign n47548 = n25410 ^ n7203 ^ 1'b0 ;
  assign n47549 = ~n47547 & n47548 ;
  assign n47550 = ~n29736 & n47549 ;
  assign n47551 = n8193 & n47550 ;
  assign n47546 = n23403 & n46898 ;
  assign n47555 = n47554 ^ n47551 ^ n47546 ;
  assign n47556 = ~n9301 & n16903 ;
  assign n47557 = ~n15129 & n47556 ;
  assign n47558 = n9463 & ~n22100 ;
  assign n47561 = n34745 ^ n9746 ^ 1'b0 ;
  assign n47562 = n12311 & n47561 ;
  assign n47563 = n1279 & n47562 ;
  assign n47564 = ~n20516 & n47563 ;
  assign n47559 = ( ~x211 & n5039 ) | ( ~x211 & n8789 ) | ( n5039 & n8789 ) ;
  assign n47560 = ~n15514 & n47559 ;
  assign n47565 = n47564 ^ n47560 ^ 1'b0 ;
  assign n47566 = n33621 ^ n20846 ^ 1'b0 ;
  assign n47567 = n47566 ^ n37324 ^ n33011 ;
  assign n47569 = ( n8919 & n11458 ) | ( n8919 & n24559 ) | ( n11458 & n24559 ) ;
  assign n47568 = n7783 & n17457 ;
  assign n47570 = n47569 ^ n47568 ^ 1'b0 ;
  assign n47571 = n47570 ^ n24006 ^ 1'b0 ;
  assign n47572 = ~n15812 & n34053 ;
  assign n47573 = n8537 & n33901 ;
  assign n47574 = n34458 ^ n19495 ^ 1'b0 ;
  assign n47575 = n6099 & n47574 ;
  assign n47576 = ( n5162 & ~n26468 ) | ( n5162 & n47575 ) | ( ~n26468 & n47575 ) ;
  assign n47578 = n15838 ^ n10357 ^ n2163 ;
  assign n47579 = n47578 ^ n10540 ^ n7912 ;
  assign n47577 = ~n14367 & n22813 ;
  assign n47580 = n47579 ^ n47577 ^ 1'b0 ;
  assign n47581 = n13027 ^ n3918 ^ n311 ;
  assign n47582 = n10958 | n15849 ;
  assign n47583 = n47581 | n47582 ;
  assign n47584 = n29080 | n33610 ;
  assign n47585 = n1922 & n47584 ;
  assign n47586 = n47585 ^ n36489 ^ 1'b0 ;
  assign n47587 = n41468 ^ n25687 ^ 1'b0 ;
  assign n47588 = n11842 ^ n1929 ^ 1'b0 ;
  assign n47589 = n43859 | n47588 ;
  assign n47590 = ( n10191 & n42313 ) | ( n10191 & ~n47589 ) | ( n42313 & ~n47589 ) ;
  assign n47591 = n22595 ^ n20493 ^ n5375 ;
  assign n47592 = ( n25315 & n42429 ) | ( n25315 & n47591 ) | ( n42429 & n47591 ) ;
  assign n47594 = n31753 & ~n45371 ;
  assign n47595 = n16825 & n47594 ;
  assign n47593 = n39301 ^ n30268 ^ n29666 ;
  assign n47596 = n47595 ^ n47593 ^ n42118 ;
  assign n47597 = n19123 ^ n13077 ^ 1'b0 ;
  assign n47598 = n969 & ~n6582 ;
  assign n47599 = n23162 & n27899 ;
  assign n47600 = n2526 & n47599 ;
  assign n47601 = n992 & n3675 ;
  assign n47602 = n18308 & ~n28875 ;
  assign n47603 = n47602 ^ n37870 ^ 1'b0 ;
  assign n47604 = n47601 & n47603 ;
  assign n47605 = n29732 ^ n7401 ^ 1'b0 ;
  assign n47606 = n18330 & n47605 ;
  assign n47607 = n32163 ^ n16752 ^ n15246 ;
  assign n47608 = ( ~n3505 & n22662 ) | ( ~n3505 & n47607 ) | ( n22662 & n47607 ) ;
  assign n47609 = ( n3677 & ~n9288 ) | ( n3677 & n17193 ) | ( ~n9288 & n17193 ) ;
  assign n47610 = ( ~n17065 & n19442 ) | ( ~n17065 & n47609 ) | ( n19442 & n47609 ) ;
  assign n47611 = n8499 & ~n26674 ;
  assign n47612 = n47611 ^ n24300 ^ 1'b0 ;
  assign n47613 = ( ~n26101 & n26143 ) | ( ~n26101 & n30874 ) | ( n26143 & n30874 ) ;
  assign n47614 = ~n47612 & n47613 ;
  assign n47617 = n29688 ^ n12478 ^ 1'b0 ;
  assign n47615 = n43673 ^ n10221 ^ 1'b0 ;
  assign n47616 = ~n21000 & n47615 ;
  assign n47618 = n47617 ^ n47616 ^ n24516 ;
  assign n47619 = ( n17178 & n19323 ) | ( n17178 & n20031 ) | ( n19323 & n20031 ) ;
  assign n47620 = n1179 & n24036 ;
  assign n47621 = n15372 & n47620 ;
  assign n47622 = n15201 ^ n5649 ^ n1753 ;
  assign n47623 = ( n1313 & n35819 ) | ( n1313 & n47622 ) | ( n35819 & n47622 ) ;
  assign n47624 = ( n41591 & n47621 ) | ( n41591 & n47623 ) | ( n47621 & n47623 ) ;
  assign n47625 = x28 & n6750 ;
  assign n47626 = ~n6750 & n47625 ;
  assign n47627 = n15092 | n22876 ;
  assign n47628 = ( n21770 & n27522 ) | ( n21770 & n47627 ) | ( n27522 & n47627 ) ;
  assign n47629 = ( ~n10608 & n26367 ) | ( ~n10608 & n47628 ) | ( n26367 & n47628 ) ;
  assign n47630 = ( n44239 & n47626 ) | ( n44239 & ~n47629 ) | ( n47626 & ~n47629 ) ;
  assign n47631 = n39319 ^ n18555 ^ n9061 ;
  assign n47632 = ( n13173 & n15055 ) | ( n13173 & ~n38712 ) | ( n15055 & ~n38712 ) ;
  assign n47633 = n44962 ^ n35731 ^ n11107 ;
  assign n47634 = n10229 ^ n471 ^ 1'b0 ;
  assign n47635 = n13000 & n47634 ;
  assign n47636 = n47635 ^ n5318 ^ n1222 ;
  assign n47637 = n15352 | n47636 ;
  assign n47638 = n11727 ^ n4196 ^ 1'b0 ;
  assign n47639 = n3314 & n47638 ;
  assign n47640 = ( n21178 & n24413 ) | ( n21178 & n47639 ) | ( n24413 & n47639 ) ;
  assign n47641 = n31657 & n47640 ;
  assign n47642 = n47641 ^ n17733 ^ 1'b0 ;
  assign n47643 = n32608 ^ n327 ^ 1'b0 ;
  assign n47644 = n47642 | n47643 ;
  assign n47649 = n13917 ^ n6411 ^ 1'b0 ;
  assign n47650 = n39647 & ~n43469 ;
  assign n47651 = n47650 ^ n40884 ^ 1'b0 ;
  assign n47652 = n47649 & n47651 ;
  assign n47645 = ~n11288 & n26333 ;
  assign n47646 = ~n20027 & n47645 ;
  assign n47647 = n21672 | n47646 ;
  assign n47648 = n25609 | n47647 ;
  assign n47653 = n47652 ^ n47648 ^ n20143 ;
  assign n47654 = n21693 ^ n16922 ^ n15655 ;
  assign n47655 = n39566 ^ n31656 ^ 1'b0 ;
  assign n47658 = n14078 ^ n12768 ^ 1'b0 ;
  assign n47659 = n1489 | n47658 ;
  assign n47656 = n20108 ^ n4821 ^ 1'b0 ;
  assign n47657 = ~n13174 & n47656 ;
  assign n47660 = n47659 ^ n47657 ^ n13393 ;
  assign n47661 = ( ~n5705 & n10753 ) | ( ~n5705 & n15124 ) | ( n10753 & n15124 ) ;
  assign n47662 = n47661 ^ n26720 ^ 1'b0 ;
  assign n47663 = ( ~n23064 & n26562 ) | ( ~n23064 & n39653 ) | ( n26562 & n39653 ) ;
  assign n47664 = ( n13664 & n20711 ) | ( n13664 & n47663 ) | ( n20711 & n47663 ) ;
  assign n47665 = n31440 | n32898 ;
  assign n47666 = n4192 & ~n47665 ;
  assign n47667 = n12960 | n47666 ;
  assign n47668 = n3164 & n45433 ;
  assign n47669 = ( n4586 & ~n16121 ) | ( n4586 & n47668 ) | ( ~n16121 & n47668 ) ;
  assign n47670 = ~n1916 & n47669 ;
  assign n47671 = ( n7817 & n11544 ) | ( n7817 & ~n15821 ) | ( n11544 & ~n15821 ) ;
  assign n47672 = n47671 ^ n15824 ^ 1'b0 ;
  assign n47673 = n30479 ^ n11380 ^ n4349 ;
  assign n47674 = n8320 & ~n15027 ;
  assign n47675 = n47673 & n47674 ;
  assign n47676 = n1385 & n14416 ;
  assign n47677 = ( n10808 & n12169 ) | ( n10808 & n47676 ) | ( n12169 & n47676 ) ;
  assign n47678 = n40306 ^ n8017 ^ 1'b0 ;
  assign n47679 = ( n5707 & n16182 ) | ( n5707 & ~n16883 ) | ( n16182 & ~n16883 ) ;
  assign n47680 = ( n11633 & n42051 ) | ( n11633 & ~n47679 ) | ( n42051 & ~n47679 ) ;
  assign n47681 = n47680 ^ n23746 ^ n509 ;
  assign n47682 = n6004 ^ n3186 ^ n1866 ;
  assign n47683 = n34420 ^ n15642 ^ n1516 ;
  assign n47684 = ( n30045 & n47682 ) | ( n30045 & n47683 ) | ( n47682 & n47683 ) ;
  assign n47685 = n1172 & ~n6000 ;
  assign n47686 = n13038 & n47685 ;
  assign n47687 = n47686 ^ n34876 ^ n19634 ;
  assign n47688 = ( ~n3655 & n11686 ) | ( ~n3655 & n33793 ) | ( n11686 & n33793 ) ;
  assign n47689 = n47688 ^ n40025 ^ n35474 ;
  assign n47690 = n8305 & n31481 ;
  assign n47691 = n38425 ^ n26294 ^ 1'b0 ;
  assign n47692 = n7902 | n47691 ;
  assign n47693 = ~n15623 & n23793 ;
  assign n47694 = n12392 | n14956 ;
  assign n47695 = n47693 | n47694 ;
  assign n47696 = ( n5882 & ~n10673 ) | ( n5882 & n34837 ) | ( ~n10673 & n34837 ) ;
  assign n47697 = n31997 ^ n2834 ^ 1'b0 ;
  assign n47698 = n16659 & n47697 ;
  assign n47699 = ~n47696 & n47698 ;
  assign n47700 = n32570 ^ n27166 ^ n8139 ;
  assign n47701 = ( n1770 & n5375 ) | ( n1770 & ~n13994 ) | ( n5375 & ~n13994 ) ;
  assign n47702 = n24988 ^ n20042 ^ 1'b0 ;
  assign n47703 = n729 & ~n25530 ;
  assign n47704 = ( ~n47701 & n47702 ) | ( ~n47701 & n47703 ) | ( n47702 & n47703 ) ;
  assign n47707 = n12504 ^ n6164 ^ 1'b0 ;
  assign n47708 = n12297 & n47707 ;
  assign n47705 = n13736 & n22747 ;
  assign n47706 = ( ~n14919 & n31168 ) | ( ~n14919 & n47705 ) | ( n31168 & n47705 ) ;
  assign n47709 = n47708 ^ n47706 ^ 1'b0 ;
  assign n47710 = n41685 & ~n46316 ;
  assign n47711 = ~n16034 & n47710 ;
  assign n47712 = n9651 & n23978 ;
  assign n47713 = n47712 ^ n17289 ^ 1'b0 ;
  assign n47714 = n14130 & n21722 ;
  assign n47715 = n47714 ^ n14748 ^ 1'b0 ;
  assign n47716 = n32949 ^ n11413 ^ 1'b0 ;
  assign n47717 = n32435 & n47716 ;
  assign n47718 = n25014 ^ n1851 ^ 1'b0 ;
  assign n47719 = n47718 ^ n22593 ^ n5975 ;
  assign n47720 = n4932 & n16525 ;
  assign n47721 = ~n17396 & n47720 ;
  assign n47722 = ( n21161 & ~n26468 ) | ( n21161 & n47721 ) | ( ~n26468 & n47721 ) ;
  assign n47723 = ( n7911 & n15056 ) | ( n7911 & ~n29530 ) | ( n15056 & ~n29530 ) ;
  assign n47724 = ( n2924 & ~n3230 ) | ( n2924 & n20585 ) | ( ~n3230 & n20585 ) ;
  assign n47725 = ( n19323 & n31998 ) | ( n19323 & ~n47724 ) | ( n31998 & ~n47724 ) ;
  assign n47726 = n38859 ^ n28106 ^ n7473 ;
  assign n47728 = ( n25348 & n30088 ) | ( n25348 & ~n34892 ) | ( n30088 & ~n34892 ) ;
  assign n47727 = n17271 ^ n14607 ^ 1'b0 ;
  assign n47729 = n47728 ^ n47727 ^ n33140 ;
  assign n47730 = ~n7880 & n8111 ;
  assign n47731 = n47730 ^ n47617 ^ 1'b0 ;
  assign n47732 = n20909 & ~n47731 ;
  assign n47733 = n47732 ^ n39609 ^ n27953 ;
  assign n47734 = ( n7817 & n18193 ) | ( n7817 & n38723 ) | ( n18193 & n38723 ) ;
  assign n47735 = n8928 & n47734 ;
  assign n47736 = ~n47733 & n47735 ;
  assign n47737 = n40202 ^ n17515 ^ n7042 ;
  assign n47738 = n47737 ^ x45 ^ 1'b0 ;
  assign n47739 = n29077 & n47738 ;
  assign n47740 = n23170 ^ n11769 ^ 1'b0 ;
  assign n47741 = ~n22302 & n33813 ;
  assign n47742 = n47741 ^ n31525 ^ 1'b0 ;
  assign n47743 = n24505 ^ n12908 ^ n5906 ;
  assign n47744 = n9713 ^ n6868 ^ n5132 ;
  assign n47745 = n7847 | n9208 ;
  assign n47746 = n47745 ^ n40978 ^ 1'b0 ;
  assign n47747 = n47744 | n47746 ;
  assign n47748 = ( n9213 & ~n47743 ) | ( n9213 & n47747 ) | ( ~n47743 & n47747 ) ;
  assign n47749 = ( n4414 & ~n22807 ) | ( n4414 & n47748 ) | ( ~n22807 & n47748 ) ;
  assign n47751 = ~n17051 & n18505 ;
  assign n47752 = n47751 ^ n15039 ^ 1'b0 ;
  assign n47750 = n32898 ^ n10972 ^ n1044 ;
  assign n47753 = n47752 ^ n47750 ^ n16730 ;
  assign n47754 = ( n8353 & n17755 ) | ( n8353 & n45687 ) | ( n17755 & n45687 ) ;
  assign n47755 = n47754 ^ n16113 ^ n6119 ;
  assign n47756 = n977 & ~n2327 ;
  assign n47757 = ( ~n9713 & n43389 ) | ( ~n9713 & n47756 ) | ( n43389 & n47756 ) ;
  assign n47758 = ( n8755 & n23869 ) | ( n8755 & n34335 ) | ( n23869 & n34335 ) ;
  assign n47760 = ( n3232 & n17054 ) | ( n3232 & n40090 ) | ( n17054 & n40090 ) ;
  assign n47761 = ( ~n9965 & n12512 ) | ( ~n9965 & n42280 ) | ( n12512 & n42280 ) ;
  assign n47762 = ( n24566 & n47760 ) | ( n24566 & n47761 ) | ( n47760 & n47761 ) ;
  assign n47759 = n4759 | n5548 ;
  assign n47763 = n47762 ^ n47759 ^ 1'b0 ;
  assign n47764 = n45541 ^ n3959 ^ 1'b0 ;
  assign n47770 = ( n6083 & n11373 ) | ( n6083 & n23183 ) | ( n11373 & n23183 ) ;
  assign n47768 = ~n13051 & n25495 ;
  assign n47769 = n31790 & n47768 ;
  assign n47765 = n17787 ^ n13351 ^ n2798 ;
  assign n47766 = n13554 ^ n1183 ^ 1'b0 ;
  assign n47767 = n47765 | n47766 ;
  assign n47771 = n47770 ^ n47769 ^ n47767 ;
  assign n47772 = n20787 | n41350 ;
  assign n47773 = n47771 | n47772 ;
  assign n47775 = n5480 ^ n3129 ^ 1'b0 ;
  assign n47774 = ~n8090 & n36744 ;
  assign n47776 = n47775 ^ n47774 ^ 1'b0 ;
  assign n47777 = ( ~n36815 & n39266 ) | ( ~n36815 & n47776 ) | ( n39266 & n47776 ) ;
  assign n47778 = n47777 ^ n20221 ^ 1'b0 ;
  assign n47779 = n20728 ^ n19801 ^ x156 ;
  assign n47780 = n47779 ^ n43234 ^ 1'b0 ;
  assign n47781 = n45494 ^ n33854 ^ n8784 ;
  assign n47782 = ( ~n5855 & n26339 ) | ( ~n5855 & n47781 ) | ( n26339 & n47781 ) ;
  assign n47783 = ( n21240 & n38162 ) | ( n21240 & n42679 ) | ( n38162 & n42679 ) ;
  assign n47784 = ~n6885 & n24671 ;
  assign n47785 = ~n9349 & n47784 ;
  assign n47786 = n20295 ^ n9788 ^ 1'b0 ;
  assign n47787 = n15550 & ~n47786 ;
  assign n47788 = n47787 ^ n25462 ^ 1'b0 ;
  assign n47789 = n41250 ^ n14057 ^ n912 ;
  assign n47790 = n10975 & n47789 ;
  assign n47791 = n47790 ^ n4439 ^ 1'b0 ;
  assign n47794 = n14902 ^ n13109 ^ 1'b0 ;
  assign n47795 = n9468 & ~n19208 ;
  assign n47796 = n47794 & n47795 ;
  assign n47797 = n47796 ^ n2106 ^ 1'b0 ;
  assign n47798 = ~n37363 & n47797 ;
  assign n47792 = n2130 | n11459 ;
  assign n47793 = n47792 ^ n30982 ^ 1'b0 ;
  assign n47799 = n47798 ^ n47793 ^ 1'b0 ;
  assign n47800 = ~n32281 & n47799 ;
  assign n47801 = n25879 ^ n25427 ^ 1'b0 ;
  assign n47802 = n46991 | n47801 ;
  assign n47803 = n43660 ^ n26349 ^ n24683 ;
  assign n47808 = n8036 & n29720 ;
  assign n47809 = n47808 ^ n21525 ^ 1'b0 ;
  assign n47804 = ~n4807 & n10327 ;
  assign n47805 = ~n1073 & n47804 ;
  assign n47806 = n47805 ^ n24384 ^ n5145 ;
  assign n47807 = ( n27587 & n32374 ) | ( n27587 & ~n47806 ) | ( n32374 & ~n47806 ) ;
  assign n47810 = n47809 ^ n47807 ^ n3187 ;
  assign n47811 = n6124 ^ n1941 ^ 1'b0 ;
  assign n47812 = n39093 & n47811 ;
  assign n47813 = ( n10214 & n19569 ) | ( n10214 & n38611 ) | ( n19569 & n38611 ) ;
  assign n47814 = n35635 ^ n21649 ^ n7177 ;
  assign n47815 = ( ~n9077 & n44417 ) | ( ~n9077 & n47814 ) | ( n44417 & n47814 ) ;
  assign n47816 = n15311 | n47815 ;
  assign n47817 = n47816 ^ n13988 ^ 1'b0 ;
  assign n47818 = n26262 ^ n19104 ^ 1'b0 ;
  assign n47819 = ~n43056 & n47818 ;
  assign n47820 = n14305 & n38691 ;
  assign n47821 = ~n17510 & n47820 ;
  assign n47822 = n35596 ^ n33218 ^ n5236 ;
  assign n47823 = ( n22532 & n25134 ) | ( n22532 & ~n47822 ) | ( n25134 & ~n47822 ) ;
  assign n47824 = n37192 ^ n33049 ^ n14673 ;
  assign n47825 = ( n2760 & n6178 ) | ( n2760 & ~n47824 ) | ( n6178 & ~n47824 ) ;
  assign n47826 = ~n4374 & n11448 ;
  assign n47827 = n47826 ^ n40061 ^ 1'b0 ;
  assign n47828 = n47827 ^ n23633 ^ 1'b0 ;
  assign n47829 = ( n9271 & n26447 ) | ( n9271 & ~n33937 ) | ( n26447 & ~n33937 ) ;
  assign n47830 = n46630 ^ n2478 ^ 1'b0 ;
  assign n47831 = n24341 & ~n47830 ;
  assign n47832 = ( ~n3798 & n43928 ) | ( ~n3798 & n47831 ) | ( n43928 & n47831 ) ;
  assign n47833 = n10599 ^ n9280 ^ n4755 ;
  assign n47834 = ( n10553 & n26183 ) | ( n10553 & n47833 ) | ( n26183 & n47833 ) ;
  assign n47835 = n32758 ^ n10802 ^ n3603 ;
  assign n47836 = n47835 ^ n5518 ^ 1'b0 ;
  assign n47837 = ~n47834 & n47836 ;
  assign n47838 = n7261 | n10214 ;
  assign n47839 = n47838 ^ n38374 ^ 1'b0 ;
  assign n47840 = ( n27465 & n31857 ) | ( n27465 & ~n47839 ) | ( n31857 & ~n47839 ) ;
  assign n47841 = ~n10989 & n47840 ;
  assign n47842 = n47841 ^ n9219 ^ 1'b0 ;
  assign n47843 = n36496 ^ n22321 ^ n9569 ;
  assign n47844 = n21001 ^ n13539 ^ 1'b0 ;
  assign n47845 = n47843 | n47844 ;
  assign n47846 = ( ~n7351 & n13317 ) | ( ~n7351 & n21578 ) | ( n13317 & n21578 ) ;
  assign n47847 = n47846 ^ n22093 ^ n20152 ;
  assign n47848 = ( n1823 & ~n19052 ) | ( n1823 & n24579 ) | ( ~n19052 & n24579 ) ;
  assign n47849 = ( n12761 & n14901 ) | ( n12761 & ~n18505 ) | ( n14901 & ~n18505 ) ;
  assign n47850 = n47849 ^ n9206 ^ n6557 ;
  assign n47851 = ( n3837 & n8816 ) | ( n3837 & ~n47850 ) | ( n8816 & ~n47850 ) ;
  assign n47852 = ~n24112 & n47851 ;
  assign n47853 = ( ~n9042 & n16811 ) | ( ~n9042 & n20339 ) | ( n16811 & n20339 ) ;
  assign n47854 = ( n9314 & n18456 ) | ( n9314 & n47853 ) | ( n18456 & n47853 ) ;
  assign n47855 = n28093 ^ n21470 ^ n7141 ;
  assign n47856 = n20553 ^ n19875 ^ n10920 ;
  assign n47857 = n25197 & ~n35070 ;
  assign n47858 = ~n32526 & n47857 ;
  assign n47859 = n1474 | n47858 ;
  assign n47860 = n47859 ^ n14466 ^ 1'b0 ;
  assign n47861 = ( n18463 & n20679 ) | ( n18463 & n22911 ) | ( n20679 & n22911 ) ;
  assign n47862 = n47861 ^ n2394 ^ 1'b0 ;
  assign n47863 = n27334 | n43906 ;
  assign n47864 = n35070 & ~n47863 ;
  assign n47866 = ( n5050 & n9329 ) | ( n5050 & ~n18088 ) | ( n9329 & ~n18088 ) ;
  assign n47865 = n27214 ^ n8998 ^ 1'b0 ;
  assign n47867 = n47866 ^ n47865 ^ n2819 ;
  assign n47868 = ( n8751 & ~n9288 ) | ( n8751 & n15719 ) | ( ~n9288 & n15719 ) ;
  assign n47869 = n47868 ^ n47442 ^ 1'b0 ;
  assign n47870 = ( n26730 & n37913 ) | ( n26730 & ~n47869 ) | ( n37913 & ~n47869 ) ;
  assign n47871 = n7984 ^ n2071 ^ 1'b0 ;
  assign n47872 = n17211 ^ n4403 ^ n1567 ;
  assign n47873 = ~n7472 & n23032 ;
  assign n47874 = n47873 ^ n29629 ^ 1'b0 ;
  assign n47875 = ~n7705 & n10945 ;
  assign n47876 = ( ~n4925 & n8003 ) | ( ~n4925 & n47875 ) | ( n8003 & n47875 ) ;
  assign n47877 = ( ~n47872 & n47874 ) | ( ~n47872 & n47876 ) | ( n47874 & n47876 ) ;
  assign n47878 = ( n4083 & n20332 ) | ( n4083 & ~n26157 ) | ( n20332 & ~n26157 ) ;
  assign n47879 = ( n7351 & n12181 ) | ( n7351 & n47878 ) | ( n12181 & n47878 ) ;
  assign n47880 = ( n13504 & ~n33534 ) | ( n13504 & n47879 ) | ( ~n33534 & n47879 ) ;
  assign n47881 = n6457 | n47880 ;
  assign n47883 = n8431 & n9050 ;
  assign n47882 = n45863 ^ n25944 ^ n6659 ;
  assign n47884 = n47883 ^ n47882 ^ n6938 ;
  assign n47885 = ( n12641 & n15950 ) | ( n12641 & ~n29004 ) | ( n15950 & ~n29004 ) ;
  assign n47886 = n35908 ^ n13886 ^ 1'b0 ;
  assign n47887 = n47885 & ~n47886 ;
  assign n47888 = n43633 ^ n26253 ^ 1'b0 ;
  assign n47889 = n6937 | n30700 ;
  assign n47890 = n42872 ^ n19477 ^ n5548 ;
  assign n47891 = n47890 ^ n43158 ^ 1'b0 ;
  assign n47892 = ( n16515 & n22353 ) | ( n16515 & n39028 ) | ( n22353 & n39028 ) ;
  assign n47893 = ~n18386 & n22545 ;
  assign n47894 = ~n6484 & n47893 ;
  assign n47895 = ( n2485 & n13356 ) | ( n2485 & ~n47894 ) | ( n13356 & ~n47894 ) ;
  assign n47896 = n34074 ^ n25574 ^ n14175 ;
  assign n47897 = n3803 | n11650 ;
  assign n47898 = n47897 ^ n27237 ^ 1'b0 ;
  assign n47899 = n12040 ^ n1544 ^ 1'b0 ;
  assign n47900 = ~n5581 & n47899 ;
  assign n47901 = n2629 & n47900 ;
  assign n47902 = n1448 & n11413 ;
  assign n47903 = x44 | n2027 ;
  assign n47904 = ( n17114 & ~n19748 ) | ( n17114 & n47903 ) | ( ~n19748 & n47903 ) ;
  assign n47905 = n10048 & n42625 ;
  assign n47906 = n14507 & n47905 ;
  assign n47907 = n17185 | n47906 ;
  assign n47908 = ( n12370 & n15470 ) | ( n12370 & ~n47103 ) | ( n15470 & ~n47103 ) ;
  assign n47909 = n28617 ^ n22807 ^ x200 ;
  assign n47910 = n14117 & n46666 ;
  assign n47914 = ( n2924 & n5828 ) | ( n2924 & n13509 ) | ( n5828 & n13509 ) ;
  assign n47911 = n4544 & ~n13245 ;
  assign n47912 = n16830 & n47911 ;
  assign n47913 = n7418 & ~n47912 ;
  assign n47915 = n47914 ^ n47913 ^ 1'b0 ;
  assign n47916 = ( ~n43201 & n44967 ) | ( ~n43201 & n47915 ) | ( n44967 & n47915 ) ;
  assign n47917 = n15877 & n16079 ;
  assign n47918 = n47917 ^ n28775 ^ 1'b0 ;
  assign n47919 = n4053 ^ n1192 ^ 1'b0 ;
  assign n47920 = n6291 & n47919 ;
  assign n47921 = n36381 ^ n11166 ^ n5393 ;
  assign n47922 = ~n42531 & n47921 ;
  assign n47923 = n14491 ^ n962 ^ 1'b0 ;
  assign n47924 = n47922 & ~n47923 ;
  assign n47925 = n47920 & ~n47924 ;
  assign n47926 = n14279 ^ n7973 ^ 1'b0 ;
  assign n47928 = ( n20215 & n21195 ) | ( n20215 & n24566 ) | ( n21195 & n24566 ) ;
  assign n47927 = n20325 & ~n21234 ;
  assign n47929 = n47928 ^ n47927 ^ 1'b0 ;
  assign n47934 = n4141 | n6877 ;
  assign n47935 = n47934 ^ n31382 ^ 1'b0 ;
  assign n47930 = n32546 ^ n32155 ^ 1'b0 ;
  assign n47931 = ~n28896 & n47930 ;
  assign n47932 = ( n3847 & ~n34605 ) | ( n3847 & n47931 ) | ( ~n34605 & n47931 ) ;
  assign n47933 = ~n14788 & n47932 ;
  assign n47936 = n47935 ^ n47933 ^ 1'b0 ;
  assign n47937 = n1892 ^ n1732 ^ 1'b0 ;
  assign n47938 = ( n10917 & ~n12510 ) | ( n10917 & n47937 ) | ( ~n12510 & n47937 ) ;
  assign n47939 = n47938 ^ n34553 ^ 1'b0 ;
  assign n47940 = n9092 ^ n2814 ^ 1'b0 ;
  assign n47941 = ~n7308 & n47940 ;
  assign n47942 = ( ~n19068 & n19328 ) | ( ~n19068 & n47941 ) | ( n19328 & n47941 ) ;
  assign n47943 = ~n1966 & n4445 ;
  assign n47944 = ( n3119 & n41782 ) | ( n3119 & n47943 ) | ( n41782 & n47943 ) ;
  assign n47945 = ~n24816 & n47944 ;
  assign n47946 = ( ~n1068 & n5202 ) | ( ~n1068 & n7942 ) | ( n5202 & n7942 ) ;
  assign n47947 = ( n750 & n38365 ) | ( n750 & n47946 ) | ( n38365 & n47946 ) ;
  assign n47948 = n28960 ^ n2353 ^ n2233 ;
  assign n47949 = n38597 & n41314 ;
  assign n47950 = ~n17129 & n47949 ;
  assign n47951 = n2146 | n42026 ;
  assign n47952 = n42044 ^ n9475 ^ n5281 ;
  assign n47953 = n47952 ^ n44112 ^ n16202 ;
  assign n47957 = n541 | n1934 ;
  assign n47958 = n1934 & ~n47957 ;
  assign n47959 = x161 & ~n47958 ;
  assign n47960 = n47958 & n47959 ;
  assign n47954 = n2441 | n14805 ;
  assign n47955 = n2441 & ~n47954 ;
  assign n47956 = n47955 ^ n30634 ^ n10015 ;
  assign n47961 = n47960 ^ n47956 ^ n37090 ;
  assign n47962 = n35134 ^ n5285 ^ 1'b0 ;
  assign n47963 = ~n12591 & n33442 ;
  assign n47964 = ~n29928 & n47963 ;
  assign n47965 = ( n47961 & ~n47962 ) | ( n47961 & n47964 ) | ( ~n47962 & n47964 ) ;
  assign n47966 = ( n662 & n3303 ) | ( n662 & ~n6490 ) | ( n3303 & ~n6490 ) ;
  assign n47967 = ( n3373 & n10022 ) | ( n3373 & n47966 ) | ( n10022 & n47966 ) ;
  assign n47968 = n47967 ^ n45671 ^ n28238 ;
  assign n47969 = n6810 & n25369 ;
  assign n47970 = ~n6956 & n9396 ;
  assign n47971 = ~n27323 & n27548 ;
  assign n47972 = n47971 ^ n719 ^ 1'b0 ;
  assign n47973 = n20109 | n47972 ;
  assign n47974 = n38146 & ~n47973 ;
  assign n47975 = n15918 ^ n5965 ^ n3377 ;
  assign n47976 = ( ~n18708 & n33092 ) | ( ~n18708 & n47975 ) | ( n33092 & n47975 ) ;
  assign n47977 = n47976 ^ n37561 ^ 1'b0 ;
  assign n47978 = n32546 | n47977 ;
  assign n47979 = ( n7133 & n42102 ) | ( n7133 & n47978 ) | ( n42102 & n47978 ) ;
  assign n47980 = n47979 ^ n26455 ^ 1'b0 ;
  assign n47981 = n23472 & ~n47980 ;
  assign n47982 = n17654 | n22353 ;
  assign n47983 = n47982 ^ n17294 ^ 1'b0 ;
  assign n47984 = n25212 & ~n31594 ;
  assign n47985 = n23858 ^ n2103 ^ 1'b0 ;
  assign n47986 = n45488 ^ n18123 ^ 1'b0 ;
  assign n47987 = n17909 ^ n14254 ^ 1'b0 ;
  assign n47988 = ~n10989 & n47987 ;
  assign n47989 = ( n8736 & ~n21290 ) | ( n8736 & n43126 ) | ( ~n21290 & n43126 ) ;
  assign n47990 = n40686 ^ n27539 ^ 1'b0 ;
  assign n47991 = ( n6702 & ~n21303 ) | ( n6702 & n24834 ) | ( ~n21303 & n24834 ) ;
  assign n47992 = n36836 ^ n35348 ^ n6540 ;
  assign n47993 = ( n11341 & n26443 ) | ( n11341 & ~n44800 ) | ( n26443 & ~n44800 ) ;
  assign n47994 = ( ~n30693 & n32538 ) | ( ~n30693 & n32946 ) | ( n32538 & n32946 ) ;
  assign n47995 = n18504 ^ n9576 ^ 1'b0 ;
  assign n47996 = n7320 | n36061 ;
  assign n47997 = n47996 ^ n19200 ^ 1'b0 ;
  assign n47998 = n35701 ^ n511 ^ 1'b0 ;
  assign n47999 = ( ~n7663 & n9963 ) | ( ~n7663 & n12066 ) | ( n9963 & n12066 ) ;
  assign n48000 = n47375 ^ n40013 ^ n12110 ;
  assign n48001 = n24611 ^ n21465 ^ 1'b0 ;
  assign n48002 = n12370 & ~n48001 ;
  assign n48003 = n48002 ^ n7655 ^ n6966 ;
  assign n48004 = n44505 ^ n41925 ^ 1'b0 ;
  assign n48005 = n7110 & ~n48004 ;
  assign n48006 = n43061 ^ n3157 ^ 1'b0 ;
  assign n48008 = n13671 ^ n11616 ^ 1'b0 ;
  assign n48009 = n3324 & n48008 ;
  assign n48007 = n4857 & ~n6517 ;
  assign n48010 = n48009 ^ n48007 ^ 1'b0 ;
  assign n48011 = n16958 | n19957 ;
  assign n48012 = n9821 | n48011 ;
  assign n48013 = n384 | n16961 ;
  assign n48014 = n29289 | n48013 ;
  assign n48015 = ( n12534 & ~n21914 ) | ( n12534 & n43038 ) | ( ~n21914 & n43038 ) ;
  assign n48016 = n16226 ^ n14008 ^ 1'b0 ;
  assign n48017 = n15136 | n48016 ;
  assign n48018 = ( n347 & n16894 ) | ( n347 & ~n48017 ) | ( n16894 & ~n48017 ) ;
  assign n48019 = n4076 | n44307 ;
  assign n48020 = n23678 ^ n4014 ^ 1'b0 ;
  assign n48021 = n29306 ^ n19519 ^ 1'b0 ;
  assign n48022 = n8589 & ~n16699 ;
  assign n48023 = ~n2884 & n48022 ;
  assign n48024 = n16610 & ~n48023 ;
  assign n48025 = n7719 & n48024 ;
  assign n48026 = n43209 ^ n7186 ^ n2998 ;
  assign n48028 = ( n20687 & n32911 ) | ( n20687 & n36107 ) | ( n32911 & n36107 ) ;
  assign n48027 = ( n6844 & n22755 ) | ( n6844 & n31071 ) | ( n22755 & n31071 ) ;
  assign n48029 = n48028 ^ n48027 ^ n32728 ;
  assign n48030 = n48029 ^ n25224 ^ n20366 ;
  assign n48031 = n14620 | n38896 ;
  assign n48032 = n24735 ^ n14611 ^ 1'b0 ;
  assign n48033 = n19474 | n48032 ;
  assign n48034 = ( n9580 & n12030 ) | ( n9580 & ~n48033 ) | ( n12030 & ~n48033 ) ;
  assign n48035 = n37692 ^ n11634 ^ n9513 ;
  assign n48036 = n34874 ^ n8308 ^ 1'b0 ;
  assign n48037 = n48035 & n48036 ;
  assign n48038 = n18932 ^ n10406 ^ 1'b0 ;
  assign n48039 = n1362 | n48038 ;
  assign n48040 = n273 | n23046 ;
  assign n48041 = n12147 & ~n48040 ;
  assign n48042 = n48041 ^ n10415 ^ n1461 ;
  assign n48043 = n35552 ^ n10584 ^ 1'b0 ;
  assign n48044 = x181 & n13479 ;
  assign n48045 = ( x149 & ~n13204 ) | ( x149 & n48044 ) | ( ~n13204 & n48044 ) ;
  assign n48049 = n16078 ^ n6135 ^ 1'b0 ;
  assign n48050 = ~n18987 & n48049 ;
  assign n48046 = n39065 ^ n21579 ^ 1'b0 ;
  assign n48047 = n5788 | n48046 ;
  assign n48048 = n29032 & ~n48047 ;
  assign n48051 = n48050 ^ n48048 ^ 1'b0 ;
  assign n48052 = n40489 ^ n22704 ^ n13212 ;
  assign n48053 = n13366 & ~n48052 ;
  assign n48054 = n48053 ^ n26212 ^ 1'b0 ;
  assign n48055 = n40828 ^ n17086 ^ 1'b0 ;
  assign n48056 = n45684 ^ n37957 ^ 1'b0 ;
  assign n48058 = n47914 ^ n14337 ^ n2780 ;
  assign n48059 = n48058 ^ n21531 ^ n5003 ;
  assign n48057 = ~n1839 & n16075 ;
  assign n48060 = n48059 ^ n48057 ^ 1'b0 ;
  assign n48061 = ( ~n14659 & n35970 ) | ( ~n14659 & n48060 ) | ( n35970 & n48060 ) ;
  assign n48062 = n7341 ^ n4315 ^ 1'b0 ;
  assign n48063 = n17386 & n48062 ;
  assign n48064 = ( n10676 & n18916 ) | ( n10676 & ~n25561 ) | ( n18916 & ~n25561 ) ;
  assign n48065 = ( n37937 & n46589 ) | ( n37937 & ~n48064 ) | ( n46589 & ~n48064 ) ;
  assign n48066 = ( ~n14032 & n21037 ) | ( ~n14032 & n48065 ) | ( n21037 & n48065 ) ;
  assign n48067 = n3333 | n8861 ;
  assign n48068 = ~n1249 & n9909 ;
  assign n48069 = n48068 ^ n15910 ^ 1'b0 ;
  assign n48070 = n6028 & n41357 ;
  assign n48071 = n48069 & n48070 ;
  assign n48072 = ~n21268 & n44206 ;
  assign n48073 = n48072 ^ n16634 ^ 1'b0 ;
  assign n48074 = ~n48071 & n48073 ;
  assign n48075 = n11880 | n12962 ;
  assign n48076 = n48075 ^ n31222 ^ 1'b0 ;
  assign n48077 = n21456 & ~n41374 ;
  assign n48078 = ~n23010 & n38005 ;
  assign n48079 = n2899 & n48078 ;
  assign n48080 = n26834 & ~n34266 ;
  assign n48081 = n13847 & ~n40970 ;
  assign n48082 = n27486 ^ n2215 ^ 1'b0 ;
  assign n48083 = ~n12350 & n48082 ;
  assign n48085 = ~n3480 & n11298 ;
  assign n48086 = n9100 & n48085 ;
  assign n48087 = n22259 | n48086 ;
  assign n48088 = n48087 ^ n15887 ^ 1'b0 ;
  assign n48084 = n27266 & ~n38677 ;
  assign n48089 = n48088 ^ n48084 ^ 1'b0 ;
  assign n48090 = ( n33177 & n48083 ) | ( n33177 & ~n48089 ) | ( n48083 & ~n48089 ) ;
  assign n48091 = x30 & n8946 ;
  assign n48092 = n48091 ^ n38292 ^ 1'b0 ;
  assign n48095 = ~n6165 & n7134 ;
  assign n48096 = n48095 ^ n5133 ^ 1'b0 ;
  assign n48097 = n43240 & ~n48096 ;
  assign n48093 = n32609 ^ n10786 ^ 1'b0 ;
  assign n48094 = ~n7610 & n48093 ;
  assign n48098 = n48097 ^ n48094 ^ 1'b0 ;
  assign n48099 = n48098 ^ n14591 ^ n12889 ;
  assign n48100 = n45270 ^ n23498 ^ n12623 ;
  assign n48101 = n36293 ^ n405 ^ 1'b0 ;
  assign n48102 = ( n37540 & ~n48100 ) | ( n37540 & n48101 ) | ( ~n48100 & n48101 ) ;
  assign n48103 = n36236 ^ n34330 ^ n18328 ;
  assign n48104 = n48103 ^ n18807 ^ 1'b0 ;
  assign n48105 = ~n11868 & n42619 ;
  assign n48106 = n48105 ^ n22773 ^ 1'b0 ;
  assign n48112 = ~n19915 & n44527 ;
  assign n48107 = n28450 ^ n21143 ^ 1'b0 ;
  assign n48108 = n48107 ^ n14626 ^ n2880 ;
  assign n48109 = ~n13250 & n48108 ;
  assign n48110 = n48109 ^ n37953 ^ n11426 ;
  assign n48111 = ~n2234 & n48110 ;
  assign n48113 = n48112 ^ n48111 ^ 1'b0 ;
  assign n48115 = ( n1192 & ~n12131 ) | ( n1192 & n24955 ) | ( ~n12131 & n24955 ) ;
  assign n48114 = n36517 & ~n45999 ;
  assign n48116 = n48115 ^ n48114 ^ 1'b0 ;
  assign n48118 = ( n10755 & n11209 ) | ( n10755 & n44356 ) | ( n11209 & n44356 ) ;
  assign n48117 = ~n4315 & n19916 ;
  assign n48119 = n48118 ^ n48117 ^ 1'b0 ;
  assign n48120 = ( n1937 & ~n8581 ) | ( n1937 & n36317 ) | ( ~n8581 & n36317 ) ;
  assign n48121 = n48120 ^ n31153 ^ n16858 ;
  assign n48122 = n16334 & n46193 ;
  assign n48123 = ( n4034 & ~n18875 ) | ( n4034 & n34387 ) | ( ~n18875 & n34387 ) ;
  assign n48124 = ( n4460 & ~n16903 ) | ( n4460 & n46129 ) | ( ~n16903 & n46129 ) ;
  assign n48125 = n3666 | n37430 ;
  assign n48126 = n31222 & ~n48125 ;
  assign n48127 = ( n353 & n39855 ) | ( n353 & ~n48126 ) | ( n39855 & ~n48126 ) ;
  assign n48128 = ( ~n18992 & n19067 ) | ( ~n18992 & n24914 ) | ( n19067 & n24914 ) ;
  assign n48129 = n18563 | n48128 ;
  assign n48130 = ~n5654 & n13523 ;
  assign n48132 = ( n8364 & ~n34300 ) | ( n8364 & n35914 ) | ( ~n34300 & n35914 ) ;
  assign n48131 = n44159 ^ n5823 ^ n3276 ;
  assign n48133 = n48132 ^ n48131 ^ n5437 ;
  assign n48134 = ~n5343 & n48133 ;
  assign n48135 = ~n48130 & n48134 ;
  assign n48136 = n34510 | n39943 ;
  assign n48137 = n48136 ^ n1593 ^ 1'b0 ;
  assign n48138 = n5225 & ~n27913 ;
  assign n48139 = n48138 ^ n9509 ^ 1'b0 ;
  assign n48140 = ( n1990 & n10689 ) | ( n1990 & n48139 ) | ( n10689 & n48139 ) ;
  assign n48141 = n18914 ^ n12062 ^ n320 ;
  assign n48145 = ( n30666 & n34998 ) | ( n30666 & n36116 ) | ( n34998 & n36116 ) ;
  assign n48143 = ~n355 & n13144 ;
  assign n48142 = n34698 ^ n15139 ^ n2545 ;
  assign n48144 = n48143 ^ n48142 ^ n12534 ;
  assign n48146 = n48145 ^ n48144 ^ n28793 ;
  assign n48147 = n25855 ^ n11830 ^ 1'b0 ;
  assign n48148 = ~n1892 & n32547 ;
  assign n48149 = ( n3290 & n19356 ) | ( n3290 & ~n24321 ) | ( n19356 & ~n24321 ) ;
  assign n48150 = ( n48147 & n48148 ) | ( n48147 & n48149 ) | ( n48148 & n48149 ) ;
  assign n48151 = ~n27389 & n33053 ;
  assign n48152 = n48151 ^ n23026 ^ 1'b0 ;
  assign n48153 = n48152 ^ n26620 ^ n13760 ;
  assign n48154 = n45924 ^ n26991 ^ n18006 ;
  assign n48155 = n8233 ^ n4344 ^ 1'b0 ;
  assign n48156 = n36101 ^ n28356 ^ n11499 ;
  assign n48157 = n38047 | n46958 ;
  assign n48158 = n48157 ^ n12125 ^ 1'b0 ;
  assign n48159 = n26295 ^ n12186 ^ 1'b0 ;
  assign n48160 = n17942 | n22696 ;
  assign n48161 = n27768 | n48160 ;
  assign n48162 = ( n34624 & ~n42285 ) | ( n34624 & n48161 ) | ( ~n42285 & n48161 ) ;
  assign n48163 = n2644 | n38238 ;
  assign n48164 = ~n18147 & n31440 ;
  assign n48165 = ( n4234 & n12419 ) | ( n4234 & n35403 ) | ( n12419 & n35403 ) ;
  assign n48166 = ~n8551 & n12885 ;
  assign n48167 = ( n3917 & ~n12764 ) | ( n3917 & n48166 ) | ( ~n12764 & n48166 ) ;
  assign n48168 = n48167 ^ n25277 ^ 1'b0 ;
  assign n48169 = n13440 ^ n10777 ^ n665 ;
  assign n48170 = ~n12427 & n48169 ;
  assign n48171 = n13461 & ~n34214 ;
  assign n48172 = n16955 & ~n33319 ;
  assign n48173 = n48172 ^ n26948 ^ 1'b0 ;
  assign n48174 = ( n17065 & ~n32737 ) | ( n17065 & n48173 ) | ( ~n32737 & n48173 ) ;
  assign n48175 = n48174 ^ n7133 ^ 1'b0 ;
  assign n48176 = n34475 | n48175 ;
  assign n48177 = n48176 ^ n11407 ^ 1'b0 ;
  assign n48178 = n15674 ^ n10330 ^ 1'b0 ;
  assign n48179 = n40946 ^ n37182 ^ 1'b0 ;
  assign n48180 = n10182 & ~n26797 ;
  assign n48181 = n48180 ^ n5212 ^ 1'b0 ;
  assign n48182 = ( n15076 & n19222 ) | ( n15076 & n27334 ) | ( n19222 & n27334 ) ;
  assign n48184 = n30223 | n37632 ;
  assign n48183 = n20079 ^ n10678 ^ n1932 ;
  assign n48185 = n48184 ^ n48183 ^ n26531 ;
  assign n48186 = ( ~n13319 & n13626 ) | ( ~n13319 & n28666 ) | ( n13626 & n28666 ) ;
  assign n48187 = ( ~n27766 & n48185 ) | ( ~n27766 & n48186 ) | ( n48185 & n48186 ) ;
  assign n48188 = n29769 ^ n8139 ^ 1'b0 ;
  assign n48189 = ( n6652 & ~n42074 ) | ( n6652 & n48188 ) | ( ~n42074 & n48188 ) ;
  assign n48190 = n38083 ^ n29475 ^ n17316 ;
  assign n48191 = ( n2640 & n13981 ) | ( n2640 & n28510 ) | ( n13981 & n28510 ) ;
  assign n48192 = n20460 & ~n40591 ;
  assign n48193 = ~n6109 & n29849 ;
  assign n48194 = n48193 ^ n32073 ^ 1'b0 ;
  assign n48195 = ~n5708 & n12813 ;
  assign n48196 = n43299 ^ n33816 ^ n17889 ;
  assign n48197 = n23576 | n48196 ;
  assign n48198 = n40841 ^ n17036 ^ 1'b0 ;
  assign n48199 = ( n16648 & n30178 ) | ( n16648 & ~n34811 ) | ( n30178 & ~n34811 ) ;
  assign n48200 = n9468 ^ n4337 ^ 1'b0 ;
  assign n48201 = n21755 & n48200 ;
  assign n48202 = n15535 & n25196 ;
  assign n48203 = ( n22660 & n29605 ) | ( n22660 & ~n48202 ) | ( n29605 & ~n48202 ) ;
  assign n48204 = ~n11051 & n25405 ;
  assign n48205 = ~n2283 & n48204 ;
  assign n48206 = n12792 ^ n538 ^ 1'b0 ;
  assign n48207 = n10845 & ~n48206 ;
  assign n48208 = n19754 ^ n13723 ^ 1'b0 ;
  assign n48209 = n48207 & ~n48208 ;
  assign n48210 = n25085 ^ n644 ^ 1'b0 ;
  assign n48213 = n6226 & ~n17661 ;
  assign n48214 = n48213 ^ n5663 ^ 1'b0 ;
  assign n48215 = ~n12434 & n48214 ;
  assign n48216 = n48215 ^ n48202 ^ n27519 ;
  assign n48211 = ( n1355 & n3996 ) | ( n1355 & ~n15714 ) | ( n3996 & ~n15714 ) ;
  assign n48212 = n20068 & n48211 ;
  assign n48217 = n48216 ^ n48212 ^ 1'b0 ;
  assign n48218 = n599 & ~n8008 ;
  assign n48219 = n12272 & n48218 ;
  assign n48220 = ( n6418 & n29281 ) | ( n6418 & ~n42887 ) | ( n29281 & ~n42887 ) ;
  assign n48221 = ( n4828 & n48219 ) | ( n4828 & n48220 ) | ( n48219 & n48220 ) ;
  assign n48222 = n48221 ^ n38310 ^ n30131 ;
  assign n48223 = n48222 ^ n28663 ^ n3556 ;
  assign n48224 = ( n26041 & ~n30798 ) | ( n26041 & n48223 ) | ( ~n30798 & n48223 ) ;
  assign n48225 = n35413 ^ n13759 ^ n5799 ;
  assign n48226 = n7504 ^ n6599 ^ n509 ;
  assign n48227 = n20313 | n48226 ;
  assign n48228 = n29058 ^ n13523 ^ n6721 ;
  assign n48229 = n48228 ^ n9092 ^ 1'b0 ;
  assign n48230 = n1470 & n25016 ;
  assign n48231 = n48230 ^ n4315 ^ 1'b0 ;
  assign n48232 = n48231 ^ n24277 ^ 1'b0 ;
  assign n48233 = n18518 ^ n12845 ^ 1'b0 ;
  assign n48234 = n48233 ^ n41045 ^ n23141 ;
  assign n48235 = n34528 ^ n24893 ^ n7029 ;
  assign n48236 = n19457 ^ n6003 ^ 1'b0 ;
  assign n48237 = n7268 & ~n48236 ;
  assign n48238 = n48237 ^ n32773 ^ n28599 ;
  assign n48239 = ( n41044 & ~n48235 ) | ( n41044 & n48238 ) | ( ~n48235 & n48238 ) ;
  assign n48240 = n3330 | n48239 ;
  assign n48241 = n48240 ^ n15479 ^ 1'b0 ;
  assign n48242 = n394 | n46185 ;
  assign n48243 = x151 & ~n48242 ;
  assign n48244 = n48243 ^ n8785 ^ 1'b0 ;
  assign n48245 = n48244 ^ n21666 ^ 1'b0 ;
  assign n48246 = ~n16632 & n48245 ;
  assign n48247 = n10822 & ~n17180 ;
  assign n48248 = n48247 ^ n17724 ^ 1'b0 ;
  assign n48249 = ( n24001 & n33842 ) | ( n24001 & ~n48248 ) | ( n33842 & ~n48248 ) ;
  assign n48250 = ( ~n5459 & n19545 ) | ( ~n5459 & n48249 ) | ( n19545 & n48249 ) ;
  assign n48251 = n25034 & n48250 ;
  assign n48252 = ~n32159 & n48251 ;
  assign n48253 = n13429 | n25652 ;
  assign n48254 = n48253 ^ n34943 ^ 1'b0 ;
  assign n48255 = ( n2967 & n11951 ) | ( n2967 & n23549 ) | ( n11951 & n23549 ) ;
  assign n48256 = n34451 & n48255 ;
  assign n48257 = n9565 & ~n28356 ;
  assign n48258 = n36564 ^ n30594 ^ 1'b0 ;
  assign n48259 = n28044 ^ n21341 ^ 1'b0 ;
  assign n48260 = n30846 ^ n12553 ^ n10349 ;
  assign n48261 = n48260 ^ n31240 ^ n2098 ;
  assign n48262 = ~n2987 & n4424 ;
  assign n48263 = n48261 & n48262 ;
  assign n48265 = n11655 & ~n40851 ;
  assign n48266 = n48265 ^ n7990 ^ 1'b0 ;
  assign n48264 = n27048 ^ n25797 ^ 1'b0 ;
  assign n48267 = n48266 ^ n48264 ^ n6969 ;
  assign n48268 = n23269 | n45449 ;
  assign n48270 = n20069 ^ n17466 ^ 1'b0 ;
  assign n48271 = n5183 & ~n48270 ;
  assign n48269 = ~n25839 & n34163 ;
  assign n48272 = n48271 ^ n48269 ^ 1'b0 ;
  assign n48273 = ( n48267 & n48268 ) | ( n48267 & ~n48272 ) | ( n48268 & ~n48272 ) ;
  assign n48274 = n48273 ^ n20021 ^ n12976 ;
  assign n48275 = n7859 & n48274 ;
  assign n48276 = n37678 & n48275 ;
  assign n48277 = n12418 & ~n32425 ;
  assign n48278 = n12136 & ~n12250 ;
  assign n48279 = n48278 ^ n33951 ^ 1'b0 ;
  assign n48280 = ( n28989 & ~n48277 ) | ( n28989 & n48279 ) | ( ~n48277 & n48279 ) ;
  assign n48281 = n1997 & n40422 ;
  assign n48282 = n48281 ^ n43486 ^ n2504 ;
  assign n48283 = ( n45435 & ~n48280 ) | ( n45435 & n48282 ) | ( ~n48280 & n48282 ) ;
  assign n48290 = n25443 ^ n4527 ^ 1'b0 ;
  assign n48291 = n38342 & ~n48290 ;
  assign n48292 = n48291 ^ n32922 ^ 1'b0 ;
  assign n48285 = n26901 & n27248 ;
  assign n48286 = n48285 ^ n39369 ^ 1'b0 ;
  assign n48287 = ( n12729 & n21261 ) | ( n12729 & n48286 ) | ( n21261 & n48286 ) ;
  assign n48288 = n23655 & n48287 ;
  assign n48289 = n48288 ^ n22736 ^ 1'b0 ;
  assign n48284 = n34178 ^ n12504 ^ n5602 ;
  assign n48293 = n48292 ^ n48289 ^ n48284 ;
  assign n48294 = ( n3801 & n9651 ) | ( n3801 & ~n11367 ) | ( n9651 & ~n11367 ) ;
  assign n48295 = ( ~n28176 & n35684 ) | ( ~n28176 & n48294 ) | ( n35684 & n48294 ) ;
  assign n48296 = n40499 ^ n38779 ^ n33276 ;
  assign n48297 = n48296 ^ n4193 ^ 1'b0 ;
  assign n48298 = ~n4315 & n6040 ;
  assign n48299 = n48298 ^ n5797 ^ 1'b0 ;
  assign n48300 = n48299 ^ n40520 ^ n36383 ;
  assign n48301 = n45978 ^ n14914 ^ 1'b0 ;
  assign n48302 = n38909 & n48301 ;
  assign n48303 = n6944 | n25499 ;
  assign n48304 = n39318 | n48303 ;
  assign n48305 = n48304 ^ n38532 ^ n15624 ;
  assign n48306 = ~n41943 & n48305 ;
  assign n48307 = n21335 & n48306 ;
  assign n48308 = n48307 ^ n43303 ^ n33472 ;
  assign n48309 = n48308 ^ n1233 ^ 1'b0 ;
  assign n48310 = n48302 & ~n48309 ;
  assign n48311 = n41375 ^ n11488 ^ 1'b0 ;
  assign n48312 = n44173 & n48311 ;
  assign n48313 = n8000 & ~n29998 ;
  assign n48314 = ~n307 & n48313 ;
  assign n48315 = ~n26571 & n31064 ;
  assign n48316 = n48315 ^ n24987 ^ 1'b0 ;
  assign n48317 = n46329 | n48316 ;
  assign n48318 = n26575 | n29040 ;
  assign n48319 = n44287 ^ n7829 ^ 1'b0 ;
  assign n48320 = n2750 & n30777 ;
  assign n48321 = n27832 ^ n16230 ^ 1'b0 ;
  assign n48322 = n2946 & n9061 ;
  assign n48323 = n27574 & n48322 ;
  assign n48324 = ( n1155 & ~n2782 ) | ( n1155 & n48323 ) | ( ~n2782 & n48323 ) ;
  assign n48325 = n38834 ^ n13722 ^ n12198 ;
  assign n48326 = n11452 & ~n42981 ;
  assign n48327 = n6404 | n18253 ;
  assign n48328 = n48327 ^ n2145 ^ 1'b0 ;
  assign n48329 = ~n2684 & n48328 ;
  assign n48330 = ~n48326 & n48329 ;
  assign n48331 = n40189 ^ n18711 ^ 1'b0 ;
  assign n48332 = n3523 | n19663 ;
  assign n48333 = n2661 | n48332 ;
  assign n48334 = n18385 ^ n17449 ^ n8544 ;
  assign n48335 = n27310 ^ n3342 ^ 1'b0 ;
  assign n48336 = n7679 & n48335 ;
  assign n48337 = n1981 & n48336 ;
  assign n48338 = ( n3958 & ~n19139 ) | ( n3958 & n48337 ) | ( ~n19139 & n48337 ) ;
  assign n48339 = n48334 & n48338 ;
  assign n48340 = ( n857 & ~n952 ) | ( n857 & n8015 ) | ( ~n952 & n8015 ) ;
  assign n48341 = ( n7097 & n33106 ) | ( n7097 & ~n34451 ) | ( n33106 & ~n34451 ) ;
  assign n48342 = ( n26045 & n29316 ) | ( n26045 & ~n33898 ) | ( n29316 & ~n33898 ) ;
  assign n48343 = n33921 ^ n12032 ^ n1264 ;
  assign n48344 = n14281 & n37273 ;
  assign n48345 = n18576 & n48344 ;
  assign n48346 = n8138 & ~n20754 ;
  assign n48347 = n48346 ^ n301 ^ 1'b0 ;
  assign n48348 = ~n1100 & n48347 ;
  assign n48349 = n37267 ^ n7874 ^ 1'b0 ;
  assign n48350 = n45198 & n48349 ;
  assign n48351 = n38736 ^ n5702 ^ 1'b0 ;
  assign n48352 = n46642 ^ n279 ^ 1'b0 ;
  assign n48353 = n33371 ^ n12008 ^ x83 ;
  assign n48354 = n8209 | n17042 ;
  assign n48355 = n40700 ^ n20234 ^ n8514 ;
  assign n48356 = ( n10072 & ~n10896 ) | ( n10072 & n28749 ) | ( ~n10896 & n28749 ) ;
  assign n48357 = ( n10132 & n11666 ) | ( n10132 & n30953 ) | ( n11666 & n30953 ) ;
  assign n48358 = n48357 ^ n12275 ^ 1'b0 ;
  assign n48359 = n48358 ^ n5042 ^ n1797 ;
  assign n48360 = n48359 ^ n7766 ^ 1'b0 ;
  assign n48362 = ( n9177 & n11894 ) | ( n9177 & n18860 ) | ( n11894 & n18860 ) ;
  assign n48361 = n6334 & n38335 ;
  assign n48363 = n48362 ^ n48361 ^ n4618 ;
  assign n48364 = ~n29939 & n45059 ;
  assign n48365 = n48364 ^ n40981 ^ 1'b0 ;
  assign n48366 = ( n14419 & n35592 ) | ( n14419 & ~n48365 ) | ( n35592 & ~n48365 ) ;
  assign n48367 = n37608 ^ n27685 ^ n25368 ;
  assign n48368 = n47537 ^ n8307 ^ 1'b0 ;
  assign n48369 = ~n4293 & n6234 ;
  assign n48370 = n48369 ^ n21581 ^ 1'b0 ;
  assign n48371 = n19521 ^ n3151 ^ 1'b0 ;
  assign n48372 = n48370 & n48371 ;
  assign n48373 = ~x158 & n48372 ;
  assign n48374 = n37007 ^ n16068 ^ n2230 ;
  assign n48375 = n48374 ^ n17560 ^ 1'b0 ;
  assign n48376 = ~n43246 & n48375 ;
  assign n48377 = n19894 | n29756 ;
  assign n48378 = n40338 | n48377 ;
  assign n48379 = n43793 ^ n37192 ^ n32748 ;
  assign n48380 = n8799 & n44889 ;
  assign n48381 = n48380 ^ n37273 ^ n5718 ;
  assign n48382 = ~n8053 & n38438 ;
  assign n48383 = n45205 ^ n33887 ^ n2138 ;
  assign n48384 = n38861 ^ n3225 ^ 1'b0 ;
  assign n48385 = ~n48351 & n48384 ;
  assign n48386 = n48385 ^ n16904 ^ n12231 ;
  assign n48387 = n25484 ^ n9568 ^ 1'b0 ;
  assign n48388 = n7952 & ~n48387 ;
  assign n48389 = n48388 ^ n39056 ^ 1'b0 ;
  assign n48390 = n36517 & ~n48389 ;
  assign n48391 = n12318 & n48390 ;
  assign n48392 = n48391 ^ n43446 ^ 1'b0 ;
  assign n48393 = ~n4988 & n16330 ;
  assign n48394 = n47724 ^ n31213 ^ 1'b0 ;
  assign n48395 = n10220 & ~n48394 ;
  assign n48396 = ( n2311 & n3034 ) | ( n2311 & ~n41724 ) | ( n3034 & ~n41724 ) ;
  assign n48397 = n21014 & n48280 ;
  assign n48398 = ( n812 & ~n2659 ) | ( n812 & n5408 ) | ( ~n2659 & n5408 ) ;
  assign n48399 = n34501 ^ n21473 ^ 1'b0 ;
  assign n48400 = n17288 ^ n9671 ^ n7393 ;
  assign n48401 = n29787 ^ n25111 ^ n3364 ;
  assign n48402 = n48401 ^ n31035 ^ 1'b0 ;
  assign n48403 = n32227 ^ n15693 ^ 1'b0 ;
  assign n48404 = n48402 | n48403 ;
  assign n48405 = n24744 | n47994 ;
  assign n48406 = n48405 ^ n275 ^ 1'b0 ;
  assign n48407 = ~n15963 & n28228 ;
  assign n48408 = n7384 & n48407 ;
  assign n48409 = ( n725 & n7554 ) | ( n725 & n21081 ) | ( n7554 & n21081 ) ;
  assign n48410 = n41091 & n48409 ;
  assign n48411 = n48410 ^ n40893 ^ 1'b0 ;
  assign n48412 = n9711 | n17326 ;
  assign n48413 = ~n16376 & n24775 ;
  assign n48414 = n48413 ^ n1343 ^ 1'b0 ;
  assign n48415 = n39382 ^ n5068 ^ 1'b0 ;
  assign n48416 = n5509 | n5581 ;
  assign n48417 = n33945 & n48416 ;
  assign n48418 = n15504 | n26834 ;
  assign n48419 = n31020 | n48418 ;
  assign n48420 = n4693 & ~n29562 ;
  assign n48421 = ~n48419 & n48420 ;
  assign n48422 = n31117 & ~n46136 ;
  assign n48423 = n48421 & n48422 ;
  assign n48427 = n2405 & ~n10001 ;
  assign n48424 = n6674 ^ n6000 ^ 1'b0 ;
  assign n48425 = ~n25881 & n48424 ;
  assign n48426 = n48425 ^ n16237 ^ 1'b0 ;
  assign n48428 = n48427 ^ n48426 ^ 1'b0 ;
  assign n48429 = n22266 & n37127 ;
  assign n48430 = n48429 ^ n36029 ^ 1'b0 ;
  assign n48431 = n7377 | n8736 ;
  assign n48432 = n9403 & ~n48431 ;
  assign n48433 = ( n31354 & ~n44078 ) | ( n31354 & n48432 ) | ( ~n44078 & n48432 ) ;
  assign n48434 = n48433 ^ n41969 ^ n28581 ;
  assign n48435 = ~n3166 & n31032 ;
  assign n48436 = n48435 ^ n10350 ^ 1'b0 ;
  assign n48437 = n44417 ^ n39438 ^ n22266 ;
  assign n48438 = n24041 ^ n1277 ^ 1'b0 ;
  assign n48439 = n3432 & n48438 ;
  assign n48440 = n48439 ^ n15792 ^ 1'b0 ;
  assign n48441 = n19159 ^ n9227 ^ 1'b0 ;
  assign n48442 = ~n48440 & n48441 ;
  assign n48443 = n41363 & n48442 ;
  assign n48444 = ( n20617 & n24838 ) | ( n20617 & n44634 ) | ( n24838 & n44634 ) ;
  assign n48445 = n41442 ^ n17930 ^ 1'b0 ;
  assign n48446 = n48445 ^ n38717 ^ n16076 ;
  assign n48447 = n9413 & ~n48446 ;
  assign n48448 = n48447 ^ n14358 ^ 1'b0 ;
  assign n48449 = ~n47304 & n48448 ;
  assign n48450 = ~n15849 & n16969 ;
  assign n48451 = ~n6937 & n48450 ;
  assign n48452 = n14797 & n48451 ;
  assign n48453 = n6676 & ~n48452 ;
  assign n48454 = n28084 & n48453 ;
  assign n48455 = n39808 ^ n4412 ^ 1'b0 ;
  assign n48456 = n40750 & ~n48455 ;
  assign n48457 = ( n1482 & n17030 ) | ( n1482 & ~n25168 ) | ( n17030 & ~n25168 ) ;
  assign n48458 = ( n19123 & n32350 ) | ( n19123 & n48457 ) | ( n32350 & n48457 ) ;
  assign n48459 = n43646 ^ n1623 ^ 1'b0 ;
  assign n48460 = ( ~n2952 & n16451 ) | ( ~n2952 & n40832 ) | ( n16451 & n40832 ) ;
  assign n48461 = ( ~n5992 & n27963 ) | ( ~n5992 & n48460 ) | ( n27963 & n48460 ) ;
  assign n48462 = ( n2337 & n34625 ) | ( n2337 & ~n48461 ) | ( n34625 & ~n48461 ) ;
  assign n48463 = n36656 ^ n25385 ^ 1'b0 ;
  assign n48464 = n29407 & n48463 ;
  assign n48465 = n48464 ^ n34673 ^ n31491 ;
  assign n48466 = ( ~n30124 & n42716 ) | ( ~n30124 & n47846 ) | ( n42716 & n47846 ) ;
  assign n48467 = n33802 & ~n41393 ;
  assign n48468 = n48467 ^ n4682 ^ 1'b0 ;
  assign n48469 = n28545 & ~n35340 ;
  assign n48470 = n48469 ^ n34669 ^ 1'b0 ;
  assign n48471 = n13848 ^ n3231 ^ n1793 ;
  assign n48472 = n14727 | n48471 ;
  assign n48473 = n8895 & ~n48472 ;
  assign n48474 = n46630 ^ n29809 ^ 1'b0 ;
  assign n48475 = n14077 & n33856 ;
  assign n48476 = n48475 ^ n2367 ^ 1'b0 ;
  assign n48477 = ( n23077 & n33387 ) | ( n23077 & n48476 ) | ( n33387 & n48476 ) ;
  assign n48478 = n44707 ^ n11579 ^ n374 ;
  assign n48479 = ( ~n17479 & n23054 ) | ( ~n17479 & n36720 ) | ( n23054 & n36720 ) ;
  assign n48480 = n4095 ^ n1190 ^ 1'b0 ;
  assign n48481 = ~n812 & n25310 ;
  assign n48482 = n24450 & n46599 ;
  assign n48483 = n2167 & ~n30474 ;
  assign n48484 = ( n1394 & ~n28777 ) | ( n1394 & n33920 ) | ( ~n28777 & n33920 ) ;
  assign n48485 = n11541 & n42578 ;
  assign n48486 = n26719 ^ n752 ^ 1'b0 ;
  assign n48487 = n8079 & n13703 ;
  assign n48488 = ~n22453 & n48487 ;
  assign n48489 = n21896 ^ n6014 ^ 1'b0 ;
  assign n48490 = n17076 | n48489 ;
  assign n48491 = n48490 ^ n4316 ^ 1'b0 ;
  assign n48492 = n17591 & ~n44770 ;
  assign n48493 = n48492 ^ n5713 ^ 1'b0 ;
  assign n48494 = n21912 & n48493 ;
  assign n48495 = ~n26910 & n48494 ;
  assign n48496 = n44872 ^ n25467 ^ n1410 ;
  assign n48497 = n48496 ^ n10717 ^ 1'b0 ;
  assign n48498 = n4750 ^ n2418 ^ 1'b0 ;
  assign n48499 = ~n10499 & n48498 ;
  assign n48500 = ( n14650 & n22525 ) | ( n14650 & n48499 ) | ( n22525 & n48499 ) ;
  assign n48501 = n23364 ^ n4830 ^ 1'b0 ;
  assign n48502 = n12591 ^ n8635 ^ 1'b0 ;
  assign n48503 = n48502 ^ n11975 ^ n5253 ;
  assign n48504 = n5800 ^ n5723 ^ n1803 ;
  assign n48505 = n15219 ^ n14523 ^ n7752 ;
  assign n48506 = ( n4203 & ~n17476 ) | ( n4203 & n48505 ) | ( ~n17476 & n48505 ) ;
  assign n48507 = ( n5385 & n48504 ) | ( n5385 & ~n48506 ) | ( n48504 & ~n48506 ) ;
  assign n48508 = n9596 | n45449 ;
  assign n48511 = ( n12781 & ~n22963 ) | ( n12781 & n40942 ) | ( ~n22963 & n40942 ) ;
  assign n48509 = n20213 ^ n7384 ^ 1'b0 ;
  assign n48510 = n43347 & ~n48509 ;
  assign n48512 = n48511 ^ n48510 ^ 1'b0 ;
  assign n48513 = n48512 ^ n36880 ^ n9325 ;
  assign n48517 = n21252 ^ n10589 ^ 1'b0 ;
  assign n48514 = ( n3992 & ~n7377 ) | ( n3992 & n43720 ) | ( ~n7377 & n43720 ) ;
  assign n48515 = ( n6094 & ~n15924 ) | ( n6094 & n27154 ) | ( ~n15924 & n27154 ) ;
  assign n48516 = ( n16283 & n48514 ) | ( n16283 & n48515 ) | ( n48514 & n48515 ) ;
  assign n48518 = n48517 ^ n48516 ^ n3863 ;
  assign n48519 = n8644 & ~n38434 ;
  assign n48522 = x52 & ~n19818 ;
  assign n48523 = ~n752 & n48522 ;
  assign n48520 = n26440 ^ n9977 ^ 1'b0 ;
  assign n48521 = n802 & ~n48520 ;
  assign n48524 = n48523 ^ n48521 ^ 1'b0 ;
  assign n48525 = n8632 & n12807 ;
  assign n48526 = n48525 ^ n12618 ^ 1'b0 ;
  assign n48527 = ~n5340 & n46674 ;
  assign n48530 = n11746 ^ n9182 ^ n910 ;
  assign n48531 = ( n25604 & n44713 ) | ( n25604 & ~n48530 ) | ( n44713 & ~n48530 ) ;
  assign n48528 = n14265 & n30107 ;
  assign n48529 = n15872 | n48528 ;
  assign n48532 = n48531 ^ n48529 ^ 1'b0 ;
  assign n48533 = n14285 ^ n13159 ^ n7250 ;
  assign n48534 = n20849 & ~n46554 ;
  assign n48536 = ~n6074 & n37515 ;
  assign n48537 = n36818 & n48536 ;
  assign n48535 = n27026 ^ n17497 ^ n1049 ;
  assign n48538 = n48537 ^ n48535 ^ n33138 ;
  assign n48539 = n8676 ^ n6484 ^ n1351 ;
  assign n48540 = ~n26455 & n37637 ;
  assign n48541 = n2110 & n41966 ;
  assign n48542 = n16306 & n26657 ;
  assign n48543 = n45690 & n48542 ;
  assign n48544 = ~n1136 & n3497 ;
  assign n48545 = n48544 ^ n11428 ^ 1'b0 ;
  assign n48546 = n8055 ^ n4413 ^ 1'b0 ;
  assign n48547 = n1455 & n48546 ;
  assign n48548 = n32661 ^ n3632 ^ 1'b0 ;
  assign n48549 = ~n6717 & n48548 ;
  assign n48550 = n29928 ^ n25162 ^ n11999 ;
  assign n48551 = n48550 ^ n22850 ^ 1'b0 ;
  assign n48552 = n8929 ^ n5192 ^ 1'b0 ;
  assign n48553 = n46670 & n48552 ;
  assign n48554 = n7621 & n8593 ;
  assign n48555 = n48554 ^ n21269 ^ 1'b0 ;
  assign n48556 = ( n3804 & n6384 ) | ( n3804 & ~n32531 ) | ( n6384 & ~n32531 ) ;
  assign n48557 = ( ~n24104 & n48555 ) | ( ~n24104 & n48556 ) | ( n48555 & n48556 ) ;
  assign n48558 = ( n1544 & n5888 ) | ( n1544 & n9204 ) | ( n5888 & n9204 ) ;
  assign n48559 = ( n8182 & n16607 ) | ( n8182 & ~n17471 ) | ( n16607 & ~n17471 ) ;
  assign n48560 = ( ~n4256 & n8336 ) | ( ~n4256 & n10625 ) | ( n8336 & n10625 ) ;
  assign n48561 = n48560 ^ n34980 ^ n15217 ;
  assign n48562 = n2882 & ~n11476 ;
  assign n48563 = ~n11595 & n48562 ;
  assign n48564 = n10782 | n29450 ;
  assign n48565 = n48563 & ~n48564 ;
  assign n48566 = n22498 ^ n6515 ^ 1'b0 ;
  assign n48567 = n37326 & ~n48566 ;
  assign n48568 = n24055 ^ n4126 ^ 1'b0 ;
  assign n48569 = n48567 & n48568 ;
  assign n48570 = n11163 ^ n1866 ^ 1'b0 ;
  assign n48571 = n48570 ^ n38229 ^ n29549 ;
  assign n48572 = ( n3818 & n29771 ) | ( n3818 & ~n48571 ) | ( n29771 & ~n48571 ) ;
  assign n48573 = n14309 | n48572 ;
  assign n48574 = n48573 ^ n48474 ^ 1'b0 ;
  assign n48575 = n18783 & ~n24663 ;
  assign n48576 = n22601 & n48575 ;
  assign n48577 = n23307 ^ n14811 ^ 1'b0 ;
  assign n48578 = n24561 & n39220 ;
  assign n48579 = ( n1820 & n46828 ) | ( n1820 & ~n48578 ) | ( n46828 & ~n48578 ) ;
  assign n48580 = ( n9479 & n10537 ) | ( n9479 & n41430 ) | ( n10537 & n41430 ) ;
  assign n48581 = n5336 & n46101 ;
  assign n48582 = ( ~n22238 & n48580 ) | ( ~n22238 & n48581 ) | ( n48580 & n48581 ) ;
  assign n48583 = n14460 & ~n16385 ;
  assign n48584 = n48583 ^ n19441 ^ n17555 ;
  assign n48585 = n17254 ^ n7668 ^ 1'b0 ;
  assign n48586 = ~n41655 & n48585 ;
  assign n48587 = ( n37562 & n38802 ) | ( n37562 & ~n48586 ) | ( n38802 & ~n48586 ) ;
  assign n48588 = n23921 ^ n12370 ^ 1'b0 ;
  assign n48589 = n22251 & ~n33892 ;
  assign n48590 = n23106 & ~n40574 ;
  assign n48593 = n1314 & n20243 ;
  assign n48591 = n24770 ^ n13396 ^ n483 ;
  assign n48592 = n44360 | n48591 ;
  assign n48594 = n48593 ^ n48592 ^ n42555 ;
  assign n48595 = ( n9162 & ~n27871 ) | ( n9162 & n38427 ) | ( ~n27871 & n38427 ) ;
  assign n48596 = ( ~n5566 & n35338 ) | ( ~n5566 & n41091 ) | ( n35338 & n41091 ) ;
  assign n48597 = n13946 ^ n6753 ^ n6305 ;
  assign n48598 = ( ~n11113 & n17800 ) | ( ~n11113 & n34535 ) | ( n17800 & n34535 ) ;
  assign n48599 = n30379 & ~n48598 ;
  assign n48600 = n1344 & n48599 ;
  assign n48601 = ( n10846 & n48597 ) | ( n10846 & ~n48600 ) | ( n48597 & ~n48600 ) ;
  assign n48602 = ~n18226 & n34475 ;
  assign n48603 = n48602 ^ n10048 ^ 1'b0 ;
  assign n48604 = n28516 & n43187 ;
  assign n48605 = n48604 ^ n25203 ^ n24285 ;
  assign n48606 = n448 | n48605 ;
  assign n48607 = n30919 & ~n48606 ;
  assign n48608 = ~n30285 & n48607 ;
  assign n48609 = n37840 ^ n2411 ^ 1'b0 ;
  assign n48610 = n24896 & ~n48609 ;
  assign n48611 = ~n8735 & n42811 ;
  assign n48612 = n48611 ^ n8606 ^ 1'b0 ;
  assign n48613 = n10482 ^ n3739 ^ 1'b0 ;
  assign n48614 = ( n12220 & n30195 ) | ( n12220 & n31826 ) | ( n30195 & n31826 ) ;
  assign n48615 = n24678 ^ n11294 ^ 1'b0 ;
  assign n48618 = n19564 ^ n3807 ^ 1'b0 ;
  assign n48616 = n5976 & n25375 ;
  assign n48617 = ( n7500 & n38630 ) | ( n7500 & n48616 ) | ( n38630 & n48616 ) ;
  assign n48619 = n48618 ^ n48617 ^ n1988 ;
  assign n48620 = n14447 ^ n8422 ^ 1'b0 ;
  assign n48621 = n42960 ^ n13022 ^ n1877 ;
  assign n48622 = n48621 ^ n27145 ^ n14150 ;
  assign n48623 = ~n27065 & n48622 ;
  assign n48624 = ~n48620 & n48623 ;
  assign n48625 = n4954 ^ n840 ^ 1'b0 ;
  assign n48626 = n909 & n48625 ;
  assign n48627 = n17393 & ~n43641 ;
  assign n48628 = ( n3370 & ~n18421 ) | ( n3370 & n48627 ) | ( ~n18421 & n48627 ) ;
  assign n48629 = n48628 ^ n40810 ^ 1'b0 ;
  assign n48630 = n48626 & ~n48629 ;
  assign n48631 = n12842 ^ n6789 ^ 1'b0 ;
  assign n48632 = ~n30635 & n48631 ;
  assign n48633 = n30042 ^ n12131 ^ 1'b0 ;
  assign n48634 = n13478 | n48633 ;
  assign n48635 = ( ~n11505 & n16125 ) | ( ~n11505 & n48634 ) | ( n16125 & n48634 ) ;
  assign n48636 = ( n5338 & n23755 ) | ( n5338 & ~n48635 ) | ( n23755 & ~n48635 ) ;
  assign n48637 = n9952 | n31624 ;
  assign n48638 = n2007 & ~n48637 ;
  assign n48639 = n48638 ^ n5881 ^ n1814 ;
  assign n48640 = n17663 ^ n10265 ^ n3972 ;
  assign n48641 = n48622 ^ n34895 ^ n17397 ;
  assign n48642 = n46449 ^ n42251 ^ n41036 ;
  assign n48643 = ( n15177 & ~n21510 ) | ( n15177 & n44550 ) | ( ~n21510 & n44550 ) ;
  assign n48644 = n48643 ^ n24235 ^ 1'b0 ;
  assign n48645 = n7464 & n29732 ;
  assign n48646 = n1578 & ~n37054 ;
  assign n48647 = n48646 ^ n1753 ^ 1'b0 ;
  assign n48648 = n40395 & ~n48647 ;
  assign n48649 = ~n10643 & n13661 ;
  assign n48650 = ( n9604 & n27555 ) | ( n9604 & n39850 ) | ( n27555 & n39850 ) ;
  assign n48651 = ( n439 & n2031 ) | ( n439 & n21169 ) | ( n2031 & n21169 ) ;
  assign n48652 = n48651 ^ n21179 ^ 1'b0 ;
  assign n48653 = n48650 & ~n48652 ;
  assign n48654 = ~n6598 & n10320 ;
  assign n48655 = n48654 ^ n33218 ^ 1'b0 ;
  assign n48656 = n32721 | n48655 ;
  assign n48657 = ( n23081 & n48653 ) | ( n23081 & ~n48656 ) | ( n48653 & ~n48656 ) ;
  assign n48658 = n46466 ^ n26141 ^ n2965 ;
  assign n48659 = ( ~n7934 & n20818 ) | ( ~n7934 & n23726 ) | ( n20818 & n23726 ) ;
  assign n48660 = ( n23551 & n48097 ) | ( n23551 & ~n48659 ) | ( n48097 & ~n48659 ) ;
  assign n48661 = ( n20077 & n27725 ) | ( n20077 & n30183 ) | ( n27725 & n30183 ) ;
  assign n48662 = n22635 ^ n1803 ^ 1'b0 ;
  assign n48663 = n33767 ^ n12984 ^ n2826 ;
  assign n48664 = n21342 & n47256 ;
  assign n48665 = ( ~n2841 & n48663 ) | ( ~n2841 & n48664 ) | ( n48663 & n48664 ) ;
  assign n48666 = n41012 ^ n38416 ^ 1'b0 ;
  assign n48669 = ( n11264 & ~n14500 ) | ( n11264 & n32105 ) | ( ~n14500 & n32105 ) ;
  assign n48667 = n13566 ^ n5690 ^ n2077 ;
  assign n48668 = n3464 | n48667 ;
  assign n48670 = n48669 ^ n48668 ^ 1'b0 ;
  assign n48671 = n15544 | n34286 ;
  assign n48672 = n34258 & ~n48671 ;
  assign n48673 = n48670 & ~n48672 ;
  assign n48674 = n40918 ^ n39831 ^ n9328 ;
  assign n48675 = n16652 | n47309 ;
  assign n48676 = n19492 & ~n48675 ;
  assign n48677 = ~n11318 & n48676 ;
  assign n48678 = n4398 & ~n25698 ;
  assign n48679 = n2600 & ~n48678 ;
  assign n48681 = ~n1438 & n21833 ;
  assign n48682 = n48681 ^ n412 ^ 1'b0 ;
  assign n48680 = n21591 ^ n20288 ^ n19435 ;
  assign n48683 = n48682 ^ n48680 ^ n10476 ;
  assign n48684 = n20073 ^ n15530 ^ 1'b0 ;
  assign n48685 = n48684 ^ n29233 ^ n2866 ;
  assign n48686 = n48685 ^ n38009 ^ n23279 ;
  assign n48687 = n46783 ^ n39960 ^ n14666 ;
  assign n48688 = n38337 ^ n9711 ^ 1'b0 ;
  assign n48689 = n46515 & ~n48688 ;
  assign n48690 = n18782 ^ n2729 ^ n534 ;
  assign n48691 = n25841 ^ n15570 ^ 1'b0 ;
  assign n48692 = n48690 & n48691 ;
  assign n48693 = n7278 & n25995 ;
  assign n48694 = ~n34376 & n48693 ;
  assign n48695 = ( n1721 & n34383 ) | ( n1721 & ~n44065 ) | ( n34383 & ~n44065 ) ;
  assign n48696 = n45270 ^ n13035 ^ n9938 ;
  assign n48697 = n48696 ^ n36437 ^ n17574 ;
  assign n48698 = ( n7235 & n15274 ) | ( n7235 & ~n28402 ) | ( n15274 & ~n28402 ) ;
  assign n48699 = n3651 | n14042 ;
  assign n48700 = n48699 ^ n1089 ^ 1'b0 ;
  assign n48701 = n48700 ^ n30917 ^ n15501 ;
  assign n48702 = n40670 ^ n17385 ^ n1969 ;
  assign n48703 = ( ~n7890 & n30962 ) | ( ~n7890 & n48702 ) | ( n30962 & n48702 ) ;
  assign n48704 = ( n18894 & ~n40970 ) | ( n18894 & n48703 ) | ( ~n40970 & n48703 ) ;
  assign n48705 = n15703 & ~n17987 ;
  assign n48706 = ( ~n15062 & n29431 ) | ( ~n15062 & n48705 ) | ( n29431 & n48705 ) ;
  assign n48707 = n7511 ^ n3189 ^ 1'b0 ;
  assign n48708 = n45971 & n48707 ;
  assign n48709 = n48351 ^ n5580 ^ 1'b0 ;
  assign n48710 = ~n10520 & n48709 ;
  assign n48711 = ~n38602 & n48710 ;
  assign n48712 = n48711 ^ n34652 ^ 1'b0 ;
  assign n48713 = n48712 ^ n37297 ^ 1'b0 ;
  assign n48714 = n43881 ^ n34538 ^ n21521 ;
  assign n48715 = x71 & n25589 ;
  assign n48716 = n15461 | n15494 ;
  assign n48717 = n48716 ^ n44159 ^ 1'b0 ;
  assign n48718 = n48717 ^ n46125 ^ x228 ;
  assign n48719 = n48718 ^ n43931 ^ n26453 ;
  assign n48720 = n16532 ^ n9205 ^ n4298 ;
  assign n48721 = n48720 ^ n35920 ^ 1'b0 ;
  assign n48722 = n11783 ^ n8135 ^ 1'b0 ;
  assign n48723 = ~n15529 & n48722 ;
  assign n48724 = n48723 ^ n11113 ^ n4467 ;
  assign n48725 = ~n22807 & n35246 ;
  assign n48726 = ~n48724 & n48725 ;
  assign n48727 = n4779 ^ n2700 ^ 1'b0 ;
  assign n48728 = n48727 ^ n40791 ^ n24324 ;
  assign n48729 = n14592 & n48728 ;
  assign n48730 = n22328 ^ n13031 ^ n11489 ;
  assign n48731 = n17941 & n48730 ;
  assign n48733 = n43250 & ~n46664 ;
  assign n48734 = n33576 & n48733 ;
  assign n48732 = ~n44441 & n48258 ;
  assign n48735 = n48734 ^ n48732 ^ 1'b0 ;
  assign n48736 = ( n18813 & n22625 ) | ( n18813 & n29239 ) | ( n22625 & n29239 ) ;
  assign n48737 = n2936 & ~n4325 ;
  assign n48738 = n48737 ^ n13877 ^ x197 ;
  assign n48739 = n48736 & n48738 ;
  assign n48740 = n24001 ^ n17178 ^ n11108 ;
  assign n48741 = n1072 | n39939 ;
  assign n48742 = n29921 & ~n48741 ;
  assign n48743 = ( n14942 & ~n34085 ) | ( n14942 & n48742 ) | ( ~n34085 & n48742 ) ;
  assign n48744 = ~n48740 & n48743 ;
  assign n48745 = n2140 | n2247 ;
  assign n48746 = n48745 ^ n8851 ^ 1'b0 ;
  assign n48747 = n48746 ^ n36998 ^ 1'b0 ;
  assign n48748 = n48744 | n48747 ;
  assign n48749 = n23446 ^ n22644 ^ n7073 ;
  assign n48752 = ( ~n911 & n9074 ) | ( ~n911 & n28416 ) | ( n9074 & n28416 ) ;
  assign n48751 = n16190 & ~n20330 ;
  assign n48753 = n48752 ^ n48751 ^ 1'b0 ;
  assign n48750 = n25538 & ~n33294 ;
  assign n48754 = n48753 ^ n48750 ^ 1'b0 ;
  assign n48755 = n48754 ^ n21561 ^ n4209 ;
  assign n48756 = n41968 ^ n26173 ^ 1'b0 ;
  assign n48757 = n7470 & ~n10498 ;
  assign n48758 = ~n48756 & n48757 ;
  assign n48759 = n48758 ^ n12524 ^ 1'b0 ;
  assign n48760 = n793 | n4373 ;
  assign n48761 = ( n12857 & ~n17140 ) | ( n12857 & n48760 ) | ( ~n17140 & n48760 ) ;
  assign n48762 = ( n5114 & n33122 ) | ( n5114 & ~n48125 ) | ( n33122 & ~n48125 ) ;
  assign n48763 = ~n32252 & n48762 ;
  assign n48764 = ( n2014 & n16635 ) | ( n2014 & n47777 ) | ( n16635 & n47777 ) ;
  assign n48765 = n39819 ^ n10546 ^ n9292 ;
  assign n48766 = n38363 ^ n19342 ^ n12102 ;
  assign n48767 = ( n29908 & ~n45116 ) | ( n29908 & n48766 ) | ( ~n45116 & n48766 ) ;
  assign n48768 = n24879 ^ n7031 ^ 1'b0 ;
  assign n48769 = n1462 & n48768 ;
  assign n48770 = n30129 ^ n11459 ^ 1'b0 ;
  assign n48771 = ( ~n32570 & n48769 ) | ( ~n32570 & n48770 ) | ( n48769 & n48770 ) ;
  assign n48772 = ~n36829 & n48771 ;
  assign n48774 = ( n3430 & n5171 ) | ( n3430 & ~n18737 ) | ( n5171 & ~n18737 ) ;
  assign n48775 = ( n3169 & n6086 ) | ( n3169 & ~n48774 ) | ( n6086 & ~n48774 ) ;
  assign n48776 = n7094 | n48775 ;
  assign n48777 = n48776 ^ n26744 ^ 1'b0 ;
  assign n48773 = ( ~n1288 & n39044 ) | ( ~n1288 & n45532 ) | ( n39044 & n45532 ) ;
  assign n48778 = n48777 ^ n48773 ^ n5217 ;
  assign n48779 = ( ~n11633 & n18015 ) | ( ~n11633 & n24537 ) | ( n18015 & n24537 ) ;
  assign n48780 = n47037 ^ n44336 ^ n9664 ;
  assign n48781 = ( n18863 & n48779 ) | ( n18863 & n48780 ) | ( n48779 & n48780 ) ;
  assign n48782 = n30931 ^ n21780 ^ 1'b0 ;
  assign n48783 = n17976 & n48782 ;
  assign n48784 = n14811 & n17081 ;
  assign n48785 = n48784 ^ n30474 ^ 1'b0 ;
  assign n48786 = n40246 ^ n22130 ^ n5760 ;
  assign n48787 = n22211 | n48786 ;
  assign n48788 = n32906 & ~n48787 ;
  assign n48789 = ~n22423 & n43572 ;
  assign n48790 = ( n1399 & ~n8677 ) | ( n1399 & n15677 ) | ( ~n8677 & n15677 ) ;
  assign n48791 = ( n1751 & n3596 ) | ( n1751 & n16500 ) | ( n3596 & n16500 ) ;
  assign n48792 = n48791 ^ n42003 ^ n13810 ;
  assign n48793 = n9605 | n19750 ;
  assign n48794 = n3413 | n48793 ;
  assign n48795 = n48794 ^ n25798 ^ 1'b0 ;
  assign n48796 = n48795 ^ n20826 ^ n13429 ;
  assign n48797 = n48796 ^ n26138 ^ n24702 ;
  assign n48798 = ( ~n17944 & n22073 ) | ( ~n17944 & n45651 ) | ( n22073 & n45651 ) ;
  assign n48799 = ( n8228 & n19074 ) | ( n8228 & n23535 ) | ( n19074 & n23535 ) ;
  assign n48800 = ~n22858 & n41816 ;
  assign n48802 = n39414 ^ n26913 ^ 1'b0 ;
  assign n48803 = ( n26151 & ~n29207 ) | ( n26151 & n48802 ) | ( ~n29207 & n48802 ) ;
  assign n48801 = n4780 & ~n20192 ;
  assign n48804 = n48803 ^ n48801 ^ 1'b0 ;
  assign n48805 = ~n16682 & n47789 ;
  assign n48806 = n39078 & n48805 ;
  assign n48807 = n36698 ^ n7551 ^ 1'b0 ;
  assign n48808 = n30522 ^ n17391 ^ 1'b0 ;
  assign n48809 = n45884 ^ n22277 ^ 1'b0 ;
  assign n48810 = ~n24661 & n48809 ;
  assign n48811 = n48810 ^ n10170 ^ n3340 ;
  assign n48812 = ( ~n6479 & n11831 ) | ( ~n6479 & n26322 ) | ( n11831 & n26322 ) ;
  assign n48813 = n36422 ^ n23895 ^ n19216 ;
  assign n48814 = n44751 ^ n40297 ^ n29067 ;
  assign n48815 = ( n2142 & ~n5638 ) | ( n2142 & n10140 ) | ( ~n5638 & n10140 ) ;
  assign n48816 = n4560 | n48815 ;
  assign n48817 = x120 | n48816 ;
  assign n48818 = n9693 & ~n28750 ;
  assign n48819 = n43886 & n48818 ;
  assign n48820 = n16279 & n35846 ;
  assign n48821 = ~n8704 & n48820 ;
  assign n48822 = ( n9231 & ~n11197 ) | ( n9231 & n46874 ) | ( ~n11197 & n46874 ) ;
  assign n48823 = ( n8813 & n18372 ) | ( n8813 & ~n48822 ) | ( n18372 & ~n48822 ) ;
  assign n48826 = n39653 ^ n32972 ^ 1'b0 ;
  assign n48824 = ( n18951 & n31529 ) | ( n18951 & ~n34121 ) | ( n31529 & ~n34121 ) ;
  assign n48825 = n1957 | n48824 ;
  assign n48827 = n48826 ^ n48825 ^ 1'b0 ;
  assign n48828 = ( n3771 & ~n40841 ) | ( n3771 & n48827 ) | ( ~n40841 & n48827 ) ;
  assign n48829 = n6026 ^ n5265 ^ 1'b0 ;
  assign n48830 = n5720 & ~n48829 ;
  assign n48831 = ( ~n28321 & n31425 ) | ( ~n28321 & n48830 ) | ( n31425 & n48830 ) ;
  assign n48832 = n15839 ^ n4642 ^ 1'b0 ;
  assign n48833 = n4767 & ~n7009 ;
  assign n48834 = ( n8447 & n15667 ) | ( n8447 & ~n48833 ) | ( n15667 & ~n48833 ) ;
  assign n48835 = n10333 & ~n24582 ;
  assign n48836 = n48835 ^ n46421 ^ 1'b0 ;
  assign n48837 = ( n4744 & n48834 ) | ( n4744 & ~n48836 ) | ( n48834 & ~n48836 ) ;
  assign n48838 = n48837 ^ n6479 ^ 1'b0 ;
  assign n48839 = n36196 ^ n11094 ^ 1'b0 ;
  assign n48840 = n29877 & ~n48839 ;
  assign n48841 = n6876 | n13152 ;
  assign n48842 = n15562 & n48841 ;
  assign n48843 = n18154 | n42043 ;
  assign n48844 = n48843 ^ n11099 ^ 1'b0 ;
  assign n48845 = ( n18818 & n25515 ) | ( n18818 & n30670 ) | ( n25515 & n30670 ) ;
  assign n48846 = n35843 | n48845 ;
  assign n48847 = n17575 ^ n8130 ^ 1'b0 ;
  assign n48848 = ( n19461 & ~n30700 ) | ( n19461 & n48847 ) | ( ~n30700 & n48847 ) ;
  assign n48849 = ~n20361 & n22962 ;
  assign n48850 = n48849 ^ n13404 ^ 1'b0 ;
  assign n48851 = ( ~n36140 & n45516 ) | ( ~n36140 & n48850 ) | ( n45516 & n48850 ) ;
  assign n48852 = n2930 & n36543 ;
  assign n48853 = n22476 ^ n20793 ^ n16208 ;
  assign n48854 = n12730 & n48853 ;
  assign n48855 = n11905 | n37449 ;
  assign n48856 = n6806 | n48855 ;
  assign n48857 = n35853 ^ n16675 ^ 1'b0 ;
  assign n48858 = n12971 | n48857 ;
  assign n48859 = n48856 & ~n48858 ;
  assign n48860 = n34887 & ~n41252 ;
  assign n48861 = n48860 ^ n16726 ^ n3437 ;
  assign n48862 = n31193 ^ n25197 ^ n25058 ;
  assign n48866 = ( n9259 & n26975 ) | ( n9259 & n29486 ) | ( n26975 & n29486 ) ;
  assign n48867 = n48866 ^ n16776 ^ n3383 ;
  assign n48868 = ~n2532 & n48867 ;
  assign n48863 = n43061 ^ n16292 ^ 1'b0 ;
  assign n48864 = n42782 | n48863 ;
  assign n48865 = ( n27979 & n40888 ) | ( n27979 & n48864 ) | ( n40888 & n48864 ) ;
  assign n48869 = n48868 ^ n48865 ^ n632 ;
  assign n48870 = n48869 ^ n33387 ^ n5420 ;
  assign n48871 = ( n9740 & n21081 ) | ( n9740 & n41761 ) | ( n21081 & n41761 ) ;
  assign n48873 = ( n2139 & n10078 ) | ( n2139 & ~n34042 ) | ( n10078 & ~n34042 ) ;
  assign n48872 = n19774 ^ n7938 ^ n1257 ;
  assign n48874 = n48873 ^ n48872 ^ n12562 ;
  assign n48875 = n46813 ^ n6287 ^ 1'b0 ;
  assign n48876 = ~n48874 & n48875 ;
  assign n48877 = n3162 | n23333 ;
  assign n48878 = n33876 & ~n48877 ;
  assign n48879 = ( n3820 & n4192 ) | ( n3820 & ~n5947 ) | ( n4192 & ~n5947 ) ;
  assign n48880 = n20579 ^ n11952 ^ 1'b0 ;
  assign n48881 = n26955 & n48880 ;
  assign n48882 = n8272 | n48881 ;
  assign n48883 = ( n7788 & n48879 ) | ( n7788 & ~n48882 ) | ( n48879 & ~n48882 ) ;
  assign n48884 = n47846 ^ n22842 ^ n11540 ;
  assign n48885 = n39051 ^ n24859 ^ n23074 ;
  assign n48886 = n5276 & ~n15314 ;
  assign n48887 = n48886 ^ n8606 ^ 1'b0 ;
  assign n48888 = ( n3566 & ~n16219 ) | ( n3566 & n48887 ) | ( ~n16219 & n48887 ) ;
  assign n48889 = n15638 ^ n12630 ^ n2722 ;
  assign n48890 = n19751 | n35807 ;
  assign n48891 = n48890 ^ n31668 ^ n20780 ;
  assign n48892 = n47962 & ~n48891 ;
  assign n48893 = n15132 ^ n793 ^ 1'b0 ;
  assign n48894 = n48893 ^ n3055 ^ n2490 ;
  assign n48895 = n14099 & ~n14559 ;
  assign n48896 = n30966 & n48895 ;
  assign n48897 = n48896 ^ n1714 ^ 1'b0 ;
  assign n48898 = n48894 & n48897 ;
  assign n48899 = n48898 ^ x153 ^ 1'b0 ;
  assign n48900 = n31932 & n48899 ;
  assign n48901 = n1216 ^ n363 ^ 1'b0 ;
  assign n48902 = ~n2407 & n48901 ;
  assign n48903 = n48902 ^ n20597 ^ n18542 ;
  assign n48904 = n45484 ^ n24434 ^ 1'b0 ;
  assign n48905 = ~n48903 & n48904 ;
  assign n48906 = n32699 ^ n28943 ^ 1'b0 ;
  assign n48907 = n48305 & ~n48906 ;
  assign n48908 = n7885 & n48907 ;
  assign n48909 = n48908 ^ n23066 ^ 1'b0 ;
  assign n48910 = n21117 & ~n23752 ;
  assign n48911 = ~n2097 & n48910 ;
  assign n48912 = n41385 ^ n29919 ^ 1'b0 ;
  assign n48913 = n47254 & n48912 ;
  assign n48914 = n27731 ^ n6588 ^ 1'b0 ;
  assign n48915 = x169 & ~n48914 ;
  assign n48916 = ~n23826 & n42184 ;
  assign n48917 = ~n48915 & n48916 ;
  assign n48918 = n48917 ^ n19875 ^ n19470 ;
  assign n48919 = ( n11197 & n25851 ) | ( n11197 & n33344 ) | ( n25851 & n33344 ) ;
  assign n48920 = n48071 ^ n44323 ^ n419 ;
  assign n48921 = n43369 ^ n28149 ^ n12080 ;
  assign n48922 = n48921 ^ n4319 ^ 1'b0 ;
  assign n48923 = ( ~n20423 & n25365 ) | ( ~n20423 & n29244 ) | ( n25365 & n29244 ) ;
  assign n48924 = n3516 | n4512 ;
  assign n48925 = n48924 ^ n10897 ^ 1'b0 ;
  assign n48926 = n2443 | n48925 ;
  assign n48927 = n23212 ^ n10327 ^ 1'b0 ;
  assign n48928 = n16333 | n30095 ;
  assign n48929 = n48927 | n48928 ;
  assign n48930 = n5566 & n20373 ;
  assign n48931 = n48930 ^ n34673 ^ 1'b0 ;
  assign n48932 = n45153 ^ n43335 ^ 1'b0 ;
  assign n48933 = ( n33668 & n45377 ) | ( n33668 & n47045 ) | ( n45377 & n47045 ) ;
  assign n48934 = ( ~n10763 & n21071 ) | ( ~n10763 & n35713 ) | ( n21071 & n35713 ) ;
  assign n48935 = ( n4379 & n19812 ) | ( n4379 & ~n48934 ) | ( n19812 & ~n48934 ) ;
  assign n48936 = n5278 & ~n48845 ;
  assign n48937 = n31017 ^ n25870 ^ n8928 ;
  assign n48938 = n48937 ^ n32446 ^ n26228 ;
  assign n48939 = n13500 & n40116 ;
  assign n48941 = n36379 ^ n21368 ^ n5228 ;
  assign n48940 = ~n11136 & n39322 ;
  assign n48942 = n48941 ^ n48940 ^ 1'b0 ;
  assign n48943 = n36594 & n45523 ;
  assign n48944 = ~x83 & n48943 ;
  assign n48945 = n37602 ^ n511 ^ 1'b0 ;
  assign n48946 = n48945 ^ n5659 ^ 1'b0 ;
  assign n48947 = n8649 & ~n47214 ;
  assign n48948 = ~n48946 & n48947 ;
  assign n48949 = n19279 ^ n3329 ^ 1'b0 ;
  assign n48950 = ~n11137 & n48949 ;
  assign n48951 = ~n6456 & n48950 ;
  assign n48952 = n19595 & n48951 ;
  assign n48953 = n43402 ^ n16372 ^ 1'b0 ;
  assign n48954 = n34273 & n48953 ;
  assign n48955 = n48954 ^ n29410 ^ 1'b0 ;
  assign n48956 = ~n32906 & n37004 ;
  assign n48957 = n48956 ^ n32620 ^ 1'b0 ;
  assign n48958 = n13526 & ~n35602 ;
  assign n48959 = ( n25583 & n48957 ) | ( n25583 & n48958 ) | ( n48957 & n48958 ) ;
  assign n48960 = ( n10647 & ~n40745 ) | ( n10647 & n48959 ) | ( ~n40745 & n48959 ) ;
  assign n48961 = n39510 ^ n18889 ^ n1367 ;
  assign n48962 = n13059 | n26336 ;
  assign n48963 = n28805 & ~n33836 ;
  assign n48964 = n48963 ^ n8447 ^ 1'b0 ;
  assign n48965 = n48964 ^ n17351 ^ 1'b0 ;
  assign n48966 = ( n3604 & n28272 ) | ( n3604 & ~n44491 ) | ( n28272 & ~n44491 ) ;
  assign n48967 = ~n27921 & n33385 ;
  assign n48968 = n10807 & ~n19796 ;
  assign n48969 = n48968 ^ n43673 ^ 1'b0 ;
  assign n48970 = n43284 ^ n12275 ^ 1'b0 ;
  assign n48971 = n48969 | n48970 ;
  assign n48972 = n32299 | n45756 ;
  assign n48973 = n21347 & ~n48972 ;
  assign n48974 = n46809 ^ n21130 ^ 1'b0 ;
  assign n48975 = n20503 & ~n48974 ;
  assign n48976 = n48975 ^ n9332 ^ 1'b0 ;
  assign n48977 = ( n24385 & ~n32298 ) | ( n24385 & n41385 ) | ( ~n32298 & n41385 ) ;
  assign n48978 = ~n32984 & n48977 ;
  assign n48979 = n22353 ^ n15716 ^ 1'b0 ;
  assign n48980 = n48979 ^ n32666 ^ n14724 ;
  assign n48981 = n10244 ^ n8570 ^ 1'b0 ;
  assign n48982 = ( ~n11206 & n13029 ) | ( ~n11206 & n48981 ) | ( n13029 & n48981 ) ;
  assign n48983 = n5421 & n9304 ;
  assign n48984 = n11903 & n48983 ;
  assign n48985 = n13630 ^ n7403 ^ 1'b0 ;
  assign n48986 = n48984 | n48985 ;
  assign n48987 = ( ~n7683 & n48982 ) | ( ~n7683 & n48986 ) | ( n48982 & n48986 ) ;
  assign n48988 = ( ~n7391 & n30886 ) | ( ~n7391 & n39004 ) | ( n30886 & n39004 ) ;
  assign n48989 = n36953 ^ n13195 ^ 1'b0 ;
  assign n48990 = n22028 ^ n13074 ^ n5388 ;
  assign n48991 = n48990 ^ n11965 ^ 1'b0 ;
  assign n48992 = n29127 | n48991 ;
  assign n48993 = n40975 ^ n37980 ^ 1'b0 ;
  assign n48994 = n42076 & n48993 ;
  assign n48995 = ( ~n40115 & n48992 ) | ( ~n40115 & n48994 ) | ( n48992 & n48994 ) ;
  assign n48996 = n16013 | n25698 ;
  assign n48997 = n38599 & ~n48996 ;
  assign n48998 = n4871 | n48997 ;
  assign n48999 = n2401 | n48998 ;
  assign n49000 = n5712 & ~n23849 ;
  assign n49001 = ~n12965 & n49000 ;
  assign n49002 = n17874 ^ n6736 ^ 1'b0 ;
  assign n49003 = n22873 ^ n1129 ^ 1'b0 ;
  assign n49004 = n49002 & ~n49003 ;
  assign n49007 = n20457 ^ n15272 ^ n3354 ;
  assign n49005 = ~n6602 & n21405 ;
  assign n49006 = ( n13354 & n24949 ) | ( n13354 & ~n49005 ) | ( n24949 & ~n49005 ) ;
  assign n49008 = n49007 ^ n49006 ^ 1'b0 ;
  assign n49009 = ~n36215 & n46588 ;
  assign n49011 = n7592 | n28440 ;
  assign n49010 = ( n18461 & ~n26285 ) | ( n18461 & n41250 ) | ( ~n26285 & n41250 ) ;
  assign n49012 = n49011 ^ n49010 ^ n9673 ;
  assign n49013 = ( n3116 & n29190 ) | ( n3116 & n32964 ) | ( n29190 & n32964 ) ;
  assign n49014 = ( n2070 & n15942 ) | ( n2070 & n38935 ) | ( n15942 & n38935 ) ;
  assign n49015 = ( n1010 & n22919 ) | ( n1010 & ~n29002 ) | ( n22919 & ~n29002 ) ;
  assign n49016 = ( n14192 & ~n23052 ) | ( n14192 & n49015 ) | ( ~n23052 & n49015 ) ;
  assign n49017 = n11044 & n41202 ;
  assign n49018 = n3154 ^ n443 ^ 1'b0 ;
  assign n49022 = n15328 ^ n12098 ^ n9396 ;
  assign n49019 = n24838 ^ n9963 ^ 1'b0 ;
  assign n49020 = ~n10180 & n13487 ;
  assign n49021 = n49019 & n49020 ;
  assign n49023 = n49022 ^ n49021 ^ n12640 ;
  assign n49024 = n22034 ^ n12614 ^ n6881 ;
  assign n49025 = n49024 ^ n28149 ^ n27605 ;
  assign n49026 = n49025 ^ n38338 ^ n355 ;
  assign n49027 = n18098 | n49026 ;
  assign n49028 = n49023 | n49027 ;
  assign n49029 = n16318 ^ n9196 ^ x154 ;
  assign n49030 = ~n8337 & n49029 ;
  assign n49031 = n18309 & ~n32635 ;
  assign n49032 = ~n733 & n25849 ;
  assign n49033 = n24199 ^ n18402 ^ n3703 ;
  assign n49034 = ( ~n16156 & n49032 ) | ( ~n16156 & n49033 ) | ( n49032 & n49033 ) ;
  assign n49035 = ( n24300 & n29224 ) | ( n24300 & n49034 ) | ( n29224 & n49034 ) ;
  assign n49036 = n46779 ^ n13484 ^ n8558 ;
  assign n49037 = n2691 & ~n49036 ;
  assign n49038 = ~n31741 & n49037 ;
  assign n49039 = n49038 ^ n28438 ^ n8587 ;
  assign n49040 = n49039 ^ n47866 ^ n42259 ;
  assign n49041 = n38711 ^ n22003 ^ n6588 ;
  assign n49042 = ( n7379 & n16250 ) | ( n7379 & n19133 ) | ( n16250 & n19133 ) ;
  assign n49043 = n6638 & ~n25506 ;
  assign n49044 = ~n13505 & n49043 ;
  assign n49045 = n36641 | n49044 ;
  assign n49046 = n49045 ^ n5840 ^ 1'b0 ;
  assign n49047 = n11455 & n30522 ;
  assign n49048 = n8083 | n23756 ;
  assign n49049 = n49047 & ~n49048 ;
  assign n49050 = n22322 | n30084 ;
  assign n49051 = n49050 ^ n42881 ^ 1'b0 ;
  assign n49052 = n37711 ^ n4145 ^ 1'b0 ;
  assign n49053 = ( n7417 & n8581 ) | ( n7417 & n49052 ) | ( n8581 & n49052 ) ;
  assign n49054 = n23176 ^ n12387 ^ 1'b0 ;
  assign n49055 = n24927 ^ n15117 ^ 1'b0 ;
  assign n49056 = n16655 & n49055 ;
  assign n49057 = ( n17195 & n36891 ) | ( n17195 & n49056 ) | ( n36891 & n49056 ) ;
  assign n49058 = ( n13427 & ~n49054 ) | ( n13427 & n49057 ) | ( ~n49054 & n49057 ) ;
  assign n49059 = ( n1255 & ~n25937 ) | ( n1255 & n29935 ) | ( ~n25937 & n29935 ) ;
  assign n49060 = n7009 ^ n5081 ^ n2962 ;
  assign n49061 = n10888 ^ n5001 ^ 1'b0 ;
  assign n49062 = n47008 ^ n13008 ^ n2595 ;
  assign n49065 = ( n22964 & ~n28803 ) | ( n22964 & n36450 ) | ( ~n28803 & n36450 ) ;
  assign n49066 = n49065 ^ n35542 ^ n28384 ;
  assign n49063 = n26168 ^ n2254 ^ 1'b0 ;
  assign n49064 = n5681 | n49063 ;
  assign n49067 = n49066 ^ n49064 ^ 1'b0 ;
  assign n49068 = ~n5624 & n38250 ;
  assign n49069 = n13093 & ~n35115 ;
  assign n49070 = n37041 ^ n20741 ^ n6806 ;
  assign n49071 = n44344 ^ n33133 ^ n16729 ;
  assign n49072 = n49071 ^ n22514 ^ n8473 ;
  assign n49073 = n6240 & ~n17110 ;
  assign n49074 = ~n2540 & n49073 ;
  assign n49075 = ( n21000 & n43700 ) | ( n21000 & n49074 ) | ( n43700 & n49074 ) ;
  assign n49076 = n49075 ^ n23861 ^ n17263 ;
  assign n49077 = n24925 ^ n20720 ^ n10514 ;
  assign n49078 = ( ~n5029 & n20533 ) | ( ~n5029 & n23484 ) | ( n20533 & n23484 ) ;
  assign n49079 = ( n2247 & ~n7531 ) | ( n2247 & n42334 ) | ( ~n7531 & n42334 ) ;
  assign n49080 = n23230 | n49079 ;
  assign n49081 = n49080 ^ n3731 ^ 1'b0 ;
  assign n49082 = n25322 ^ n1816 ^ 1'b0 ;
  assign n49083 = ~n4664 & n49082 ;
  assign n49084 = ( n11178 & n40602 ) | ( n11178 & ~n49083 ) | ( n40602 & ~n49083 ) ;
  assign n49085 = n15193 & ~n16948 ;
  assign n49086 = n41712 & n49085 ;
  assign n49087 = n46718 & ~n49086 ;
  assign n49088 = ~n49084 & n49087 ;
  assign n49089 = n42221 ^ n33938 ^ n9025 ;
  assign n49090 = n27434 ^ n16221 ^ n12240 ;
  assign n49091 = n6529 | n39278 ;
  assign n49092 = n49091 ^ n12475 ^ n9159 ;
  assign n49093 = n31113 ^ n27666 ^ 1'b0 ;
  assign n49094 = n20506 | n49093 ;
  assign n49095 = n1276 & ~n49094 ;
  assign n49096 = n49095 ^ n12220 ^ n7881 ;
  assign n49097 = ( n9717 & n13356 ) | ( n9717 & n13671 ) | ( n13356 & n13671 ) ;
  assign n49098 = n49097 ^ n29173 ^ n3403 ;
  assign n49099 = n16082 ^ n7016 ^ 1'b0 ;
  assign n49100 = n4041 | n49099 ;
  assign n49101 = n1063 | n40502 ;
  assign n49102 = n33134 ^ n29809 ^ 1'b0 ;
  assign n49103 = n37210 & ~n49102 ;
  assign n49104 = n28679 ^ n15168 ^ 1'b0 ;
  assign n49105 = n11627 & n15829 ;
  assign n49106 = n49105 ^ n11643 ^ 1'b0 ;
  assign n49107 = n49106 ^ n22687 ^ n19355 ;
  assign n49108 = n8952 & ~n31555 ;
  assign n49109 = n26369 ^ n21503 ^ 1'b0 ;
  assign n49120 = n20214 ^ n6196 ^ n5595 ;
  assign n49121 = n49120 ^ n15414 ^ 1'b0 ;
  assign n49112 = n5733 | n35309 ;
  assign n49113 = n1288 | n49112 ;
  assign n49110 = n18838 ^ n17980 ^ n4819 ;
  assign n49111 = ( n3968 & n6625 ) | ( n3968 & ~n49110 ) | ( n6625 & ~n49110 ) ;
  assign n49114 = n49113 ^ n49111 ^ n47787 ;
  assign n49115 = ( n800 & n26196 ) | ( n800 & n49114 ) | ( n26196 & n49114 ) ;
  assign n49116 = n40439 ^ n17231 ^ n4930 ;
  assign n49117 = n39440 ^ n10367 ^ 1'b0 ;
  assign n49118 = n39041 & ~n49117 ;
  assign n49119 = ( n49115 & n49116 ) | ( n49115 & ~n49118 ) | ( n49116 & ~n49118 ) ;
  assign n49122 = n49121 ^ n49119 ^ n4097 ;
  assign n49123 = n25916 & ~n36648 ;
  assign n49124 = n19441 ^ n5949 ^ 1'b0 ;
  assign n49125 = n20206 | n46827 ;
  assign n49129 = n37649 ^ n34256 ^ n26342 ;
  assign n49126 = n12292 & n21050 ;
  assign n49127 = n49126 ^ n17365 ^ 1'b0 ;
  assign n49128 = n27832 & n49127 ;
  assign n49130 = n49129 ^ n49128 ^ 1'b0 ;
  assign n49131 = ( ~n11926 & n40192 ) | ( ~n11926 & n45028 ) | ( n40192 & n45028 ) ;
  assign n49132 = ( n10644 & n14310 ) | ( n10644 & n15084 ) | ( n14310 & n15084 ) ;
  assign n49133 = n33913 & ~n34973 ;
  assign n49134 = ~n4161 & n49133 ;
  assign n49135 = n49134 ^ n42359 ^ n13926 ;
  assign n49136 = ( n4878 & ~n9157 ) | ( n4878 & n11830 ) | ( ~n9157 & n11830 ) ;
  assign n49137 = n34961 ^ n33207 ^ 1'b0 ;
  assign n49138 = ( ~n4327 & n26963 ) | ( ~n4327 & n37972 ) | ( n26963 & n37972 ) ;
  assign n49139 = ~n32321 & n49138 ;
  assign n49140 = n32647 & n49139 ;
  assign n49141 = n20289 | n21033 ;
  assign n49142 = n29525 | n49141 ;
  assign n49143 = n49142 ^ n13142 ^ 1'b0 ;
  assign n49144 = ~n36813 & n42988 ;
  assign n49145 = n10667 & n49144 ;
  assign n49146 = n49145 ^ n19122 ^ 1'b0 ;
  assign n49147 = n19889 | n25416 ;
  assign n49148 = n723 | n19762 ;
  assign n49149 = ( ~n13204 & n14149 ) | ( ~n13204 & n49148 ) | ( n14149 & n49148 ) ;
  assign n49150 = n40664 ^ n8995 ^ n6181 ;
  assign n49151 = n5637 | n19895 ;
  assign n49152 = n49151 ^ n21310 ^ 1'b0 ;
  assign n49154 = ( n2765 & n8756 ) | ( n2765 & ~n21399 ) | ( n8756 & ~n21399 ) ;
  assign n49153 = n9635 ^ n2985 ^ 1'b0 ;
  assign n49155 = n49154 ^ n49153 ^ n44090 ;
  assign n49156 = ~n20623 & n20660 ;
  assign n49157 = ~n4829 & n37150 ;
  assign n49158 = ( n39708 & n49156 ) | ( n39708 & ~n49157 ) | ( n49156 & ~n49157 ) ;
  assign n49159 = ( ~n1786 & n32989 ) | ( ~n1786 & n39363 ) | ( n32989 & n39363 ) ;
  assign n49160 = n24958 ^ n11346 ^ 1'b0 ;
  assign n49161 = ~n49159 & n49160 ;
  assign n49162 = ( n35749 & ~n45362 ) | ( n35749 & n49161 ) | ( ~n45362 & n49161 ) ;
  assign n49163 = n11384 & n40561 ;
  assign n49164 = ~n49162 & n49163 ;
  assign n49165 = n7694 & n27248 ;
  assign n49166 = n49165 ^ n9061 ^ 1'b0 ;
  assign n49167 = n43417 ^ n8658 ^ 1'b0 ;
  assign n49168 = n35927 ^ n19106 ^ n10288 ;
  assign n49169 = ~n30866 & n49168 ;
  assign n49170 = n49169 ^ n16266 ^ n2991 ;
  assign n49171 = n49170 ^ n19667 ^ 1'b0 ;
  assign n49172 = n25738 ^ n6072 ^ x110 ;
  assign n49173 = ( n5620 & ~n8537 ) | ( n5620 & n29544 ) | ( ~n8537 & n29544 ) ;
  assign n49174 = n45187 ^ n43408 ^ 1'b0 ;
  assign n49175 = n3339 & n27306 ;
  assign n49176 = ~n3620 & n31959 ;
  assign n49177 = ~n11255 & n45006 ;
  assign n49178 = n49177 ^ n24005 ^ 1'b0 ;
  assign n49179 = n8423 & ~n10015 ;
  assign n49180 = ( n3440 & ~n17449 ) | ( n3440 & n33425 ) | ( ~n17449 & n33425 ) ;
  assign n49181 = n49180 ^ n25645 ^ 1'b0 ;
  assign n49182 = n49179 & n49181 ;
  assign n49183 = n16664 ^ n7141 ^ 1'b0 ;
  assign n49184 = n1662 | n49183 ;
  assign n49185 = n18513 ^ n16719 ^ 1'b0 ;
  assign n49186 = n17076 | n49185 ;
  assign n49187 = n22201 ^ n14060 ^ n10769 ;
  assign n49188 = n1216 & ~n13802 ;
  assign n49189 = n5809 & n49188 ;
  assign n49190 = n49189 ^ n30750 ^ n21047 ;
  assign n49191 = n46918 ^ n32908 ^ n14994 ;
  assign n49192 = n49191 ^ n24539 ^ n19056 ;
  assign n49193 = n44777 ^ n43244 ^ n4122 ;
  assign n49194 = n12783 & n42568 ;
  assign n49195 = n6799 | n17706 ;
  assign n49196 = n49194 & ~n49195 ;
  assign n49197 = n49196 ^ n7069 ^ 1'b0 ;
  assign n49198 = ( n4412 & ~n19655 ) | ( n4412 & n27700 ) | ( ~n19655 & n27700 ) ;
  assign n49199 = ( n5556 & n13109 ) | ( n5556 & ~n36422 ) | ( n13109 & ~n36422 ) ;
  assign n49200 = n26535 | n49199 ;
  assign n49201 = n30180 ^ n19913 ^ n14870 ;
  assign n49202 = n29888 & n49201 ;
  assign n49203 = n32040 ^ n17687 ^ n8182 ;
  assign n49204 = ~n17942 & n24580 ;
  assign n49205 = ~n49203 & n49204 ;
  assign n49206 = ~n11922 & n16297 ;
  assign n49207 = ~n30876 & n49206 ;
  assign n49208 = ( ~n7184 & n40646 ) | ( ~n7184 & n49207 ) | ( n40646 & n49207 ) ;
  assign n49209 = n22147 ^ n20135 ^ n6671 ;
  assign n49210 = ( n478 & n31552 ) | ( n478 & n49209 ) | ( n31552 & n49209 ) ;
  assign n49212 = n13502 ^ n10146 ^ 1'b0 ;
  assign n49211 = ( n1102 & n6497 ) | ( n1102 & n24860 ) | ( n6497 & n24860 ) ;
  assign n49213 = n49212 ^ n49211 ^ n17990 ;
  assign n49214 = n30248 ^ n27131 ^ n1856 ;
  assign n49215 = n49214 ^ n29733 ^ 1'b0 ;
  assign n49216 = ( n2080 & ~n6216 ) | ( n2080 & n40253 ) | ( ~n6216 & n40253 ) ;
  assign n49217 = ( n7498 & n19333 ) | ( n7498 & ~n31124 ) | ( n19333 & ~n31124 ) ;
  assign n49218 = n13877 | n27691 ;
  assign n49219 = n3305 & ~n49218 ;
  assign n49222 = n46478 ^ n5475 ^ 1'b0 ;
  assign n49223 = n31896 & n49222 ;
  assign n49224 = n11120 & n49223 ;
  assign n49225 = ~n8656 & n49224 ;
  assign n49220 = ~n13528 & n45341 ;
  assign n49221 = n49220 ^ n16791 ^ n2641 ;
  assign n49226 = n49225 ^ n49221 ^ n30194 ;
  assign n49227 = n49226 ^ n48990 ^ n40473 ;
  assign n49228 = ( n5681 & n19353 ) | ( n5681 & ~n25248 ) | ( n19353 & ~n25248 ) ;
  assign n49229 = n9892 | n40435 ;
  assign n49230 = n49229 ^ n48221 ^ 1'b0 ;
  assign n49231 = n31834 ^ n22135 ^ n4477 ;
  assign n49232 = ( ~n7636 & n36168 ) | ( ~n7636 & n46790 ) | ( n36168 & n46790 ) ;
  assign n49236 = n35961 ^ n18505 ^ n6971 ;
  assign n49233 = n19168 ^ n9775 ^ n6966 ;
  assign n49234 = n49233 ^ n18288 ^ n11378 ;
  assign n49235 = n13807 | n49234 ;
  assign n49237 = n49236 ^ n49235 ^ 1'b0 ;
  assign n49238 = n49232 & n49237 ;
  assign n49239 = ( n10887 & n14859 ) | ( n10887 & ~n37223 ) | ( n14859 & ~n37223 ) ;
  assign n49241 = n8594 | n16923 ;
  assign n49242 = n49241 ^ n39342 ^ 1'b0 ;
  assign n49243 = n49242 ^ n48616 ^ n36730 ;
  assign n49240 = ~n13251 & n28855 ;
  assign n49244 = n49243 ^ n49240 ^ 1'b0 ;
  assign n49245 = ~n20705 & n41217 ;
  assign n49246 = n36263 & n49245 ;
  assign n49247 = n46961 ^ n28241 ^ 1'b0 ;
  assign n49248 = ( x195 & n5548 ) | ( x195 & ~n16742 ) | ( n5548 & ~n16742 ) ;
  assign n49249 = n14297 & ~n27074 ;
  assign n49250 = ( ~n37176 & n49248 ) | ( ~n37176 & n49249 ) | ( n49248 & n49249 ) ;
  assign n49251 = n32028 ^ n20425 ^ n2853 ;
  assign n49252 = n49251 ^ n41017 ^ n26680 ;
  assign n49253 = n49252 ^ n17440 ^ n15575 ;
  assign n49254 = n30801 & ~n32589 ;
  assign n49261 = ( n3534 & n18442 ) | ( n3534 & ~n24802 ) | ( n18442 & ~n24802 ) ;
  assign n49259 = n14373 & ~n17592 ;
  assign n49260 = ~n24873 & n49259 ;
  assign n49262 = n49261 ^ n49260 ^ 1'b0 ;
  assign n49255 = n17661 ^ n11858 ^ n7630 ;
  assign n49256 = n4653 | n21773 ;
  assign n49257 = n49256 ^ n33417 ^ 1'b0 ;
  assign n49258 = ( n39720 & n49255 ) | ( n39720 & n49257 ) | ( n49255 & n49257 ) ;
  assign n49263 = n49262 ^ n49258 ^ 1'b0 ;
  assign n49264 = n6838 | n29180 ;
  assign n49265 = n49264 ^ n4741 ^ 1'b0 ;
  assign n49266 = n13221 | n44938 ;
  assign n49267 = ~n19798 & n35340 ;
  assign n49270 = ~n2357 & n8819 ;
  assign n49268 = n2267 & ~n19299 ;
  assign n49269 = n49268 ^ n2243 ^ 1'b0 ;
  assign n49271 = n49270 ^ n49269 ^ n5204 ;
  assign n49272 = ~n14630 & n23168 ;
  assign n49273 = ~n6769 & n49272 ;
  assign n49274 = n48872 & ~n49273 ;
  assign n49275 = ( n6598 & n10259 ) | ( n6598 & n41048 ) | ( n10259 & n41048 ) ;
  assign n49276 = n30306 ^ n3200 ^ 1'b0 ;
  assign n49277 = n34176 & ~n49276 ;
  assign n49278 = ~n7739 & n13438 ;
  assign n49279 = n49278 ^ n8666 ^ 1'b0 ;
  assign n49280 = n20964 & n23038 ;
  assign n49281 = ( ~n3196 & n35886 ) | ( ~n3196 & n37428 ) | ( n35886 & n37428 ) ;
  assign n49282 = n49281 ^ n40412 ^ n26878 ;
  assign n49283 = n46036 ^ n36633 ^ n8290 ;
  assign n49284 = ( n4463 & ~n30170 ) | ( n4463 & n35946 ) | ( ~n30170 & n35946 ) ;
  assign n49285 = ( n11512 & ~n13238 ) | ( n11512 & n15323 ) | ( ~n13238 & n15323 ) ;
  assign n49286 = ( n24193 & ~n40013 ) | ( n24193 & n49285 ) | ( ~n40013 & n49285 ) ;
  assign n49287 = n624 | n6825 ;
  assign n49288 = n49287 ^ n1003 ^ 1'b0 ;
  assign n49293 = n6765 & ~n18910 ;
  assign n49289 = n46772 ^ n46127 ^ n19600 ;
  assign n49290 = n29350 ^ n12361 ^ 1'b0 ;
  assign n49291 = n2771 | n49290 ;
  assign n49292 = ( n4965 & n49289 ) | ( n4965 & n49291 ) | ( n49289 & n49291 ) ;
  assign n49294 = n49293 ^ n49292 ^ n6796 ;
  assign n49295 = n49288 | n49294 ;
  assign n49296 = n32020 ^ n8701 ^ 1'b0 ;
  assign n49297 = n22668 & ~n49296 ;
  assign n49298 = n49297 ^ n26363 ^ 1'b0 ;
  assign n49299 = n21754 & n40940 ;
  assign n49300 = n49299 ^ n26174 ^ 1'b0 ;
  assign n49301 = n16512 ^ n2325 ^ 1'b0 ;
  assign n49302 = n39894 ^ n35756 ^ 1'b0 ;
  assign n49303 = n36858 & ~n49302 ;
  assign n49304 = n49301 & n49303 ;
  assign n49305 = ( x62 & ~n10433 ) | ( x62 & n19359 ) | ( ~n10433 & n19359 ) ;
  assign n49306 = ( n34665 & ~n36242 ) | ( n34665 & n49305 ) | ( ~n36242 & n49305 ) ;
  assign n49307 = ( n16233 & ~n42783 ) | ( n16233 & n45965 ) | ( ~n42783 & n45965 ) ;
  assign n49308 = n30777 ^ n25424 ^ n2309 ;
  assign n49309 = n6688 | n15087 ;
  assign n49310 = n12196 ^ n4294 ^ 1'b0 ;
  assign n49311 = ~n42931 & n49310 ;
  assign n49312 = n3593 & ~n16677 ;
  assign n49313 = n49312 ^ n26090 ^ 1'b0 ;
  assign n49314 = n23127 ^ n10055 ^ 1'b0 ;
  assign n49315 = n49313 & n49314 ;
  assign n49316 = ~n19489 & n27174 ;
  assign n49317 = ~n23994 & n49316 ;
  assign n49318 = n6616 & ~n14991 ;
  assign n49319 = ~n26140 & n49318 ;
  assign n49323 = n16961 ^ n13274 ^ n2451 ;
  assign n49320 = n8718 | n20109 ;
  assign n49321 = n49320 ^ n914 ^ 1'b0 ;
  assign n49322 = n49321 ^ n7080 ^ 1'b0 ;
  assign n49324 = n49323 ^ n49322 ^ n12982 ;
  assign n49325 = ( n8917 & n23576 ) | ( n8917 & ~n31020 ) | ( n23576 & ~n31020 ) ;
  assign n49326 = ( ~n44736 & n48296 ) | ( ~n44736 & n49325 ) | ( n48296 & n49325 ) ;
  assign n49329 = n1760 & n3717 ;
  assign n49330 = n49329 ^ n2391 ^ 1'b0 ;
  assign n49327 = n9667 & ~n13552 ;
  assign n49328 = n49327 ^ n1588 ^ 1'b0 ;
  assign n49331 = n49330 ^ n49328 ^ 1'b0 ;
  assign n49332 = ~n5548 & n30476 ;
  assign n49333 = ~n49331 & n49332 ;
  assign n49334 = n49333 ^ n38666 ^ 1'b0 ;
  assign n49335 = n28694 ^ n27886 ^ n15859 ;
  assign n49336 = n28430 ^ n15700 ^ n4990 ;
  assign n49337 = ~n26129 & n32993 ;
  assign n49338 = n34637 & n49337 ;
  assign n49339 = n49336 | n49338 ;
  assign n49340 = n13674 & ~n32368 ;
  assign n49341 = n9620 & n49340 ;
  assign n49342 = ~n8218 & n25789 ;
  assign n49343 = ~n6246 & n49342 ;
  assign n49344 = n5497 & ~n49343 ;
  assign n49345 = n39101 ^ n3959 ^ 1'b0 ;
  assign n49346 = n47878 ^ n34387 ^ n30625 ;
  assign n49347 = n6903 | n7063 ;
  assign n49348 = n16682 ^ n3178 ^ 1'b0 ;
  assign n49349 = n49348 ^ n24461 ^ n880 ;
  assign n49350 = ( n5265 & n13537 ) | ( n5265 & ~n42709 ) | ( n13537 & ~n42709 ) ;
  assign n49351 = n37395 ^ n15767 ^ 1'b0 ;
  assign n49352 = n2104 & n49351 ;
  assign n49353 = n49352 ^ n25114 ^ n11689 ;
  assign n49354 = n14649 | n49353 ;
  assign n49355 = n30336 ^ n5197 ^ 1'b0 ;
  assign n49356 = n18157 ^ n15566 ^ n13869 ;
  assign n49357 = n16944 ^ n4020 ^ n1478 ;
  assign n49358 = n9947 ^ n6998 ^ 1'b0 ;
  assign n49359 = n49357 & n49358 ;
  assign n49360 = n49359 ^ n39573 ^ 1'b0 ;
  assign n49361 = n3790 & ~n49360 ;
  assign n49362 = n49361 ^ n41208 ^ n17658 ;
  assign n49363 = ( n16250 & n24776 ) | ( n16250 & n35461 ) | ( n24776 & n35461 ) ;
  assign n49364 = n44013 ^ n40165 ^ n35442 ;
  assign n49365 = n31613 ^ n28518 ^ 1'b0 ;
  assign n49366 = ( ~n30671 & n46214 ) | ( ~n30671 & n49365 ) | ( n46214 & n49365 ) ;
  assign n49368 = ( n857 & n1961 ) | ( n857 & n6486 ) | ( n1961 & n6486 ) ;
  assign n49367 = ~n10896 & n13473 ;
  assign n49369 = n49368 ^ n49367 ^ 1'b0 ;
  assign n49370 = ~n15650 & n49369 ;
  assign n49371 = n7359 | n14649 ;
  assign n49372 = n49371 ^ n2597 ^ 1'b0 ;
  assign n49374 = n9625 ^ n4723 ^ 1'b0 ;
  assign n49373 = n22121 & n34998 ;
  assign n49375 = n49374 ^ n49373 ^ 1'b0 ;
  assign n49380 = n29839 ^ n10625 ^ 1'b0 ;
  assign n49381 = n10526 & n49380 ;
  assign n49382 = n49381 ^ n30607 ^ 1'b0 ;
  assign n49376 = ( n8589 & n12990 ) | ( n8589 & ~n25585 ) | ( n12990 & ~n25585 ) ;
  assign n49377 = n8790 & n17807 ;
  assign n49378 = ( n44515 & n49376 ) | ( n44515 & n49377 ) | ( n49376 & n49377 ) ;
  assign n49379 = ~n46283 & n49378 ;
  assign n49383 = n49382 ^ n49379 ^ 1'b0 ;
  assign n49384 = ( n9698 & n24442 ) | ( n9698 & ~n49383 ) | ( n24442 & ~n49383 ) ;
  assign n49385 = n32458 ^ n7186 ^ 1'b0 ;
  assign n49386 = n43869 ^ n1155 ^ 1'b0 ;
  assign n49387 = ( n33587 & n39649 ) | ( n33587 & ~n49386 ) | ( n39649 & ~n49386 ) ;
  assign n49388 = ~n14485 & n14891 ;
  assign n49389 = n31902 ^ n25162 ^ n18973 ;
  assign n49390 = ( n19336 & ~n38604 ) | ( n19336 & n49389 ) | ( ~n38604 & n49389 ) ;
  assign n49391 = n1885 & n17785 ;
  assign n49392 = n27310 & n49391 ;
  assign n49393 = n49392 ^ n25875 ^ 1'b0 ;
  assign n49394 = ( n49388 & ~n49390 ) | ( n49388 & n49393 ) | ( ~n49390 & n49393 ) ;
  assign n49395 = ( n11642 & ~n25160 ) | ( n11642 & n26636 ) | ( ~n25160 & n26636 ) ;
  assign n49396 = n26310 & n35010 ;
  assign n49397 = n474 & ~n23329 ;
  assign n49398 = n49397 ^ n10753 ^ 1'b0 ;
  assign n49399 = ~n9214 & n43389 ;
  assign n49400 = n49399 ^ n5346 ^ 1'b0 ;
  assign n49401 = ~n17983 & n25203 ;
  assign n49402 = n35276 | n49401 ;
  assign n49403 = n8750 & n22985 ;
  assign n49404 = n32754 ^ n18320 ^ 1'b0 ;
  assign n49405 = n1589 & ~n2530 ;
  assign n49406 = n49405 ^ n23617 ^ 1'b0 ;
  assign n49407 = n49406 ^ n10937 ^ 1'b0 ;
  assign n49408 = ( ~n49403 & n49404 ) | ( ~n49403 & n49407 ) | ( n49404 & n49407 ) ;
  assign n49409 = n2030 | n40912 ;
  assign n49410 = n49409 ^ n45293 ^ n3520 ;
  assign n49411 = ~n1828 & n20480 ;
  assign n49412 = n49411 ^ n9711 ^ 1'b0 ;
  assign n49413 = n49412 ^ n27105 ^ n9921 ;
  assign n49414 = n34437 ^ n28767 ^ n16282 ;
  assign n49415 = n11353 | n16118 ;
  assign n49416 = n10835 ^ n6017 ^ 1'b0 ;
  assign n49417 = n9373 & n49416 ;
  assign n49418 = n17809 | n30456 ;
  assign n49419 = n49417 | n49418 ;
  assign n49420 = n2804 | n39592 ;
  assign n49421 = n7077 & ~n49420 ;
  assign n49422 = n49421 ^ n11422 ^ 1'b0 ;
  assign n49423 = n19735 | n46159 ;
  assign n49424 = n20325 ^ n5183 ^ 1'b0 ;
  assign n49425 = ~n49423 & n49424 ;
  assign n49426 = n8819 | n43771 ;
  assign n49427 = n49426 ^ n30134 ^ 1'b0 ;
  assign n49428 = n34408 ^ n32273 ^ n16019 ;
  assign n49429 = n35746 ^ n31268 ^ n14288 ;
  assign n49430 = n49429 ^ n35523 ^ n25961 ;
  assign n49431 = n22184 ^ n18072 ^ n3269 ;
  assign n49432 = n37322 ^ n8482 ^ 1'b0 ;
  assign n49433 = n44904 & n49432 ;
  assign n49434 = n49433 ^ n45029 ^ n25318 ;
  assign n49435 = n13440 | n32229 ;
  assign n49436 = n11492 & ~n49435 ;
  assign n49437 = n40825 ^ n26925 ^ n24013 ;
  assign n49438 = n18798 | n48945 ;
  assign n49439 = n6793 ^ n4494 ^ 1'b0 ;
  assign n49440 = n26154 ^ n21215 ^ x29 ;
  assign n49441 = n49440 ^ n22502 ^ n6015 ;
  assign n49442 = ~n17983 & n23399 ;
  assign n49443 = ~n49441 & n49442 ;
  assign n49444 = n13438 & n19083 ;
  assign n49445 = n13804 & ~n26433 ;
  assign n49447 = ~n6301 & n11223 ;
  assign n49446 = n29094 & ~n38811 ;
  assign n49448 = n49447 ^ n49446 ^ 1'b0 ;
  assign n49449 = ( ~n1598 & n13374 ) | ( ~n1598 & n29740 ) | ( n13374 & n29740 ) ;
  assign n49450 = n25030 ^ n13134 ^ n8380 ;
  assign n49451 = ( n8177 & ~n15694 ) | ( n8177 & n16928 ) | ( ~n15694 & n16928 ) ;
  assign n49452 = ( n8191 & n17076 ) | ( n8191 & n49451 ) | ( n17076 & n49451 ) ;
  assign n49453 = ( n32069 & n40298 ) | ( n32069 & ~n41892 ) | ( n40298 & ~n41892 ) ;
  assign n49454 = ~n5755 & n49453 ;
  assign n49455 = n49454 ^ n33232 ^ 1'b0 ;
  assign n49456 = n49455 ^ n31570 ^ x227 ;
  assign n49457 = n16225 & ~n49456 ;
  assign n49458 = n33000 ^ n31067 ^ 1'b0 ;
  assign n49459 = n6237 | n49458 ;
  assign n49460 = n49459 ^ n6560 ^ x216 ;
  assign n49461 = ~n1022 & n11917 ;
  assign n49462 = ~n49460 & n49461 ;
  assign n49463 = n49462 ^ n14465 ^ 1'b0 ;
  assign n49464 = n8083 | n31983 ;
  assign n49465 = n49464 ^ n7407 ^ 1'b0 ;
  assign n49466 = n8182 ^ n5022 ^ 1'b0 ;
  assign n49467 = n17496 & n49466 ;
  assign n49468 = n39050 ^ n36207 ^ 1'b0 ;
  assign n49469 = n35760 & ~n49468 ;
  assign n49470 = ~n21476 & n24484 ;
  assign n49471 = ( n26228 & n42039 ) | ( n26228 & n49234 ) | ( n42039 & n49234 ) ;
  assign n49472 = n38536 ^ n30483 ^ n17547 ;
  assign n49473 = n20408 ^ n7798 ^ n1572 ;
  assign n49474 = n49473 ^ n40908 ^ n9761 ;
  assign n49475 = n32283 ^ n2945 ^ 1'b0 ;
  assign n49476 = n675 & n49475 ;
  assign n49477 = n21093 & ~n49476 ;
  assign n49478 = ( n8864 & n11343 ) | ( n8864 & ~n49477 ) | ( n11343 & ~n49477 ) ;
  assign n49479 = n49478 ^ n10735 ^ 1'b0 ;
  assign n49481 = n28160 ^ n20551 ^ 1'b0 ;
  assign n49480 = n10565 & n42612 ;
  assign n49482 = n49481 ^ n49480 ^ 1'b0 ;
  assign n49483 = n2475 | n42301 ;
  assign n49484 = ( ~n5772 & n21133 ) | ( ~n5772 & n21887 ) | ( n21133 & n21887 ) ;
  assign n49485 = n48103 & n49484 ;
  assign n49486 = n10244 & ~n44665 ;
  assign n49487 = ( n6616 & n21542 ) | ( n6616 & ~n49486 ) | ( n21542 & ~n49486 ) ;
  assign n49488 = n2132 & n38597 ;
  assign n49489 = n49488 ^ n5815 ^ n5653 ;
  assign n49490 = n14443 ^ n10336 ^ n8966 ;
  assign n49491 = n49490 ^ n34882 ^ n7868 ;
  assign n49492 = n8111 & ~n45208 ;
  assign n49493 = n49492 ^ n8721 ^ 1'b0 ;
  assign n49494 = n13484 & n49493 ;
  assign n49495 = n3709 & ~n24181 ;
  assign n49496 = n49495 ^ n18502 ^ 1'b0 ;
  assign n49497 = n49496 ^ n11493 ^ 1'b0 ;
  assign n49499 = n15202 ^ n11063 ^ 1'b0 ;
  assign n49500 = n12873 & n49499 ;
  assign n49498 = ( n34538 & ~n37196 ) | ( n34538 & n49194 ) | ( ~n37196 & n49194 ) ;
  assign n49501 = n49500 ^ n49498 ^ n23735 ;
  assign n49502 = ( n16119 & ~n49497 ) | ( n16119 & n49501 ) | ( ~n49497 & n49501 ) ;
  assign n49503 = ~n3050 & n15864 ;
  assign n49504 = n33010 & n49503 ;
  assign n49505 = ( n7128 & n49502 ) | ( n7128 & ~n49504 ) | ( n49502 & ~n49504 ) ;
  assign n49506 = n46673 ^ n24898 ^ n8612 ;
  assign n49507 = n39133 ^ n12321 ^ 1'b0 ;
  assign n49508 = n20010 ^ n11305 ^ n2773 ;
  assign n49509 = n40105 ^ n31457 ^ 1'b0 ;
  assign n49510 = n49508 | n49509 ;
  assign n49511 = n4249 & n4733 ;
  assign n49512 = n26285 | n49511 ;
  assign n49513 = n49510 & ~n49512 ;
  assign n49514 = n20192 | n21668 ;
  assign n49515 = n21421 | n49514 ;
  assign n49516 = n32067 ^ n29570 ^ n26733 ;
  assign n49517 = n31654 & n49516 ;
  assign n49518 = ( n1534 & n7646 ) | ( n1534 & n25187 ) | ( n7646 & n25187 ) ;
  assign n49519 = ( n10415 & n27759 ) | ( n10415 & ~n49518 ) | ( n27759 & ~n49518 ) ;
  assign n49520 = ( n1548 & n5715 ) | ( n1548 & ~n14870 ) | ( n5715 & ~n14870 ) ;
  assign n49521 = ~n1427 & n8966 ;
  assign n49522 = n9406 & ~n18823 ;
  assign n49523 = n49522 ^ n9242 ^ 1'b0 ;
  assign n49524 = n40675 ^ n6250 ^ n5242 ;
  assign n49525 = ( ~n17205 & n49523 ) | ( ~n17205 & n49524 ) | ( n49523 & n49524 ) ;
  assign n49526 = n43738 ^ n41207 ^ 1'b0 ;
  assign n49527 = n9814 ^ x46 ^ 1'b0 ;
  assign n49528 = n49526 & n49527 ;
  assign n49529 = ~n21911 & n35617 ;
  assign n49530 = n4837 & n22962 ;
  assign n49531 = ( ~n36717 & n41109 ) | ( ~n36717 & n49530 ) | ( n41109 & n49530 ) ;
  assign n49532 = n3588 | n25943 ;
  assign n49533 = n49532 ^ n26486 ^ 1'b0 ;
  assign n49534 = n49533 ^ n47544 ^ n46512 ;
  assign n49535 = n44010 ^ n38757 ^ n5733 ;
  assign n49536 = ( ~n684 & n44996 ) | ( ~n684 & n47868 ) | ( n44996 & n47868 ) ;
  assign n49537 = n49536 ^ n32956 ^ n18912 ;
  assign n49538 = n3068 & n23503 ;
  assign n49539 = n49538 ^ n29983 ^ n1553 ;
  assign n49540 = n49539 ^ n21170 ^ n6990 ;
  assign n49541 = ~n1461 & n3636 ;
  assign n49542 = ~n21446 & n49541 ;
  assign n49543 = ( n15700 & n22570 ) | ( n15700 & n26039 ) | ( n22570 & n26039 ) ;
  assign n49544 = n3885 | n49543 ;
  assign n49545 = n49544 ^ n20473 ^ 1'b0 ;
  assign n49546 = n33511 | n49471 ;
  assign n49547 = n47301 ^ n33540 ^ 1'b0 ;
  assign n49548 = n45898 & ~n49547 ;
  assign n49549 = ( n3199 & n30206 ) | ( n3199 & n31937 ) | ( n30206 & n31937 ) ;
  assign n49552 = ~n8171 & n30957 ;
  assign n49550 = ~n7301 & n47701 ;
  assign n49551 = n49550 ^ n3248 ^ 1'b0 ;
  assign n49553 = n49552 ^ n49551 ^ n31811 ;
  assign n49554 = ( ~n4746 & n34778 ) | ( ~n4746 & n46442 ) | ( n34778 & n46442 ) ;
  assign n49555 = ( n12544 & ~n29548 ) | ( n12544 & n39068 ) | ( ~n29548 & n39068 ) ;
  assign n49556 = n49376 ^ n21669 ^ 1'b0 ;
  assign n49557 = n36082 ^ n30034 ^ n14259 ;
  assign n49558 = ( n1881 & n9192 ) | ( n1881 & n13500 ) | ( n9192 & n13500 ) ;
  assign n49559 = n2387 & n13161 ;
  assign n49560 = ~n49558 & n49559 ;
  assign n49561 = ~n3740 & n22428 ;
  assign n49562 = n49561 ^ n18651 ^ 1'b0 ;
  assign n49563 = ( n4194 & n5387 ) | ( n4194 & ~n6396 ) | ( n5387 & ~n6396 ) ;
  assign n49564 = ( ~n10918 & n18087 ) | ( ~n10918 & n49563 ) | ( n18087 & n49563 ) ;
  assign n49565 = n49564 ^ n26077 ^ 1'b0 ;
  assign n49566 = n9433 & ~n25792 ;
  assign n49567 = n5836 & n49566 ;
  assign n49568 = n49567 ^ n20656 ^ n20512 ;
  assign n49570 = n26133 ^ n11436 ^ n6683 ;
  assign n49569 = n24434 ^ n2718 ^ 1'b0 ;
  assign n49571 = n49570 ^ n49569 ^ n24859 ;
  assign n49572 = ( n13122 & n18818 ) | ( n13122 & n22604 ) | ( n18818 & n22604 ) ;
  assign n49573 = ( n3011 & n4475 ) | ( n3011 & n4582 ) | ( n4475 & n4582 ) ;
  assign n49574 = n49573 ^ n22951 ^ n887 ;
  assign n49575 = n49574 ^ n41997 ^ n3596 ;
  assign n49576 = n9622 ^ n9595 ^ 1'b0 ;
  assign n49577 = n9584 & n49576 ;
  assign n49578 = ( n1508 & n6726 ) | ( n1508 & n49577 ) | ( n6726 & n49577 ) ;
  assign n49579 = ( n26424 & ~n44186 ) | ( n26424 & n47026 ) | ( ~n44186 & n47026 ) ;
  assign n49580 = n49579 ^ n29745 ^ n13195 ;
  assign n49581 = n49580 ^ n38330 ^ 1'b0 ;
  assign n49582 = n36365 & n49581 ;
  assign n49583 = n41011 ^ n3615 ^ 1'b0 ;
  assign n49584 = ~n1150 & n49583 ;
  assign n49586 = ~n3937 & n37021 ;
  assign n49585 = n18310 & ~n20942 ;
  assign n49587 = n49586 ^ n49585 ^ 1'b0 ;
  assign n49588 = ( n2150 & n10665 ) | ( n2150 & ~n30245 ) | ( n10665 & ~n30245 ) ;
  assign n49589 = ( ~n7806 & n27443 ) | ( ~n7806 & n49588 ) | ( n27443 & n49588 ) ;
  assign n49590 = ( n20886 & n31055 ) | ( n20886 & ~n49589 ) | ( n31055 & ~n49589 ) ;
  assign n49592 = n18430 ^ n9126 ^ n1930 ;
  assign n49591 = ~n24058 & n33459 ;
  assign n49593 = n49592 ^ n49591 ^ 1'b0 ;
  assign n49594 = ( n26339 & n46796 ) | ( n26339 & ~n49593 ) | ( n46796 & ~n49593 ) ;
  assign n49596 = ( x119 & ~n4067 ) | ( x119 & n28462 ) | ( ~n4067 & n28462 ) ;
  assign n49595 = n17843 ^ n1573 ^ 1'b0 ;
  assign n49597 = n49596 ^ n49595 ^ n22032 ;
  assign n49598 = ( n16321 & ~n17650 ) | ( n16321 & n21582 ) | ( ~n17650 & n21582 ) ;
  assign n49599 = n49598 ^ n13469 ^ n5164 ;
  assign n49600 = n44838 ^ n3425 ^ 1'b0 ;
  assign n49601 = n19697 | n49600 ;
  assign n49602 = n10238 | n44510 ;
  assign n49603 = n49602 ^ n44321 ^ 1'b0 ;
  assign n49609 = n4938 & ~n15151 ;
  assign n49610 = ~n11559 & n49609 ;
  assign n49604 = n27305 ^ n24003 ^ n1834 ;
  assign n49605 = ( ~n24008 & n27140 ) | ( ~n24008 & n49604 ) | ( n27140 & n49604 ) ;
  assign n49606 = n7514 | n49605 ;
  assign n49607 = n9338 | n49606 ;
  assign n49608 = n7566 & n49607 ;
  assign n49611 = n49610 ^ n49608 ^ 1'b0 ;
  assign n49612 = ( n13149 & n49603 ) | ( n13149 & n49611 ) | ( n49603 & n49611 ) ;
  assign n49613 = n10926 & ~n45395 ;
  assign n49614 = n12218 ^ n8163 ^ 1'b0 ;
  assign n49615 = ~n21795 & n49614 ;
  assign n49616 = ( n24493 & n28155 ) | ( n24493 & n49615 ) | ( n28155 & n49615 ) ;
  assign n49617 = n16267 ^ n1412 ^ 1'b0 ;
  assign n49618 = n3814 & ~n8563 ;
  assign n49619 = ~n9212 & n49618 ;
  assign n49620 = n8999 | n10676 ;
  assign n49621 = n13799 & n49620 ;
  assign n49622 = n49619 & n49621 ;
  assign n49623 = n49622 ^ n25499 ^ 1'b0 ;
  assign n49624 = n42033 ^ n5645 ^ 1'b0 ;
  assign n49625 = ~n17433 & n49624 ;
  assign n49626 = ( ~n6162 & n16255 ) | ( ~n6162 & n49625 ) | ( n16255 & n49625 ) ;
  assign n49627 = n3620 | n12605 ;
  assign n49628 = n49627 ^ n7362 ^ 1'b0 ;
  assign n49629 = n38250 ^ n21572 ^ 1'b0 ;
  assign n49630 = n8672 & n49629 ;
  assign n49631 = n12534 & ~n39162 ;
  assign n49632 = ~n12237 & n49631 ;
  assign n49633 = n47042 ^ n13099 ^ 1'b0 ;
  assign n49634 = n1145 | n42388 ;
  assign n49635 = ~n12930 & n26253 ;
  assign n49636 = ~n49634 & n49635 ;
  assign n49637 = n31160 & n34619 ;
  assign n49638 = ( ~n10567 & n42910 ) | ( ~n10567 & n49637 ) | ( n42910 & n49637 ) ;
  assign n49639 = n12607 ^ n8354 ^ n5543 ;
  assign n49640 = n11633 ^ n8604 ^ 1'b0 ;
  assign n49642 = x86 & ~n14101 ;
  assign n49643 = n49642 ^ n15225 ^ 1'b0 ;
  assign n49641 = n32679 ^ n22922 ^ n2787 ;
  assign n49644 = n49643 ^ n49641 ^ n19080 ;
  assign n49646 = x240 & n22003 ;
  assign n49647 = n49646 ^ n9742 ^ 1'b0 ;
  assign n49645 = n567 & ~n7022 ;
  assign n49648 = n49647 ^ n49645 ^ 1'b0 ;
  assign n49649 = n2680 & n36851 ;
  assign n49650 = n19067 ^ n16645 ^ n3179 ;
  assign n49651 = ( x180 & n1614 ) | ( x180 & ~n25776 ) | ( n1614 & ~n25776 ) ;
  assign n49652 = n49651 ^ n16905 ^ n6521 ;
  assign n49653 = ( n12890 & n43522 ) | ( n12890 & n49652 ) | ( n43522 & n49652 ) ;
  assign n49654 = n32777 ^ n31071 ^ n7795 ;
  assign n49655 = n39843 ^ n8458 ^ 1'b0 ;
  assign n49656 = ~n1162 & n49655 ;
  assign n49657 = n24026 | n49656 ;
  assign n49658 = n45877 | n49657 ;
  assign n49659 = ( n1749 & ~n22970 ) | ( n1749 & n49658 ) | ( ~n22970 & n49658 ) ;
  assign n49660 = n31966 ^ n30692 ^ 1'b0 ;
  assign n49661 = n25403 | n32580 ;
  assign n49662 = n18193 | n49661 ;
  assign n49663 = n49662 ^ n34619 ^ n5598 ;
  assign n49664 = n49331 ^ n35023 ^ 1'b0 ;
  assign n49665 = n10185 | n49664 ;
  assign n49666 = n21610 ^ n14042 ^ n11386 ;
  assign n49667 = n19056 ^ n6131 ^ 1'b0 ;
  assign n49668 = n49666 | n49667 ;
  assign n49669 = ~n6479 & n19342 ;
  assign n49670 = ~n19342 & n49669 ;
  assign n49671 = n29320 ^ n21295 ^ n17826 ;
  assign n49672 = ( n43411 & ~n49670 ) | ( n43411 & n49671 ) | ( ~n49670 & n49671 ) ;
  assign n49673 = n49672 ^ n24253 ^ n16242 ;
  assign n49674 = n25884 ^ n7805 ^ 1'b0 ;
  assign n49675 = n11572 & n49674 ;
  assign n49676 = n47214 | n49675 ;
  assign n49677 = n17908 ^ n6864 ^ 1'b0 ;
  assign n49678 = n23168 & n49677 ;
  assign n49679 = ( n6522 & n45221 ) | ( n6522 & ~n49678 ) | ( n45221 & ~n49678 ) ;
  assign n49680 = ~n4789 & n49679 ;
  assign n49681 = n36946 ^ n13851 ^ 1'b0 ;
  assign n49682 = ( n25468 & ~n30271 ) | ( n25468 & n33767 ) | ( ~n30271 & n33767 ) ;
  assign n49683 = n9288 & ~n26997 ;
  assign n49684 = n22853 & n42988 ;
  assign n49685 = n3679 & n35823 ;
  assign n49686 = ~n24588 & n25684 ;
  assign n49687 = ~n5917 & n49686 ;
  assign n49688 = ~n1894 & n18359 ;
  assign n49689 = ~n19627 & n23918 ;
  assign n49690 = ~n18309 & n49689 ;
  assign n49691 = n9980 ^ n4038 ^ 1'b0 ;
  assign n49692 = ( n592 & n49690 ) | ( n592 & n49691 ) | ( n49690 & n49691 ) ;
  assign n49693 = n39137 ^ n4630 ^ 1'b0 ;
  assign n49694 = n48268 ^ n4819 ^ 1'b0 ;
  assign n49695 = n45785 ^ n3256 ^ x31 ;
  assign n49696 = ( n8943 & n49694 ) | ( n8943 & ~n49695 ) | ( n49694 & ~n49695 ) ;
  assign n49697 = n49696 ^ n45101 ^ n32389 ;
  assign n49698 = ( n26346 & ~n27231 ) | ( n26346 & n47542 ) | ( ~n27231 & n47542 ) ;
  assign n49699 = n49698 ^ n2584 ^ 1'b0 ;
  assign n49700 = ~n6334 & n49699 ;
  assign n49701 = n29232 ^ n24946 ^ n6982 ;
  assign n49702 = ~n547 & n23041 ;
  assign n49703 = ~n49701 & n49702 ;
  assign n49704 = n17237 ^ n3196 ^ 1'b0 ;
  assign n49705 = n24239 & n49704 ;
  assign n49706 = n2226 & n49705 ;
  assign n49707 = ~n40216 & n49706 ;
  assign n49708 = ( n10261 & ~n10277 ) | ( n10261 & n21326 ) | ( ~n10277 & n21326 ) ;
  assign n49709 = n34718 ^ n32653 ^ n11259 ;
  assign n49710 = n26561 ^ n23615 ^ n15854 ;
  assign n49711 = n37752 | n49710 ;
  assign n49712 = n15180 ^ n12661 ^ n5504 ;
  assign n49715 = n10305 | n21455 ;
  assign n49716 = n13057 & n49715 ;
  assign n49717 = n49716 ^ n44010 ^ 1'b0 ;
  assign n49713 = n27171 ^ n2603 ^ 1'b0 ;
  assign n49714 = n41461 & ~n49713 ;
  assign n49718 = n49717 ^ n49714 ^ n36926 ;
  assign n49719 = n4865 | n7138 ;
  assign n49720 = n29699 & ~n49719 ;
  assign n49721 = n9643 ^ n1688 ^ 1'b0 ;
  assign n49722 = ~n49720 & n49721 ;
  assign n49723 = n49508 ^ x102 ^ 1'b0 ;
  assign n49724 = n3411 | n4334 ;
  assign n49725 = n11858 ^ n1028 ^ 1'b0 ;
  assign n49726 = n49724 | n49725 ;
  assign n49727 = n27810 ^ n10138 ^ 1'b0 ;
  assign n49728 = n11876 | n49727 ;
  assign n49729 = n582 & ~n43211 ;
  assign n49730 = n22638 & ~n24144 ;
  assign n49731 = n49730 ^ n23120 ^ n18374 ;
  assign n49732 = n49731 ^ n39318 ^ n11885 ;
  assign n49733 = n46241 ^ n34614 ^ 1'b0 ;
  assign n49737 = n19117 ^ n15551 ^ n4844 ;
  assign n49738 = ( n6357 & n27434 ) | ( n6357 & n49737 ) | ( n27434 & n49737 ) ;
  assign n49739 = ( n37353 & ~n42993 ) | ( n37353 & n49738 ) | ( ~n42993 & n49738 ) ;
  assign n49734 = ~n10219 & n10779 ;
  assign n49735 = n49734 ^ n14804 ^ 1'b0 ;
  assign n49736 = n49735 ^ n19369 ^ 1'b0 ;
  assign n49740 = n49739 ^ n49736 ^ n12753 ;
  assign n49741 = n28409 ^ n27316 ^ n16137 ;
  assign n49742 = ( ~n17352 & n30332 ) | ( ~n17352 & n49741 ) | ( n30332 & n49741 ) ;
  assign n49743 = n14222 ^ n5681 ^ 1'b0 ;
  assign n49744 = ~n12684 & n49743 ;
  assign n49745 = n11806 & n49744 ;
  assign n49746 = n49745 ^ n40458 ^ 1'b0 ;
  assign n49747 = n29674 ^ n2983 ^ 1'b0 ;
  assign n49748 = ( n36338 & n37262 ) | ( n36338 & n39156 ) | ( n37262 & n39156 ) ;
  assign n49749 = ( n2273 & n23633 ) | ( n2273 & ~n24374 ) | ( n23633 & ~n24374 ) ;
  assign n49750 = n46459 ^ n26032 ^ n9948 ;
  assign n49751 = ~n26275 & n39978 ;
  assign n49752 = n6040 ^ n1155 ^ 1'b0 ;
  assign n49753 = n22453 & ~n49752 ;
  assign n49754 = n33469 ^ n7285 ^ 1'b0 ;
  assign n49755 = n18759 ^ n399 ^ 1'b0 ;
  assign n49756 = n17164 | n49755 ;
  assign n49757 = n44653 ^ n475 ^ 1'b0 ;
  assign n49758 = n5213 & ~n32684 ;
  assign n49759 = ~n5994 & n49758 ;
  assign n49760 = n19714 | n49759 ;
  assign n49761 = ( n7990 & n49757 ) | ( n7990 & ~n49760 ) | ( n49757 & ~n49760 ) ;
  assign n49762 = ( ~n8753 & n24579 ) | ( ~n8753 & n34653 ) | ( n24579 & n34653 ) ;
  assign n49763 = ( n24112 & ~n48758 ) | ( n24112 & n49762 ) | ( ~n48758 & n49762 ) ;
  assign n49764 = n8356 & n10129 ;
  assign n49765 = ~n27500 & n49764 ;
  assign n49766 = ( ~n7061 & n27457 ) | ( ~n7061 & n49765 ) | ( n27457 & n49765 ) ;
  assign n49767 = n10916 & ~n18583 ;
  assign n49768 = n49767 ^ n10405 ^ 1'b0 ;
  assign n49769 = n49768 ^ n7774 ^ n5608 ;
  assign n49770 = n42780 ^ n42312 ^ n18883 ;
  assign n49771 = n7700 ^ n3400 ^ 1'b0 ;
  assign n49772 = n27548 & n49746 ;
  assign n49773 = n49772 ^ n40731 ^ 1'b0 ;
  assign n49774 = n46890 ^ n8743 ^ 1'b0 ;
  assign n49775 = n265 & ~n49774 ;
  assign n49776 = ~n18968 & n49775 ;
  assign n49777 = ~n3044 & n49776 ;
  assign n49778 = n17221 ^ n11842 ^ n8942 ;
  assign n49779 = x121 & n22662 ;
  assign n49780 = n49779 ^ n17947 ^ 1'b0 ;
  assign n49781 = ( n4471 & ~n34133 ) | ( n4471 & n49780 ) | ( ~n34133 & n49780 ) ;
  assign n49782 = ~n42626 & n49781 ;
  assign n49783 = n49778 & n49782 ;
  assign n49784 = n15772 ^ n12229 ^ 1'b0 ;
  assign n49785 = n3943 | n49784 ;
  assign n49786 = n20062 & ~n49785 ;
  assign n49787 = ( n26342 & n35338 ) | ( n26342 & n49786 ) | ( n35338 & n49786 ) ;
  assign n49788 = n37932 ^ n31330 ^ 1'b0 ;
  assign n49789 = n47794 ^ n16496 ^ 1'b0 ;
  assign n49790 = ~n6083 & n8478 ;
  assign n49791 = ~n17152 & n49790 ;
  assign n49792 = n49791 ^ n37095 ^ n28855 ;
  assign n49793 = ( n31756 & ~n49789 ) | ( n31756 & n49792 ) | ( ~n49789 & n49792 ) ;
  assign n49794 = n1785 ^ n547 ^ 1'b0 ;
  assign n49795 = n31077 ^ n17889 ^ n6388 ;
  assign n49796 = ( ~n7094 & n12623 ) | ( ~n7094 & n30874 ) | ( n12623 & n30874 ) ;
  assign n49797 = n23323 & ~n49796 ;
  assign n49798 = ~n48777 & n49797 ;
  assign n49799 = n49798 ^ n11013 ^ 1'b0 ;
  assign n49800 = n5437 & n49799 ;
  assign n49801 = n509 | n49800 ;
  assign n49802 = n47394 ^ n26738 ^ 1'b0 ;
  assign n49803 = n48211 & n49802 ;
  assign n49804 = n21910 & n44502 ;
  assign n49805 = n13345 | n24915 ;
  assign n49806 = n49805 ^ n19193 ^ n932 ;
  assign n49807 = n12873 & n49806 ;
  assign n49808 = n28888 | n44368 ;
  assign n49809 = n49808 ^ n12919 ^ 1'b0 ;
  assign n49811 = n8216 ^ n7658 ^ n6681 ;
  assign n49812 = ( n11490 & n26771 ) | ( n11490 & n49811 ) | ( n26771 & n49811 ) ;
  assign n49813 = n26033 & n49812 ;
  assign n49814 = n33046 & n49813 ;
  assign n49815 = n49814 ^ n26525 ^ 1'b0 ;
  assign n49810 = n9505 & ~n9998 ;
  assign n49816 = n49815 ^ n49810 ^ n34098 ;
  assign n49817 = n47869 ^ n28556 ^ n15302 ;
  assign n49818 = n20340 ^ n17798 ^ n13875 ;
  assign n49819 = n49818 ^ n34074 ^ n12829 ;
  assign n49820 = n49819 ^ n37984 ^ n18487 ;
  assign n49821 = n49820 ^ n15282 ^ n873 ;
  assign n49822 = ( n6701 & n24488 ) | ( n6701 & n49651 ) | ( n24488 & n49651 ) ;
  assign n49823 = ( n15083 & n22218 ) | ( n15083 & n49822 ) | ( n22218 & n49822 ) ;
  assign n49825 = n29446 ^ n12897 ^ n1105 ;
  assign n49824 = ( n15035 & ~n18763 ) | ( n15035 & n19158 ) | ( ~n18763 & n19158 ) ;
  assign n49826 = n49825 ^ n49824 ^ 1'b0 ;
  assign n49827 = n31937 & n46120 ;
  assign n49828 = n27953 & n49827 ;
  assign n49829 = ~n12945 & n14385 ;
  assign n49830 = ~n8915 & n49829 ;
  assign n49831 = ~n5380 & n37439 ;
  assign n49832 = n23700 ^ n18478 ^ 1'b0 ;
  assign n49833 = n49032 & n49832 ;
  assign n49834 = n20994 ^ n1152 ^ 1'b0 ;
  assign n49835 = n49833 | n49834 ;
  assign n49836 = n34592 ^ n16913 ^ 1'b0 ;
  assign n49837 = n14394 ^ n11304 ^ 1'b0 ;
  assign n49838 = n49837 ^ n27552 ^ n1681 ;
  assign n49839 = n49838 ^ n38966 ^ n3211 ;
  assign n49840 = n38475 ^ n10048 ^ 1'b0 ;
  assign n49841 = n6353 & ~n49840 ;
  assign n49842 = n49841 ^ n11499 ^ n8730 ;
  assign n49843 = n23660 ^ n19172 ^ n509 ;
  assign n49844 = ~n35891 & n49843 ;
  assign n49845 = n49844 ^ n17010 ^ 1'b0 ;
  assign n49846 = ( ~n1317 & n16839 ) | ( ~n1317 & n49845 ) | ( n16839 & n49845 ) ;
  assign n49847 = n36744 ^ n9331 ^ n6945 ;
  assign n49848 = ( ~n10945 & n30998 ) | ( ~n10945 & n49847 ) | ( n30998 & n49847 ) ;
  assign n49849 = n41470 ^ n36176 ^ 1'b0 ;
  assign n49850 = ( n13574 & n31932 ) | ( n13574 & n49849 ) | ( n31932 & n49849 ) ;
  assign n49851 = n35945 ^ n14700 ^ n1384 ;
  assign n49852 = n3024 | n43238 ;
  assign n49853 = n49851 & ~n49852 ;
  assign n49854 = n17130 | n44564 ;
  assign n49855 = n11220 & ~n48845 ;
  assign n49856 = n49855 ^ n26443 ^ n6862 ;
  assign n49857 = n42028 ^ n17372 ^ n1372 ;
  assign n49858 = ( ~n1969 & n2592 ) | ( ~n1969 & n26135 ) | ( n2592 & n26135 ) ;
  assign n49859 = n30937 ^ n30053 ^ n16347 ;
  assign n49860 = ~n18434 & n41785 ;
  assign n49861 = ~n19840 & n34300 ;
  assign n49862 = n49429 & n49861 ;
  assign n49863 = ~n6762 & n11730 ;
  assign n49864 = n49863 ^ n8780 ^ 1'b0 ;
  assign n49865 = n46398 ^ n28913 ^ 1'b0 ;
  assign n49866 = n37880 & ~n49865 ;
  assign n49867 = n29960 ^ n22529 ^ 1'b0 ;
  assign n49868 = n49866 & n49867 ;
  assign n49869 = n19897 | n29114 ;
  assign n49870 = n49869 ^ n5990 ^ 1'b0 ;
  assign n49871 = ( ~n22119 & n26415 ) | ( ~n22119 & n49870 ) | ( n26415 & n49870 ) ;
  assign n49872 = ( n10494 & n20529 ) | ( n10494 & ~n20915 ) | ( n20529 & ~n20915 ) ;
  assign n49873 = n17606 ^ n10980 ^ 1'b0 ;
  assign n49874 = n2267 & ~n49873 ;
  assign n49875 = n49874 ^ n21431 ^ n6829 ;
  assign n49876 = n7709 ^ n7401 ^ 1'b0 ;
  assign n49877 = n49876 ^ n15263 ^ n13865 ;
  assign n49878 = ( ~n437 & n8772 ) | ( ~n437 & n49877 ) | ( n8772 & n49877 ) ;
  assign n49879 = n41582 ^ n31895 ^ n1031 ;
  assign n49880 = n49879 ^ n22003 ^ n15414 ;
  assign n49881 = ( n7364 & n49878 ) | ( n7364 & n49880 ) | ( n49878 & n49880 ) ;
  assign n49882 = n49881 ^ n15953 ^ n7867 ;
  assign n49883 = ~n27104 & n44264 ;
  assign n49884 = n13843 & n49811 ;
  assign n49885 = n49883 & n49884 ;
  assign n49886 = n9219 | n22236 ;
  assign n49887 = n37554 | n49886 ;
  assign n49888 = n11582 | n14972 ;
  assign n49889 = n49888 ^ n34969 ^ 1'b0 ;
  assign n49890 = n49889 ^ n21409 ^ n17735 ;
  assign n49891 = ( n36703 & ~n42494 ) | ( n36703 & n49890 ) | ( ~n42494 & n49890 ) ;
  assign n49892 = n49891 ^ n26207 ^ 1'b0 ;
  assign n49893 = n47701 ^ n32288 ^ 1'b0 ;
  assign n49894 = x173 & ~n28469 ;
  assign n49895 = ~n25540 & n49894 ;
  assign n49896 = n49895 ^ n31369 ^ n23948 ;
  assign n49897 = n49896 ^ n34683 ^ n18167 ;
  assign n49898 = n49897 ^ n38160 ^ n27686 ;
  assign n49899 = n9694 ^ n8944 ^ 1'b0 ;
  assign n49900 = n31551 ^ n4245 ^ n4077 ;
  assign n49901 = n49900 ^ n24751 ^ 1'b0 ;
  assign n49902 = n14591 & n49901 ;
  assign n49903 = n16481 & n31185 ;
  assign n49904 = n49903 ^ n4122 ^ 1'b0 ;
  assign n49905 = n23452 ^ n10862 ^ n8067 ;
  assign n49906 = ( ~n49902 & n49904 ) | ( ~n49902 & n49905 ) | ( n49904 & n49905 ) ;
  assign n49907 = n23429 | n46111 ;
  assign n49908 = ( n7453 & n16667 ) | ( n7453 & ~n17770 ) | ( n16667 & ~n17770 ) ;
  assign n49909 = ( n19624 & ~n24656 ) | ( n19624 & n49908 ) | ( ~n24656 & n49908 ) ;
  assign n49910 = n30332 ^ n18235 ^ 1'b0 ;
  assign n49911 = n48266 | n49910 ;
  assign n49914 = n18147 ^ n14285 ^ n4038 ;
  assign n49912 = n8935 | n11183 ;
  assign n49913 = n24509 & ~n49912 ;
  assign n49915 = n49914 ^ n49913 ^ 1'b0 ;
  assign n49916 = n47899 ^ n8299 ^ 1'b0 ;
  assign n49917 = n45230 ^ n26056 ^ 1'b0 ;
  assign n49918 = n4848 | n49917 ;
  assign n49919 = ( ~n32098 & n49916 ) | ( ~n32098 & n49918 ) | ( n49916 & n49918 ) ;
  assign n49920 = n7174 & ~n48504 ;
  assign n49921 = n49920 ^ n16935 ^ n5720 ;
  assign n49922 = ( n14049 & n28149 ) | ( n14049 & ~n48248 ) | ( n28149 & ~n48248 ) ;
  assign n49923 = ( n5725 & n16892 ) | ( n5725 & ~n26431 ) | ( n16892 & ~n26431 ) ;
  assign n49924 = ( n15066 & ~n49922 ) | ( n15066 & n49923 ) | ( ~n49922 & n49923 ) ;
  assign n49931 = n42288 ^ n31815 ^ 1'b0 ;
  assign n49932 = n49931 ^ n3339 ^ n918 ;
  assign n49933 = n49932 ^ n37760 ^ n5549 ;
  assign n49934 = n21028 | n49933 ;
  assign n49927 = n27337 & n40583 ;
  assign n49926 = n12604 & n26975 ;
  assign n49928 = n49927 ^ n49926 ^ 1'b0 ;
  assign n49925 = ( ~n16286 & n42637 ) | ( ~n16286 & n47701 ) | ( n42637 & n47701 ) ;
  assign n49929 = n49928 ^ n49925 ^ n5809 ;
  assign n49930 = n49929 ^ n36101 ^ n32803 ;
  assign n49935 = n49934 ^ n49930 ^ n20990 ;
  assign n49936 = ( n26241 & n35348 ) | ( n26241 & ~n49935 ) | ( n35348 & ~n49935 ) ;
  assign n49937 = ( x225 & ~n4636 ) | ( x225 & n5643 ) | ( ~n4636 & n5643 ) ;
  assign n49938 = n49937 ^ n7470 ^ 1'b0 ;
  assign n49939 = n17479 | n21234 ;
  assign n49940 = ~n17696 & n31043 ;
  assign n49942 = ( ~n1885 & n15833 ) | ( ~n1885 & n27894 ) | ( n15833 & n27894 ) ;
  assign n49941 = n37642 & n43687 ;
  assign n49943 = n49942 ^ n49941 ^ 1'b0 ;
  assign n49944 = n37004 ^ n34946 ^ 1'b0 ;
  assign n49945 = x205 & ~n40158 ;
  assign n49946 = ( ~n13216 & n38838 ) | ( ~n13216 & n49945 ) | ( n38838 & n49945 ) ;
  assign n49947 = ( x132 & n17935 ) | ( x132 & ~n49946 ) | ( n17935 & ~n49946 ) ;
  assign n49948 = ( n9132 & ~n14051 ) | ( n9132 & n33176 ) | ( ~n14051 & n33176 ) ;
  assign n49949 = n47868 ^ n16578 ^ n8772 ;
  assign n49950 = ( ~n46441 & n49948 ) | ( ~n46441 & n49949 ) | ( n49948 & n49949 ) ;
  assign n49951 = n48493 ^ n47730 ^ n15442 ;
  assign n49952 = n46012 ^ n3684 ^ 1'b0 ;
  assign n49953 = n15259 | n18022 ;
  assign n49954 = n1940 | n49953 ;
  assign n49955 = n49954 ^ n20015 ^ n2300 ;
  assign n49956 = n7421 & n45563 ;
  assign n49957 = n10679 & ~n49956 ;
  assign n49958 = n37957 ^ n6410 ^ 1'b0 ;
  assign n49959 = n10941 ^ n10033 ^ 1'b0 ;
  assign n49960 = ~n49958 & n49959 ;
  assign n49961 = n33354 ^ n12566 ^ 1'b0 ;
  assign n49962 = ~n5623 & n49961 ;
  assign n49963 = x100 & n18229 ;
  assign n49964 = ~n11341 & n49963 ;
  assign n49965 = ( n2976 & ~n8689 ) | ( n2976 & n23100 ) | ( ~n8689 & n23100 ) ;
  assign n49966 = n12740 ^ n3117 ^ 1'b0 ;
  assign n49967 = ~n28450 & n49966 ;
  assign n49968 = ( n18276 & n49965 ) | ( n18276 & n49967 ) | ( n49965 & n49967 ) ;
  assign n49969 = ( n18698 & n41138 ) | ( n18698 & ~n49968 ) | ( n41138 & ~n49968 ) ;
  assign n49970 = n49969 ^ n26230 ^ 1'b0 ;
  assign n49971 = n49964 & n49970 ;
  assign n49972 = n7494 ^ x220 ^ 1'b0 ;
  assign n49973 = n9452 & n49972 ;
  assign n49975 = n15655 & n20741 ;
  assign n49974 = n14093 & ~n24124 ;
  assign n49976 = n49975 ^ n49974 ^ 1'b0 ;
  assign n49977 = n49976 ^ n43396 ^ 1'b0 ;
  assign n49978 = ( n15845 & ~n28027 ) | ( n15845 & n30883 ) | ( ~n28027 & n30883 ) ;
  assign n49979 = ( n2026 & ~n36717 ) | ( n2026 & n49978 ) | ( ~n36717 & n49978 ) ;
  assign n49980 = ( n1254 & ~n21432 ) | ( n1254 & n29972 ) | ( ~n21432 & n29972 ) ;
  assign n49981 = n6464 & ~n12714 ;
  assign n49982 = ~n26073 & n49981 ;
  assign n49983 = ~n6370 & n27120 ;
  assign n49984 = n49982 & n49983 ;
  assign n49985 = n49980 | n49984 ;
  assign n49986 = n10390 ^ n7788 ^ 1'b0 ;
  assign n49987 = n49986 ^ n18348 ^ n3426 ;
  assign n49988 = n37220 & n46166 ;
  assign n49989 = ~x207 & n41801 ;
  assign n49990 = n22323 & ~n49989 ;
  assign n49991 = n1669 & n24174 ;
  assign n49992 = ( n23798 & n29932 ) | ( n23798 & ~n36082 ) | ( n29932 & ~n36082 ) ;
  assign n49993 = ~n26313 & n49992 ;
  assign n49994 = ~n49991 & n49993 ;
  assign n49995 = ~n16333 & n35880 ;
  assign n49996 = n49995 ^ n37155 ^ n3951 ;
  assign n49997 = n11043 ^ n11006 ^ n1367 ;
  assign n49998 = ~n17788 & n49997 ;
  assign n49999 = n49998 ^ n12970 ^ n7265 ;
  assign n50000 = n15934 ^ n15683 ^ 1'b0 ;
  assign n50001 = n50000 ^ n48743 ^ n30217 ;
  assign n50002 = n4426 & ~n11488 ;
  assign n50003 = n50002 ^ n1572 ^ 1'b0 ;
  assign n50004 = ( ~n5905 & n43595 ) | ( ~n5905 & n50003 ) | ( n43595 & n50003 ) ;
  assign n50005 = n7381 ^ n4253 ^ 1'b0 ;
  assign n50006 = n33548 ^ n33079 ^ n15436 ;
  assign n50007 = n45135 & n50006 ;
  assign n50008 = n50007 ^ n13176 ^ 1'b0 ;
  assign n50009 = n18640 & ~n20055 ;
  assign n50010 = ~n32680 & n50009 ;
  assign n50011 = n23965 & ~n45388 ;
  assign n50012 = n50010 & n50011 ;
  assign n50013 = n50012 ^ n10842 ^ 1'b0 ;
  assign n50014 = n19911 ^ n5752 ^ 1'b0 ;
  assign n50016 = n11585 & n41582 ;
  assign n50017 = n16475 & n50016 ;
  assign n50018 = n23279 & n50017 ;
  assign n50015 = n4753 | n22925 ;
  assign n50019 = n50018 ^ n50015 ^ 1'b0 ;
  assign n50020 = n10093 ^ n7492 ^ 1'b0 ;
  assign n50021 = ~n20357 & n50020 ;
  assign n50022 = n50021 ^ n43343 ^ n13590 ;
  assign n50023 = n50022 ^ n627 ^ 1'b0 ;
  assign n50024 = n38342 ^ n14096 ^ 1'b0 ;
  assign n50025 = n30766 ^ n16914 ^ x59 ;
  assign n50026 = ~n19848 & n25798 ;
  assign n50027 = ~n40141 & n50026 ;
  assign n50028 = n50027 ^ n13851 ^ n8413 ;
  assign n50029 = n36861 ^ n28365 ^ 1'b0 ;
  assign n50030 = ( ~n2809 & n2986 ) | ( ~n2809 & n21227 ) | ( n2986 & n21227 ) ;
  assign n50031 = n50030 ^ n49655 ^ 1'b0 ;
  assign n50032 = n28578 & n38105 ;
  assign n50033 = n50032 ^ n19324 ^ 1'b0 ;
  assign n50034 = n19888 & ~n30009 ;
  assign n50035 = n2558 & n50034 ;
  assign n50036 = n666 & n20909 ;
  assign n50037 = n50036 ^ n15742 ^ 1'b0 ;
  assign n50038 = ~n27069 & n48289 ;
  assign n50039 = ~n22723 & n50038 ;
  assign n50040 = n11857 & n50039 ;
  assign n50041 = n30323 ^ n1950 ^ 1'b0 ;
  assign n50043 = n8651 ^ n7908 ^ n2070 ;
  assign n50042 = n11806 & ~n37322 ;
  assign n50044 = n50043 ^ n50042 ^ 1'b0 ;
  assign n50045 = ( n1927 & n8636 ) | ( n1927 & ~n17627 ) | ( n8636 & ~n17627 ) ;
  assign n50046 = n20265 ^ n12416 ^ n10758 ;
  assign n50047 = ~n6787 & n38242 ;
  assign n50048 = ( n12301 & n38202 ) | ( n12301 & ~n40287 ) | ( n38202 & ~n40287 ) ;
  assign n50049 = ( n2260 & n5231 ) | ( n2260 & ~n7226 ) | ( n5231 & ~n7226 ) ;
  assign n50050 = n50049 ^ n38232 ^ n20669 ;
  assign n50051 = n26393 | n28769 ;
  assign n50052 = n48512 ^ n18684 ^ 1'b0 ;
  assign n50053 = n7501 ^ n5104 ^ n494 ;
  assign n50054 = n622 & ~n50053 ;
  assign n50055 = n23824 ^ n20987 ^ n2924 ;
  assign n50056 = n26967 ^ n5086 ^ 1'b0 ;
  assign n50057 = ~n2841 & n20238 ;
  assign n50058 = n50057 ^ n23813 ^ 1'b0 ;
  assign n50059 = n50058 ^ n48853 ^ n47885 ;
  assign n50060 = n5911 ^ n2968 ^ 1'b0 ;
  assign n50061 = ~n2412 & n50060 ;
  assign n50062 = n50061 ^ n43790 ^ n26217 ;
  assign n50063 = n31625 ^ n4662 ^ n2796 ;
  assign n50064 = n3529 & ~n50063 ;
  assign n50065 = ~n17971 & n50064 ;
  assign n50066 = ~n25090 & n30570 ;
  assign n50067 = n50066 ^ n38584 ^ 1'b0 ;
  assign n50068 = n10366 | n11615 ;
  assign n50069 = n50068 ^ n880 ^ 1'b0 ;
  assign n50070 = ~n8416 & n13374 ;
  assign n50071 = n26636 & n50070 ;
  assign n50072 = n3792 | n50071 ;
  assign n50073 = ( n16800 & n48977 ) | ( n16800 & n50072 ) | ( n48977 & n50072 ) ;
  assign n50074 = n21342 ^ n14524 ^ 1'b0 ;
  assign n50075 = ~n31618 & n50074 ;
  assign n50076 = ~n37782 & n49377 ;
  assign n50077 = n50076 ^ n29237 ^ 1'b0 ;
  assign n50078 = n50077 ^ n2873 ^ 1'b0 ;
  assign n50079 = n50075 & n50078 ;
  assign n50080 = n5569 & ~n9643 ;
  assign n50081 = n9793 & n50080 ;
  assign n50082 = ( n10009 & n25691 ) | ( n10009 & n50081 ) | ( n25691 & n50081 ) ;
  assign n50083 = n50079 & ~n50082 ;
  assign n50087 = ~n4706 & n27009 ;
  assign n50088 = n50087 ^ n19014 ^ n2503 ;
  assign n50084 = n24146 ^ n12602 ^ n3437 ;
  assign n50085 = ( ~n12037 & n13584 ) | ( ~n12037 & n50084 ) | ( n13584 & n50084 ) ;
  assign n50086 = n50085 ^ n40093 ^ n8536 ;
  assign n50089 = n50088 ^ n50086 ^ n27248 ;
  assign n50090 = n28790 ^ n26044 ^ 1'b0 ;
  assign n50091 = n30379 ^ n19171 ^ 1'b0 ;
  assign n50092 = n50091 ^ n37502 ^ n1666 ;
  assign n50097 = n24380 | n45553 ;
  assign n50093 = n10233 ^ n3811 ^ 1'b0 ;
  assign n50094 = n15221 & n50093 ;
  assign n50095 = n50094 ^ n9919 ^ n1380 ;
  assign n50096 = n46063 & n50095 ;
  assign n50098 = n50097 ^ n50096 ^ 1'b0 ;
  assign n50099 = n28350 & ~n39579 ;
  assign n50100 = n12967 ^ n7601 ^ 1'b0 ;
  assign n50101 = ~n50099 & n50100 ;
  assign n50102 = n29851 & n46681 ;
  assign n50105 = n27880 ^ n15359 ^ 1'b0 ;
  assign n50103 = n7098 & n14735 ;
  assign n50104 = n7812 & n50103 ;
  assign n50106 = n50105 ^ n50104 ^ n29570 ;
  assign n50107 = n19685 | n24470 ;
  assign n50109 = ~n1826 & n3873 ;
  assign n50110 = ~n4204 & n50109 ;
  assign n50108 = n7942 & ~n25157 ;
  assign n50111 = n50110 ^ n50108 ^ 1'b0 ;
  assign n50112 = ~n13224 & n50111 ;
  assign n50116 = n16080 ^ n6848 ^ 1'b0 ;
  assign n50113 = ( n14318 & ~n34468 ) | ( n14318 & n39004 ) | ( ~n34468 & n39004 ) ;
  assign n50114 = ( n15140 & n17599 ) | ( n15140 & n50113 ) | ( n17599 & n50113 ) ;
  assign n50115 = n50114 ^ n36848 ^ n784 ;
  assign n50117 = n50116 ^ n50115 ^ n13031 ;
  assign n50118 = n30315 & ~n49365 ;
  assign n50119 = n50118 ^ n27222 ^ n6297 ;
  assign n50120 = n684 & ~n2418 ;
  assign n50121 = ~n3955 & n50120 ;
  assign n50122 = n24891 ^ n6940 ^ 1'b0 ;
  assign n50123 = n42225 | n50122 ;
  assign n50124 = ( n15004 & ~n50121 ) | ( n15004 & n50123 ) | ( ~n50121 & n50123 ) ;
  assign n50125 = ~n14279 & n22758 ;
  assign n50126 = n50115 & n50125 ;
  assign n50127 = ( n9115 & ~n10092 ) | ( n9115 & n35062 ) | ( ~n10092 & n35062 ) ;
  assign n50128 = n42253 ^ n36444 ^ 1'b0 ;
  assign n50129 = n50127 & n50128 ;
  assign n50130 = n4754 ^ x222 ^ 1'b0 ;
  assign n50131 = n44054 & ~n50130 ;
  assign n50132 = n14941 & n50131 ;
  assign n50133 = ( n9497 & n48824 ) | ( n9497 & n50132 ) | ( n48824 & n50132 ) ;
  assign n50134 = ( n6027 & ~n6414 ) | ( n6027 & n50133 ) | ( ~n6414 & n50133 ) ;
  assign n50135 = n23437 ^ x173 ^ 1'b0 ;
  assign n50136 = ( n5443 & n11858 ) | ( n5443 & ~n50135 ) | ( n11858 & ~n50135 ) ;
  assign n50138 = n47070 ^ n28512 ^ n12097 ;
  assign n50137 = n48598 ^ n20923 ^ n4198 ;
  assign n50139 = n50138 ^ n50137 ^ x83 ;
  assign n50140 = ( n43640 & ~n50136 ) | ( n43640 & n50139 ) | ( ~n50136 & n50139 ) ;
  assign n50141 = n20665 ^ n15296 ^ n10232 ;
  assign n50142 = ( n1620 & n16895 ) | ( n1620 & n49111 ) | ( n16895 & n49111 ) ;
  assign n50143 = ( n1303 & n6753 ) | ( n1303 & ~n30008 ) | ( n6753 & ~n30008 ) ;
  assign n50145 = ( n16877 & ~n19393 ) | ( n16877 & n26255 ) | ( ~n19393 & n26255 ) ;
  assign n50144 = n30894 | n45192 ;
  assign n50146 = n50145 ^ n50144 ^ n32762 ;
  assign n50147 = n50146 ^ n46249 ^ n2614 ;
  assign n50148 = n33033 | n42971 ;
  assign n50149 = n20973 ^ n19068 ^ 1'b0 ;
  assign n50150 = n17657 & ~n41044 ;
  assign n50151 = ~n30428 & n50150 ;
  assign n50153 = ( n27844 & n34811 ) | ( n27844 & ~n35608 ) | ( n34811 & ~n35608 ) ;
  assign n50154 = n50153 ^ n8417 ^ n4367 ;
  assign n50152 = n14300 & ~n46250 ;
  assign n50155 = n50154 ^ n50152 ^ 1'b0 ;
  assign n50156 = n41998 ^ n4559 ^ 1'b0 ;
  assign n50157 = ( n39430 & n40959 ) | ( n39430 & ~n50156 ) | ( n40959 & ~n50156 ) ;
  assign n50158 = ( n1355 & ~n7616 ) | ( n1355 & n29771 ) | ( ~n7616 & n29771 ) ;
  assign n50159 = n3505 | n10917 ;
  assign n50160 = n50159 ^ n34029 ^ n1941 ;
  assign n50161 = n34410 ^ n8861 ^ n7607 ;
  assign n50162 = n50161 ^ n23023 ^ 1'b0 ;
  assign n50164 = ( n6786 & ~n20720 ) | ( n6786 & n36476 ) | ( ~n20720 & n36476 ) ;
  assign n50163 = n11095 ^ n10939 ^ 1'b0 ;
  assign n50165 = n50164 ^ n50163 ^ n11239 ;
  assign n50166 = n1378 & ~n1942 ;
  assign n50167 = ( ~n17853 & n21711 ) | ( ~n17853 & n50166 ) | ( n21711 & n50166 ) ;
  assign n50168 = ~n50165 & n50167 ;
  assign n50169 = n30537 & ~n50168 ;
  assign n50170 = n49890 ^ n8217 ^ n6840 ;
  assign n50171 = n26627 ^ n2209 ^ 1'b0 ;
  assign n50172 = ( n16914 & n21800 ) | ( n16914 & ~n25157 ) | ( n21800 & ~n25157 ) ;
  assign n50173 = n23377 | n50172 ;
  assign n50174 = n14228 ^ n7931 ^ 1'b0 ;
  assign n50175 = n39420 | n50174 ;
  assign n50176 = n26044 ^ n580 ^ 1'b0 ;
  assign n50177 = n50176 ^ n30719 ^ n14723 ;
  assign n50178 = ~n46487 & n50177 ;
  assign n50179 = n35546 & ~n44634 ;
  assign n50180 = ( n7377 & n17125 ) | ( n7377 & n50179 ) | ( n17125 & n50179 ) ;
  assign n50181 = ( n4078 & n8821 ) | ( n4078 & ~n33364 ) | ( n8821 & ~n33364 ) ;
  assign n50182 = ( n20559 & n37784 ) | ( n20559 & ~n50181 ) | ( n37784 & ~n50181 ) ;
  assign n50183 = n30766 ^ n10916 ^ 1'b0 ;
  assign n50184 = ~n15211 & n50183 ;
  assign n50185 = ( n14455 & n26679 ) | ( n14455 & n50184 ) | ( n26679 & n50184 ) ;
  assign n50186 = n49273 ^ n46550 ^ n11343 ;
  assign n50187 = x93 & n4240 ;
  assign n50188 = ~n31615 & n39758 ;
  assign n50189 = n10659 | n50188 ;
  assign n50190 = n50189 ^ n12244 ^ n7895 ;
  assign n50191 = n14531 & n48676 ;
  assign n50192 = n9329 & ~n19991 ;
  assign n50193 = ~n25875 & n50192 ;
  assign n50194 = n37345 ^ n34706 ^ n30483 ;
  assign n50195 = n50194 ^ n41765 ^ n35908 ;
  assign n50196 = ~n15542 & n41915 ;
  assign n50197 = ( n8071 & n31802 ) | ( n8071 & n50196 ) | ( n31802 & n50196 ) ;
  assign n50198 = n35297 ^ n3084 ^ n2999 ;
  assign n50199 = n50198 ^ n42689 ^ 1'b0 ;
  assign n50200 = n14324 & ~n50199 ;
  assign n50201 = ( n11668 & ~n14232 ) | ( n11668 & n50200 ) | ( ~n14232 & n50200 ) ;
  assign n50204 = n20627 ^ n7588 ^ 1'b0 ;
  assign n50202 = n17748 | n20698 ;
  assign n50203 = n50202 ^ n37813 ^ 1'b0 ;
  assign n50205 = n50204 ^ n50203 ^ n8560 ;
  assign n50208 = n35616 ^ n16675 ^ n6114 ;
  assign n50206 = n8986 & ~n9900 ;
  assign n50207 = n50206 ^ n14481 ^ n11784 ;
  assign n50209 = n50208 ^ n50207 ^ n14595 ;
  assign n50211 = n6728 ^ n3754 ^ 1'b0 ;
  assign n50212 = n26714 ^ n7070 ^ 1'b0 ;
  assign n50213 = ( n10152 & ~n11221 ) | ( n10152 & n50212 ) | ( ~n11221 & n50212 ) ;
  assign n50214 = ( n7503 & n50211 ) | ( n7503 & ~n50213 ) | ( n50211 & ~n50213 ) ;
  assign n50210 = n20614 & ~n25514 ;
  assign n50215 = n50214 ^ n50210 ^ 1'b0 ;
  assign n50216 = n9064 | n12453 ;
  assign n50217 = n50216 ^ n8704 ^ 1'b0 ;
  assign n50218 = n12941 & n50217 ;
  assign n50219 = ~x46 & n50218 ;
  assign n50220 = n4662 & ~n30527 ;
  assign n50221 = n20780 & n50220 ;
  assign n50222 = n28682 ^ n7286 ^ 1'b0 ;
  assign n50223 = ( n1722 & ~n40727 ) | ( n1722 & n50222 ) | ( ~n40727 & n50222 ) ;
  assign n50224 = n30635 & ~n50223 ;
  assign n50225 = n50224 ^ n47793 ^ 1'b0 ;
  assign n50226 = n40195 ^ n23390 ^ n10043 ;
  assign n50227 = n31417 ^ n5793 ^ 1'b0 ;
  assign n50228 = n25149 & n50227 ;
  assign n50229 = n50228 ^ n6091 ^ 1'b0 ;
  assign n50230 = n10289 | n15765 ;
  assign n50231 = n9275 | n50230 ;
  assign n50232 = n50231 ^ n17061 ^ 1'b0 ;
  assign n50233 = n50232 ^ n6114 ^ 1'b0 ;
  assign n50234 = n27664 ^ n17415 ^ n4980 ;
  assign n50235 = ~n29663 & n44713 ;
  assign n50236 = ( n11680 & ~n22479 ) | ( n11680 & n35560 ) | ( ~n22479 & n35560 ) ;
  assign n50237 = n50236 ^ n12024 ^ 1'b0 ;
  assign n50238 = n40822 ^ n1915 ^ 1'b0 ;
  assign n50239 = ~n5974 & n50238 ;
  assign n50240 = n27394 & n47262 ;
  assign n50241 = n50240 ^ n29509 ^ 1'b0 ;
  assign n50242 = n13405 & ~n42392 ;
  assign n50243 = n37686 & n50242 ;
  assign n50244 = n36576 ^ n24483 ^ 1'b0 ;
  assign n50245 = n50243 | n50244 ;
  assign n50246 = n14686 ^ n7772 ^ 1'b0 ;
  assign n50247 = ( n3262 & n24851 ) | ( n3262 & ~n50246 ) | ( n24851 & ~n50246 ) ;
  assign n50248 = ( n14904 & ~n18789 ) | ( n14904 & n40574 ) | ( ~n18789 & n40574 ) ;
  assign n50249 = ( n3942 & ~n17936 ) | ( n3942 & n50248 ) | ( ~n17936 & n50248 ) ;
  assign n50250 = ( n15855 & ~n23644 ) | ( n15855 & n27719 ) | ( ~n23644 & n27719 ) ;
  assign n50251 = n32444 ^ n6178 ^ n5643 ;
  assign n50252 = n50251 ^ n28233 ^ n2588 ;
  assign n50253 = ~n3219 & n31604 ;
  assign n50254 = n50253 ^ n2349 ^ 1'b0 ;
  assign n50255 = n45415 ^ n44014 ^ n25740 ;
  assign n50256 = ( n50252 & ~n50254 ) | ( n50252 & n50255 ) | ( ~n50254 & n50255 ) ;
  assign n50257 = n32253 ^ n5300 ^ 1'b0 ;
  assign n50258 = n50257 ^ n32011 ^ n13333 ;
  assign n50259 = n24671 ^ n13918 ^ n10942 ;
  assign n50260 = n32899 ^ n16667 ^ n4051 ;
  assign n50261 = ( n20024 & n36270 ) | ( n20024 & n50260 ) | ( n36270 & n50260 ) ;
  assign n50262 = n10429 & n37866 ;
  assign n50263 = ~n50261 & n50262 ;
  assign n50264 = n3535 & n15442 ;
  assign n50265 = n48981 & n50264 ;
  assign n50266 = ( ~n10318 & n20491 ) | ( ~n10318 & n50265 ) | ( n20491 & n50265 ) ;
  assign n50267 = n50266 ^ n23859 ^ 1'b0 ;
  assign n50268 = n50267 ^ n16541 ^ 1'b0 ;
  assign n50269 = n7665 | n50268 ;
  assign n50270 = ~n31491 & n50269 ;
  assign n50271 = ~n22595 & n50270 ;
  assign n50272 = n47343 ^ n38914 ^ 1'b0 ;
  assign n50273 = ~n8107 & n23064 ;
  assign n50274 = ~n40785 & n50273 ;
  assign n50275 = n50274 ^ n45028 ^ 1'b0 ;
  assign n50278 = ( n19803 & ~n29618 ) | ( n19803 & n32556 ) | ( ~n29618 & n32556 ) ;
  assign n50279 = n17627 & n22690 ;
  assign n50280 = ~n50278 & n50279 ;
  assign n50276 = n23961 ^ n3765 ^ 1'b0 ;
  assign n50277 = n9538 | n50276 ;
  assign n50281 = n50280 ^ n50277 ^ 1'b0 ;
  assign n50282 = ( n20652 & ~n21665 ) | ( n20652 & n36489 ) | ( ~n21665 & n36489 ) ;
  assign n50283 = n19038 & ~n21132 ;
  assign n50284 = ~n2965 & n41594 ;
  assign n50285 = n50284 ^ n38056 ^ 1'b0 ;
  assign n50286 = n19618 & n50285 ;
  assign n50287 = ~n50283 & n50286 ;
  assign n50288 = n50287 ^ n46890 ^ n3056 ;
  assign n50289 = ( n27076 & ~n50282 ) | ( n27076 & n50288 ) | ( ~n50282 & n50288 ) ;
  assign n50290 = n6204 ^ n4618 ^ 1'b0 ;
  assign n50291 = n14285 & ~n50290 ;
  assign n50292 = n50291 ^ n32079 ^ n1271 ;
  assign n50293 = n46050 & n49695 ;
  assign n50294 = n50293 ^ n12875 ^ n10536 ;
  assign n50295 = n6749 & ~n10987 ;
  assign n50296 = ( n7900 & n27658 ) | ( n7900 & ~n32052 ) | ( n27658 & ~n32052 ) ;
  assign n50297 = n29432 & n45352 ;
  assign n50298 = n42808 ^ n32763 ^ 1'b0 ;
  assign n50299 = n30787 ^ n21403 ^ n13804 ;
  assign n50300 = n298 & ~n50299 ;
  assign n50301 = ( n2940 & n11706 ) | ( n2940 & ~n18518 ) | ( n11706 & ~n18518 ) ;
  assign n50302 = n46314 ^ n12912 ^ 1'b0 ;
  assign n50303 = n50301 & n50302 ;
  assign n50304 = ~n36886 & n42176 ;
  assign n50305 = n8113 & n14294 ;
  assign n50306 = n50305 ^ n1647 ^ 1'b0 ;
  assign n50307 = n50306 ^ n17246 ^ 1'b0 ;
  assign n50308 = n32288 ^ n26661 ^ n8745 ;
  assign n50309 = ( n6138 & n49110 ) | ( n6138 & ~n50308 ) | ( n49110 & ~n50308 ) ;
  assign n50310 = ( n883 & n34952 ) | ( n883 & ~n43586 ) | ( n34952 & ~n43586 ) ;
  assign n50311 = n16630 ^ n7695 ^ 1'b0 ;
  assign n50312 = ( n8861 & n21644 ) | ( n8861 & n50311 ) | ( n21644 & n50311 ) ;
  assign n50313 = n37357 ^ n36836 ^ n30805 ;
  assign n50314 = n46783 ^ n1732 ^ 1'b0 ;
  assign n50315 = n4523 & n50314 ;
  assign n50316 = n15010 & n38352 ;
  assign n50317 = n50316 ^ n9570 ^ 1'b0 ;
  assign n50318 = n41918 ^ n18319 ^ 1'b0 ;
  assign n50319 = ~n50317 & n50318 ;
  assign n50320 = ~n4360 & n39388 ;
  assign n50321 = n29686 & ~n34718 ;
  assign n50322 = ~n50320 & n50321 ;
  assign n50323 = ( n11751 & ~n15959 ) | ( n11751 & n33901 ) | ( ~n15959 & n33901 ) ;
  assign n50324 = n29261 & n37652 ;
  assign n50325 = ( n4709 & ~n16030 ) | ( n4709 & n30707 ) | ( ~n16030 & n30707 ) ;
  assign n50326 = n27394 & n50325 ;
  assign n50327 = n43084 ^ n25598 ^ 1'b0 ;
  assign n50328 = n27995 & ~n50327 ;
  assign n50330 = n16433 ^ n1055 ^ 1'b0 ;
  assign n50329 = ( n2344 & n5693 ) | ( n2344 & n5934 ) | ( n5693 & n5934 ) ;
  assign n50331 = n50330 ^ n50329 ^ n7812 ;
  assign n50332 = n6080 | n10485 ;
  assign n50333 = n1331 | n50332 ;
  assign n50334 = ( n10830 & n50331 ) | ( n10830 & ~n50333 ) | ( n50331 & ~n50333 ) ;
  assign n50335 = n1293 | n15169 ;
  assign n50336 = ( n23663 & n28252 ) | ( n23663 & n50335 ) | ( n28252 & n50335 ) ;
  assign n50337 = n50336 ^ n31033 ^ n17185 ;
  assign n50338 = n50337 ^ n35894 ^ n32999 ;
  assign n50339 = n5411 & ~n38002 ;
  assign n50340 = n50339 ^ n9240 ^ 1'b0 ;
  assign n50341 = n19768 & ~n32617 ;
  assign n50342 = n50341 ^ n14341 ^ 1'b0 ;
  assign n50343 = n42610 ^ n30243 ^ 1'b0 ;
  assign n50344 = n15714 | n50343 ;
  assign n50346 = n37208 ^ n7694 ^ n2069 ;
  assign n50345 = n4011 | n42447 ;
  assign n50347 = n50346 ^ n50345 ^ 1'b0 ;
  assign n50348 = ( n26526 & n42661 ) | ( n26526 & n50347 ) | ( n42661 & n50347 ) ;
  assign n50349 = n42725 ^ n24517 ^ n16763 ;
  assign n50350 = ~n16040 & n30877 ;
  assign n50351 = ( n9010 & n14108 ) | ( n9010 & n26707 ) | ( n14108 & n26707 ) ;
  assign n50352 = n14079 ^ n6959 ^ 1'b0 ;
  assign n50353 = n45718 & n50352 ;
  assign n50354 = ( n47131 & ~n50351 ) | ( n47131 & n50353 ) | ( ~n50351 & n50353 ) ;
  assign n50355 = n29150 ^ n24047 ^ 1'b0 ;
  assign n50356 = ~n11656 & n50355 ;
  assign n50357 = ~n3579 & n50356 ;
  assign n50358 = n6097 | n18018 ;
  assign n50359 = ( x228 & ~n1920 ) | ( x228 & n50358 ) | ( ~n1920 & n50358 ) ;
  assign n50360 = n23823 | n50359 ;
  assign n50361 = n27541 ^ n16002 ^ 1'b0 ;
  assign n50362 = n2410 | n25375 ;
  assign n50363 = n11185 & ~n50362 ;
  assign n50364 = ~n10383 & n34444 ;
  assign n50368 = ( n9816 & n16939 ) | ( n9816 & ~n24967 ) | ( n16939 & ~n24967 ) ;
  assign n50369 = n50368 ^ n39877 ^ n18861 ;
  assign n50365 = ( n5435 & ~n6648 ) | ( n5435 & n11952 ) | ( ~n6648 & n11952 ) ;
  assign n50366 = ~n26941 & n50365 ;
  assign n50367 = n50366 ^ n23829 ^ 1'b0 ;
  assign n50370 = n50369 ^ n50367 ^ n49737 ;
  assign n50371 = n36478 ^ n15033 ^ n11542 ;
  assign n50372 = n47102 ^ n9655 ^ 1'b0 ;
  assign n50373 = n11091 & ~n33269 ;
  assign n50374 = n42648 ^ n9644 ^ n5068 ;
  assign n50375 = n47549 & ~n50374 ;
  assign n50376 = ( ~n14454 & n50373 ) | ( ~n14454 & n50375 ) | ( n50373 & n50375 ) ;
  assign n50377 = x9 & n15206 ;
  assign n50378 = n9542 & n50377 ;
  assign n50379 = n16962 ^ n11777 ^ 1'b0 ;
  assign n50380 = n50378 & ~n50379 ;
  assign n50381 = ( n3798 & n4956 ) | ( n3798 & ~n30795 ) | ( n4956 & ~n30795 ) ;
  assign n50382 = ( n29562 & n50380 ) | ( n29562 & n50381 ) | ( n50380 & n50381 ) ;
  assign n50383 = n40422 ^ n6360 ^ 1'b0 ;
  assign n50384 = ~n28231 & n50383 ;
  assign n50385 = n50384 ^ n24826 ^ n3358 ;
  assign n50386 = n6246 & ~n50385 ;
  assign n50387 = n13736 ^ n12593 ^ 1'b0 ;
  assign n50388 = n46038 | n50387 ;
  assign n50392 = n9311 & ~n47627 ;
  assign n50393 = n2001 & n50392 ;
  assign n50394 = n50393 ^ n1681 ^ 1'b0 ;
  assign n50389 = n23038 ^ n9341 ^ n3373 ;
  assign n50390 = ( ~n8790 & n24148 ) | ( ~n8790 & n50389 ) | ( n24148 & n50389 ) ;
  assign n50391 = n9632 | n50390 ;
  assign n50395 = n50394 ^ n50391 ^ 1'b0 ;
  assign n50396 = n1404 & n48271 ;
  assign n50397 = n50396 ^ n39949 ^ 1'b0 ;
  assign n50398 = ~n28848 & n50397 ;
  assign n50399 = n50398 ^ n33867 ^ n10888 ;
  assign n50400 = n50399 ^ n1772 ^ 1'b0 ;
  assign n50401 = ~n42032 & n50400 ;
  assign n50402 = n31858 & n32981 ;
  assign n50403 = ( n21753 & n29090 ) | ( n21753 & ~n32143 ) | ( n29090 & ~n32143 ) ;
  assign n50404 = n14933 & ~n47526 ;
  assign n50405 = n50404 ^ n11733 ^ 1'b0 ;
  assign n50406 = n48071 ^ n471 ^ 1'b0 ;
  assign n50407 = n13729 ^ n10836 ^ n10553 ;
  assign n50408 = n26106 ^ n21809 ^ 1'b0 ;
  assign n50409 = n31144 ^ n21036 ^ n20136 ;
  assign n50410 = n38337 & ~n50409 ;
  assign n50411 = n50410 ^ n6206 ^ 1'b0 ;
  assign n50412 = n33143 ^ n10413 ^ 1'b0 ;
  assign n50413 = n14842 | n50412 ;
  assign n50414 = n50413 ^ n8193 ^ 1'b0 ;
  assign n50415 = x53 & n4405 ;
  assign n50416 = ~n14797 & n25650 ;
  assign n50417 = n50416 ^ n26780 ^ n11617 ;
  assign n50419 = n3994 ^ n748 ^ 1'b0 ;
  assign n50420 = ~n27989 & n50419 ;
  assign n50418 = n23327 ^ n12202 ^ 1'b0 ;
  assign n50421 = n50420 ^ n50418 ^ n13347 ;
  assign n50422 = n2184 & ~n2866 ;
  assign n50423 = n50422 ^ n37223 ^ 1'b0 ;
  assign n50424 = ( ~n33218 & n39399 ) | ( ~n33218 & n50423 ) | ( n39399 & n50423 ) ;
  assign n50425 = n23025 & ~n41870 ;
  assign n50426 = n50425 ^ n10781 ^ 1'b0 ;
  assign n50427 = ~n19331 & n50426 ;
  assign n50428 = ~n18007 & n50427 ;
  assign n50429 = n10872 & ~n16552 ;
  assign n50430 = n14165 & ~n50429 ;
  assign n50431 = n50428 | n50430 ;
  assign n50432 = n14645 ^ n14228 ^ n306 ;
  assign n50433 = n28840 ^ n15495 ^ n1305 ;
  assign n50434 = ( n10346 & ~n17115 ) | ( n10346 & n50433 ) | ( ~n17115 & n50433 ) ;
  assign n50435 = n48896 ^ n20047 ^ 1'b0 ;
  assign n50436 = n32966 ^ n18462 ^ 1'b0 ;
  assign n50437 = n781 | n50436 ;
  assign n50438 = n16560 ^ n8927 ^ 1'b0 ;
  assign n50439 = ~n26854 & n50438 ;
  assign n50440 = n23767 & n25837 ;
  assign n50441 = n39530 & n50440 ;
  assign n50442 = ( n826 & n14207 ) | ( n826 & ~n50441 ) | ( n14207 & ~n50441 ) ;
  assign n50443 = ~n27794 & n45565 ;
  assign n50444 = n14503 ^ n12540 ^ 1'b0 ;
  assign n50445 = n2552 & n50444 ;
  assign n50446 = ~n16486 & n50445 ;
  assign n50447 = n50446 ^ n8379 ^ 1'b0 ;
  assign n50448 = ( n3019 & ~n5665 ) | ( n3019 & n9212 ) | ( ~n5665 & n9212 ) ;
  assign n50449 = ( n1927 & n42316 ) | ( n1927 & n50448 ) | ( n42316 & n50448 ) ;
  assign n50450 = n28499 ^ n16762 ^ 1'b0 ;
  assign n50451 = n50450 ^ n1065 ^ n494 ;
  assign n50452 = ( n4184 & ~n4624 ) | ( n4184 & n4889 ) | ( ~n4624 & n4889 ) ;
  assign n50453 = n50451 & ~n50452 ;
  assign n50454 = ( n4939 & n10541 ) | ( n4939 & ~n50453 ) | ( n10541 & ~n50453 ) ;
  assign n50455 = n50454 ^ n42993 ^ n3352 ;
  assign n50456 = n31844 ^ n3937 ^ 1'b0 ;
  assign n50457 = n22283 ^ n16850 ^ 1'b0 ;
  assign n50458 = n43126 & n50457 ;
  assign n50459 = n6618 & ~n47852 ;
  assign n50460 = n31092 & n50459 ;
  assign n50462 = n47228 ^ n16349 ^ 1'b0 ;
  assign n50463 = ( n3994 & ~n6332 ) | ( n3994 & n50462 ) | ( ~n6332 & n50462 ) ;
  assign n50461 = n6980 & ~n8935 ;
  assign n50464 = n50463 ^ n50461 ^ 1'b0 ;
  assign n50465 = n31996 & n46563 ;
  assign n50466 = n14552 & ~n29854 ;
  assign n50467 = n50466 ^ n47518 ^ n35460 ;
  assign n50468 = n21990 ^ x77 ^ 1'b0 ;
  assign n50469 = ( n9704 & ~n48401 ) | ( n9704 & n50468 ) | ( ~n48401 & n50468 ) ;
  assign n50470 = n50469 ^ n49986 ^ n35807 ;
  assign n50471 = n26769 ^ n7596 ^ 1'b0 ;
  assign n50472 = n34424 & n35669 ;
  assign n50473 = n44756 & n50472 ;
  assign n50474 = ( n15990 & ~n20972 ) | ( n15990 & n30428 ) | ( ~n20972 & n30428 ) ;
  assign n50475 = ( n4103 & ~n34154 ) | ( n4103 & n50474 ) | ( ~n34154 & n50474 ) ;
  assign n50476 = n25098 & ~n50475 ;
  assign n50477 = ~n11035 & n50476 ;
  assign n50478 = ~n7138 & n27724 ;
  assign n50479 = ~n28363 & n43335 ;
  assign n50480 = ~n19604 & n25571 ;
  assign n50481 = n17855 & n50480 ;
  assign n50483 = n14381 ^ n12840 ^ 1'b0 ;
  assign n50484 = ~n9624 & n16737 ;
  assign n50485 = ~n50483 & n50484 ;
  assign n50486 = ( n7354 & ~n15831 ) | ( n7354 & n50485 ) | ( ~n15831 & n50485 ) ;
  assign n50482 = n4331 | n28388 ;
  assign n50487 = n50486 ^ n50482 ^ 1'b0 ;
  assign n50491 = ( n23376 & n33744 ) | ( n23376 & ~n34802 ) | ( n33744 & ~n34802 ) ;
  assign n50488 = n16103 | n24146 ;
  assign n50489 = n28829 | n50488 ;
  assign n50490 = n17963 & ~n50489 ;
  assign n50492 = n50491 ^ n50490 ^ 1'b0 ;
  assign n50493 = ( ~n9974 & n27550 ) | ( ~n9974 & n50492 ) | ( n27550 & n50492 ) ;
  assign n50494 = n41267 ^ n14908 ^ n5799 ;
  assign n50495 = ~n34808 & n50494 ;
  assign n50496 = n24594 ^ n5521 ^ 1'b0 ;
  assign n50497 = n20210 & n50496 ;
  assign n50498 = n50497 ^ n46518 ^ 1'b0 ;
  assign n50499 = n31888 ^ n12089 ^ n5974 ;
  assign n50500 = n50499 ^ n7859 ^ n5300 ;
  assign n50501 = ~n5054 & n40095 ;
  assign n50502 = n3480 & n50501 ;
  assign n50503 = ~n3306 & n6522 ;
  assign n50504 = n50503 ^ n7425 ^ 1'b0 ;
  assign n50505 = n50504 ^ n25598 ^ n2907 ;
  assign n50506 = n23380 & n50505 ;
  assign n50510 = n36792 ^ n26507 ^ n26431 ;
  assign n50511 = n10307 & n50510 ;
  assign n50512 = n40092 & n50511 ;
  assign n50513 = ~n28038 & n50512 ;
  assign n50507 = ( n13682 & ~n24005 ) | ( n13682 & n48200 ) | ( ~n24005 & n48200 ) ;
  assign n50508 = ( ~n8880 & n17690 ) | ( ~n8880 & n50507 ) | ( n17690 & n50507 ) ;
  assign n50509 = n15701 | n50508 ;
  assign n50514 = n50513 ^ n50509 ^ 1'b0 ;
  assign n50515 = n14269 ^ n3107 ^ 1'b0 ;
  assign n50516 = ~n32227 & n50515 ;
  assign n50517 = n1653 ^ n947 ^ 1'b0 ;
  assign n50518 = ( n1288 & ~n25998 ) | ( n1288 & n50517 ) | ( ~n25998 & n50517 ) ;
  assign n50519 = n50518 ^ n4735 ^ 1'b0 ;
  assign n50520 = n29148 & n30428 ;
  assign n50521 = n36564 ^ n36092 ^ 1'b0 ;
  assign n50522 = n23776 & ~n50521 ;
  assign n50523 = ( ~n4480 & n17013 ) | ( ~n4480 & n50522 ) | ( n17013 & n50522 ) ;
  assign n50526 = n31071 ^ n9750 ^ n8980 ;
  assign n50524 = n18477 & ~n33320 ;
  assign n50525 = n16135 & n50524 ;
  assign n50527 = n50526 ^ n50525 ^ n15978 ;
  assign n50528 = n9626 | n22514 ;
  assign n50529 = n50379 & ~n50528 ;
  assign n50530 = n11896 ^ n10555 ^ n1476 ;
  assign n50531 = ( n10505 & n50529 ) | ( n10505 & ~n50530 ) | ( n50529 & ~n50530 ) ;
  assign n50532 = n21264 ^ n12409 ^ n12093 ;
  assign n50533 = n19194 | n50532 ;
  assign n50534 = n50533 ^ n16655 ^ 1'b0 ;
  assign n50535 = ( n1708 & n17198 ) | ( n1708 & ~n42867 ) | ( n17198 & ~n42867 ) ;
  assign n50536 = n17211 & ~n50535 ;
  assign n50537 = n41504 & n50536 ;
  assign n50538 = n38264 & n39035 ;
  assign n50539 = ~n35747 & n50538 ;
  assign n50540 = n28388 ^ n24083 ^ 1'b0 ;
  assign n50541 = n7316 & n50540 ;
  assign n50542 = n42356 & n50541 ;
  assign n50543 = n50542 ^ n40311 ^ 1'b0 ;
  assign n50544 = ( n521 & ~n7243 ) | ( n521 & n13680 ) | ( ~n7243 & n13680 ) ;
  assign n50545 = ~n15489 & n19647 ;
  assign n50546 = n2827 | n22078 ;
  assign n50547 = ( n9291 & n25030 ) | ( n9291 & n50546 ) | ( n25030 & n50546 ) ;
  assign n50548 = ~n1026 & n4187 ;
  assign n50549 = ( n1904 & n29096 ) | ( n1904 & ~n50548 ) | ( n29096 & ~n50548 ) ;
  assign n50550 = n2951 & ~n6744 ;
  assign n50551 = ~n2951 & n50550 ;
  assign n50552 = n50551 ^ n34940 ^ n32857 ;
  assign n50553 = n3535 & n16110 ;
  assign n50554 = n16746 ^ n9358 ^ 1'b0 ;
  assign n50555 = n41017 ^ n22813 ^ 1'b0 ;
  assign n50556 = n13272 & ~n50555 ;
  assign n50557 = n19119 ^ n17332 ^ 1'b0 ;
  assign n50558 = n15855 & n25061 ;
  assign n50559 = ~n2316 & n50558 ;
  assign n50560 = n22983 & n34419 ;
  assign n50561 = n50560 ^ n17720 ^ n14614 ;
  assign n50562 = ( ~n11359 & n11916 ) | ( ~n11359 & n40426 ) | ( n11916 & n40426 ) ;
  assign n50563 = n3738 ^ n2073 ^ n1668 ;
  assign n50564 = n50563 ^ n41621 ^ n7664 ;
  assign n50565 = ~n6773 & n50564 ;
  assign n50566 = n50565 ^ n26339 ^ 1'b0 ;
  assign n50567 = ( n18201 & n42363 ) | ( n18201 & n50566 ) | ( n42363 & n50566 ) ;
  assign n50568 = ( n11527 & n13277 ) | ( n11527 & ~n33112 ) | ( n13277 & ~n33112 ) ;
  assign n50569 = ( n7553 & n9727 ) | ( n7553 & ~n14854 ) | ( n9727 & ~n14854 ) ;
  assign n50570 = n50569 ^ n19323 ^ 1'b0 ;
  assign n50571 = n49876 ^ n49500 ^ n33314 ;
  assign n50572 = n34701 | n41369 ;
  assign n50573 = n6105 | n50572 ;
  assign n50574 = n33655 ^ n8856 ^ 1'b0 ;
  assign n50575 = ~n23796 & n50574 ;
  assign n50576 = n25247 ^ n11283 ^ 1'b0 ;
  assign n50577 = n13639 | n50576 ;
  assign n50579 = ( n8486 & n16039 ) | ( n8486 & n28611 ) | ( n16039 & n28611 ) ;
  assign n50578 = n23244 & n31108 ;
  assign n50580 = n50579 ^ n50578 ^ 1'b0 ;
  assign n50581 = n1309 & ~n22645 ;
  assign n50582 = ~n1307 & n50581 ;
  assign n50583 = n50582 ^ n34528 ^ n13165 ;
  assign n50584 = n20168 | n50583 ;
  assign n50585 = ( ~n4994 & n9730 ) | ( ~n4994 & n13069 ) | ( n9730 & n13069 ) ;
  assign n50586 = n4613 & n7776 ;
  assign n50587 = ~n6213 & n50586 ;
  assign n50588 = n18015 | n50587 ;
  assign n50589 = n23014 & ~n50588 ;
  assign n50590 = n23785 & ~n50589 ;
  assign n50591 = n50590 ^ n3777 ^ 1'b0 ;
  assign n50592 = ( ~n38635 & n49368 ) | ( ~n38635 & n50591 ) | ( n49368 & n50591 ) ;
  assign n50593 = n25937 ^ n332 ^ 1'b0 ;
  assign n50594 = n50593 ^ n24617 ^ n20889 ;
  assign n50595 = ( n971 & n2638 ) | ( n971 & ~n42020 ) | ( n2638 & ~n42020 ) ;
  assign n50596 = n6406 ^ n3193 ^ n280 ;
  assign n50597 = n29814 & ~n50596 ;
  assign n50598 = n8666 & ~n10269 ;
  assign n50599 = n19868 & n50598 ;
  assign n50600 = n12756 | n50599 ;
  assign n50601 = n50597 & ~n50600 ;
  assign n50602 = n12498 | n33301 ;
  assign n50603 = n8536 | n50602 ;
  assign n50604 = n40343 ^ n15546 ^ 1'b0 ;
  assign n50605 = n50603 & ~n50604 ;
  assign n50606 = n14962 & n30552 ;
  assign n50607 = ~n50605 & n50606 ;
  assign n50608 = ~n6428 & n24008 ;
  assign n50609 = n21108 & n50608 ;
  assign n50610 = n3337 & ~n50517 ;
  assign n50611 = ( n2390 & ~n8354 ) | ( n2390 & n50610 ) | ( ~n8354 & n50610 ) ;
  assign n50612 = n50049 ^ n8267 ^ n3149 ;
  assign n50613 = n50612 ^ n38979 ^ n35231 ;
  assign n50614 = n1103 & ~n16417 ;
  assign n50615 = ( n3348 & ~n4902 ) | ( n3348 & n50614 ) | ( ~n4902 & n50614 ) ;
  assign n50616 = ( ~n21820 & n30788 ) | ( ~n21820 & n49543 ) | ( n30788 & n49543 ) ;
  assign n50617 = n41037 ^ n6877 ^ 1'b0 ;
  assign n50618 = n27419 & ~n50617 ;
  assign n50619 = ~n5066 & n41555 ;
  assign n50620 = n31125 & n50619 ;
  assign n50621 = ~n28205 & n33957 ;
  assign n50622 = ~n26493 & n50621 ;
  assign n50623 = n32256 ^ n30971 ^ n9286 ;
  assign n50624 = ( n8109 & n10022 ) | ( n8109 & ~n42638 ) | ( n10022 & ~n42638 ) ;
  assign n50625 = n50624 ^ n21316 ^ n9781 ;
  assign n50626 = n14842 ^ n8656 ^ n1275 ;
  assign n50627 = ( n11269 & ~n18939 ) | ( n11269 & n50626 ) | ( ~n18939 & n50626 ) ;
  assign n50628 = n42725 ^ n892 ^ 1'b0 ;
  assign n50629 = ~n10943 & n20059 ;
  assign n50630 = n50629 ^ n42190 ^ n12895 ;
  assign n50631 = n36149 ^ n22156 ^ 1'b0 ;
  assign n50632 = n3213 & ~n50631 ;
  assign n50633 = n50632 ^ n50283 ^ n21178 ;
  assign n50635 = n37347 ^ n16045 ^ 1'b0 ;
  assign n50636 = n7663 & ~n50635 ;
  assign n50634 = n14914 & n48295 ;
  assign n50637 = n50636 ^ n50634 ^ 1'b0 ;
  assign n50638 = ( n7274 & n11554 ) | ( n7274 & n30111 ) | ( n11554 & n30111 ) ;
  assign n50639 = n22127 & n50638 ;
  assign n50640 = ~n24425 & n50639 ;
  assign n50641 = n50640 ^ n12131 ^ 1'b0 ;
  assign n50642 = ~n18194 & n21112 ;
  assign n50643 = n50641 & n50642 ;
  assign n50644 = n12353 & n46093 ;
  assign n50645 = n7241 & n50644 ;
  assign n50646 = n21626 | n25329 ;
  assign n50647 = ( n12429 & n13232 ) | ( n12429 & ~n45194 ) | ( n13232 & ~n45194 ) ;
  assign n50648 = ~n26834 & n34170 ;
  assign n50649 = n50648 ^ n40064 ^ n29241 ;
  assign n50650 = ~n280 & n28366 ;
  assign n50651 = ~n5362 & n50650 ;
  assign n50652 = ( n2497 & n2885 ) | ( n2497 & ~n50651 ) | ( n2885 & ~n50651 ) ;
  assign n50653 = ( n5686 & n32854 ) | ( n5686 & n35317 ) | ( n32854 & n35317 ) ;
  assign n50654 = n23868 ^ n3559 ^ 1'b0 ;
  assign n50655 = n29056 ^ n5755 ^ 1'b0 ;
  assign n50656 = n17782 & n50655 ;
  assign n50657 = n28141 & ~n33001 ;
  assign n50658 = ~n50656 & n50657 ;
  assign n50659 = n9008 ^ n4199 ^ 1'b0 ;
  assign n50660 = ~n25058 & n50659 ;
  assign n50661 = n50660 ^ n46368 ^ n26076 ;
  assign n50662 = n50661 ^ n48852 ^ 1'b0 ;
  assign n50663 = n4859 & ~n50662 ;
  assign n50664 = ~n29091 & n30946 ;
  assign n50665 = ( ~n32575 & n35325 ) | ( ~n32575 & n50664 ) | ( n35325 & n50664 ) ;
  assign n50666 = ~n8018 & n50665 ;
  assign n50667 = n43720 ^ n39137 ^ n8299 ;
  assign n50674 = ~n5383 & n29019 ;
  assign n50675 = n50674 ^ n5998 ^ 1'b0 ;
  assign n50672 = ~n11948 & n14033 ;
  assign n50669 = n42368 ^ n20371 ^ 1'b0 ;
  assign n50670 = n7974 & ~n50669 ;
  assign n50671 = n50670 ^ n11793 ^ n6712 ;
  assign n50673 = n50672 ^ n50671 ^ n8770 ;
  assign n50668 = ( ~n15491 & n44768 ) | ( ~n15491 & n45819 ) | ( n44768 & n45819 ) ;
  assign n50676 = n50675 ^ n50673 ^ n50668 ;
  assign n50677 = ~n7108 & n23703 ;
  assign n50678 = n50677 ^ n43912 ^ n25331 ;
  assign n50679 = n46676 ^ n25502 ^ n11038 ;
  assign n50680 = ~n7092 & n27156 ;
  assign n50681 = n50680 ^ n20449 ^ 1'b0 ;
  assign n50682 = n16654 ^ n5599 ^ 1'b0 ;
  assign n50683 = n737 & n50682 ;
  assign n50684 = ( n17546 & ~n46920 ) | ( n17546 & n50683 ) | ( ~n46920 & n50683 ) ;
  assign n50685 = ~n41684 & n50684 ;
  assign n50686 = n7979 ^ n4566 ^ 1'b0 ;
  assign n50687 = n30375 & n50686 ;
  assign n50689 = n26621 ^ n12935 ^ 1'b0 ;
  assign n50690 = n4228 & n8588 ;
  assign n50691 = n50689 & n50690 ;
  assign n50688 = n16339 ^ n14478 ^ x243 ;
  assign n50692 = n50691 ^ n50688 ^ 1'b0 ;
  assign n50693 = n29121 & ~n29530 ;
  assign n50694 = n50693 ^ n8356 ^ 1'b0 ;
  assign n50695 = ( n5519 & ~n21809 ) | ( n5519 & n48046 ) | ( ~n21809 & n48046 ) ;
  assign n50696 = n50694 & n50695 ;
  assign n50697 = n6145 | n12122 ;
  assign n50698 = n41367 | n50697 ;
  assign n50699 = n17286 & ~n18048 ;
  assign n50700 = ( n13502 & ~n16866 ) | ( n13502 & n50699 ) | ( ~n16866 & n50699 ) ;
  assign n50701 = n10593 ^ n10223 ^ 1'b0 ;
  assign n50702 = n13196 & n17981 ;
  assign n50703 = n50702 ^ n3360 ^ 1'b0 ;
  assign n50704 = x95 & n33442 ;
  assign n50705 = n38918 & n50704 ;
  assign n50706 = n22094 | n44103 ;
  assign n50707 = n1239 | n50706 ;
  assign n50709 = n5444 ^ n657 ^ 1'b0 ;
  assign n50708 = n20529 ^ n7612 ^ 1'b0 ;
  assign n50710 = n50709 ^ n50708 ^ x16 ;
  assign n50711 = ~n35454 & n48096 ;
  assign n50712 = ~n50710 & n50711 ;
  assign n50713 = n19559 ^ n11301 ^ n3554 ;
  assign n50714 = ( n1995 & n40801 ) | ( n1995 & ~n50713 ) | ( n40801 & ~n50713 ) ;
  assign n50715 = n29019 ^ n20360 ^ 1'b0 ;
  assign n50716 = n21258 & ~n50715 ;
  assign n50717 = ~n11629 & n33537 ;
  assign n50718 = n50717 ^ n22473 ^ 1'b0 ;
  assign n50719 = n50716 & ~n50718 ;
  assign n50720 = n50719 ^ n38350 ^ 1'b0 ;
  assign n50721 = ( n31737 & ~n50714 ) | ( n31737 & n50720 ) | ( ~n50714 & n50720 ) ;
  assign n50722 = n29651 ^ n18201 ^ n8970 ;
  assign n50724 = n27497 ^ n20067 ^ 1'b0 ;
  assign n50723 = ( n3002 & n11553 ) | ( n3002 & ~n32133 ) | ( n11553 & ~n32133 ) ;
  assign n50725 = n50724 ^ n50723 ^ n23132 ;
  assign n50726 = n50725 ^ n967 ^ 1'b0 ;
  assign n50727 = n15217 & ~n50726 ;
  assign n50728 = ( n16577 & ~n50722 ) | ( n16577 & n50727 ) | ( ~n50722 & n50727 ) ;
  assign n50729 = n24144 ^ n13451 ^ 1'b0 ;
  assign n50730 = n50729 ^ n16968 ^ n13618 ;
  assign n50731 = ~n19077 & n40317 ;
  assign n50732 = n20562 & n28751 ;
  assign n50733 = n2965 & n50732 ;
  assign n50734 = ( ~n11106 & n30791 ) | ( ~n11106 & n50733 ) | ( n30791 & n50733 ) ;
  assign n50735 = ( ~n19208 & n27721 ) | ( ~n19208 & n50587 ) | ( n27721 & n50587 ) ;
  assign n50736 = ( x88 & ~n3301 ) | ( x88 & n39109 ) | ( ~n3301 & n39109 ) ;
  assign n50737 = n31342 | n50736 ;
  assign n50738 = n50737 ^ x75 ^ 1'b0 ;
  assign n50739 = ( ~n1432 & n31172 ) | ( ~n1432 & n50738 ) | ( n31172 & n50738 ) ;
  assign n50740 = ( ~n1858 & n9037 ) | ( ~n1858 & n14423 ) | ( n9037 & n14423 ) ;
  assign n50741 = n50739 & n50740 ;
  assign n50742 = n25964 ^ n10609 ^ 1'b0 ;
  assign n50743 = n4661 & ~n9785 ;
  assign n50744 = n29086 & n50743 ;
  assign n50745 = n50744 ^ n3010 ^ 1'b0 ;
  assign n50746 = n27029 & ~n35839 ;
  assign n50747 = n10585 | n50746 ;
  assign n50748 = ( n11585 & ~n45352 ) | ( n11585 & n48060 ) | ( ~n45352 & n48060 ) ;
  assign n50749 = n40463 | n42632 ;
  assign n50750 = n2422 & ~n25306 ;
  assign n50751 = ( n3163 & n50560 ) | ( n3163 & n50750 ) | ( n50560 & n50750 ) ;
  assign n50752 = n11704 ^ n5419 ^ n4344 ;
  assign n50753 = x85 & ~n28827 ;
  assign n50754 = n40903 | n44737 ;
  assign n50755 = n20768 & n40908 ;
  assign n50756 = n26542 | n50755 ;
  assign n50757 = n50756 ^ n49655 ^ 1'b0 ;
  assign n50758 = n17094 | n27835 ;
  assign n50759 = n4249 | n50758 ;
  assign n50760 = n33259 ^ n25723 ^ n1558 ;
  assign n50761 = n29604 ^ n8411 ^ 1'b0 ;
  assign n50762 = ( n22054 & ~n39257 ) | ( n22054 & n50761 ) | ( ~n39257 & n50761 ) ;
  assign n50763 = ~n20892 & n29955 ;
  assign n50764 = ( n18119 & ~n29855 ) | ( n18119 & n30010 ) | ( ~n29855 & n30010 ) ;
  assign n50765 = ~n41785 & n46875 ;
  assign n50766 = n37770 & ~n39114 ;
  assign n50767 = n43417 & n50766 ;
  assign n50768 = n8287 | n46127 ;
  assign n50769 = x220 | n50768 ;
  assign n50770 = n22396 | n39169 ;
  assign n50771 = n6606 ^ n4101 ^ n2260 ;
  assign n50772 = n43220 & n50771 ;
  assign n50773 = ~n50770 & n50772 ;
  assign n50774 = n50773 ^ n15850 ^ n14311 ;
  assign n50781 = n11186 ^ n10495 ^ 1'b0 ;
  assign n50782 = n3756 | n50781 ;
  assign n50783 = n50782 ^ n45910 ^ n17865 ;
  assign n50776 = n27453 ^ n5200 ^ 1'b0 ;
  assign n50777 = ~n30946 & n50776 ;
  assign n50778 = n26507 ^ n19995 ^ 1'b0 ;
  assign n50779 = ( ~n18950 & n50777 ) | ( ~n18950 & n50778 ) | ( n50777 & n50778 ) ;
  assign n50780 = ~n44344 & n50779 ;
  assign n50775 = ( n6173 & n16935 ) | ( n6173 & n27849 ) | ( n16935 & n27849 ) ;
  assign n50784 = n50783 ^ n50780 ^ n50775 ;
  assign n50785 = n24810 ^ n3583 ^ n327 ;
  assign n50786 = ( n26244 & ~n49157 ) | ( n26244 & n50785 ) | ( ~n49157 & n50785 ) ;
  assign n50787 = n23896 ^ n15579 ^ n10544 ;
  assign n50788 = n17737 ^ n7974 ^ 1'b0 ;
  assign n50789 = ( n29035 & n33758 ) | ( n29035 & n50788 ) | ( n33758 & n50788 ) ;
  assign n50790 = ~n19585 & n34932 ;
  assign n50791 = n47442 & ~n50790 ;
  assign n50792 = n1239 & ~n40293 ;
  assign n50793 = n11018 & n50792 ;
  assign n50794 = n24288 ^ n19077 ^ 1'b0 ;
  assign n50795 = n50794 ^ n48850 ^ 1'b0 ;
  assign n50796 = ~n3666 & n50795 ;
  assign n50797 = n45399 & n50796 ;
  assign n50798 = n12747 ^ n8371 ^ 1'b0 ;
  assign n50799 = n41114 & n48708 ;
  assign n50800 = n50798 & n50799 ;
  assign n50801 = n31417 & n43310 ;
  assign n50802 = n50801 ^ n49243 ^ 1'b0 ;
  assign n50803 = n9765 & ~n50535 ;
  assign n50804 = n24206 ^ n22421 ^ 1'b0 ;
  assign n50805 = n20835 ^ n1154 ^ 1'b0 ;
  assign n50806 = ( n1264 & n50804 ) | ( n1264 & ~n50805 ) | ( n50804 & ~n50805 ) ;
  assign n50807 = n47026 ^ n39767 ^ n2933 ;
  assign n50808 = ( n4706 & n19257 ) | ( n4706 & n50807 ) | ( n19257 & n50807 ) ;
  assign n50809 = n25288 ^ n18096 ^ n10116 ;
  assign n50810 = n50809 ^ n25290 ^ n9946 ;
  assign n50811 = n12478 ^ n1431 ^ 1'b0 ;
  assign n50812 = n9117 & ~n14960 ;
  assign n50813 = n50811 & n50812 ;
  assign n50814 = n40851 ^ n17922 ^ n7084 ;
  assign n50815 = n50813 & ~n50814 ;
  assign n50816 = n2417 & n4373 ;
  assign n50817 = n50816 ^ n6494 ^ 1'b0 ;
  assign n50818 = ( n9552 & ~n45316 ) | ( n9552 & n50817 ) | ( ~n45316 & n50817 ) ;
  assign n50819 = n19473 & n44142 ;
  assign n50820 = n50819 ^ n4100 ^ 1'b0 ;
  assign n50822 = n6269 | n28007 ;
  assign n50823 = n13806 | n50822 ;
  assign n50824 = n35156 & n50823 ;
  assign n50825 = ~n22229 & n50824 ;
  assign n50821 = n3394 & n18828 ;
  assign n50826 = n50825 ^ n50821 ^ 1'b0 ;
  assign n50827 = n5869 & ~n19823 ;
  assign n50828 = n12621 & n50827 ;
  assign n50829 = n17640 ^ n7919 ^ 1'b0 ;
  assign n50830 = ~n50828 & n50829 ;
  assign n50831 = n50830 ^ n1268 ^ 1'b0 ;
  assign n50832 = n45687 ^ n28019 ^ n3366 ;
  assign n50833 = n25964 | n48937 ;
  assign n50834 = n2623 & n50833 ;
  assign n50835 = n17677 ^ n4222 ^ 1'b0 ;
  assign n50836 = ~n46772 & n50835 ;
  assign n50837 = ( n10176 & n24106 ) | ( n10176 & ~n50836 ) | ( n24106 & ~n50836 ) ;
  assign n50838 = n23442 & ~n45013 ;
  assign n50839 = n50838 ^ n8847 ^ 1'b0 ;
  assign n50843 = ( n22396 & ~n27670 ) | ( n22396 & n46571 ) | ( ~n27670 & n46571 ) ;
  assign n50841 = n28522 ^ n19144 ^ x18 ;
  assign n50840 = n16480 | n18944 ;
  assign n50842 = n50841 ^ n50840 ^ 1'b0 ;
  assign n50844 = n50843 ^ n50842 ^ n48833 ;
  assign n50845 = n49189 ^ n5066 ^ 1'b0 ;
  assign n50846 = n16231 & n50845 ;
  assign n50847 = ~n2707 & n43538 ;
  assign n50848 = n50847 ^ n1261 ^ 1'b0 ;
  assign n50849 = n40385 & n50261 ;
  assign n50850 = ~n12072 & n50849 ;
  assign n50851 = n47152 ^ n6318 ^ 1'b0 ;
  assign n50852 = n23978 | n42920 ;
  assign n50853 = ( n6196 & n25408 ) | ( n6196 & ~n41836 ) | ( n25408 & ~n41836 ) ;
  assign n50854 = n9200 & n10101 ;
  assign n50855 = ~n2935 & n50854 ;
  assign n50856 = ( n6057 & n50853 ) | ( n6057 & ~n50855 ) | ( n50853 & ~n50855 ) ;
  assign n50858 = ( ~n7049 & n21133 ) | ( ~n7049 & n33319 ) | ( n21133 & n33319 ) ;
  assign n50859 = n50858 ^ n38612 ^ 1'b0 ;
  assign n50857 = ~n31213 & n31594 ;
  assign n50860 = n50859 ^ n50857 ^ n31688 ;
  assign n50865 = n21761 & n35109 ;
  assign n50864 = n5276 | n23340 ;
  assign n50862 = n32400 ^ n21160 ^ n14337 ;
  assign n50861 = ( n13813 & n39731 ) | ( n13813 & n41560 ) | ( n39731 & n41560 ) ;
  assign n50863 = n50862 ^ n50861 ^ n15586 ;
  assign n50866 = n50865 ^ n50864 ^ n50863 ;
  assign n50867 = ( ~n21956 & n36835 ) | ( ~n21956 & n42940 ) | ( n36835 & n42940 ) ;
  assign n50871 = n8030 & ~n12261 ;
  assign n50870 = n21864 ^ n14118 ^ 1'b0 ;
  assign n50868 = n23320 ^ n16777 ^ 1'b0 ;
  assign n50869 = n29348 | n50868 ;
  assign n50872 = n50871 ^ n50870 ^ n50869 ;
  assign n50873 = ( n9019 & n34250 ) | ( n9019 & n48083 ) | ( n34250 & n48083 ) ;
  assign n50874 = n50873 ^ n37220 ^ n690 ;
  assign n50875 = n50874 ^ n10960 ^ 1'b0 ;
  assign n50876 = n20663 & n50875 ;
  assign n50877 = ~n21505 & n35251 ;
  assign n50878 = n43585 & ~n50877 ;
  assign n50879 = n50878 ^ n26433 ^ 1'b0 ;
  assign n50880 = n42562 ^ n18353 ^ 1'b0 ;
  assign n50881 = n45774 & n50880 ;
  assign n50882 = n19626 & n50881 ;
  assign n50883 = n19705 ^ n15244 ^ n12616 ;
  assign n50884 = n27185 ^ n24064 ^ n1989 ;
  assign n50885 = ( ~n4756 & n16842 ) | ( ~n4756 & n50884 ) | ( n16842 & n50884 ) ;
  assign n50886 = ( ~n1307 & n5634 ) | ( ~n1307 & n19352 ) | ( n5634 & n19352 ) ;
  assign n50890 = n17635 ^ n14541 ^ 1'b0 ;
  assign n50887 = n7258 | n21292 ;
  assign n50888 = ( n6177 & n15004 ) | ( n6177 & n43610 ) | ( n15004 & n43610 ) ;
  assign n50889 = n50887 & ~n50888 ;
  assign n50891 = n50890 ^ n50889 ^ 1'b0 ;
  assign n50892 = ~n8533 & n40082 ;
  assign n50893 = ( ~n2800 & n32392 ) | ( ~n2800 & n50892 ) | ( n32392 & n50892 ) ;
  assign n50894 = n50893 ^ n46365 ^ n32809 ;
  assign n50895 = n41560 ^ n26135 ^ n24002 ;
  assign n50896 = ~n6744 & n19233 ;
  assign n50897 = n50896 ^ n1428 ^ 1'b0 ;
  assign n50898 = n16828 & n50897 ;
  assign n50899 = n12239 & n50898 ;
  assign n50900 = n50899 ^ n13384 ^ 1'b0 ;
  assign n50901 = n15962 & ~n50900 ;
  assign n50902 = ( n24139 & ~n50895 ) | ( n24139 & n50901 ) | ( ~n50895 & n50901 ) ;
  assign n50903 = n31968 & n34436 ;
  assign n50904 = n20419 & n50903 ;
  assign n50905 = n19283 ^ n4106 ^ 1'b0 ;
  assign n50906 = ~n9142 & n13760 ;
  assign n50907 = ~n3911 & n17307 ;
  assign n50908 = n50907 ^ n10692 ^ 1'b0 ;
  assign n50909 = n6982 ^ n1418 ^ 1'b0 ;
  assign n50910 = n35710 ^ n9386 ^ 1'b0 ;
  assign n50911 = n50910 ^ n38319 ^ n24626 ;
  assign n50912 = ( n9043 & n46411 ) | ( n9043 & n50911 ) | ( n46411 & n50911 ) ;
  assign n50913 = n21961 ^ n12326 ^ 1'b0 ;
  assign n50914 = ( n10057 & n28220 ) | ( n10057 & n50913 ) | ( n28220 & n50913 ) ;
  assign n50915 = ( n14161 & n42753 ) | ( n14161 & n50914 ) | ( n42753 & n50914 ) ;
  assign n50916 = ( ~n10732 & n27449 ) | ( ~n10732 & n46058 ) | ( n27449 & n46058 ) ;
  assign n50919 = ~n25303 & n34640 ;
  assign n50917 = n40941 ^ n19267 ^ 1'b0 ;
  assign n50918 = x100 & ~n50917 ;
  assign n50920 = n50919 ^ n50918 ^ 1'b0 ;
  assign n50921 = n19800 ^ n7598 ^ 1'b0 ;
  assign n50922 = n20249 & ~n38048 ;
  assign n50923 = n6615 | n21357 ;
  assign n50924 = n18846 | n50923 ;
  assign n50925 = n16515 & n22348 ;
  assign n50926 = n2546 & n50925 ;
  assign n50927 = n6501 & n16580 ;
  assign n50928 = n17517 & ~n38811 ;
  assign n50929 = n50928 ^ n33048 ^ 1'b0 ;
  assign n50930 = n50929 ^ n37846 ^ n25186 ;
  assign n50931 = ( n9566 & n10038 ) | ( n9566 & n30326 ) | ( n10038 & n30326 ) ;
  assign n50932 = ( ~n3677 & n12411 ) | ( ~n3677 & n20008 ) | ( n12411 & n20008 ) ;
  assign n50933 = n1978 & n50932 ;
  assign n50934 = n2512 | n10344 ;
  assign n50935 = n20331 & ~n50934 ;
  assign n50936 = ( n7111 & n18521 ) | ( n7111 & ~n19028 ) | ( n18521 & ~n19028 ) ;
  assign n50937 = n50936 ^ n39697 ^ 1'b0 ;
  assign n50938 = n6692 & n50937 ;
  assign n50939 = n50938 ^ n20449 ^ 1'b0 ;
  assign n50944 = n35612 ^ n18014 ^ 1'b0 ;
  assign n50940 = n14952 & n26290 ;
  assign n50941 = ~n17914 & n50940 ;
  assign n50942 = n22799 ^ n20168 ^ n14427 ;
  assign n50943 = n50941 | n50942 ;
  assign n50945 = n50944 ^ n50943 ^ 1'b0 ;
  assign n50948 = ( n1572 & n8462 ) | ( n1572 & ~n33344 ) | ( n8462 & ~n33344 ) ;
  assign n50947 = n23524 | n26232 ;
  assign n50949 = n50948 ^ n50947 ^ 1'b0 ;
  assign n50946 = n31946 ^ n30788 ^ n1257 ;
  assign n50950 = n50949 ^ n50946 ^ n9437 ;
  assign n50951 = n50950 ^ n6982 ^ 1'b0 ;
  assign n50952 = n47198 & ~n50951 ;
  assign n50953 = ~n3999 & n20748 ;
  assign n50954 = n35348 & n50953 ;
  assign n50955 = ( n22028 & n46829 ) | ( n22028 & ~n50954 ) | ( n46829 & ~n50954 ) ;
  assign n50956 = n36106 ^ n8477 ^ 1'b0 ;
  assign n50957 = ~n43704 & n50956 ;
  assign n50958 = n50957 ^ n23501 ^ n1278 ;
  assign n50959 = n394 & ~n50958 ;
  assign n50960 = ( n20761 & n22434 ) | ( n20761 & n43281 ) | ( n22434 & n43281 ) ;
  assign n50963 = n19245 ^ n4662 ^ n3598 ;
  assign n50964 = n9587 | n50963 ;
  assign n50965 = n38152 | n50964 ;
  assign n50961 = ~n652 & n24925 ;
  assign n50962 = n50961 ^ n30801 ^ 1'b0 ;
  assign n50966 = n50965 ^ n50962 ^ n9535 ;
  assign n50967 = ( n15934 & n20932 ) | ( n15934 & n49075 ) | ( n20932 & n49075 ) ;
  assign n50968 = n735 & ~n29293 ;
  assign n50969 = n30067 & n50968 ;
  assign n50970 = n42322 & n50969 ;
  assign n50971 = n25564 & ~n41757 ;
  assign n50972 = ~n2591 & n33459 ;
  assign n50973 = n50972 ^ n31114 ^ n12280 ;
  assign n50974 = ( n2142 & ~n28411 ) | ( n2142 & n31799 ) | ( ~n28411 & n31799 ) ;
  assign n50975 = n50974 ^ n28382 ^ n21606 ;
  assign n50976 = n27015 ^ n7365 ^ n1150 ;
  assign n50977 = n5205 & ~n45247 ;
  assign n50978 = ( n15876 & n28537 ) | ( n15876 & n50977 ) | ( n28537 & n50977 ) ;
  assign n50979 = n48872 ^ n28152 ^ n26139 ;
  assign n50980 = n37861 ^ n22845 ^ n9780 ;
  assign n50981 = n32941 & ~n50980 ;
  assign n50982 = ( n569 & n21342 ) | ( n569 & ~n21822 ) | ( n21342 & ~n21822 ) ;
  assign n50983 = ~n15718 & n50982 ;
  assign n50984 = n25396 | n27070 ;
  assign n50985 = n50984 ^ n44462 ^ 1'b0 ;
  assign n50986 = n23385 ^ n3111 ^ 1'b0 ;
  assign n50987 = n29294 & ~n50986 ;
  assign n50988 = n50987 ^ n29614 ^ 1'b0 ;
  assign n50989 = ~n7542 & n19436 ;
  assign n50990 = n32665 & n50989 ;
  assign n50991 = n50990 ^ n47081 ^ n42625 ;
  assign n50992 = n7846 | n20113 ;
  assign n50993 = n36035 ^ n30307 ^ n3740 ;
  assign n50994 = ( ~n4038 & n18560 ) | ( ~n4038 & n50993 ) | ( n18560 & n50993 ) ;
  assign n50995 = n9121 & n50994 ;
  assign n50996 = n25081 & n41608 ;
  assign n50997 = n50996 ^ n17861 ^ 1'b0 ;
  assign n50998 = n50997 ^ n48822 ^ n20662 ;
  assign n50999 = n30139 ^ n26188 ^ n14046 ;
  assign n51000 = n46999 ^ n10433 ^ 1'b0 ;
  assign n51001 = n16528 | n51000 ;
  assign n51002 = n51001 ^ n27514 ^ n1276 ;
  assign n51003 = n12551 ^ n9556 ^ n9271 ;
  assign n51004 = n21151 | n51003 ;
  assign n51005 = n24855 ^ n1336 ^ 1'b0 ;
  assign n51006 = n29314 | n51005 ;
  assign n51007 = n51006 ^ n27028 ^ 1'b0 ;
  assign n51008 = n8188 | n51007 ;
  assign n51009 = ~n12838 & n37672 ;
  assign n51010 = n51008 & n51009 ;
  assign n51011 = n3854 ^ n2110 ^ 1'b0 ;
  assign n51012 = ~n47899 & n51011 ;
  assign n51013 = ( n28543 & ~n39883 ) | ( n28543 & n41019 ) | ( ~n39883 & n41019 ) ;
  assign n51014 = n47835 ^ n33932 ^ n2602 ;
  assign n51015 = n11146 & ~n24480 ;
  assign n51016 = n1551 & ~n31701 ;
  assign n51017 = n2210 ^ n935 ^ 1'b0 ;
  assign n51018 = n34952 | n51017 ;
  assign n51019 = n16367 & n24104 ;
  assign n51020 = n36814 ^ n14820 ^ n6314 ;
  assign n51021 = n51020 ^ n9505 ^ n9406 ;
  assign n51023 = n8863 & n35417 ;
  assign n51022 = n6560 | n9003 ;
  assign n51024 = n51023 ^ n51022 ^ 1'b0 ;
  assign n51025 = ( n51019 & ~n51021 ) | ( n51019 & n51024 ) | ( ~n51021 & n51024 ) ;
  assign n51026 = n20691 & n33927 ;
  assign n51027 = ~n12673 & n51026 ;
  assign n51028 = ( n14004 & n16242 ) | ( n14004 & ~n16424 ) | ( n16242 & ~n16424 ) ;
  assign n51029 = n51028 ^ n6611 ^ n2984 ;
  assign n51030 = n2688 & n15349 ;
  assign n51031 = n51030 ^ x187 ^ 1'b0 ;
  assign n51032 = n41700 | n51031 ;
  assign n51033 = n51029 | n51032 ;
  assign n51034 = n20894 ^ n6328 ^ 1'b0 ;
  assign n51035 = n41298 & n51034 ;
  assign n51036 = n15526 ^ n9654 ^ x13 ;
  assign n51037 = n17501 ^ n16411 ^ 1'b0 ;
  assign n51038 = n51036 & n51037 ;
  assign n51039 = ( ~n5544 & n12825 ) | ( ~n5544 & n18386 ) | ( n12825 & n18386 ) ;
  assign n51040 = ( n10077 & n18455 ) | ( n10077 & ~n51039 ) | ( n18455 & ~n51039 ) ;
  assign n51041 = ( n1706 & n5954 ) | ( n1706 & n25378 ) | ( n5954 & n25378 ) ;
  assign n51042 = ( n13253 & ~n20232 ) | ( n13253 & n30123 ) | ( ~n20232 & n30123 ) ;
  assign n51043 = n4587 & n23238 ;
  assign n51044 = ( ~n51041 & n51042 ) | ( ~n51041 & n51043 ) | ( n51042 & n51043 ) ;
  assign n51045 = n5648 & ~n51044 ;
  assign n51046 = n23317 & ~n50854 ;
  assign n51047 = n4468 | n51046 ;
  assign n51048 = n26343 & ~n51047 ;
  assign n51049 = ~n33687 & n51048 ;
  assign n51050 = n22532 ^ n13290 ^ 1'b0 ;
  assign n51051 = n8301 & n8465 ;
  assign n51052 = n51051 ^ n16247 ^ 1'b0 ;
  assign n51053 = n51052 ^ n3193 ^ 1'b0 ;
  assign n51054 = n47640 ^ n44094 ^ 1'b0 ;
  assign n51055 = n51054 ^ n8903 ^ 1'b0 ;
  assign n51056 = n42384 ^ n12208 ^ 1'b0 ;
  assign n51057 = ~n697 & n51056 ;
  assign n51058 = n15121 ^ n12952 ^ 1'b0 ;
  assign n51059 = n18560 | n51058 ;
  assign n51060 = ( n8917 & n24262 ) | ( n8917 & n27032 ) | ( n24262 & n27032 ) ;
  assign n51061 = n46555 ^ x208 ^ 1'b0 ;
  assign n51062 = n11467 ^ n5216 ^ 1'b0 ;
  assign n51063 = ( n38500 & n46478 ) | ( n38500 & ~n51062 ) | ( n46478 & ~n51062 ) ;
  assign n51064 = ( n1489 & n18310 ) | ( n1489 & n51063 ) | ( n18310 & n51063 ) ;
  assign n51065 = n15678 | n51064 ;
  assign n51066 = n23802 ^ n21154 ^ x117 ;
  assign n51067 = ( n18430 & ~n39188 ) | ( n18430 & n51066 ) | ( ~n39188 & n51066 ) ;
  assign n51068 = ( n3596 & ~n13791 ) | ( n3596 & n19937 ) | ( ~n13791 & n19937 ) ;
  assign n51069 = ~n31468 & n36564 ;
  assign n51070 = ( n31409 & n51068 ) | ( n31409 & n51069 ) | ( n51068 & n51069 ) ;
  assign n51071 = n24253 ^ n21326 ^ 1'b0 ;
  assign n51072 = n34832 & ~n51071 ;
  assign n51073 = n6665 & ~n41654 ;
  assign n51074 = n51073 ^ n20102 ^ 1'b0 ;
  assign n51075 = n2010 | n15897 ;
  assign n51076 = ( n4946 & n12739 ) | ( n4946 & ~n45570 ) | ( n12739 & ~n45570 ) ;
  assign n51077 = n1473 & n29966 ;
  assign n51078 = n51076 & n51077 ;
  assign n51080 = n21778 ^ n10429 ^ x84 ;
  assign n51081 = n51080 ^ n25845 ^ n4032 ;
  assign n51082 = n31775 & n51081 ;
  assign n51079 = n26684 ^ n3875 ^ 1'b0 ;
  assign n51083 = n51082 ^ n51079 ^ n39754 ;
  assign n51084 = n34382 ^ n25967 ^ 1'b0 ;
  assign n51085 = n13556 & n51084 ;
  assign n51086 = n7995 & ~n28761 ;
  assign n51087 = n46043 ^ n21132 ^ 1'b0 ;
  assign n51088 = ( ~n2318 & n51086 ) | ( ~n2318 & n51087 ) | ( n51086 & n51087 ) ;
  assign n51089 = n7381 & ~n50794 ;
  assign n51090 = ( n28934 & n44478 ) | ( n28934 & ~n51089 ) | ( n44478 & ~n51089 ) ;
  assign n51091 = ( ~n19368 & n20227 ) | ( ~n19368 & n51090 ) | ( n20227 & n51090 ) ;
  assign n51092 = ( n1783 & ~n12431 ) | ( n1783 & n22729 ) | ( ~n12431 & n22729 ) ;
  assign n51093 = n995 & ~n24750 ;
  assign n51094 = n51092 & n51093 ;
  assign n51095 = n37067 ^ n16233 ^ 1'b0 ;
  assign n51096 = n18328 & n51095 ;
  assign n51097 = ( n16119 & n19356 ) | ( n16119 & n24168 ) | ( n19356 & n24168 ) ;
  assign n51098 = n51097 ^ n38697 ^ n32646 ;
  assign n51099 = n1656 & n51098 ;
  assign n51100 = n8564 & n51099 ;
  assign n51101 = n15312 & ~n21190 ;
  assign n51102 = n51101 ^ n15036 ^ 1'b0 ;
  assign n51103 = n36531 ^ n2948 ^ 1'b0 ;
  assign n51104 = n44744 & ~n51103 ;
  assign n51105 = n22010 ^ n20724 ^ n13345 ;
  assign n51106 = n51105 ^ n7782 ^ 1'b0 ;
  assign n51107 = n11474 | n36953 ;
  assign n51108 = n3408 | n51107 ;
  assign n51109 = n28144 & ~n51108 ;
  assign n51110 = n17713 ^ n10220 ^ 1'b0 ;
  assign n51111 = n51109 | n51110 ;
  assign n51112 = n51111 ^ n48380 ^ n15155 ;
  assign n51113 = n18215 & ~n43011 ;
  assign n51114 = n12850 & ~n51113 ;
  assign n51115 = ( n6864 & ~n20338 ) | ( n6864 & n21217 ) | ( ~n20338 & n21217 ) ;
  assign n51116 = ( n6193 & n23540 ) | ( n6193 & n51115 ) | ( n23540 & n51115 ) ;
  assign n51117 = n36449 ^ n11716 ^ 1'b0 ;
  assign n51118 = n47899 ^ n13803 ^ n10824 ;
  assign n51119 = n19258 ^ n19247 ^ 1'b0 ;
  assign n51120 = n36754 ^ n29044 ^ n18201 ;
  assign n51121 = n2145 & n8599 ;
  assign n51122 = n51121 ^ n38438 ^ 1'b0 ;
  assign n51123 = ~n25274 & n51122 ;
  assign n51124 = n51123 ^ n28909 ^ 1'b0 ;
  assign n51125 = ~n51120 & n51124 ;
  assign n51126 = n35414 ^ n2610 ^ 1'b0 ;
  assign n51128 = ~n12456 & n15793 ;
  assign n51127 = n2806 & ~n16391 ;
  assign n51129 = n51128 ^ n51127 ^ 1'b0 ;
  assign n51130 = ( n24693 & n39782 ) | ( n24693 & n51129 ) | ( n39782 & n51129 ) ;
  assign n51131 = n40704 ^ n38880 ^ n25956 ;
  assign n51132 = n26716 & n38365 ;
  assign n51133 = n51132 ^ n16153 ^ 1'b0 ;
  assign n51134 = n51133 ^ n37802 ^ n8842 ;
  assign n51135 = n9051 & n29709 ;
  assign n51136 = ~n24266 & n51135 ;
  assign n51137 = n45244 | n51136 ;
  assign n51138 = ~n12515 & n20429 ;
  assign n51140 = ( n7133 & ~n23066 ) | ( n7133 & n42843 ) | ( ~n23066 & n42843 ) ;
  assign n51141 = n51140 ^ n16538 ^ n4822 ;
  assign n51139 = ~n9425 & n24612 ;
  assign n51142 = n51141 ^ n51139 ^ 1'b0 ;
  assign n51143 = n22390 & ~n29360 ;
  assign n51144 = ~n21320 & n37575 ;
  assign n51145 = n14902 & n51144 ;
  assign n51146 = n46977 ^ n37644 ^ n33229 ;
  assign n51147 = n25326 & ~n31957 ;
  assign n51148 = n45461 ^ n21041 ^ 1'b0 ;
  assign n51149 = n21014 ^ n14271 ^ n8659 ;
  assign n51150 = n6737 | n13969 ;
  assign n51151 = ( n5883 & ~n16679 ) | ( n5883 & n36370 ) | ( ~n16679 & n36370 ) ;
  assign n51152 = n51151 ^ n11840 ^ 1'b0 ;
  assign n51153 = ~n16962 & n45464 ;
  assign n51154 = n51153 ^ n46320 ^ 1'b0 ;
  assign n51155 = ~n626 & n51154 ;
  assign n51156 = n12676 & n31633 ;
  assign n51157 = n34753 ^ n15767 ^ n10918 ;
  assign n51158 = ~n1230 & n25185 ;
  assign n51161 = n3501 & ~n4115 ;
  assign n51162 = n17264 | n51161 ;
  assign n51159 = ~n5342 & n10196 ;
  assign n51160 = n37677 & n51159 ;
  assign n51163 = n51162 ^ n51160 ^ n1225 ;
  assign n51164 = n41235 ^ n37828 ^ n14172 ;
  assign n51165 = n51164 ^ n36578 ^ n2404 ;
  assign n51166 = n40234 ^ n15960 ^ 1'b0 ;
  assign n51167 = ( n18404 & n45540 ) | ( n18404 & ~n51166 ) | ( n45540 & ~n51166 ) ;
  assign n51168 = n2773 | n13345 ;
  assign n51169 = n51168 ^ n10521 ^ 1'b0 ;
  assign n51170 = n51169 ^ n45563 ^ 1'b0 ;
  assign n51171 = ~n37074 & n51170 ;
  assign n51172 = n26991 ^ n26595 ^ 1'b0 ;
  assign n51173 = n22035 & ~n51172 ;
  assign n51174 = n50167 ^ n38049 ^ 1'b0 ;
  assign n51175 = ~n15499 & n35396 ;
  assign n51176 = ~n51174 & n51175 ;
  assign n51177 = n39428 | n47394 ;
  assign n51178 = n51177 ^ n49765 ^ 1'b0 ;
  assign n51179 = n20136 ^ n14102 ^ 1'b0 ;
  assign n51180 = ( n4539 & n12855 ) | ( n4539 & n13810 ) | ( n12855 & n13810 ) ;
  assign n51181 = n51180 ^ n28466 ^ n13148 ;
  assign n51182 = ( n20831 & ~n39046 ) | ( n20831 & n51181 ) | ( ~n39046 & n51181 ) ;
  assign n51183 = n40347 & ~n51182 ;
  assign n51184 = ~n51179 & n51183 ;
  assign n51185 = ( n6642 & n15390 ) | ( n6642 & ~n15622 ) | ( n15390 & ~n15622 ) ;
  assign n51186 = n39032 ^ n6923 ^ 1'b0 ;
  assign n51187 = ~n16054 & n51186 ;
  assign n51188 = ~n20160 & n51187 ;
  assign n51189 = ( n2530 & n5177 ) | ( n2530 & n10327 ) | ( n5177 & n10327 ) ;
  assign n51190 = ( x52 & n9546 ) | ( x52 & ~n51189 ) | ( n9546 & ~n51189 ) ;
  assign n51191 = ( n51185 & n51188 ) | ( n51185 & ~n51190 ) | ( n51188 & ~n51190 ) ;
  assign n51192 = n34163 | n45555 ;
  assign n51193 = n50353 ^ n36881 ^ n5835 ;
  assign n51194 = ~n14140 & n20511 ;
  assign n51195 = ( n23578 & n43994 ) | ( n23578 & ~n51194 ) | ( n43994 & ~n51194 ) ;
  assign n51196 = n27795 ^ n26795 ^ 1'b0 ;
  assign n51197 = n37340 & ~n51196 ;
  assign n51198 = n7256 ^ n2195 ^ 1'b0 ;
  assign n51199 = n51198 ^ n28694 ^ 1'b0 ;
  assign n51200 = n16936 | n51199 ;
  assign n51201 = n44491 ^ n30307 ^ n13813 ;
  assign n51202 = ~n34869 & n51201 ;
  assign n51203 = n29519 | n32992 ;
  assign n51204 = n51203 ^ n30677 ^ 1'b0 ;
  assign n51205 = n29642 ^ n16739 ^ n3408 ;
  assign n51206 = n51205 ^ n27201 ^ n11886 ;
  assign n51207 = n7815 | n27610 ;
  assign n51208 = n51207 ^ n48305 ^ 1'b0 ;
  assign n51209 = ( ~n12516 & n20962 ) | ( ~n12516 & n51208 ) | ( n20962 & n51208 ) ;
  assign n51210 = n10223 | n33606 ;
  assign n51211 = n39080 ^ n3358 ^ 1'b0 ;
  assign n51212 = ~n2932 & n8877 ;
  assign n51213 = n51212 ^ n14801 ^ 1'b0 ;
  assign n51214 = ( n7490 & n21093 ) | ( n7490 & ~n51213 ) | ( n21093 & ~n51213 ) ;
  assign n51216 = ( n6208 & n8671 ) | ( n6208 & ~n27437 ) | ( n8671 & ~n27437 ) ;
  assign n51215 = n39448 ^ n17822 ^ n10391 ;
  assign n51217 = n51216 ^ n51215 ^ n49913 ;
  assign n51218 = ~n32501 & n41358 ;
  assign n51219 = n36372 & n51218 ;
  assign n51222 = n11986 & n38000 ;
  assign n51220 = n15542 ^ x102 ^ 1'b0 ;
  assign n51221 = ~n5140 & n51220 ;
  assign n51223 = n51222 ^ n51221 ^ 1'b0 ;
  assign n51224 = n42540 ^ n21930 ^ 1'b0 ;
  assign n51225 = n12653 | n51224 ;
  assign n51226 = n21694 ^ n9263 ^ n6239 ;
  assign n51227 = ( ~n4263 & n32242 ) | ( ~n4263 & n51226 ) | ( n32242 & n51226 ) ;
  assign n51228 = ( n9963 & n11924 ) | ( n9963 & ~n20938 ) | ( n11924 & ~n20938 ) ;
  assign n51229 = n29036 ^ n6647 ^ 1'b0 ;
  assign n51230 = n565 | n20447 ;
  assign n51231 = n51230 ^ n35870 ^ 1'b0 ;
  assign n51232 = ~n1428 & n6611 ;
  assign n51233 = n51232 ^ n41374 ^ n16161 ;
  assign n51234 = ( n6072 & n51231 ) | ( n6072 & ~n51233 ) | ( n51231 & ~n51233 ) ;
  assign n51235 = ( n16706 & n33619 ) | ( n16706 & n43222 ) | ( n33619 & n43222 ) ;
  assign n51236 = n5739 | n16103 ;
  assign n51237 = n8572 & n9205 ;
  assign n51238 = ~n8420 & n51237 ;
  assign n51239 = ( ~n2680 & n4965 ) | ( ~n2680 & n38427 ) | ( n4965 & n38427 ) ;
  assign n51240 = ~n37752 & n51239 ;
  assign n51241 = n51238 & n51240 ;
  assign n51242 = n1826 | n38287 ;
  assign n51243 = n47109 & ~n51242 ;
  assign n51248 = ( n7137 & n17451 ) | ( n7137 & n20583 ) | ( n17451 & n20583 ) ;
  assign n51249 = n20023 & ~n51248 ;
  assign n51250 = n19492 & n51249 ;
  assign n51244 = n36449 ^ n9146 ^ 1'b0 ;
  assign n51245 = ~n27033 & n51244 ;
  assign n51246 = n51245 ^ n16857 ^ n10948 ;
  assign n51247 = n5514 | n51246 ;
  assign n51251 = n51250 ^ n51247 ^ 1'b0 ;
  assign n51252 = n6317 & ~n9457 ;
  assign n51253 = n51252 ^ n15059 ^ 1'b0 ;
  assign n51254 = n51253 ^ n28788 ^ n6711 ;
  assign n51255 = x144 & ~n3307 ;
  assign n51256 = n51255 ^ n2162 ^ 1'b0 ;
  assign n51257 = n51256 ^ n45466 ^ n4348 ;
  assign n51258 = ( n6015 & n15104 ) | ( n6015 & n39938 ) | ( n15104 & n39938 ) ;
  assign n51259 = n48118 ^ n23034 ^ n5152 ;
  assign n51260 = ( n17245 & n24770 ) | ( n17245 & n43701 ) | ( n24770 & n43701 ) ;
  assign n51261 = n28372 ^ n26847 ^ n11197 ;
  assign n51262 = n2834 ^ n999 ^ 1'b0 ;
  assign n51263 = n51262 ^ n35244 ^ 1'b0 ;
  assign n51264 = n43675 & n51263 ;
  assign n51265 = ( ~n1802 & n4283 ) | ( ~n1802 & n12285 ) | ( n4283 & n12285 ) ;
  assign n51266 = n47976 ^ n16119 ^ 1'b0 ;
  assign n51267 = n51265 & ~n51266 ;
  assign n51268 = n5069 & n45905 ;
  assign n51269 = ( n10935 & n22473 ) | ( n10935 & ~n28078 ) | ( n22473 & ~n28078 ) ;
  assign n51270 = ( n4782 & ~n25338 ) | ( n4782 & n32322 ) | ( ~n25338 & n32322 ) ;
  assign n51271 = n20873 ^ n20147 ^ 1'b0 ;
  assign n51272 = n40902 & n51271 ;
  assign n51273 = ( ~n7443 & n13529 ) | ( ~n7443 & n51272 ) | ( n13529 & n51272 ) ;
  assign n51274 = n51270 | n51273 ;
  assign n51275 = ( n12442 & n14619 ) | ( n12442 & n19190 ) | ( n14619 & n19190 ) ;
  assign n51276 = n14789 ^ n12451 ^ n8876 ;
  assign n51277 = ( n38987 & ~n47846 ) | ( n38987 & n51276 ) | ( ~n47846 & n51276 ) ;
  assign n51278 = n5695 & n24578 ;
  assign n51279 = n51278 ^ n21119 ^ 1'b0 ;
  assign n51280 = ( ~n8086 & n45687 ) | ( ~n8086 & n51279 ) | ( n45687 & n51279 ) ;
  assign n51281 = n51280 ^ n27922 ^ 1'b0 ;
  assign n51282 = ( ~n25199 & n28492 ) | ( ~n25199 & n51021 ) | ( n28492 & n51021 ) ;
  assign n51283 = n40090 ^ n403 ^ 1'b0 ;
  assign n51284 = n51283 ^ n25973 ^ n25061 ;
  assign n51285 = n51284 ^ n6261 ^ 1'b0 ;
  assign n51286 = n21576 & n51285 ;
  assign n51287 = n28764 ^ n20212 ^ 1'b0 ;
  assign n51288 = n30457 | n51287 ;
  assign n51289 = ( n18020 & n19913 ) | ( n18020 & ~n43720 ) | ( n19913 & ~n43720 ) ;
  assign n51290 = n21268 ^ n16773 ^ n9595 ;
  assign n51291 = n51290 ^ n46900 ^ n14380 ;
  assign n51292 = n23449 | n51291 ;
  assign n51293 = n51289 | n51292 ;
  assign n51294 = n7616 | n10953 ;
  assign n51295 = n51294 ^ n7612 ^ 1'b0 ;
  assign n51296 = n15687 & ~n20887 ;
  assign n51297 = n36095 & n51296 ;
  assign n51298 = n1387 | n51297 ;
  assign n51299 = n51298 ^ n49404 ^ 1'b0 ;
  assign n51300 = n51299 ^ n38987 ^ 1'b0 ;
  assign n51301 = n44352 & n51300 ;
  assign n51302 = n7359 | n23200 ;
  assign n51303 = n46661 | n51302 ;
  assign n51304 = n51303 ^ n26285 ^ 1'b0 ;
  assign n51308 = ( n2555 & ~n10582 ) | ( n2555 & n22505 ) | ( ~n10582 & n22505 ) ;
  assign n51307 = n37297 ^ n17261 ^ n2791 ;
  assign n51309 = n51308 ^ n51307 ^ n5853 ;
  assign n51305 = n23381 & ~n26093 ;
  assign n51306 = ~n28365 & n51305 ;
  assign n51310 = n51309 ^ n51306 ^ 1'b0 ;
  assign n51311 = n38024 ^ n16249 ^ n15163 ;
  assign n51312 = n49997 ^ n20034 ^ 1'b0 ;
  assign n51313 = ( n4601 & ~n46212 ) | ( n4601 & n51312 ) | ( ~n46212 & n51312 ) ;
  assign n51314 = n43073 ^ n31807 ^ 1'b0 ;
  assign n51315 = n29914 ^ n9781 ^ 1'b0 ;
  assign n51316 = n7157 & n29227 ;
  assign n51317 = n51316 ^ n26363 ^ 1'b0 ;
  assign n51318 = n29966 ^ n10539 ^ 1'b0 ;
  assign n51319 = ( n1481 & n5258 ) | ( n1481 & ~n14568 ) | ( n5258 & ~n14568 ) ;
  assign n51320 = n51319 ^ n23858 ^ n9139 ;
  assign n51321 = n51318 & ~n51320 ;
  assign n51324 = n6372 | n13144 ;
  assign n51325 = n3860 & ~n51324 ;
  assign n51322 = n2748 | n9179 ;
  assign n51323 = n51322 ^ n32570 ^ n17093 ;
  assign n51326 = n51325 ^ n51323 ^ n1606 ;
  assign n51327 = n15360 & ~n27628 ;
  assign n51328 = n45866 ^ n43023 ^ n16760 ;
  assign n51329 = n24275 ^ n10372 ^ n6718 ;
  assign n51330 = n22205 | n42242 ;
  assign n51331 = n51330 ^ n8955 ^ 1'b0 ;
  assign n51332 = ( ~n12446 & n51329 ) | ( ~n12446 & n51331 ) | ( n51329 & n51331 ) ;
  assign n51333 = ( n11009 & n21165 ) | ( n11009 & ~n51332 ) | ( n21165 & ~n51332 ) ;
  assign n51334 = n10550 & ~n46963 ;
  assign n51335 = n28241 & n51334 ;
  assign n51336 = n15284 | n45771 ;
  assign n51337 = n51336 ^ n22781 ^ 1'b0 ;
  assign n51338 = n2766 & ~n47895 ;
  assign n51339 = n2207 | n12714 ;
  assign n51340 = n1166 | n51339 ;
  assign n51341 = n17922 | n51340 ;
  assign n51342 = ( n9526 & n20031 ) | ( n9526 & n43430 ) | ( n20031 & n43430 ) ;
  assign n51343 = n3499 & ~n35868 ;
  assign n51344 = ~n2452 & n3234 ;
  assign n51345 = ( n9756 & n25303 ) | ( n9756 & ~n35618 ) | ( n25303 & ~n35618 ) ;
  assign n51348 = n43317 ^ n2176 ^ 1'b0 ;
  assign n51346 = ~n20114 & n33067 ;
  assign n51347 = n24265 & n51346 ;
  assign n51349 = n51348 ^ n51347 ^ n50396 ;
  assign n51350 = n16864 & ~n34694 ;
  assign n51351 = n1942 & n51350 ;
  assign n51352 = n43511 | n50632 ;
  assign n51353 = n1753 & n18644 ;
  assign n51354 = n3668 & ~n51353 ;
  assign n51355 = n17196 | n51354 ;
  assign n51356 = n18377 | n51355 ;
  assign n51357 = ( ~n6855 & n47157 ) | ( ~n6855 & n49619 ) | ( n47157 & n49619 ) ;
  assign n51358 = n11104 | n51357 ;
  assign n51359 = n51358 ^ n12162 ^ 1'b0 ;
  assign n51360 = n51359 ^ n48266 ^ 1'b0 ;
  assign n51361 = n34413 & ~n51360 ;
  assign n51362 = ~n51356 & n51361 ;
  assign n51363 = n894 & ~n51253 ;
  assign n51364 = n51363 ^ n27954 ^ 1'b0 ;
  assign n51365 = ( n15090 & n42604 ) | ( n15090 & ~n51364 ) | ( n42604 & ~n51364 ) ;
  assign n51366 = n29582 ^ n10345 ^ 1'b0 ;
  assign n51367 = n47578 ^ n29965 ^ 1'b0 ;
  assign n51371 = n10817 ^ n8254 ^ 1'b0 ;
  assign n51368 = n14770 ^ n7644 ^ 1'b0 ;
  assign n51369 = n33157 & ~n51368 ;
  assign n51370 = n51369 ^ n13978 ^ n6227 ;
  assign n51372 = n51371 ^ n51370 ^ n7821 ;
  assign n51373 = n29272 ^ n19133 ^ n7696 ;
  assign n51374 = n30078 | n34644 ;
  assign n51375 = ( n12695 & ~n29371 ) | ( n12695 & n51374 ) | ( ~n29371 & n51374 ) ;
  assign n51376 = ( ~x19 & n10641 ) | ( ~x19 & n14006 ) | ( n10641 & n14006 ) ;
  assign n51377 = n51376 ^ n49149 ^ 1'b0 ;
  assign n51378 = n25107 & ~n51377 ;
  assign n51379 = ~n6523 & n51173 ;
  assign n51380 = n51379 ^ n20404 ^ 1'b0 ;
  assign n51381 = ( ~n14070 & n28228 ) | ( ~n14070 & n36191 ) | ( n28228 & n36191 ) ;
  assign n51382 = n15284 ^ n8820 ^ 1'b0 ;
  assign n51383 = x63 & ~n51382 ;
  assign n51384 = n51383 ^ n27848 ^ n23135 ;
  assign n51385 = n6529 | n39776 ;
  assign n51386 = ( n17669 & ~n33177 ) | ( n17669 & n43045 ) | ( ~n33177 & n43045 ) ;
  assign n51389 = n20519 & n22703 ;
  assign n51390 = n51389 ^ n37227 ^ 1'b0 ;
  assign n51387 = n17297 ^ n13867 ^ n3612 ;
  assign n51388 = ( n20432 & n29112 ) | ( n20432 & ~n51387 ) | ( n29112 & ~n51387 ) ;
  assign n51391 = n51390 ^ n51388 ^ n7456 ;
  assign n51392 = ~n27904 & n34146 ;
  assign n51393 = n343 & n19390 ;
  assign n51394 = ~n17023 & n51393 ;
  assign n51395 = n22248 | n32193 ;
  assign n51396 = n21352 & n38353 ;
  assign n51397 = n18090 ^ n11849 ^ 1'b0 ;
  assign n51398 = ~n3831 & n51397 ;
  assign n51399 = n425 & n51398 ;
  assign n51400 = ~n7008 & n51399 ;
  assign n51401 = n28078 ^ n21099 ^ n16496 ;
  assign n51402 = n39381 ^ x254 ^ 1'b0 ;
  assign n51403 = ( ~n10928 & n46211 ) | ( ~n10928 & n51402 ) | ( n46211 & n51402 ) ;
  assign n51404 = n20774 ^ n6878 ^ 1'b0 ;
  assign n51405 = n10561 ^ n7379 ^ 1'b0 ;
  assign n51406 = n51405 ^ n14216 ^ n6312 ;
  assign n51407 = n51406 ^ n13611 ^ n1304 ;
  assign n51408 = ( n9491 & n10943 ) | ( n9491 & n51407 ) | ( n10943 & n51407 ) ;
  assign n51409 = ( n21755 & ~n23144 ) | ( n21755 & n51408 ) | ( ~n23144 & n51408 ) ;
  assign n51410 = n41742 ^ n18360 ^ 1'b0 ;
  assign n51411 = n42931 ^ n6813 ^ 1'b0 ;
  assign n51412 = n4633 & ~n51411 ;
  assign n51413 = ( n32672 & n51410 ) | ( n32672 & ~n51412 ) | ( n51410 & ~n51412 ) ;
  assign n51414 = n42709 & ~n51413 ;
  assign n51415 = n46929 ^ n44302 ^ n28513 ;
  assign n51416 = n49388 ^ n4619 ^ 1'b0 ;
  assign n51417 = n32575 & ~n51416 ;
  assign n51418 = ( n7892 & ~n11961 ) | ( n7892 & n16182 ) | ( ~n11961 & n16182 ) ;
  assign n51419 = n51418 ^ n29237 ^ 1'b0 ;
  assign n51420 = n12178 | n51419 ;
  assign n51421 = n28584 ^ n7827 ^ 1'b0 ;
  assign n51422 = n721 & n5846 ;
  assign n51423 = ~n6255 & n51422 ;
  assign n51424 = n51423 ^ n3895 ^ 1'b0 ;
  assign n51425 = n11349 | n51424 ;
  assign n51426 = n7350 & n24862 ;
  assign n51427 = n40314 ^ n20284 ^ 1'b0 ;
  assign n51428 = n51426 & n51427 ;
  assign n51429 = n8922 ^ n6450 ^ 1'b0 ;
  assign n51430 = ( ~n8983 & n36270 ) | ( ~n8983 & n48093 ) | ( n36270 & n48093 ) ;
  assign n51432 = n22337 & n34470 ;
  assign n51433 = ( n17343 & ~n19084 ) | ( n17343 & n51432 ) | ( ~n19084 & n51432 ) ;
  assign n51431 = n19569 | n23240 ;
  assign n51434 = n51433 ^ n51431 ^ 1'b0 ;
  assign n51435 = n51434 ^ n30355 ^ 1'b0 ;
  assign n51436 = n1421 | n51435 ;
  assign n51437 = n9433 & n15736 ;
  assign n51438 = ~n5132 & n51437 ;
  assign n51439 = ( n16784 & n39710 ) | ( n16784 & ~n51438 ) | ( n39710 & ~n51438 ) ;
  assign n51440 = ( n1848 & ~n15154 ) | ( n1848 & n51439 ) | ( ~n15154 & n51439 ) ;
  assign n51441 = n47846 ^ n10760 ^ n10236 ;
  assign n51442 = n51441 ^ n32240 ^ n6880 ;
  assign n51443 = n4322 & n8400 ;
  assign n51444 = n9444 & n51443 ;
  assign n51445 = n2700 | n13822 ;
  assign n51446 = n51445 ^ n2397 ^ 1'b0 ;
  assign n51447 = ( n51081 & ~n51444 ) | ( n51081 & n51446 ) | ( ~n51444 & n51446 ) ;
  assign n51448 = n51447 ^ n29023 ^ 1'b0 ;
  assign n51449 = n47728 ^ n14665 ^ n4988 ;
  assign n51450 = n51449 ^ n28957 ^ 1'b0 ;
  assign n51451 = n704 | n33778 ;
  assign n51452 = n25944 | n47967 ;
  assign n51453 = n51452 ^ n35466 ^ 1'b0 ;
  assign n51454 = ( n17815 & ~n35488 ) | ( n17815 & n51453 ) | ( ~n35488 & n51453 ) ;
  assign n51455 = n26208 ^ n20197 ^ 1'b0 ;
  assign n51456 = n51454 | n51455 ;
  assign n51457 = n36851 ^ n26786 ^ n21691 ;
  assign n51458 = n51457 ^ n3979 ^ n3031 ;
  assign n51459 = n42718 | n51458 ;
  assign n51460 = n16354 ^ n2923 ^ n632 ;
  assign n51461 = ( n18441 & n51322 ) | ( n18441 & ~n51460 ) | ( n51322 & ~n51460 ) ;
  assign n51462 = n51461 ^ n33557 ^ 1'b0 ;
  assign n51463 = x54 & n51462 ;
  assign n51464 = n51463 ^ n18447 ^ n4176 ;
  assign n51465 = n10252 | n18917 ;
  assign n51466 = ( n4696 & n20279 ) | ( n4696 & ~n51465 ) | ( n20279 & ~n51465 ) ;
  assign n51467 = ~n19969 & n32709 ;
  assign n51468 = n32273 ^ n9785 ^ n4141 ;
  assign n51469 = n18544 | n31083 ;
  assign n51470 = ( n11261 & n51468 ) | ( n11261 & ~n51469 ) | ( n51468 & ~n51469 ) ;
  assign n51471 = ~n51467 & n51470 ;
  assign n51472 = n44774 ^ n6240 ^ 1'b0 ;
  assign n51475 = n40472 ^ n18103 ^ n13870 ;
  assign n51473 = n3025 & ~n9286 ;
  assign n51474 = n51473 ^ n14223 ^ 1'b0 ;
  assign n51476 = n51475 ^ n51474 ^ n17098 ;
  assign n51477 = n51476 ^ n2246 ^ 1'b0 ;
  assign n51478 = n50452 ^ n36340 ^ n33098 ;
  assign n51479 = n51478 ^ n9294 ^ 1'b0 ;
  assign n51480 = n38968 | n51479 ;
  assign n51481 = n51480 ^ n29304 ^ 1'b0 ;
  assign n51482 = n37444 ^ n31035 ^ n23680 ;
  assign n51483 = n2370 & n51482 ;
  assign n51484 = n51483 ^ n3245 ^ 1'b0 ;
  assign n51485 = ( n6997 & n22250 ) | ( n6997 & ~n51484 ) | ( n22250 & ~n51484 ) ;
  assign n51486 = ( n18194 & n18734 ) | ( n18194 & ~n20234 ) | ( n18734 & ~n20234 ) ;
  assign n51487 = n41989 ^ n15318 ^ 1'b0 ;
  assign n51489 = n32333 ^ n5281 ^ 1'b0 ;
  assign n51490 = ( ~n3242 & n15966 ) | ( ~n3242 & n51489 ) | ( n15966 & n51489 ) ;
  assign n51488 = n33292 ^ n32861 ^ 1'b0 ;
  assign n51491 = n51490 ^ n51488 ^ 1'b0 ;
  assign n51492 = n4861 ^ n1563 ^ 1'b0 ;
  assign n51493 = n51492 ^ n22192 ^ 1'b0 ;
  assign n51494 = n34432 ^ n28742 ^ 1'b0 ;
  assign n51495 = n15641 & ~n29304 ;
  assign n51496 = ~n1643 & n18276 ;
  assign n51497 = n26247 ^ n7365 ^ 1'b0 ;
  assign n51498 = n51496 & n51497 ;
  assign n51499 = ( ~n3340 & n11583 ) | ( ~n3340 & n25325 ) | ( n11583 & n25325 ) ;
  assign n51500 = n16149 & n51499 ;
  assign n51501 = n51500 ^ n7201 ^ n4208 ;
  assign n51502 = n19334 & ~n20281 ;
  assign n51503 = n17855 | n21099 ;
  assign n51504 = n51503 ^ n15632 ^ 1'b0 ;
  assign n51505 = n5723 & n51504 ;
  assign n51506 = ( n43719 & n51502 ) | ( n43719 & ~n51505 ) | ( n51502 & ~n51505 ) ;
  assign n51507 = n2858 & ~n5348 ;
  assign n51508 = ( n19777 & n50268 ) | ( n19777 & n51507 ) | ( n50268 & n51507 ) ;
  assign n51510 = n18484 & ~n49033 ;
  assign n51509 = n30700 ^ n17635 ^ n14202 ;
  assign n51511 = n51510 ^ n51509 ^ n18980 ;
  assign n51512 = n51511 ^ n34081 ^ 1'b0 ;
  assign n51513 = n38648 ^ n36712 ^ n33475 ;
  assign n51514 = n30577 ^ n8526 ^ 1'b0 ;
  assign n51515 = n50836 ^ n20267 ^ n18050 ;
  assign n51516 = n51515 ^ n10243 ^ 1'b0 ;
  assign n51517 = n13114 ^ n5606 ^ 1'b0 ;
  assign n51519 = n5905 & n8649 ;
  assign n51520 = n51519 ^ n21890 ^ 1'b0 ;
  assign n51518 = n18712 & n27849 ;
  assign n51521 = n51520 ^ n51518 ^ n45537 ;
  assign n51522 = ( n32984 & ~n51517 ) | ( n32984 & n51521 ) | ( ~n51517 & n51521 ) ;
  assign n51523 = ( ~n10445 & n10986 ) | ( ~n10445 & n21990 ) | ( n10986 & n21990 ) ;
  assign n51524 = ( ~n1288 & n7561 ) | ( ~n1288 & n37824 ) | ( n7561 & n37824 ) ;
  assign n51525 = ( n795 & ~n10208 ) | ( n795 & n18505 ) | ( ~n10208 & n18505 ) ;
  assign n51526 = ( ~n12811 & n14555 ) | ( ~n12811 & n51525 ) | ( n14555 & n51525 ) ;
  assign n51527 = n1783 | n27393 ;
  assign n51528 = n37673 & ~n51527 ;
  assign n51529 = ( n5297 & ~n51526 ) | ( n5297 & n51528 ) | ( ~n51526 & n51528 ) ;
  assign n51531 = n4338 | n11003 ;
  assign n51532 = n14054 & ~n51531 ;
  assign n51530 = n2070 & n40189 ;
  assign n51533 = n51532 ^ n51530 ^ n29004 ;
  assign n51534 = ( n3618 & n6064 ) | ( n3618 & ~n10573 ) | ( n6064 & ~n10573 ) ;
  assign n51535 = n51534 ^ n11617 ^ n9505 ;
  assign n51536 = ( n1753 & n24455 ) | ( n1753 & n27610 ) | ( n24455 & n27610 ) ;
  assign n51537 = n13675 & ~n51536 ;
  assign n51538 = n18184 & n51537 ;
  assign n51539 = n1831 & ~n47852 ;
  assign n51540 = ~n6049 & n51539 ;
  assign n51545 = n14300 ^ n7880 ^ 1'b0 ;
  assign n51546 = n3375 & n51545 ;
  assign n51541 = n21216 & n31460 ;
  assign n51542 = n51541 ^ n14414 ^ 1'b0 ;
  assign n51543 = n20206 | n51542 ;
  assign n51544 = n4045 | n51543 ;
  assign n51547 = n51546 ^ n51544 ^ 1'b0 ;
  assign n51548 = n6913 | n23776 ;
  assign n51549 = n51548 ^ n33543 ^ 1'b0 ;
  assign n51550 = n42434 ^ n29263 ^ n19250 ;
  assign n51551 = n44096 ^ n43501 ^ 1'b0 ;
  assign n51552 = n36406 ^ n35200 ^ 1'b0 ;
  assign n51553 = n29169 ^ n4359 ^ 1'b0 ;
  assign n51554 = n41130 ^ n12753 ^ n8565 ;
  assign n51555 = n49257 & n51554 ;
  assign n51556 = n43602 ^ n31663 ^ n3355 ;
  assign n51557 = ( n9848 & n23346 ) | ( n9848 & n51556 ) | ( n23346 & n51556 ) ;
  assign n51558 = n1230 & ~n19104 ;
  assign n51559 = n12087 | n51558 ;
  assign n51560 = n25754 & ~n51559 ;
  assign n51561 = n21404 | n49364 ;
  assign n51562 = n50518 | n51561 ;
  assign n51563 = n15990 | n23474 ;
  assign n51564 = n51563 ^ n3466 ^ 1'b0 ;
  assign n51565 = ~n6775 & n7697 ;
  assign n51566 = n51565 ^ n9406 ^ 1'b0 ;
  assign n51567 = n27248 ^ n12664 ^ 1'b0 ;
  assign n51568 = n19036 ^ x227 ^ 1'b0 ;
  assign n51569 = n25652 ^ n9656 ^ 1'b0 ;
  assign n51570 = ~n51568 & n51569 ;
  assign n51571 = ( n8484 & ~n39519 ) | ( n8484 & n51570 ) | ( ~n39519 & n51570 ) ;
  assign n51574 = n16935 ^ n12710 ^ 1'b0 ;
  assign n51572 = n1305 & ~n5059 ;
  assign n51573 = ( n7056 & n19009 ) | ( n7056 & n51572 ) | ( n19009 & n51572 ) ;
  assign n51575 = n51574 ^ n51573 ^ n25061 ;
  assign n51576 = n36042 ^ n8481 ^ n2375 ;
  assign n51577 = n51576 ^ n18476 ^ n17543 ;
  assign n51578 = n47151 ^ n42015 ^ 1'b0 ;
  assign n51579 = ( n11381 & n16424 ) | ( n11381 & n23450 ) | ( n16424 & n23450 ) ;
  assign n51580 = n47051 ^ n6601 ^ n3348 ;
  assign n51581 = ( n48139 & n51579 ) | ( n48139 & n51580 ) | ( n51579 & n51580 ) ;
  assign n51582 = n29107 ^ n8218 ^ 1'b0 ;
  assign n51583 = n23524 | n47345 ;
  assign n51584 = n22150 & n39598 ;
  assign n51585 = n40705 ^ n18527 ^ n5342 ;
  assign n51586 = n27401 ^ n17127 ^ 1'b0 ;
  assign n51587 = ( n5617 & n35709 ) | ( n5617 & n41782 ) | ( n35709 & n41782 ) ;
  assign n51588 = ( n2359 & ~n24157 ) | ( n2359 & n51587 ) | ( ~n24157 & n51587 ) ;
  assign n51589 = ( n22566 & ~n39665 ) | ( n22566 & n51588 ) | ( ~n39665 & n51588 ) ;
  assign n51590 = ~n10625 & n51589 ;
  assign n51591 = n48586 ^ n22758 ^ 1'b0 ;
  assign n51592 = ( n5773 & n7558 ) | ( n5773 & n20763 ) | ( n7558 & n20763 ) ;
  assign n51593 = n39007 ^ n13711 ^ 1'b0 ;
  assign n51594 = ( ~n23192 & n51592 ) | ( ~n23192 & n51593 ) | ( n51592 & n51593 ) ;
  assign n51595 = n24906 ^ n12413 ^ n3230 ;
  assign n51596 = n3249 & n51595 ;
  assign n51597 = n51596 ^ n15132 ^ 1'b0 ;
  assign n51598 = n8491 & n48571 ;
  assign n51599 = n51598 ^ n7836 ^ 1'b0 ;
  assign n51603 = n3067 & n21864 ;
  assign n51604 = n11416 & n51603 ;
  assign n51605 = n1721 ^ n1506 ^ 1'b0 ;
  assign n51606 = ~n51604 & n51605 ;
  assign n51607 = ( ~n10488 & n14789 ) | ( ~n10488 & n51606 ) | ( n14789 & n51606 ) ;
  assign n51602 = n18531 ^ n11681 ^ n4375 ;
  assign n51608 = n51607 ^ n51602 ^ 1'b0 ;
  assign n51600 = ~n17356 & n45866 ;
  assign n51601 = n22178 | n51600 ;
  assign n51609 = n51608 ^ n51601 ^ 1'b0 ;
  assign n51611 = n3981 & ~n37067 ;
  assign n51610 = ( n10782 & n22494 ) | ( n10782 & ~n45640 ) | ( n22494 & ~n45640 ) ;
  assign n51612 = n51611 ^ n51610 ^ n31286 ;
  assign n51613 = n20125 & ~n51612 ;
  assign n51614 = n51613 ^ n24427 ^ 1'b0 ;
  assign n51615 = n21199 | n23129 ;
  assign n51616 = n16770 & n51615 ;
  assign n51617 = n17504 & ~n51616 ;
  assign n51618 = n6724 & ~n51617 ;
  assign n51619 = ( n7884 & n18911 ) | ( n7884 & n44054 ) | ( n18911 & n44054 ) ;
  assign n51620 = n51619 ^ n25641 ^ n7492 ;
  assign n51621 = n30764 ^ n11708 ^ n11417 ;
  assign n51622 = ~n17180 & n29964 ;
  assign n51623 = n12382 & n12472 ;
  assign n51624 = n51623 ^ n15802 ^ 1'b0 ;
  assign n51625 = n51624 ^ n43624 ^ n14975 ;
  assign n51626 = ( n24522 & n51622 ) | ( n24522 & ~n51625 ) | ( n51622 & ~n51625 ) ;
  assign n51634 = n20772 ^ n16403 ^ 1'b0 ;
  assign n51627 = n43720 ^ n32128 ^ 1'b0 ;
  assign n51628 = ~n23013 & n42850 ;
  assign n51629 = n51628 ^ n21566 ^ 1'b0 ;
  assign n51630 = n41875 ^ n16438 ^ 1'b0 ;
  assign n51631 = n51629 & n51630 ;
  assign n51632 = ( n7429 & ~n51627 ) | ( n7429 & n51631 ) | ( ~n51627 & n51631 ) ;
  assign n51633 = n51632 ^ n36121 ^ n32447 ;
  assign n51635 = n51634 ^ n51633 ^ n29987 ;
  assign n51636 = n5115 ^ n3446 ^ 1'b0 ;
  assign n51637 = n9246 & ~n40306 ;
  assign n51638 = ~n10317 & n51637 ;
  assign n51639 = n39016 ^ n11572 ^ 1'b0 ;
  assign n51640 = ~n16347 & n51639 ;
  assign n51641 = n20163 & n29970 ;
  assign n51642 = ~n17433 & n31083 ;
  assign n51643 = ( ~n40158 & n46875 ) | ( ~n40158 & n51520 ) | ( n46875 & n51520 ) ;
  assign n51644 = ( n3250 & ~n8030 ) | ( n3250 & n47333 ) | ( ~n8030 & n47333 ) ;
  assign n51645 = n45335 ^ n23301 ^ n21063 ;
  assign n51646 = n6728 | n32149 ;
  assign n51647 = n4063 & n45905 ;
  assign n51648 = n25274 ^ n23630 ^ 1'b0 ;
  assign n51649 = n3563 | n24684 ;
  assign n51650 = n35534 & ~n51649 ;
  assign n51651 = n36423 ^ n7851 ^ n5427 ;
  assign n51652 = ~n11893 & n35988 ;
  assign n51653 = n51652 ^ n34448 ^ 1'b0 ;
  assign n51654 = n23125 ^ n19035 ^ 1'b0 ;
  assign n51655 = n51654 ^ n17400 ^ n13531 ;
  assign n51656 = ( n7326 & ~n11730 ) | ( n7326 & n39782 ) | ( ~n11730 & n39782 ) ;
  assign n51657 = ~n42151 & n44340 ;
  assign n51658 = n51657 ^ n12036 ^ n10749 ;
  assign n51659 = ~n3400 & n15167 ;
  assign n51660 = n26697 | n35314 ;
  assign n51661 = n8428 | n51660 ;
  assign n51662 = n48937 & ~n51661 ;
  assign n51663 = n24232 ^ n12972 ^ n6120 ;
  assign n51664 = n39280 & ~n51663 ;
  assign n51665 = n51664 ^ n842 ^ 1'b0 ;
  assign n51666 = n30670 ^ n22676 ^ n3353 ;
  assign n51667 = ~n4568 & n35228 ;
  assign n51668 = n5902 ^ n3899 ^ n3504 ;
  assign n51669 = n51668 ^ n10337 ^ n10308 ;
  assign n51670 = n51669 ^ n46145 ^ n29432 ;
  assign n51671 = ( n9346 & n13849 ) | ( n9346 & n27559 ) | ( n13849 & n27559 ) ;
  assign n51672 = n51671 ^ n31118 ^ n4770 ;
  assign n51673 = n27574 ^ n16917 ^ n10083 ;
  assign n51674 = n51673 ^ n30529 ^ n19163 ;
  assign n51675 = ( ~n3201 & n30240 ) | ( ~n3201 & n51674 ) | ( n30240 & n51674 ) ;
  assign n51676 = n6685 ^ n5578 ^ n2254 ;
  assign n51677 = n51676 ^ n13801 ^ 1'b0 ;
  assign n51678 = n26585 & ~n51677 ;
  assign n51679 = n19840 | n51678 ;
  assign n51680 = ( n1266 & n10611 ) | ( n1266 & ~n20506 ) | ( n10611 & ~n20506 ) ;
  assign n51681 = ~n33214 & n51680 ;
  assign n51682 = n4095 & ~n21617 ;
  assign n51683 = n51682 ^ n49735 ^ 1'b0 ;
  assign n51684 = n25281 ^ n12249 ^ x186 ;
  assign n51685 = n6314 ^ n3532 ^ n882 ;
  assign n51686 = n51685 ^ n38788 ^ n36086 ;
  assign n51687 = ( n38580 & ~n51684 ) | ( n38580 & n51686 ) | ( ~n51684 & n51686 ) ;
  assign n51688 = n24764 & ~n28902 ;
  assign n51689 = n51688 ^ n5522 ^ 1'b0 ;
  assign n51690 = ( n648 & n1927 ) | ( n648 & ~n51689 ) | ( n1927 & ~n51689 ) ;
  assign n51691 = n28552 ^ n12042 ^ 1'b0 ;
  assign n51692 = n3287 & ~n24382 ;
  assign n51693 = ( n24266 & ~n35269 ) | ( n24266 & n51692 ) | ( ~n35269 & n51692 ) ;
  assign n51694 = n37267 ^ n8519 ^ n2555 ;
  assign n51695 = ( ~n2840 & n32290 ) | ( ~n2840 & n51694 ) | ( n32290 & n51694 ) ;
  assign n51696 = n40090 ^ n14942 ^ 1'b0 ;
  assign n51697 = n27392 ^ n11564 ^ 1'b0 ;
  assign n51698 = n36854 ^ n25522 ^ n14266 ;
  assign n51699 = n21132 ^ n9192 ^ n9073 ;
  assign n51700 = n51699 ^ n18270 ^ 1'b0 ;
  assign n51701 = n51698 & n51700 ;
  assign n51703 = n21910 ^ n16292 ^ 1'b0 ;
  assign n51704 = n6826 & n51703 ;
  assign n51705 = ( ~x219 & n8111 ) | ( ~x219 & n45429 ) | ( n8111 & n45429 ) ;
  assign n51706 = n20673 ^ n4721 ^ 1'b0 ;
  assign n51707 = n1753 | n51706 ;
  assign n51708 = n51707 ^ n34343 ^ 1'b0 ;
  assign n51709 = ( n6215 & ~n51705 ) | ( n6215 & n51708 ) | ( ~n51705 & n51708 ) ;
  assign n51710 = ( n31236 & ~n51704 ) | ( n31236 & n51709 ) | ( ~n51704 & n51709 ) ;
  assign n51702 = n528 & n18155 ;
  assign n51711 = n51710 ^ n51702 ^ 1'b0 ;
  assign n51712 = n48308 ^ n7846 ^ 1'b0 ;
  assign n51713 = n6903 | n39519 ;
  assign n51714 = n31895 ^ n24875 ^ n1722 ;
  assign n51715 = ( n25961 & ~n37363 ) | ( n25961 & n40364 ) | ( ~n37363 & n40364 ) ;
  assign n51716 = n41268 ^ n39051 ^ n28258 ;
  assign n51717 = n18057 ^ n12773 ^ 1'b0 ;
  assign n51718 = ~n9227 & n51717 ;
  assign n51719 = ~n1544 & n21148 ;
  assign n51720 = ~n51718 & n51719 ;
  assign n51721 = n5464 & ~n33401 ;
  assign n51722 = n26958 ^ n19840 ^ n3111 ;
  assign n51723 = n31876 & n51722 ;
  assign n51724 = n40897 ^ n13860 ^ n8743 ;
  assign n51725 = n51511 ^ n51198 ^ 1'b0 ;
  assign n51726 = n38914 ^ n25416 ^ n17880 ;
  assign n51727 = ( x182 & n21647 ) | ( x182 & ~n34011 ) | ( n21647 & ~n34011 ) ;
  assign n51728 = n7024 & n17626 ;
  assign n51729 = n3885 & n51728 ;
  assign n51730 = n36931 | n51729 ;
  assign n51731 = n1502 & ~n51730 ;
  assign n51732 = n51731 ^ n43108 ^ n22843 ;
  assign n51733 = ( n4131 & ~n12171 ) | ( n4131 & n20100 ) | ( ~n12171 & n20100 ) ;
  assign n51734 = ~n514 & n17578 ;
  assign n51735 = n51733 & n51734 ;
  assign n51736 = n16488 & ~n51735 ;
  assign n51737 = ( n5505 & n7487 ) | ( n5505 & n45508 ) | ( n7487 & n45508 ) ;
  assign n51738 = n40613 | n51737 ;
  assign n51739 = n37505 | n51738 ;
  assign n51740 = n1974 & n20537 ;
  assign n51741 = ( n4601 & ~n4924 ) | ( n4601 & n21115 ) | ( ~n4924 & n21115 ) ;
  assign n51742 = n8127 | n16233 ;
  assign n51743 = n31888 ^ n5500 ^ 1'b0 ;
  assign n51744 = ~n51742 & n51743 ;
  assign n51745 = n8422 ^ n8245 ^ 1'b0 ;
  assign n51746 = ( n12534 & n23827 ) | ( n12534 & ~n51745 ) | ( n23827 & ~n51745 ) ;
  assign n51747 = n27015 | n35592 ;
  assign n51748 = ( ~n9952 & n51746 ) | ( ~n9952 & n51747 ) | ( n51746 & n51747 ) ;
  assign n51749 = n15431 ^ n5976 ^ 1'b0 ;
  assign n51750 = ~n10114 & n11508 ;
  assign n51751 = n44364 ^ n34177 ^ n14394 ;
  assign n51752 = n3549 & ~n51751 ;
  assign n51753 = ~n51750 & n51752 ;
  assign n51754 = ( n23796 & n51749 ) | ( n23796 & n51753 ) | ( n51749 & n51753 ) ;
  assign n51755 = ( ~n32144 & n45716 ) | ( ~n32144 & n50942 ) | ( n45716 & n50942 ) ;
  assign n51756 = n34116 ^ n6160 ^ n1072 ;
  assign n51757 = n51756 ^ n50485 ^ n44743 ;
  assign n51758 = n28307 | n37191 ;
  assign n51759 = n2583 | n51758 ;
  assign n51760 = n51759 ^ n22883 ^ 1'b0 ;
  assign n51761 = n39815 ^ n29027 ^ n5412 ;
  assign n51762 = ( n13891 & n14734 ) | ( n13891 & n50306 ) | ( n14734 & n50306 ) ;
  assign n51763 = ( n11238 & ~n14545 ) | ( n11238 & n51762 ) | ( ~n14545 & n51762 ) ;
  assign n51764 = n51761 | n51763 ;
  assign n51765 = n40501 ^ n36153 ^ 1'b0 ;
  assign n51766 = ( n2354 & ~n10840 ) | ( n2354 & n47127 ) | ( ~n10840 & n47127 ) ;
  assign n51767 = n21914 ^ n14279 ^ x113 ;
  assign n51768 = n24522 ^ n22843 ^ n18716 ;
  assign n51770 = n8827 ^ n3382 ^ 1'b0 ;
  assign n51771 = n829 & n51770 ;
  assign n51769 = ( n16603 & ~n34573 ) | ( n16603 & n36404 ) | ( ~n34573 & n36404 ) ;
  assign n51772 = n51771 ^ n51769 ^ 1'b0 ;
  assign n51773 = ( n13739 & ~n39648 ) | ( n13739 & n51772 ) | ( ~n39648 & n51772 ) ;
  assign n51774 = n33152 ^ n2123 ^ 1'b0 ;
  assign n51775 = ( n25050 & n30562 ) | ( n25050 & ~n46507 ) | ( n30562 & ~n46507 ) ;
  assign n51776 = n33765 & n51775 ;
  assign n51777 = n14809 & n41759 ;
  assign n51778 = n15621 & n51777 ;
  assign n51779 = n16243 & n22064 ;
  assign n51780 = n51778 | n51779 ;
  assign n51781 = ~n6130 & n10742 ;
  assign n51782 = n49145 & n51781 ;
  assign n51783 = n36881 ^ n11255 ^ 1'b0 ;
  assign n51784 = n19354 & n41746 ;
  assign n51785 = n51784 ^ n1859 ^ 1'b0 ;
  assign n51786 = n33569 ^ n28912 ^ n13804 ;
  assign n51787 = ~n39078 & n51786 ;
  assign n51788 = n51787 ^ n36361 ^ 1'b0 ;
  assign n51789 = ( ~n11395 & n51785 ) | ( ~n11395 & n51788 ) | ( n51785 & n51788 ) ;
  assign n51790 = ( n10214 & ~n22404 ) | ( n10214 & n51789 ) | ( ~n22404 & n51789 ) ;
  assign n51791 = n49705 ^ n24714 ^ 1'b0 ;
  assign n51794 = n14438 & n20895 ;
  assign n51793 = n40591 ^ n34422 ^ 1'b0 ;
  assign n51792 = ( n19378 & n30964 ) | ( n19378 & n38351 ) | ( n30964 & n38351 ) ;
  assign n51795 = n51794 ^ n51793 ^ n51792 ;
  assign n51796 = ( n8847 & ~n21448 ) | ( n8847 & n49810 ) | ( ~n21448 & n49810 ) ;
  assign n51797 = ~n9083 & n14291 ;
  assign n51798 = n51797 ^ n29632 ^ 1'b0 ;
  assign n51799 = ( n4495 & n5788 ) | ( n4495 & ~n22473 ) | ( n5788 & ~n22473 ) ;
  assign n51800 = n30677 | n51799 ;
  assign n51801 = n51800 ^ n19453 ^ 1'b0 ;
  assign n51802 = n45399 ^ n1303 ^ n981 ;
  assign n51803 = n1906 & ~n51802 ;
  assign n51804 = ~n40443 & n51803 ;
  assign n51805 = n28212 ^ n21742 ^ 1'b0 ;
  assign n51806 = n3982 | n51805 ;
  assign n51807 = n12460 | n14860 ;
  assign n51808 = n40618 ^ n35053 ^ n21801 ;
  assign n51809 = ( n14497 & ~n19291 ) | ( n14497 & n36007 ) | ( ~n19291 & n36007 ) ;
  assign n51810 = n10572 & ~n51809 ;
  assign n51811 = n11430 & n51810 ;
  assign n51812 = ( ~n6926 & n10808 ) | ( ~n6926 & n51811 ) | ( n10808 & n51811 ) ;
  assign n51813 = n42765 ^ n35697 ^ n14574 ;
  assign n51814 = ( ~n17898 & n29432 ) | ( ~n17898 & n51813 ) | ( n29432 & n51813 ) ;
  assign n51819 = n20970 & ~n37513 ;
  assign n51820 = n51819 ^ n2900 ^ 1'b0 ;
  assign n51818 = n27544 ^ n19350 ^ n16028 ;
  assign n51816 = n8219 & ~n34107 ;
  assign n51815 = ( n2835 & ~n14379 ) | ( n2835 & n20767 ) | ( ~n14379 & n20767 ) ;
  assign n51817 = n51816 ^ n51815 ^ n14875 ;
  assign n51821 = n51820 ^ n51818 ^ n51817 ;
  assign n51822 = ( n4051 & n32144 ) | ( n4051 & n34244 ) | ( n32144 & n34244 ) ;
  assign n51823 = n46188 ^ n1451 ^ 1'b0 ;
  assign n51824 = ( n7085 & n7139 ) | ( n7085 & n51823 ) | ( n7139 & n51823 ) ;
  assign n51825 = n38641 & n51824 ;
  assign n51826 = n51825 ^ n47938 ^ 1'b0 ;
  assign n51828 = ( x2 & n5186 ) | ( x2 & ~n27600 ) | ( n5186 & ~n27600 ) ;
  assign n51827 = ~n5502 & n41031 ;
  assign n51829 = n51828 ^ n51827 ^ 1'b0 ;
  assign n51830 = ( n643 & n1547 ) | ( n643 & ~n9685 ) | ( n1547 & ~n9685 ) ;
  assign n51831 = n51830 ^ n286 ^ 1'b0 ;
  assign n51832 = n51831 ^ n51257 ^ 1'b0 ;
  assign n51833 = n34975 & n51832 ;
  assign n51834 = n34107 ^ n5557 ^ 1'b0 ;
  assign n51835 = n7438 & ~n51834 ;
  assign n51836 = n19703 ^ n9597 ^ n3991 ;
  assign n51837 = n51836 ^ n857 ^ 1'b0 ;
  assign n51838 = n3309 | n51837 ;
  assign n51839 = ( n6351 & ~n51276 ) | ( n6351 & n51838 ) | ( ~n51276 & n51838 ) ;
  assign n51842 = n10540 ^ n5244 ^ 1'b0 ;
  assign n51843 = n46426 & n51842 ;
  assign n51840 = ~n1647 & n49870 ;
  assign n51841 = ~n50761 & n51840 ;
  assign n51844 = n51843 ^ n51841 ^ n15935 ;
  assign n51845 = n666 & ~n19187 ;
  assign n51846 = n51845 ^ n14860 ^ 1'b0 ;
  assign n51847 = ( n11968 & n16829 ) | ( n11968 & ~n51846 ) | ( n16829 & ~n51846 ) ;
  assign n51848 = n50165 ^ n49460 ^ x184 ;
  assign n51849 = n47330 ^ n27453 ^ n3678 ;
  assign n51850 = ( n19894 & n20588 ) | ( n19894 & ~n50097 ) | ( n20588 & ~n50097 ) ;
  assign n51851 = n1725 ^ x63 ^ 1'b0 ;
  assign n51852 = n43391 & n51851 ;
  assign n51853 = ~n4733 & n51852 ;
  assign n51854 = ~n9022 & n51853 ;
  assign n51855 = n16708 ^ n1837 ^ 1'b0 ;
  assign n51856 = ~n32425 & n51855 ;
  assign n51857 = n24683 & ~n47676 ;
  assign n51858 = n51857 ^ n38884 ^ 1'b0 ;
  assign n51859 = n51856 & ~n51858 ;
  assign n51860 = n41623 ^ n6747 ^ 1'b0 ;
  assign n51861 = n4066 & n51860 ;
  assign n51862 = ( n4714 & n11970 ) | ( n4714 & ~n18615 ) | ( n11970 & ~n18615 ) ;
  assign n51863 = ( n20017 & n21840 ) | ( n20017 & n33404 ) | ( n21840 & n33404 ) ;
  assign n51864 = ( ~n3634 & n18294 ) | ( ~n3634 & n22889 ) | ( n18294 & n22889 ) ;
  assign n51865 = n51864 ^ n41775 ^ n12697 ;
  assign n51866 = ~n690 & n51865 ;
  assign n51867 = ~n17313 & n37602 ;
  assign n51868 = n21987 ^ n11322 ^ n939 ;
  assign n51869 = ( n5031 & ~n38631 ) | ( n5031 & n51868 ) | ( ~n38631 & n51868 ) ;
  assign n51870 = n10890 & n16955 ;
  assign n51871 = n29746 & n51870 ;
  assign n51872 = n26507 ^ n23656 ^ n3511 ;
  assign n51873 = n16431 ^ n15319 ^ 1'b0 ;
  assign n51874 = n51872 | n51873 ;
  assign n51875 = n16546 ^ n5322 ^ x128 ;
  assign n51876 = n51875 ^ n24068 ^ 1'b0 ;
  assign n51877 = n7358 | n51876 ;
  assign n51878 = n11585 & n33395 ;
  assign n51879 = n51878 ^ n23001 ^ 1'b0 ;
  assign n51880 = n32907 ^ n22525 ^ 1'b0 ;
  assign n51881 = n38744 ^ n20232 ^ n13346 ;
  assign n51882 = n45561 ^ n25715 ^ 1'b0 ;
  assign n51883 = ( ~n43457 & n51881 ) | ( ~n43457 & n51882 ) | ( n51881 & n51882 ) ;
  assign n51884 = n45305 ^ n28584 ^ n20657 ;
  assign n51885 = n34466 ^ n3449 ^ 1'b0 ;
  assign n51886 = ~n28346 & n38418 ;
  assign n51887 = n51886 ^ n43040 ^ n40732 ;
  assign n51888 = n12388 | n13320 ;
  assign n51889 = n51888 ^ n4784 ^ 1'b0 ;
  assign n51890 = ~n8049 & n15548 ;
  assign n51891 = ~n10080 & n51890 ;
  assign n51892 = ~n7665 & n42532 ;
  assign n51894 = n12407 & n40395 ;
  assign n51895 = n51894 ^ n17663 ^ 1'b0 ;
  assign n51893 = ~n7830 & n35710 ;
  assign n51896 = n51895 ^ n51893 ^ 1'b0 ;
  assign n51897 = n23732 ^ n1203 ^ 1'b0 ;
  assign n51898 = n21609 & ~n51897 ;
  assign n51899 = ( n6345 & ~n8553 ) | ( n6345 & n51898 ) | ( ~n8553 & n51898 ) ;
  assign n51900 = ( n24364 & n40632 ) | ( n24364 & n51899 ) | ( n40632 & n51899 ) ;
  assign n51901 = ( n2835 & n18456 ) | ( n2835 & ~n38132 ) | ( n18456 & ~n38132 ) ;
  assign n51902 = n16290 ^ n14832 ^ n10690 ;
  assign n51903 = n33294 ^ n31033 ^ n18226 ;
  assign n51904 = ( n38533 & ~n51902 ) | ( n38533 & n51903 ) | ( ~n51902 & n51903 ) ;
  assign n51905 = n39948 & n50006 ;
  assign n51906 = ~n6355 & n51905 ;
  assign n51907 = ( ~n43358 & n49378 ) | ( ~n43358 & n51906 ) | ( n49378 & n51906 ) ;
  assign n51908 = ~n4961 & n22041 ;
  assign n51909 = ( n13298 & n30295 ) | ( n13298 & n45550 ) | ( n30295 & n45550 ) ;
  assign n51910 = n3221 ^ n386 ^ 1'b0 ;
  assign n51911 = ~n12362 & n51910 ;
  assign n51912 = ~n17130 & n51911 ;
  assign n51913 = n39523 & n51912 ;
  assign n51915 = n30318 ^ n24360 ^ n13618 ;
  assign n51914 = ~n5440 & n51439 ;
  assign n51916 = n51915 ^ n51914 ^ 1'b0 ;
  assign n51917 = n17594 ^ n739 ^ 1'b0 ;
  assign n51918 = n51917 ^ n38500 ^ n15357 ;
  assign n51919 = n9328 ^ n2234 ^ 1'b0 ;
  assign n51920 = ( n21200 & n50137 ) | ( n21200 & n51919 ) | ( n50137 & n51919 ) ;
  assign n51921 = n9438 ^ n7677 ^ 1'b0 ;
  assign n51922 = ( n32469 & n37092 ) | ( n32469 & ~n51921 ) | ( n37092 & ~n51921 ) ;
  assign n51923 = ~n7355 & n41473 ;
  assign n51924 = n48873 ^ n36772 ^ n14109 ;
  assign n51925 = n12504 & n27976 ;
  assign n51926 = n51925 ^ n50077 ^ n12036 ;
  assign n51927 = ( n7541 & n19281 ) | ( n7541 & n19507 ) | ( n19281 & n19507 ) ;
  assign n51928 = n51927 ^ n35866 ^ 1'b0 ;
  assign n51929 = n1081 & ~n51928 ;
  assign n51930 = n40281 ^ n24362 ^ 1'b0 ;
  assign n51931 = n21537 & ~n51930 ;
  assign n51932 = n37868 ^ n1779 ^ 1'b0 ;
  assign n51933 = ~n21362 & n51932 ;
  assign n51934 = ( n4245 & n18648 ) | ( n4245 & n45551 ) | ( n18648 & n45551 ) ;
  assign n51935 = ( n11204 & n39575 ) | ( n11204 & ~n51934 ) | ( n39575 & ~n51934 ) ;
  assign n51936 = ( n2605 & ~n4933 ) | ( n2605 & n15012 ) | ( ~n4933 & n15012 ) ;
  assign n51937 = ( ~n13544 & n39320 ) | ( ~n13544 & n51936 ) | ( n39320 & n51936 ) ;
  assign n51938 = n24549 ^ n5400 ^ n3370 ;
  assign n51939 = n34273 & n51938 ;
  assign n51940 = n51939 ^ n49331 ^ n35611 ;
  assign n51941 = n33044 ^ n18441 ^ n12338 ;
  assign n51942 = n2816 ^ n518 ^ 1'b0 ;
  assign n51943 = n51942 ^ n37930 ^ n9035 ;
  assign n51944 = n24104 ^ n23630 ^ n10760 ;
  assign n51945 = ( ~x249 & n24518 ) | ( ~x249 & n51944 ) | ( n24518 & n51944 ) ;
  assign n51946 = n8199 ^ n7610 ^ n585 ;
  assign n51947 = n51946 ^ n7379 ^ 1'b0 ;
  assign n51948 = ( n35789 & n51945 ) | ( n35789 & ~n51947 ) | ( n51945 & ~n51947 ) ;
  assign n51949 = ( n2208 & n10616 ) | ( n2208 & n51948 ) | ( n10616 & n51948 ) ;
  assign n51950 = n33430 & n38751 ;
  assign n51951 = ~n35988 & n51950 ;
  assign n51952 = n36191 ^ n27578 ^ n18379 ;
  assign n51953 = n37668 ^ n18917 ^ 1'b0 ;
  assign n51954 = ~n22019 & n51953 ;
  assign n51955 = ( ~n30053 & n51952 ) | ( ~n30053 & n51954 ) | ( n51952 & n51954 ) ;
  assign n51956 = ( n35833 & n37443 ) | ( n35833 & n51955 ) | ( n37443 & n51955 ) ;
  assign n51957 = n6763 & ~n51956 ;
  assign n51958 = n19859 | n27086 ;
  assign n51959 = ( n10195 & n30053 ) | ( n10195 & ~n30807 ) | ( n30053 & ~n30807 ) ;
  assign n51960 = ( n34808 & n42186 ) | ( n34808 & n51959 ) | ( n42186 & n51959 ) ;
  assign n51961 = ( n5905 & n8344 ) | ( n5905 & ~n15679 ) | ( n8344 & ~n15679 ) ;
  assign n51962 = n1670 & n4319 ;
  assign n51963 = n6245 & n26283 ;
  assign n51964 = n6749 | n28309 ;
  assign n51965 = n9865 & ~n51964 ;
  assign n51966 = n20464 & ~n28933 ;
  assign n51967 = n3834 & n49818 ;
  assign n51968 = n18965 & n51967 ;
  assign n51969 = n38160 & n51968 ;
  assign n51970 = n25763 ^ n20027 ^ n14189 ;
  assign n51971 = ( n4047 & ~n12181 ) | ( n4047 & n12916 ) | ( ~n12181 & n12916 ) ;
  assign n51972 = ( ~n11343 & n31999 ) | ( ~n11343 & n51971 ) | ( n31999 & n51971 ) ;
  assign n51973 = ~n744 & n7372 ;
  assign n51974 = n51973 ^ n4967 ^ 1'b0 ;
  assign n51975 = n8546 & n51974 ;
  assign n51976 = ( n5984 & ~n9526 ) | ( n5984 & n16586 ) | ( ~n9526 & n16586 ) ;
  assign n51977 = ( ~n17294 & n41276 ) | ( ~n17294 & n51976 ) | ( n41276 & n51976 ) ;
  assign n51978 = n37967 ^ n20957 ^ n16216 ;
  assign n51979 = n6662 ^ n2629 ^ 1'b0 ;
  assign n51980 = n13667 | n51979 ;
  assign n51981 = n51980 ^ n40965 ^ n6072 ;
  assign n51982 = n51944 ^ n34007 ^ n6376 ;
  assign n51983 = n51982 ^ n39205 ^ 1'b0 ;
  assign n51984 = n51983 ^ n35442 ^ 1'b0 ;
  assign n51985 = n5839 ^ n1753 ^ 1'b0 ;
  assign n51986 = n10763 | n49652 ;
  assign n51987 = n35882 & ~n51986 ;
  assign n51988 = n40433 ^ n27504 ^ n2790 ;
  assign n51989 = ( n6849 & n12750 ) | ( n6849 & ~n14261 ) | ( n12750 & ~n14261 ) ;
  assign n51990 = n15288 ^ n5692 ^ n3735 ;
  assign n51991 = n51990 ^ n18717 ^ 1'b0 ;
  assign n51992 = n15137 & ~n26037 ;
  assign n51993 = n51991 & n51992 ;
  assign n51994 = n47912 ^ n42741 ^ n5832 ;
  assign n51995 = n51993 & n51994 ;
  assign n51996 = n47770 ^ n35053 ^ n3854 ;
  assign n51997 = n51996 ^ n33977 ^ n5914 ;
  assign n51998 = n40909 ^ n15855 ^ 1'b0 ;
  assign n51999 = n31347 ^ n15792 ^ n6334 ;
  assign n52000 = x240 & ~n10856 ;
  assign n52001 = n3310 & n52000 ;
  assign n52002 = n7004 ^ n3592 ^ 1'b0 ;
  assign n52003 = n27486 & n52002 ;
  assign n52004 = n22624 & ~n52003 ;
  assign n52005 = n51877 ^ n28005 ^ 1'b0 ;
  assign n52006 = n4946 | n25843 ;
  assign n52007 = n52006 ^ n4983 ^ 1'b0 ;
  assign n52008 = n30750 ^ n4713 ^ n735 ;
  assign n52009 = n12641 ^ n785 ^ 1'b0 ;
  assign n52010 = n14412 & n52009 ;
  assign n52011 = n52010 ^ n9716 ^ n831 ;
  assign n52012 = ( ~n1943 & n32147 ) | ( ~n1943 & n34791 ) | ( n32147 & n34791 ) ;
  assign n52013 = n16019 ^ n12916 ^ n6200 ;
  assign n52014 = n16225 ^ n15488 ^ n758 ;
  assign n52015 = ( n31349 & n52013 ) | ( n31349 & n52014 ) | ( n52013 & n52014 ) ;
  assign n52016 = ( n885 & n15472 ) | ( n885 & ~n42971 ) | ( n15472 & ~n42971 ) ;
  assign n52017 = ( ~n4300 & n10456 ) | ( ~n4300 & n16400 ) | ( n10456 & n16400 ) ;
  assign n52018 = n1845 | n12449 ;
  assign n52019 = n52018 ^ n3204 ^ 1'b0 ;
  assign n52020 = n4164 ^ n1373 ^ 1'b0 ;
  assign n52021 = n33490 | n52020 ;
  assign n52022 = ( ~n21904 & n23038 ) | ( ~n21904 & n37223 ) | ( n23038 & n37223 ) ;
  assign n52023 = ( n282 & n9656 ) | ( n282 & n37485 ) | ( n9656 & n37485 ) ;
  assign n52024 = n52023 ^ n40202 ^ n18353 ;
  assign n52025 = ( ~n704 & n52022 ) | ( ~n704 & n52024 ) | ( n52022 & n52024 ) ;
  assign n52026 = n22682 ^ n12219 ^ n9490 ;
  assign n52027 = n11429 ^ n7990 ^ 1'b0 ;
  assign n52028 = ( n8175 & ~n8550 ) | ( n8175 & n52027 ) | ( ~n8550 & n52027 ) ;
  assign n52029 = n51189 ^ n33274 ^ n24266 ;
  assign n52030 = n52029 ^ n800 ^ 1'b0 ;
  assign n52031 = n1319 & n9752 ;
  assign n52032 = n15568 ^ n6660 ^ 1'b0 ;
  assign n52033 = n52031 | n52032 ;
  assign n52034 = ( n6324 & ~n29067 ) | ( n6324 & n52033 ) | ( ~n29067 & n52033 ) ;
  assign n52035 = ( x229 & n52030 ) | ( x229 & ~n52034 ) | ( n52030 & ~n52034 ) ;
  assign n52036 = n1588 ^ n962 ^ 1'b0 ;
  assign n52037 = ( n22878 & n50895 ) | ( n22878 & ~n52036 ) | ( n50895 & ~n52036 ) ;
  assign n52038 = n14868 & n52037 ;
  assign n52039 = n28996 ^ n21653 ^ x13 ;
  assign n52040 = ( n34050 & ~n40579 ) | ( n34050 & n52039 ) | ( ~n40579 & n52039 ) ;
  assign n52041 = n7217 ^ n6731 ^ n5595 ;
  assign n52042 = n52041 ^ n18001 ^ 1'b0 ;
  assign n52043 = n40602 ^ n35820 ^ n35414 ;
  assign n52044 = ~n15055 & n52043 ;
  assign n52045 = n52044 ^ n29059 ^ 1'b0 ;
  assign n52046 = n7546 | n18072 ;
  assign n52047 = n3339 | n52046 ;
  assign n52048 = n9235 ^ n1627 ^ n1272 ;
  assign n52049 = ~n37271 & n52048 ;
  assign n52050 = ( ~n9581 & n42533 ) | ( ~n9581 & n52049 ) | ( n42533 & n52049 ) ;
  assign n52051 = ( ~n27132 & n52047 ) | ( ~n27132 & n52050 ) | ( n52047 & n52050 ) ;
  assign n52052 = n2840 | n27389 ;
  assign n52053 = n52051 & ~n52052 ;
  assign n52054 = n3439 & ~n12896 ;
  assign n52055 = n52054 ^ n15689 ^ 1'b0 ;
  assign n52056 = n52055 ^ n18558 ^ n1649 ;
  assign n52057 = ~n37459 & n52056 ;
  assign n52058 = n52057 ^ n46862 ^ 1'b0 ;
  assign n52059 = n52058 ^ n20574 ^ n19155 ;
  assign n52060 = n33865 ^ n2947 ^ 1'b0 ;
  assign n52061 = n52060 ^ n44713 ^ n5601 ;
  assign n52062 = ( n12099 & n29923 ) | ( n12099 & n52061 ) | ( n29923 & n52061 ) ;
  assign n52063 = ~n36846 & n40695 ;
  assign n52064 = n24095 ^ n8374 ^ n471 ;
  assign n52065 = ( n11885 & ~n29427 ) | ( n11885 & n52064 ) | ( ~n29427 & n52064 ) ;
  assign n52069 = n12826 ^ n890 ^ 1'b0 ;
  assign n52068 = n458 | n35895 ;
  assign n52070 = n52069 ^ n52068 ^ 1'b0 ;
  assign n52066 = ( n12178 & n18513 ) | ( n12178 & n26677 ) | ( n18513 & n26677 ) ;
  assign n52067 = n52066 ^ n44817 ^ n33915 ;
  assign n52071 = n52070 ^ n52067 ^ n5696 ;
  assign n52072 = n52071 ^ n50099 ^ n3226 ;
  assign n52073 = ( ~n23545 & n38964 ) | ( ~n23545 & n39610 ) | ( n38964 & n39610 ) ;
  assign n52074 = n38499 | n43197 ;
  assign n52075 = n52074 ^ n27746 ^ 1'b0 ;
  assign n52076 = n34177 ^ n20936 ^ n7827 ;
  assign n52077 = n52076 ^ n26450 ^ 1'b0 ;
  assign n52078 = n8538 & n52077 ;
  assign n52079 = n25503 & n52078 ;
  assign n52080 = n52079 ^ n11367 ^ 1'b0 ;
  assign n52081 = n31823 & n52080 ;
  assign n52082 = ~n15801 & n46571 ;
  assign n52083 = n52082 ^ n11341 ^ 1'b0 ;
  assign n52084 = n17844 ^ n4825 ^ 1'b0 ;
  assign n52085 = n12970 & ~n52084 ;
  assign n52087 = n17488 ^ n3427 ^ n2052 ;
  assign n52086 = n26833 ^ x156 ^ 1'b0 ;
  assign n52088 = n52087 ^ n52086 ^ 1'b0 ;
  assign n52089 = n3965 & n31213 ;
  assign n52090 = n7483 | n52089 ;
  assign n52091 = ( n9697 & n10702 ) | ( n9697 & n32296 ) | ( n10702 & n32296 ) ;
  assign n52092 = n13548 ^ n8946 ^ 1'b0 ;
  assign n52093 = n52092 ^ n30444 ^ n1331 ;
  assign n52094 = n675 & n23967 ;
  assign n52095 = n25610 & n52094 ;
  assign n52096 = ( n23926 & n37357 ) | ( n23926 & n52095 ) | ( n37357 & n52095 ) ;
  assign n52097 = n8553 & ~n34265 ;
  assign n52098 = n52097 ^ n43519 ^ 1'b0 ;
  assign n52099 = n16930 ^ n9641 ^ n5566 ;
  assign n52100 = ~n3838 & n52099 ;
  assign n52101 = n37649 & n50716 ;
  assign n52102 = ~n40686 & n52101 ;
  assign n52103 = n52102 ^ n712 ^ 1'b0 ;
  assign n52104 = ~n8290 & n52103 ;
  assign n52105 = n41760 ^ n13130 ^ n6107 ;
  assign n52106 = n31649 ^ n4248 ^ 1'b0 ;
  assign n52107 = n52105 & ~n52106 ;
  assign n52108 = n20124 ^ n13380 ^ 1'b0 ;
  assign n52109 = n8676 | n52108 ;
  assign n52110 = n52109 ^ n11523 ^ n2602 ;
  assign n52113 = ( n18471 & ~n34077 ) | ( n18471 & n39437 ) | ( ~n34077 & n39437 ) ;
  assign n52114 = ( n12902 & n33323 ) | ( n12902 & n52113 ) | ( n33323 & n52113 ) ;
  assign n52112 = n22064 ^ n18625 ^ n8426 ;
  assign n52111 = n8419 & n11572 ;
  assign n52115 = n52114 ^ n52112 ^ n52111 ;
  assign n52116 = ( n6962 & n43633 ) | ( n6962 & ~n44744 ) | ( n43633 & ~n44744 ) ;
  assign n52117 = n18481 ^ n2114 ^ n1034 ;
  assign n52118 = n2768 | n52117 ;
  assign n52119 = ( n3606 & n12275 ) | ( n3606 & ~n26141 ) | ( n12275 & ~n26141 ) ;
  assign n52120 = ( n11658 & n37476 ) | ( n11658 & ~n52119 ) | ( n37476 & ~n52119 ) ;
  assign n52121 = ( n1967 & n35840 ) | ( n1967 & n52120 ) | ( n35840 & n52120 ) ;
  assign n52122 = ( n3107 & n23102 ) | ( n3107 & ~n25048 ) | ( n23102 & ~n25048 ) ;
  assign n52123 = n30297 | n52122 ;
  assign n52124 = n10007 ^ n8667 ^ x192 ;
  assign n52125 = ( n11197 & n16242 ) | ( n11197 & n52124 ) | ( n16242 & n52124 ) ;
  assign n52126 = n11048 & n52125 ;
  assign n52127 = n52126 ^ n25794 ^ n19491 ;
  assign n52128 = n26629 | n52127 ;
  assign n52129 = n52128 ^ n7073 ^ 1'b0 ;
  assign n52130 = ~n1399 & n40907 ;
  assign n52131 = n10654 & n52130 ;
  assign n52134 = n37251 ^ n11685 ^ n5170 ;
  assign n52132 = ~n34929 & n45291 ;
  assign n52133 = n15609 & n52132 ;
  assign n52135 = n52134 ^ n52133 ^ 1'b0 ;
  assign n52136 = n7926 | n22525 ;
  assign n52137 = n24140 & ~n52136 ;
  assign n52138 = n24084 ^ n14539 ^ n3490 ;
  assign n52139 = n39665 ^ n10131 ^ 1'b0 ;
  assign n52140 = n14958 | n52139 ;
  assign n52141 = n42826 ^ n25018 ^ 1'b0 ;
  assign n52142 = ( n11727 & n52140 ) | ( n11727 & ~n52141 ) | ( n52140 & ~n52141 ) ;
  assign n52152 = ( ~n5708 & n12275 ) | ( ~n5708 & n13066 ) | ( n12275 & n13066 ) ;
  assign n52150 = n26253 ^ n7080 ^ 1'b0 ;
  assign n52151 = n47151 & n52150 ;
  assign n52143 = n10340 ^ n9697 ^ 1'b0 ;
  assign n52145 = n28403 ^ n13123 ^ n6919 ;
  assign n52144 = n13232 | n22608 ;
  assign n52146 = n52145 ^ n52144 ^ 1'b0 ;
  assign n52147 = n15450 & n52146 ;
  assign n52148 = ( n19200 & n52143 ) | ( n19200 & n52147 ) | ( n52143 & n52147 ) ;
  assign n52149 = n52148 ^ n5327 ^ 1'b0 ;
  assign n52153 = n52152 ^ n52151 ^ n52149 ;
  assign n52155 = n28595 ^ n22807 ^ n6270 ;
  assign n52154 = n18328 ^ n9443 ^ n5664 ;
  assign n52156 = n52155 ^ n52154 ^ n19989 ;
  assign n52157 = n31731 ^ n27033 ^ 1'b0 ;
  assign n52158 = ~n2686 & n52157 ;
  assign n52159 = ( n7503 & n16093 ) | ( n7503 & n52158 ) | ( n16093 & n52158 ) ;
  assign n52160 = n52159 ^ n38039 ^ n12996 ;
  assign n52161 = ( n4360 & ~n12891 ) | ( n4360 & n42555 ) | ( ~n12891 & n42555 ) ;
  assign n52162 = n46891 ^ n37729 ^ 1'b0 ;
  assign n52163 = ~n8398 & n52162 ;
  assign n52164 = n52163 ^ n16199 ^ n15139 ;
  assign n52165 = ~n8327 & n52164 ;
  assign n52166 = n9577 & ~n10804 ;
  assign n52167 = n52166 ^ n42169 ^ 1'b0 ;
  assign n52170 = ( n3040 & n4145 ) | ( n3040 & ~n7809 ) | ( n4145 & ~n7809 ) ;
  assign n52169 = ( n2648 & n7630 ) | ( n2648 & n16055 ) | ( n7630 & n16055 ) ;
  assign n52171 = n52170 ^ n52169 ^ 1'b0 ;
  assign n52168 = n5810 | n21863 ;
  assign n52172 = n52171 ^ n52168 ^ 1'b0 ;
  assign n52173 = n24174 ^ n4662 ^ 1'b0 ;
  assign n52174 = n27647 | n52173 ;
  assign n52175 = ( ~n17942 & n36961 ) | ( ~n17942 & n52174 ) | ( n36961 & n52174 ) ;
  assign n52176 = n52175 ^ n37128 ^ n13802 ;
  assign n52180 = n18971 ^ n11301 ^ n2705 ;
  assign n52177 = n29543 ^ n18121 ^ 1'b0 ;
  assign n52178 = n35681 ^ n7365 ^ 1'b0 ;
  assign n52179 = n52177 & ~n52178 ;
  assign n52181 = n52180 ^ n52179 ^ n25638 ;
  assign n52182 = ~n7660 & n27845 ;
  assign n52183 = n28046 ^ n25416 ^ 1'b0 ;
  assign n52184 = n27426 & n52183 ;
  assign n52185 = n40695 ^ n31317 ^ n8173 ;
  assign n52186 = ~n3841 & n30475 ;
  assign n52187 = n12310 & n52186 ;
  assign n52188 = n52187 ^ n13465 ^ n1462 ;
  assign n52189 = n19828 & ~n37786 ;
  assign n52190 = n24351 ^ n12262 ^ 1'b0 ;
  assign n52191 = n27193 & n52190 ;
  assign n52192 = n22332 ^ n8309 ^ 1'b0 ;
  assign n52193 = n52191 | n52192 ;
  assign n52194 = ~n6566 & n52193 ;
  assign n52195 = n52194 ^ n7044 ^ 1'b0 ;
  assign n52196 = n6511 | n36195 ;
  assign n52197 = n12409 ^ n8368 ^ 1'b0 ;
  assign n52198 = n8773 | n52197 ;
  assign n52199 = ( n580 & n16239 ) | ( n580 & ~n18623 ) | ( n16239 & ~n18623 ) ;
  assign n52200 = n4298 ^ n3860 ^ 1'b0 ;
  assign n52201 = n38258 ^ n6947 ^ 1'b0 ;
  assign n52202 = n1845 | n52201 ;
  assign n52203 = n52202 ^ n10263 ^ 1'b0 ;
  assign n52204 = n43481 ^ n37159 ^ n14370 ;
  assign n52205 = n52204 ^ n31249 ^ n2349 ;
  assign n52206 = ( ~n6362 & n35415 ) | ( ~n6362 & n36758 ) | ( n35415 & n36758 ) ;
  assign n52207 = n42927 ^ n36201 ^ n3398 ;
  assign n52208 = n11861 ^ n7173 ^ x199 ;
  assign n52209 = n52208 ^ n42631 ^ 1'b0 ;
  assign n52210 = n8957 & n52209 ;
  assign n52215 = ( n9216 & n12237 ) | ( n9216 & n23054 ) | ( n12237 & n23054 ) ;
  assign n52214 = n2775 | n50329 ;
  assign n52216 = n52215 ^ n52214 ^ 1'b0 ;
  assign n52211 = n36311 ^ n22274 ^ n20147 ;
  assign n52212 = ~n9974 & n52211 ;
  assign n52213 = n51163 & n52212 ;
  assign n52217 = n52216 ^ n52213 ^ 1'b0 ;
  assign n52218 = n31895 ^ n20167 ^ n4638 ;
  assign n52219 = ~n16168 & n52218 ;
  assign n52220 = n52219 ^ n32565 ^ 1'b0 ;
  assign n52221 = n52220 ^ n15009 ^ n3865 ;
  assign n52222 = n31035 ^ n27567 ^ n27109 ;
  assign n52223 = ( n6083 & n18690 ) | ( n6083 & ~n52222 ) | ( n18690 & ~n52222 ) ;
  assign n52224 = ( n2087 & n21658 ) | ( n2087 & ~n51256 ) | ( n21658 & ~n51256 ) ;
  assign n52225 = ( n15084 & n43009 ) | ( n15084 & ~n52224 ) | ( n43009 & ~n52224 ) ;
  assign n52226 = n17566 ^ n17023 ^ n14593 ;
  assign n52227 = n51108 ^ n41142 ^ n21528 ;
  assign n52228 = n25736 | n51041 ;
  assign n52229 = n52228 ^ n1450 ^ 1'b0 ;
  assign n52230 = n52229 ^ n24352 ^ n721 ;
  assign n52231 = ( n6874 & n16121 ) | ( n6874 & ~n16715 ) | ( n16121 & ~n16715 ) ;
  assign n52232 = ~n21423 & n52231 ;
  assign n52233 = n52232 ^ n12534 ^ 1'b0 ;
  assign n52234 = n18073 & ~n49744 ;
  assign n52235 = ~n48746 & n52234 ;
  assign n52236 = n52233 & n52235 ;
  assign n52237 = n8183 & ~n52236 ;
  assign n52238 = ~n23040 & n43989 ;
  assign n52239 = n40154 & n52238 ;
  assign n52240 = n39035 & ~n52239 ;
  assign n52241 = n52240 ^ n48233 ^ 1'b0 ;
  assign n52242 = n52241 ^ n37144 ^ n33198 ;
  assign n52243 = n29040 ^ n688 ^ 1'b0 ;
  assign n52244 = n52242 & ~n52243 ;
  assign n52245 = n7254 & n12740 ;
  assign n52246 = n11071 & n52245 ;
  assign n52247 = n52246 ^ n51354 ^ 1'b0 ;
  assign n52248 = n414 & n30105 ;
  assign n52249 = n52248 ^ n3591 ^ 1'b0 ;
  assign n52250 = n8139 & n52249 ;
  assign n52251 = ~n23499 & n52250 ;
  assign n52252 = ~n52247 & n52251 ;
  assign n52253 = n1495 & n17514 ;
  assign n52257 = n13442 ^ n13353 ^ n7073 ;
  assign n52254 = n9363 ^ n4773 ^ 1'b0 ;
  assign n52255 = n8927 & n26621 ;
  assign n52256 = n52254 & n52255 ;
  assign n52258 = n52257 ^ n52256 ^ n34959 ;
  assign n52259 = n52258 ^ n43063 ^ n7771 ;
  assign n52260 = n38528 & ~n48101 ;
  assign n52261 = ( n6045 & ~n20313 ) | ( n6045 & n34694 ) | ( ~n20313 & n34694 ) ;
  assign n52262 = ( n15121 & ~n27356 ) | ( n15121 & n30361 ) | ( ~n27356 & n30361 ) ;
  assign n52263 = ( n2617 & ~n38345 ) | ( n2617 & n52262 ) | ( ~n38345 & n52262 ) ;
  assign n52264 = n30998 ^ n8992 ^ 1'b0 ;
  assign n52265 = n32907 & n50716 ;
  assign n52266 = n52265 ^ n1760 ^ 1'b0 ;
  assign n52267 = n30420 ^ n18571 ^ 1'b0 ;
  assign n52268 = ~n26545 & n52267 ;
  assign n52269 = ~n8964 & n42689 ;
  assign n52270 = n52269 ^ n33337 ^ n10182 ;
  assign n52271 = n52270 ^ n918 ^ 1'b0 ;
  assign n52273 = n23906 & ~n26158 ;
  assign n52274 = n52273 ^ n26113 ^ 1'b0 ;
  assign n52272 = ~x55 & n13954 ;
  assign n52275 = n52274 ^ n52272 ^ 1'b0 ;
  assign n52276 = n19347 & n28752 ;
  assign n52277 = n52276 ^ n8705 ^ 1'b0 ;
  assign n52278 = n52277 ^ n39794 ^ n32540 ;
  assign n52279 = ( ~n6166 & n32498 ) | ( ~n6166 & n33177 ) | ( n32498 & n33177 ) ;
  assign n52280 = ~n33269 & n42872 ;
  assign n52281 = n26372 & n52280 ;
  assign n52282 = ( n49890 & n52279 ) | ( n49890 & ~n52281 ) | ( n52279 & ~n52281 ) ;
  assign n52283 = n36071 ^ n812 ^ 1'b0 ;
  assign n52284 = ( ~n23240 & n30127 ) | ( ~n23240 & n52283 ) | ( n30127 & n52283 ) ;
  assign n52285 = n48803 ^ n48284 ^ 1'b0 ;
  assign n52286 = n41374 ^ n28024 ^ n3992 ;
  assign n52287 = ~n10099 & n25189 ;
  assign n52288 = ~n52177 & n52287 ;
  assign n52289 = ( n4594 & n9027 ) | ( n4594 & ~n52288 ) | ( n9027 & ~n52288 ) ;
  assign n52290 = n22747 | n32137 ;
  assign n52291 = n11968 & ~n52290 ;
  assign n52292 = ~n6439 & n29970 ;
  assign n52293 = n52292 ^ n35445 ^ 1'b0 ;
  assign n52294 = ~n7726 & n50217 ;
  assign n52295 = n52294 ^ n32496 ^ 1'b0 ;
  assign n52296 = n20304 & ~n29699 ;
  assign n52297 = n52296 ^ n8088 ^ n4480 ;
  assign n52298 = ( ~n4985 & n7822 ) | ( ~n4985 & n36756 ) | ( n7822 & n36756 ) ;
  assign n52299 = n356 & ~n15504 ;
  assign n52300 = ~n477 & n52299 ;
  assign n52301 = ( n17553 & n44845 ) | ( n17553 & n52300 ) | ( n44845 & n52300 ) ;
  assign n52302 = n43747 ^ n12825 ^ n6406 ;
  assign n52303 = ( n4975 & n45551 ) | ( n4975 & ~n52302 ) | ( n45551 & ~n52302 ) ;
  assign n52304 = n38802 ^ n38419 ^ n29898 ;
  assign n52305 = n7543 & n22154 ;
  assign n52306 = n52305 ^ n13792 ^ 1'b0 ;
  assign n52307 = n16800 | n51868 ;
  assign n52308 = n40011 & ~n52307 ;
  assign n52309 = n40288 ^ n15370 ^ 1'b0 ;
  assign n52310 = n22313 ^ n2907 ^ 1'b0 ;
  assign n52311 = n52310 ^ n48881 ^ 1'b0 ;
  assign n52312 = n770 & ~n38188 ;
  assign n52313 = ( n44800 & n51454 ) | ( n44800 & ~n52312 ) | ( n51454 & ~n52312 ) ;
  assign n52314 = n51868 ^ n46963 ^ n1924 ;
  assign n52315 = n20098 & n52314 ;
  assign n52316 = n25324 ^ n6503 ^ 1'b0 ;
  assign n52317 = ( n22339 & n29691 ) | ( n22339 & ~n52316 ) | ( n29691 & ~n52316 ) ;
  assign n52318 = n52317 ^ n18384 ^ n9487 ;
  assign n52319 = n46040 ^ n43604 ^ n684 ;
  assign n52320 = ( n5189 & n8391 ) | ( n5189 & ~n10363 ) | ( n8391 & ~n10363 ) ;
  assign n52321 = ( n939 & n2040 ) | ( n939 & ~n52320 ) | ( n2040 & ~n52320 ) ;
  assign n52322 = ( n6541 & ~n21358 ) | ( n6541 & n52321 ) | ( ~n21358 & n52321 ) ;
  assign n52323 = n52322 ^ n17081 ^ n1395 ;
  assign n52324 = n52323 ^ n32108 ^ 1'b0 ;
  assign n52325 = n22150 ^ n12763 ^ 1'b0 ;
  assign n52326 = n32040 | n52325 ;
  assign n52327 = n36171 ^ n32226 ^ 1'b0 ;
  assign n52328 = n27457 ^ n24079 ^ 1'b0 ;
  assign n52329 = n38453 & n52328 ;
  assign n52330 = n24152 ^ n14032 ^ 1'b0 ;
  assign n52331 = n41527 & ~n48964 ;
  assign n52332 = ( n2924 & n22886 ) | ( n2924 & ~n33003 ) | ( n22886 & ~n33003 ) ;
  assign n52333 = ( n20984 & ~n26414 ) | ( n20984 & n33881 ) | ( ~n26414 & n33881 ) ;
  assign n52334 = ( n45111 & ~n52332 ) | ( n45111 & n52333 ) | ( ~n52332 & n52333 ) ;
  assign n52341 = n8664 & ~n26887 ;
  assign n52342 = n52341 ^ n12834 ^ 1'b0 ;
  assign n52338 = n15168 | n16317 ;
  assign n52339 = n403 | n52338 ;
  assign n52335 = ( ~n6873 & n12924 ) | ( ~n6873 & n13916 ) | ( n12924 & n13916 ) ;
  assign n52336 = n52335 ^ n20728 ^ n8857 ;
  assign n52337 = ~n15671 & n52336 ;
  assign n52340 = n52339 ^ n52337 ^ 1'b0 ;
  assign n52343 = n52342 ^ n52340 ^ n23106 ;
  assign n52344 = n7517 | n18352 ;
  assign n52345 = n52344 ^ n46337 ^ 1'b0 ;
  assign n52346 = n52345 ^ n21494 ^ 1'b0 ;
  assign n52347 = n50172 & ~n52346 ;
  assign n52348 = n5284 & ~n52347 ;
  assign n52349 = n1421 | n26352 ;
  assign n52350 = ( n11801 & n21635 ) | ( n11801 & ~n52349 ) | ( n21635 & ~n52349 ) ;
  assign n52351 = n37440 ^ n29217 ^ n11376 ;
  assign n52352 = n9234 & n42039 ;
  assign n52353 = n7679 & n35218 ;
  assign n52354 = n52353 ^ n25690 ^ 1'b0 ;
  assign n52355 = n7721 & n43315 ;
  assign n52356 = n46331 ^ n10895 ^ 1'b0 ;
  assign n52357 = ~n34424 & n52356 ;
  assign n52358 = n6879 ^ n2644 ^ 1'b0 ;
  assign n52359 = n1185 | n52358 ;
  assign n52360 = n22150 ^ n13163 ^ 1'b0 ;
  assign n52361 = n52359 | n52360 ;
  assign n52362 = n46804 ^ n46796 ^ n5740 ;
  assign n52363 = ~n10284 & n26168 ;
  assign n52364 = ( ~n12621 & n36451 ) | ( ~n12621 & n52363 ) | ( n36451 & n52363 ) ;
  assign n52365 = n11477 & ~n21174 ;
  assign n52366 = n10766 | n33176 ;
  assign n52367 = n52366 ^ n25248 ^ 1'b0 ;
  assign n52368 = n52367 ^ n34822 ^ n2178 ;
  assign n52369 = n52368 ^ n12110 ^ n9836 ;
  assign n52370 = n4365 & n37430 ;
  assign n52371 = n52369 & n52370 ;
  assign n52372 = ( ~n52333 & n52365 ) | ( ~n52333 & n52371 ) | ( n52365 & n52371 ) ;
  assign n52373 = ( n3962 & n11656 ) | ( n3962 & ~n21227 ) | ( n11656 & ~n21227 ) ;
  assign n52374 = ( n14837 & n35403 ) | ( n14837 & n52373 ) | ( n35403 & n52373 ) ;
  assign n52375 = ( n11735 & ~n11956 ) | ( n11735 & n26703 ) | ( ~n11956 & n26703 ) ;
  assign n52376 = n27797 ^ n17851 ^ n5720 ;
  assign n52377 = n28004 ^ n12609 ^ 1'b0 ;
  assign n52378 = n3248 & n52377 ;
  assign n52379 = n25787 | n52378 ;
  assign n52380 = n52379 ^ n25645 ^ 1'b0 ;
  assign n52381 = n9036 & ~n13651 ;
  assign n52382 = n387 & n52381 ;
  assign n52383 = n17769 ^ n388 ^ 1'b0 ;
  assign n52385 = ( n2615 & n18101 ) | ( n2615 & n25404 ) | ( n18101 & n25404 ) ;
  assign n52386 = n27762 | n52385 ;
  assign n52387 = n26636 & ~n52386 ;
  assign n52384 = ~n8560 & n18521 ;
  assign n52388 = n52387 ^ n52384 ^ n21122 ;
  assign n52389 = n25335 ^ n20194 ^ 1'b0 ;
  assign n52390 = n15579 & ~n52389 ;
  assign n52391 = ( n28902 & ~n36006 ) | ( n28902 & n52390 ) | ( ~n36006 & n52390 ) ;
  assign n52392 = n35484 & ~n52211 ;
  assign n52393 = n21014 ^ n2459 ^ 1'b0 ;
  assign n52394 = n52393 ^ n46933 ^ n6989 ;
  assign n52395 = ( n6536 & ~n11824 ) | ( n6536 & n52394 ) | ( ~n11824 & n52394 ) ;
  assign n52396 = n22834 ^ n14061 ^ 1'b0 ;
  assign n52397 = n9973 ^ n3064 ^ 1'b0 ;
  assign n52398 = ~n6789 & n47702 ;
  assign n52399 = ~n37937 & n52398 ;
  assign n52400 = ~n1809 & n14169 ;
  assign n52401 = n52400 ^ n12018 ^ 1'b0 ;
  assign n52402 = n44145 ^ n33904 ^ n22183 ;
  assign n52403 = n52401 | n52402 ;
  assign n52404 = n39016 ^ n2340 ^ 1'b0 ;
  assign n52405 = n14690 | n52404 ;
  assign n52406 = ( ~n8459 & n13318 ) | ( ~n8459 & n16890 ) | ( n13318 & n16890 ) ;
  assign n52407 = ( n2504 & ~n38846 ) | ( n2504 & n39522 ) | ( ~n38846 & n39522 ) ;
  assign n52408 = n14975 ^ n6219 ^ n4295 ;
  assign n52409 = n15444 ^ n12302 ^ 1'b0 ;
  assign n52410 = n8139 & n52409 ;
  assign n52411 = n35006 & ~n52410 ;
  assign n52412 = n40417 ^ n8820 ^ 1'b0 ;
  assign n52413 = n21036 ^ n7253 ^ n6170 ;
  assign n52414 = n44349 | n52413 ;
  assign n52415 = n16722 | n52414 ;
  assign n52416 = n11802 & n36531 ;
  assign n52417 = n52416 ^ n9279 ^ 1'b0 ;
  assign n52418 = n6486 & n52417 ;
  assign n52419 = n26134 & n52418 ;
  assign n52420 = ~n10922 & n46921 ;
  assign n52421 = n52420 ^ n10482 ^ 1'b0 ;
  assign n52422 = n28886 ^ n5850 ^ 1'b0 ;
  assign n52423 = n30433 & n52422 ;
  assign n52424 = n11875 & n49386 ;
  assign n52425 = n52424 ^ n1850 ^ n826 ;
  assign n52426 = n50936 ^ n21582 ^ n2314 ;
  assign n52427 = n10335 ^ n8667 ^ n2780 ;
  assign n52429 = ~n11732 & n43153 ;
  assign n52430 = ~n49002 & n52429 ;
  assign n52428 = n15742 & ~n19791 ;
  assign n52431 = n52430 ^ n52428 ^ n22053 ;
  assign n52432 = ( n14994 & n19175 ) | ( n14994 & ~n28993 ) | ( n19175 & ~n28993 ) ;
  assign n52433 = n38741 ^ n23260 ^ 1'b0 ;
  assign n52434 = n52432 | n52433 ;
  assign n52439 = n7477 & ~n44527 ;
  assign n52435 = n24820 & n29827 ;
  assign n52436 = n7198 & ~n30480 ;
  assign n52437 = n52435 & n52436 ;
  assign n52438 = n42437 | n52437 ;
  assign n52440 = n52439 ^ n52438 ^ 1'b0 ;
  assign n52441 = n50647 ^ n48512 ^ 1'b0 ;
  assign n52442 = n46616 & ~n52441 ;
  assign n52443 = n280 | n49726 ;
  assign n52446 = n22757 ^ n19172 ^ 1'b0 ;
  assign n52444 = n41477 ^ n10173 ^ 1'b0 ;
  assign n52445 = n52444 ^ n27200 ^ n6388 ;
  assign n52447 = n52446 ^ n52445 ^ n11532 ;
  assign n52448 = ( n1550 & n49199 ) | ( n1550 & ~n52447 ) | ( n49199 & ~n52447 ) ;
  assign n52449 = ( n2062 & n31472 ) | ( n2062 & n31890 ) | ( n31472 & n31890 ) ;
  assign n52450 = n45861 ^ n20690 ^ 1'b0 ;
  assign n52451 = n1680 & ~n52450 ;
  assign n52452 = ( n11729 & n22414 ) | ( n11729 & ~n52451 ) | ( n22414 & ~n52451 ) ;
  assign n52453 = n40670 ^ n6101 ^ 1'b0 ;
  assign n52454 = n19083 ^ n13715 ^ n4169 ;
  assign n52455 = ( ~n2935 & n24290 ) | ( ~n2935 & n30744 ) | ( n24290 & n30744 ) ;
  assign n52456 = ( ~n11371 & n20379 ) | ( ~n11371 & n52455 ) | ( n20379 & n52455 ) ;
  assign n52457 = n52456 ^ n33870 ^ n24454 ;
  assign n52458 = n34694 ^ n3651 ^ 1'b0 ;
  assign n52459 = ~n52457 & n52458 ;
  assign n52460 = n10792 & n17156 ;
  assign n52461 = n52460 ^ n16712 ^ n6259 ;
  assign n52462 = ( n43359 & n52459 ) | ( n43359 & ~n52461 ) | ( n52459 & ~n52461 ) ;
  assign n52463 = ( ~n268 & n5665 ) | ( ~n268 & n15981 ) | ( n5665 & n15981 ) ;
  assign n52464 = n28237 ^ n6559 ^ n353 ;
  assign n52465 = n36891 & n52464 ;
  assign n52466 = ~n52463 & n52465 ;
  assign n52467 = n6741 ^ n5542 ^ 1'b0 ;
  assign n52468 = n1003 & n22437 ;
  assign n52469 = n4222 & n18239 ;
  assign n52474 = n849 & ~n5149 ;
  assign n52472 = n25960 ^ n23908 ^ n8990 ;
  assign n52470 = n16222 ^ n1527 ^ 1'b0 ;
  assign n52471 = n20143 & n52470 ;
  assign n52473 = n52472 ^ n52471 ^ n1098 ;
  assign n52475 = n52474 ^ n52473 ^ n5208 ;
  assign n52476 = n10300 ^ n8397 ^ 1'b0 ;
  assign n52477 = n35470 | n52476 ;
  assign n52478 = n52477 ^ n43937 ^ n15899 ;
  assign n52479 = ( n32931 & n48953 ) | ( n32931 & n49615 ) | ( n48953 & n49615 ) ;
  assign n52483 = ~n4216 & n19371 ;
  assign n52484 = n8988 & n52483 ;
  assign n52485 = n52484 ^ n49903 ^ n9758 ;
  assign n52482 = n8084 ^ n6918 ^ n3863 ;
  assign n52480 = n13399 ^ n3562 ^ 1'b0 ;
  assign n52481 = n10136 & n52480 ;
  assign n52486 = n52485 ^ n52482 ^ n52481 ;
  assign n52487 = n20507 | n21344 ;
  assign n52488 = n43611 ^ n17602 ^ 1'b0 ;
  assign n52489 = n3164 | n44030 ;
  assign n52490 = n20766 & ~n52489 ;
  assign n52491 = n22618 ^ n5026 ^ 1'b0 ;
  assign n52492 = n2606 & ~n52491 ;
  assign n52493 = n52492 ^ n20088 ^ 1'b0 ;
  assign n52494 = n49261 ^ n24040 ^ n17426 ;
  assign n52495 = n34009 ^ n26415 ^ n5515 ;
  assign n52496 = n5675 | n31931 ;
  assign n52497 = ( n41063 & n43054 ) | ( n41063 & ~n52496 ) | ( n43054 & ~n52496 ) ;
  assign n52498 = n39809 ^ n21240 ^ n15752 ;
  assign n52499 = ( n24703 & ~n28225 ) | ( n24703 & n52498 ) | ( ~n28225 & n52498 ) ;
  assign n52500 = n21770 ^ n18607 ^ 1'b0 ;
  assign n52501 = n37615 | n52500 ;
  assign n52502 = n28308 ^ n14358 ^ 1'b0 ;
  assign n52503 = ( ~n32409 & n52501 ) | ( ~n32409 & n52502 ) | ( n52501 & n52502 ) ;
  assign n52504 = n32638 | n45340 ;
  assign n52505 = n8156 | n52504 ;
  assign n52506 = n9108 & n23900 ;
  assign n52507 = n52506 ^ n28750 ^ 1'b0 ;
  assign n52508 = n19804 & n36385 ;
  assign n52509 = ( n30007 & ~n34216 ) | ( n30007 & n48957 ) | ( ~n34216 & n48957 ) ;
  assign n52512 = n39510 ^ n38105 ^ n24843 ;
  assign n52511 = ( n1257 & n16054 ) | ( n1257 & ~n21588 ) | ( n16054 & ~n21588 ) ;
  assign n52510 = ( n4716 & n7926 ) | ( n4716 & n19807 ) | ( n7926 & n19807 ) ;
  assign n52513 = n52512 ^ n52511 ^ n52510 ;
  assign n52514 = ~n6674 & n8777 ;
  assign n52515 = n52514 ^ n4450 ^ 1'b0 ;
  assign n52516 = ( n2892 & n17123 ) | ( n2892 & ~n17221 ) | ( n17123 & ~n17221 ) ;
  assign n52517 = ( n3587 & ~n52515 ) | ( n3587 & n52516 ) | ( ~n52515 & n52516 ) ;
  assign n52518 = n2785 & n22868 ;
  assign n52519 = n52518 ^ n6390 ^ 1'b0 ;
  assign n52520 = n52519 ^ n49508 ^ n43341 ;
  assign n52521 = ( ~n1632 & n11598 ) | ( ~n1632 & n24375 ) | ( n11598 & n24375 ) ;
  assign n52522 = n2546 | n52521 ;
  assign n52523 = ( n5236 & ~n42990 ) | ( n5236 & n51089 ) | ( ~n42990 & n51089 ) ;
  assign n52524 = n19197 ^ n5303 ^ 1'b0 ;
  assign n52525 = n52523 | n52524 ;
  assign n52527 = ~n8393 & n24182 ;
  assign n52528 = ~n10582 & n52527 ;
  assign n52529 = n52528 ^ n29085 ^ 1'b0 ;
  assign n52530 = ~n12709 & n52529 ;
  assign n52526 = ~n16920 & n38790 ;
  assign n52531 = n52530 ^ n52526 ^ n42653 ;
  assign n52532 = n17385 & ~n52531 ;
  assign n52533 = n32299 | n41596 ;
  assign n52534 = n9604 & n11157 ;
  assign n52535 = n52534 ^ n34443 ^ 1'b0 ;
  assign n52536 = ( ~n36539 & n41170 ) | ( ~n36539 & n52535 ) | ( n41170 & n52535 ) ;
  assign n52537 = n52536 ^ n36314 ^ n3760 ;
  assign n52538 = n11122 ^ n1545 ^ 1'b0 ;
  assign n52539 = n18813 ^ n2633 ^ 1'b0 ;
  assign n52540 = n23668 & n24810 ;
  assign n52541 = n4080 & n28301 ;
  assign n52542 = n52541 ^ n8928 ^ 1'b0 ;
  assign n52543 = ( n15889 & n29251 ) | ( n15889 & n52542 ) | ( n29251 & n52542 ) ;
  assign n52544 = n11178 & n52543 ;
  assign n52545 = n18035 ^ n5081 ^ 1'b0 ;
  assign n52546 = ~n1681 & n52545 ;
  assign n52547 = n31176 ^ n12219 ^ n11891 ;
  assign n52548 = n12812 | n52547 ;
  assign n52549 = n42105 ^ n3605 ^ 1'b0 ;
  assign n52550 = n898 & n31071 ;
  assign n52551 = n52550 ^ n11593 ^ n7695 ;
  assign n52552 = n36085 ^ n9932 ^ 1'b0 ;
  assign n52553 = n40199 | n51718 ;
  assign n52559 = n15556 & ~n33206 ;
  assign n52560 = n52559 ^ n698 ^ 1'b0 ;
  assign n52557 = ~n8130 & n31305 ;
  assign n52558 = ~x72 & n52557 ;
  assign n52561 = n52560 ^ n52558 ^ n16528 ;
  assign n52554 = n26712 & ~n41622 ;
  assign n52555 = ~n3532 & n52554 ;
  assign n52556 = n52555 ^ n49476 ^ n30390 ;
  assign n52562 = n52561 ^ n52556 ^ n42020 ;
  assign n52563 = ( ~n4475 & n29077 ) | ( ~n4475 & n52562 ) | ( n29077 & n52562 ) ;
  assign n52564 = n20976 ^ n2523 ^ 1'b0 ;
  assign n52565 = n315 | n52564 ;
  assign n52566 = n52565 ^ n27531 ^ 1'b0 ;
  assign n52567 = n52070 & ~n52566 ;
  assign n52568 = n27505 ^ n7473 ^ 1'b0 ;
  assign n52569 = n8066 & ~n52568 ;
  assign n52570 = ( ~n2882 & n4342 ) | ( ~n2882 & n17852 ) | ( n4342 & n17852 ) ;
  assign n52571 = n52570 ^ n5928 ^ 1'b0 ;
  assign n52572 = x6 & n52571 ;
  assign n52573 = n39947 ^ n29317 ^ n17598 ;
  assign n52574 = n30412 & n32579 ;
  assign n52575 = n52573 & n52574 ;
  assign n52576 = x64 ^ x55 ^ 1'b0 ;
  assign n52577 = n10395 ^ n3136 ^ 1'b0 ;
  assign n52578 = ( n24505 & ~n25414 ) | ( n24505 & n52577 ) | ( ~n25414 & n52577 ) ;
  assign n52579 = n52578 ^ n652 ^ 1'b0 ;
  assign n52580 = ( ~n27302 & n41404 ) | ( ~n27302 & n52579 ) | ( n41404 & n52579 ) ;
  assign n52583 = n6786 & n16095 ;
  assign n52584 = n8205 & n52583 ;
  assign n52581 = n23515 ^ n19766 ^ 1'b0 ;
  assign n52582 = ~n26866 & n52581 ;
  assign n52585 = n52584 ^ n52582 ^ n32809 ;
  assign n52586 = n24064 & ~n37673 ;
  assign n52587 = n52586 ^ n9630 ^ n6479 ;
  assign n52588 = n18679 | n34959 ;
  assign n52589 = ~n1897 & n28431 ;
  assign n52590 = n52589 ^ n2765 ^ 1'b0 ;
  assign n52591 = ( ~n16504 & n52588 ) | ( ~n16504 & n52590 ) | ( n52588 & n52590 ) ;
  assign n52592 = n18033 ^ n12407 ^ 1'b0 ;
  assign n52593 = n23650 | n52592 ;
  assign n52594 = n52593 ^ n47542 ^ n16350 ;
  assign n52595 = n34331 ^ n30364 ^ 1'b0 ;
  assign n52596 = n50811 | n52595 ;
  assign n52597 = n8424 & ~n23549 ;
  assign n52598 = n3596 & n4975 ;
  assign n52599 = n52598 ^ n11435 ^ 1'b0 ;
  assign n52600 = n1317 & n3967 ;
  assign n52601 = n15518 & n52600 ;
  assign n52602 = n52601 ^ n14477 ^ n13546 ;
  assign n52603 = n38774 & n52602 ;
  assign n52604 = n35850 & n52603 ;
  assign n52605 = n34899 ^ n2310 ^ 1'b0 ;
  assign n52606 = n26390 ^ n17884 ^ n10226 ;
  assign n52607 = ( n5098 & n20531 ) | ( n5098 & n52606 ) | ( n20531 & n52606 ) ;
  assign n52608 = n42462 ^ n23839 ^ x186 ;
  assign n52609 = n7839 ^ n477 ^ 1'b0 ;
  assign n52610 = ( n5353 & n44239 ) | ( n5353 & ~n52609 ) | ( n44239 & ~n52609 ) ;
  assign n52611 = n22845 ^ n13590 ^ 1'b0 ;
  assign n52612 = n23001 & n24928 ;
  assign n52613 = n16607 & n41170 ;
  assign n52614 = n52613 ^ n29020 ^ 1'b0 ;
  assign n52615 = n2857 ^ n2642 ^ 1'b0 ;
  assign n52616 = n16730 & n52615 ;
  assign n52617 = ~n3670 & n7473 ;
  assign n52618 = n902 & ~n15509 ;
  assign n52619 = ~n13917 & n52618 ;
  assign n52621 = ( n2592 & n40756 ) | ( n2592 & n51492 ) | ( n40756 & n51492 ) ;
  assign n52622 = ( n9730 & n32932 ) | ( n9730 & ~n52621 ) | ( n32932 & ~n52621 ) ;
  assign n52620 = n9673 & n15298 ;
  assign n52623 = n52622 ^ n52620 ^ 1'b0 ;
  assign n52624 = ~n52619 & n52623 ;
  assign n52625 = ( n27275 & n52617 ) | ( n27275 & n52624 ) | ( n52617 & n52624 ) ;
  assign n52626 = n38832 ^ n5412 ^ 1'b0 ;
  assign n52627 = ~n19797 & n28604 ;
  assign n52628 = ~n929 & n52627 ;
  assign n52629 = ( n2526 & n10243 ) | ( n2526 & n52628 ) | ( n10243 & n52628 ) ;
  assign n52630 = n34849 | n52629 ;
  assign n52631 = n45834 & ~n52630 ;
  assign n52632 = ( ~n9390 & n52626 ) | ( ~n9390 & n52631 ) | ( n52626 & n52631 ) ;
  assign n52633 = n26417 ^ n18578 ^ 1'b0 ;
  assign n52634 = n20987 & ~n52633 ;
  assign n52635 = n47025 ^ n25481 ^ n14721 ;
  assign n52636 = ( n10474 & n19242 ) | ( n10474 & n52635 ) | ( n19242 & n52635 ) ;
  assign n52638 = n1612 ^ n601 ^ 1'b0 ;
  assign n52639 = n52066 | n52638 ;
  assign n52637 = n21415 ^ n16580 ^ 1'b0 ;
  assign n52640 = n52639 ^ n52637 ^ n11400 ;
  assign n52641 = ( n1346 & n52636 ) | ( n1346 & n52640 ) | ( n52636 & n52640 ) ;
  assign n52642 = ( ~n31339 & n38859 ) | ( ~n31339 & n42186 ) | ( n38859 & n42186 ) ;
  assign n52643 = n49023 | n52642 ;
  assign n52644 = ( n3002 & n15794 ) | ( n3002 & ~n52643 ) | ( n15794 & ~n52643 ) ;
  assign n52645 = ( ~n14567 & n30852 ) | ( ~n14567 & n36294 ) | ( n30852 & n36294 ) ;
  assign n52646 = n7843 ^ n6010 ^ n303 ;
  assign n52647 = ~n8873 & n52646 ;
  assign n52648 = n31417 ^ n2036 ^ 1'b0 ;
  assign n52649 = n34370 | n52648 ;
  assign n52650 = n6201 ^ n2180 ^ 1'b0 ;
  assign n52651 = ~n52649 & n52650 ;
  assign n52652 = n52651 ^ n2847 ^ 1'b0 ;
  assign n52653 = n14347 & ~n52652 ;
  assign n52654 = n23700 ^ n21419 ^ n19590 ;
  assign n52655 = n52654 ^ n35564 ^ 1'b0 ;
  assign n52656 = n52653 & ~n52655 ;
  assign n52657 = ( n3090 & n9581 ) | ( n3090 & ~n23431 ) | ( n9581 & ~n23431 ) ;
  assign n52658 = ~n18755 & n52657 ;
  assign n52659 = ( n4166 & n39792 ) | ( n4166 & ~n39819 ) | ( n39792 & ~n39819 ) ;
  assign n52660 = n33482 | n52659 ;
  assign n52661 = n50038 & n51875 ;
  assign n52662 = n10077 & ~n14992 ;
  assign n52663 = ( ~n3627 & n45279 ) | ( ~n3627 & n52662 ) | ( n45279 & n52662 ) ;
  assign n52664 = n780 & n2943 ;
  assign n52665 = n20149 & n52664 ;
  assign n52666 = ( n4975 & n23512 ) | ( n4975 & ~n37027 ) | ( n23512 & ~n37027 ) ;
  assign n52667 = ( n26076 & n30541 ) | ( n26076 & n52666 ) | ( n30541 & n52666 ) ;
  assign n52668 = ( ~n12302 & n15207 ) | ( ~n12302 & n45174 ) | ( n15207 & n45174 ) ;
  assign n52669 = n27099 | n52668 ;
  assign n52670 = n27093 ^ n20930 ^ 1'b0 ;
  assign n52671 = n7923 & n11089 ;
  assign n52672 = n52671 ^ n9766 ^ 1'b0 ;
  assign n52673 = n490 | n8214 ;
  assign n52674 = ( ~n47475 & n52672 ) | ( ~n47475 & n52673 ) | ( n52672 & n52673 ) ;
  assign n52675 = n7878 & n10495 ;
  assign n52676 = n52675 ^ n2329 ^ 1'b0 ;
  assign n52677 = n18337 ^ n5343 ^ 1'b0 ;
  assign n52678 = n52676 & n52677 ;
  assign n52679 = n27944 ^ n4018 ^ x174 ;
  assign n52680 = n52678 | n52679 ;
  assign n52681 = n32728 ^ n4283 ^ 1'b0 ;
  assign n52682 = ~n15637 & n52681 ;
  assign n52683 = n52682 ^ n49610 ^ n11463 ;
  assign n52684 = n52683 ^ n888 ^ 1'b0 ;
  assign n52685 = n8718 | n52684 ;
  assign n52686 = n52685 ^ n12066 ^ 1'b0 ;
  assign n52688 = ~n8460 & n16944 ;
  assign n52687 = n2109 & ~n16279 ;
  assign n52689 = n52688 ^ n52687 ^ 1'b0 ;
  assign n52690 = n49671 ^ n19450 ^ 1'b0 ;
  assign n52691 = n52689 | n52690 ;
  assign n52692 = n35892 ^ n7906 ^ n1572 ;
  assign n52693 = ~n11376 & n35370 ;
  assign n52694 = ( n7483 & n8376 ) | ( n7483 & n42749 ) | ( n8376 & n42749 ) ;
  assign n52695 = n10949 & n20267 ;
  assign n52696 = ~n1680 & n52695 ;
  assign n52697 = ( ~n52693 & n52694 ) | ( ~n52693 & n52696 ) | ( n52694 & n52696 ) ;
  assign n52698 = ( n1941 & n3775 ) | ( n1941 & n37840 ) | ( n3775 & n37840 ) ;
  assign n52699 = ( n12019 & ~n29575 ) | ( n12019 & n52698 ) | ( ~n29575 & n52698 ) ;
  assign n52700 = n52699 ^ n27254 ^ n12899 ;
  assign n52707 = n5855 & ~n13578 ;
  assign n52708 = n11948 ^ n9964 ^ 1'b0 ;
  assign n52709 = ( n14474 & n52707 ) | ( n14474 & n52708 ) | ( n52707 & n52708 ) ;
  assign n52703 = n21258 ^ n6860 ^ n6803 ;
  assign n52701 = ~n10797 & n29261 ;
  assign n52702 = n35406 & n52701 ;
  assign n52704 = n52703 ^ n52702 ^ 1'b0 ;
  assign n52705 = n2754 & ~n52704 ;
  assign n52706 = ~n3713 & n52705 ;
  assign n52710 = n52709 ^ n52706 ^ n51606 ;
  assign n52711 = n7217 | n20650 ;
  assign n52712 = n44556 ^ n18120 ^ n644 ;
  assign n52713 = n52712 ^ n9125 ^ n5574 ;
  assign n52714 = n16594 & n36603 ;
  assign n52715 = n52714 ^ n44713 ^ n20942 ;
  assign n52716 = ~n50471 & n52715 ;
  assign n52717 = n52716 ^ n51220 ^ 1'b0 ;
  assign n52718 = ~n5979 & n43137 ;
  assign n52719 = n46174 ^ n22449 ^ n4556 ;
  assign n52720 = n22079 | n27005 ;
  assign n52721 = n36496 | n52720 ;
  assign n52722 = n52721 ^ n21791 ^ 1'b0 ;
  assign n52723 = n8743 & ~n52722 ;
  assign n52724 = n38049 ^ n7759 ^ 1'b0 ;
  assign n52725 = ( n11016 & n16063 ) | ( n11016 & n23976 ) | ( n16063 & n23976 ) ;
  assign n52726 = ~n37181 & n52725 ;
  assign n52727 = n34926 & n52726 ;
  assign n52728 = n52727 ^ n504 ^ 1'b0 ;
  assign n52729 = n52728 ^ n46162 ^ n2866 ;
  assign n52730 = ( n19121 & n20000 ) | ( n19121 & n46411 ) | ( n20000 & n46411 ) ;
  assign n52731 = n25134 ^ n23590 ^ n8155 ;
  assign n52732 = ( n2083 & ~n52730 ) | ( n2083 & n52731 ) | ( ~n52730 & n52731 ) ;
  assign n52733 = n12133 ^ n1792 ^ 1'b0 ;
  assign n52734 = n3067 | n51390 ;
  assign n52735 = n707 | n25693 ;
  assign n52736 = n52735 ^ n11614 ^ 1'b0 ;
  assign n52737 = ~n6635 & n10903 ;
  assign n52738 = n52736 & n52737 ;
  assign n52739 = n11970 & ~n24084 ;
  assign n52740 = n12769 & n52739 ;
  assign n52741 = ~n9431 & n37116 ;
  assign n52742 = n29274 & n52741 ;
  assign n52743 = ( n14840 & n38428 ) | ( n14840 & n47701 ) | ( n38428 & n47701 ) ;
  assign n52744 = n52743 ^ n33697 ^ n11904 ;
  assign n52745 = n5048 & ~n19754 ;
  assign n52746 = n52745 ^ n29931 ^ 1'b0 ;
  assign n52747 = ( n15568 & n21348 ) | ( n15568 & ~n52746 ) | ( n21348 & ~n52746 ) ;
  assign n52748 = n8294 ^ n4071 ^ 1'b0 ;
  assign n52749 = n17490 & n51607 ;
  assign n52750 = ~n43187 & n52749 ;
  assign n52751 = ~n28001 & n52750 ;
  assign n52752 = n31945 ^ n1668 ^ 1'b0 ;
  assign n52753 = n19350 & n52752 ;
  assign n52754 = ( ~n17790 & n31005 ) | ( ~n17790 & n52753 ) | ( n31005 & n52753 ) ;
  assign n52755 = n33881 ^ n30984 ^ n9650 ;
  assign n52756 = n26769 ^ n14539 ^ 1'b0 ;
  assign n52757 = n26744 | n52756 ;
  assign n52758 = n41586 & ~n52757 ;
  assign n52759 = ( n685 & ~n13154 ) | ( n685 & n26636 ) | ( ~n13154 & n26636 ) ;
  assign n52760 = n52759 ^ n34648 ^ n18587 ;
  assign n52761 = n52760 ^ n35145 ^ 1'b0 ;
  assign n52762 = ~n16798 & n52761 ;
  assign n52763 = ( ~n1673 & n32661 ) | ( ~n1673 & n39014 ) | ( n32661 & n39014 ) ;
  assign n52764 = ~n3557 & n8686 ;
  assign n52765 = n52764 ^ n38859 ^ n26481 ;
  assign n52766 = n8256 | n10057 ;
  assign n52767 = n17976 | n34965 ;
  assign n52768 = n10905 ^ n5793 ^ 1'b0 ;
  assign n52769 = ( ~n25349 & n52767 ) | ( ~n25349 & n52768 ) | ( n52767 & n52768 ) ;
  assign n52770 = n30045 ^ n6728 ^ 1'b0 ;
  assign n52771 = n52770 ^ n41132 ^ n27029 ;
  assign n52772 = n565 & ~n48041 ;
  assign n52773 = n28477 ^ n2214 ^ 1'b0 ;
  assign n52774 = n38493 | n52773 ;
  assign n52775 = n52774 ^ n15359 ^ 1'b0 ;
  assign n52776 = n29808 | n52775 ;
  assign n52777 = ~n10892 & n11552 ;
  assign n52778 = n12817 & n52777 ;
  assign n52779 = n37622 | n52778 ;
  assign n52780 = n17156 ^ n7007 ^ 1'b0 ;
  assign n52781 = ~n20784 & n46345 ;
  assign n52782 = n52781 ^ n1646 ^ 1'b0 ;
  assign n52783 = n52782 ^ n27218 ^ n21793 ;
  assign n52784 = n50086 ^ n17761 ^ 1'b0 ;
  assign n52785 = ( n5370 & n21211 ) | ( n5370 & ~n49251 ) | ( n21211 & ~n49251 ) ;
  assign n52786 = ( ~n7927 & n12206 ) | ( ~n7927 & n52785 ) | ( n12206 & n52785 ) ;
  assign n52787 = n38515 ^ n7922 ^ 1'b0 ;
  assign n52788 = n42173 ^ n19170 ^ n2545 ;
  assign n52789 = n10807 & ~n13070 ;
  assign n52790 = n52789 ^ n4141 ^ 1'b0 ;
  assign n52791 = n18791 | n52790 ;
  assign n52792 = n52791 ^ n24508 ^ 1'b0 ;
  assign n52793 = ~n13892 & n18062 ;
  assign n52794 = n10675 & n52793 ;
  assign n52795 = n808 & n18818 ;
  assign n52796 = ~n17058 & n52795 ;
  assign n52797 = n10922 ^ n7671 ^ 1'b0 ;
  assign n52798 = n25931 | n52797 ;
  assign n52799 = n35043 ^ n30529 ^ n1582 ;
  assign n52800 = n13613 & ~n52799 ;
  assign n52801 = n52798 & n52800 ;
  assign n52803 = ( n2605 & n37999 ) | ( n2605 & ~n40828 ) | ( n37999 & ~n40828 ) ;
  assign n52802 = n25775 ^ n17101 ^ 1'b0 ;
  assign n52804 = n52803 ^ n52802 ^ n8272 ;
  assign n52805 = ~n3324 & n18658 ;
  assign n52806 = n52805 ^ n7089 ^ 1'b0 ;
  assign n52807 = ( n6320 & n52804 ) | ( n6320 & n52806 ) | ( n52804 & n52806 ) ;
  assign n52808 = n30370 & n43128 ;
  assign n52809 = n52808 ^ n23026 ^ n13215 ;
  assign n52810 = n2409 & ~n5970 ;
  assign n52811 = ( n3274 & ~n13574 ) | ( n3274 & n52810 ) | ( ~n13574 & n52810 ) ;
  assign n52812 = n20217 & n52811 ;
  assign n52813 = n36346 & ~n52812 ;
  assign n52814 = n44446 ^ n30388 ^ n5228 ;
  assign n52815 = n52171 ^ n4650 ^ 1'b0 ;
  assign n52816 = n31245 & ~n52815 ;
  assign n52817 = ( n14751 & n16634 ) | ( n14751 & ~n26059 ) | ( n16634 & ~n26059 ) ;
  assign n52818 = n52817 ^ n28545 ^ n16957 ;
  assign n52819 = ( ~n2895 & n14744 ) | ( ~n2895 & n20066 ) | ( n14744 & n20066 ) ;
  assign n52820 = n6647 & ~n52819 ;
  assign n52821 = ~n25957 & n52820 ;
  assign n52822 = n44886 ^ n42426 ^ n37635 ;
  assign n52823 = n10091 & n52822 ;
  assign n52824 = n52823 ^ n38533 ^ 1'b0 ;
  assign n52825 = ~n15501 & n42186 ;
  assign n52826 = ~n22414 & n52825 ;
  assign n52827 = ~n30116 & n49280 ;
  assign n52828 = ~n23242 & n52827 ;
  assign n52829 = ( n1946 & ~n4686 ) | ( n1946 & n41011 ) | ( ~n4686 & n41011 ) ;
  assign n52830 = n52829 ^ n39996 ^ n34768 ;
  assign n52831 = ( n2066 & n2252 ) | ( n2066 & n11915 ) | ( n2252 & n11915 ) ;
  assign n52832 = n8087 & ~n34732 ;
  assign n52833 = ( n18314 & n52831 ) | ( n18314 & ~n52832 ) | ( n52831 & ~n52832 ) ;
  assign n52834 = n35096 ^ n3441 ^ 1'b0 ;
  assign n52835 = ~n17391 & n52834 ;
  assign n52836 = n2724 & n45150 ;
  assign n52837 = ~n52835 & n52836 ;
  assign n52838 = ( n5611 & ~n52833 ) | ( n5611 & n52837 ) | ( ~n52833 & n52837 ) ;
  assign n52839 = n11160 | n21590 ;
  assign n52840 = n52839 ^ n27489 ^ n21970 ;
  assign n52841 = ( n4155 & ~n31340 ) | ( n4155 & n52840 ) | ( ~n31340 & n52840 ) ;
  assign n52842 = n5930 | n25484 ;
  assign n52843 = ( n502 & n4666 ) | ( n502 & ~n13583 ) | ( n4666 & ~n13583 ) ;
  assign n52844 = ( n27953 & ~n46258 ) | ( n27953 & n52843 ) | ( ~n46258 & n52843 ) ;
  assign n52845 = n52844 ^ n16588 ^ 1'b0 ;
  assign n52846 = n28179 ^ n13718 ^ n12076 ;
  assign n52847 = n52846 ^ n16560 ^ n12562 ;
  assign n52848 = n4070 & ~n25541 ;
  assign n52849 = n18955 & ~n48882 ;
  assign n52850 = n52848 & n52849 ;
  assign n52851 = ( ~n20135 & n40963 ) | ( ~n20135 & n47175 ) | ( n40963 & n47175 ) ;
  assign n52852 = ~n16953 & n52851 ;
  assign n52853 = n52852 ^ n2120 ^ 1'b0 ;
  assign n52854 = n25650 ^ n6359 ^ 1'b0 ;
  assign n52855 = n13043 & n21338 ;
  assign n52856 = ~n19290 & n52855 ;
  assign n52857 = ( n5710 & n16616 ) | ( n5710 & ~n24621 ) | ( n16616 & ~n24621 ) ;
  assign n52858 = ( n5613 & ~n33621 ) | ( n5613 & n52857 ) | ( ~n33621 & n52857 ) ;
  assign n52859 = n22394 & ~n52858 ;
  assign n52860 = n52859 ^ n52371 ^ 1'b0 ;
  assign n52863 = x72 & n1544 ;
  assign n52864 = n22250 & n52863 ;
  assign n52861 = ~n5501 & n16128 ;
  assign n52862 = ~n15232 & n52861 ;
  assign n52865 = n52864 ^ n52862 ^ n38872 ;
  assign n52866 = n36592 ^ n10656 ^ 1'b0 ;
  assign n52867 = n18304 | n52866 ;
  assign n52868 = ( n3199 & n28139 ) | ( n3199 & n52867 ) | ( n28139 & n52867 ) ;
  assign n52869 = ( n1072 & n36882 ) | ( n1072 & ~n52868 ) | ( n36882 & ~n52868 ) ;
  assign n52870 = n14416 ^ n13645 ^ 1'b0 ;
  assign n52871 = ~n29769 & n52870 ;
  assign n52872 = n52871 ^ n16483 ^ n14870 ;
  assign n52873 = n35835 ^ n24901 ^ n2967 ;
  assign n52874 = ~n14425 & n17115 ;
  assign n52875 = n10039 | n52874 ;
  assign n52876 = n37543 ^ n6755 ^ 1'b0 ;
  assign n52877 = ~n37139 & n51941 ;
  assign n52878 = ~n14977 & n52877 ;
  assign n52879 = n6020 | n40189 ;
  assign n52880 = n34318 | n52879 ;
  assign n52881 = n5218 | n49151 ;
  assign n52882 = n51902 | n52881 ;
  assign n52883 = n47851 & n52882 ;
  assign n52884 = n29562 ^ n17255 ^ 1'b0 ;
  assign n52885 = n50010 ^ n21919 ^ 1'b0 ;
  assign n52886 = ( n3422 & n4500 ) | ( n3422 & n13099 ) | ( n4500 & n13099 ) ;
  assign n52887 = ( n14583 & n15498 ) | ( n14583 & n52886 ) | ( n15498 & n52886 ) ;
  assign n52888 = n6642 | n8428 ;
  assign n52889 = n17602 & ~n52888 ;
  assign n52890 = n12465 ^ n6185 ^ 1'b0 ;
  assign n52891 = ~n12227 & n52890 ;
  assign n52892 = ( n11772 & n52889 ) | ( n11772 & n52891 ) | ( n52889 & n52891 ) ;
  assign n52893 = ( ~n3826 & n19611 ) | ( ~n3826 & n20499 ) | ( n19611 & n20499 ) ;
  assign n52894 = n2851 & ~n52893 ;
  assign n52895 = ~n14629 & n52894 ;
  assign n52896 = n24919 ^ n12046 ^ n3613 ;
  assign n52897 = ( n15018 & n52895 ) | ( n15018 & ~n52896 ) | ( n52895 & ~n52896 ) ;
  assign n52898 = n25928 & ~n27671 ;
  assign n52899 = n52898 ^ n14603 ^ 1'b0 ;
  assign n52900 = n15655 ^ n15144 ^ 1'b0 ;
  assign n52901 = n52899 | n52900 ;
  assign n52902 = ~n12237 & n46908 ;
  assign n52903 = n25079 ^ n15328 ^ 1'b0 ;
  assign n52904 = ~n33174 & n52903 ;
  assign n52905 = n18316 & n30623 ;
  assign n52906 = n52905 ^ n52221 ^ 1'b0 ;
  assign n52907 = ~n28462 & n52906 ;
  assign n52908 = ( ~x229 & n824 ) | ( ~x229 & n29696 ) | ( n824 & n29696 ) ;
  assign n52909 = n6701 & ~n12735 ;
  assign n52910 = ( ~n2357 & n7463 ) | ( ~n2357 & n51309 ) | ( n7463 & n51309 ) ;
  assign n52911 = ( n1005 & n52909 ) | ( n1005 & n52910 ) | ( n52909 & n52910 ) ;
  assign n52912 = ( n18675 & n44207 ) | ( n18675 & ~n45358 ) | ( n44207 & ~n45358 ) ;
  assign n52913 = n39459 ^ n2027 ^ 1'b0 ;
  assign n52914 = n17283 | n52913 ;
  assign n52915 = ( n10249 & n17600 ) | ( n10249 & n52914 ) | ( n17600 & n52914 ) ;
  assign n52917 = n10884 & ~n25488 ;
  assign n52918 = ~n23589 & n52917 ;
  assign n52919 = n52918 ^ n36058 ^ n7228 ;
  assign n52916 = ( n1481 & n11526 ) | ( n1481 & n18936 ) | ( n11526 & n18936 ) ;
  assign n52920 = n52919 ^ n52916 ^ n9944 ;
  assign n52921 = n37100 & ~n37795 ;
  assign n52922 = ~n2569 & n52921 ;
  assign n52923 = n40862 ^ n9120 ^ 1'b0 ;
  assign n52924 = n14181 & ~n52923 ;
  assign n52925 = ( n8654 & n11364 ) | ( n8654 & ~n13634 ) | ( n11364 & ~n13634 ) ;
  assign n52926 = n16462 ^ n11589 ^ n6127 ;
  assign n52927 = ( n35047 & n39418 ) | ( n35047 & n52926 ) | ( n39418 & n52926 ) ;
  assign n52928 = n14804 | n52927 ;
  assign n52929 = n52925 | n52928 ;
  assign n52930 = n5202 | n7597 ;
  assign n52931 = n52930 ^ n1163 ^ 1'b0 ;
  assign n52932 = n10009 & ~n18821 ;
  assign n52934 = n6076 | n14215 ;
  assign n52935 = n4333 & ~n52934 ;
  assign n52933 = ( x184 & n18229 ) | ( x184 & ~n34346 ) | ( n18229 & ~n34346 ) ;
  assign n52936 = n52935 ^ n52933 ^ n1318 ;
  assign n52937 = n18304 & ~n52936 ;
  assign n52938 = n44882 ^ n15137 ^ n12408 ;
  assign n52939 = n8260 | n11106 ;
  assign n52940 = n52939 ^ n30372 ^ 1'b0 ;
  assign n52941 = n7556 & ~n35916 ;
  assign n52942 = n52940 & n52941 ;
  assign n52943 = ~n3182 & n52942 ;
  assign n52944 = n23997 ^ n23549 ^ 1'b0 ;
  assign n52945 = ~n1211 & n52944 ;
  assign n52946 = n5629 & n14319 ;
  assign n52947 = ( n15174 & ~n52945 ) | ( n15174 & n52946 ) | ( ~n52945 & n52946 ) ;
  assign n52948 = n45986 ^ n8333 ^ 1'b0 ;
  assign n52949 = ~n10884 & n52948 ;
  assign n52950 = ( n30022 & ~n51054 ) | ( n30022 & n52949 ) | ( ~n51054 & n52949 ) ;
  assign n52951 = n6418 & ~n16284 ;
  assign n52952 = ~n10505 & n52951 ;
  assign n52953 = n1623 & n32184 ;
  assign n52954 = n52953 ^ n12235 ^ 1'b0 ;
  assign n52955 = n33776 & n38876 ;
  assign n52956 = n25009 ^ n12801 ^ 1'b0 ;
  assign n52957 = n21572 & ~n52956 ;
  assign n52958 = n49336 ^ n28019 ^ 1'b0 ;
  assign n52959 = n52254 ^ n24409 ^ n7178 ;
  assign n52960 = n20654 ^ n4087 ^ n1893 ;
  assign n52961 = n16022 ^ n6399 ^ 1'b0 ;
  assign n52962 = ( n750 & ~n13656 ) | ( n750 & n52961 ) | ( ~n13656 & n52961 ) ;
  assign n52963 = n27032 ^ n24667 ^ 1'b0 ;
  assign n52964 = n52963 ^ n23307 ^ n21926 ;
  assign n52965 = ( n12799 & ~n42876 ) | ( n12799 & n51245 ) | ( ~n42876 & n51245 ) ;
  assign n52966 = n38192 | n43896 ;
  assign n52967 = n52966 ^ n18567 ^ 1'b0 ;
  assign n52968 = n660 | n7596 ;
  assign n52969 = n9108 | n52968 ;
  assign n52970 = n52969 ^ n27619 ^ 1'b0 ;
  assign n52971 = n9857 & n52970 ;
  assign n52972 = ~n6989 & n42409 ;
  assign n52973 = n52972 ^ n11798 ^ 1'b0 ;
  assign n52974 = ( n5835 & n10423 ) | ( n5835 & n52973 ) | ( n10423 & n52973 ) ;
  assign n52975 = n21802 | n25738 ;
  assign n52976 = n52975 ^ n22170 ^ 1'b0 ;
  assign n52977 = ( n29003 & ~n31037 ) | ( n29003 & n52976 ) | ( ~n31037 & n52976 ) ;
  assign n52978 = n41652 & ~n49009 ;
  assign n52979 = ~n21853 & n52978 ;
  assign n52980 = ( ~n20331 & n51370 ) | ( ~n20331 & n52979 ) | ( n51370 & n52979 ) ;
  assign n52981 = n13696 & ~n24489 ;
  assign n52982 = n32765 ^ n26981 ^ n24385 ;
  assign n52983 = ( n29883 & n34270 ) | ( n29883 & n52982 ) | ( n34270 & n52982 ) ;
  assign n52984 = n5471 ^ n1746 ^ 1'b0 ;
  assign n52985 = ~n28734 & n52984 ;
  assign n52986 = ~n20546 & n52985 ;
  assign n52987 = n14476 ^ n11054 ^ 1'b0 ;
  assign n52988 = n1284 | n14781 ;
  assign n52989 = n42251 & ~n52988 ;
  assign n52990 = n13004 & n52989 ;
  assign n52991 = n29173 ^ n17230 ^ n2539 ;
  assign n52992 = n31477 ^ n21401 ^ 1'b0 ;
  assign n52993 = n10469 ^ n9832 ^ n6160 ;
  assign n52994 = n52993 ^ n47695 ^ n42286 ;
  assign n52995 = ( n980 & ~n1039 ) | ( n980 & n3006 ) | ( ~n1039 & n3006 ) ;
  assign n52996 = n52995 ^ n41482 ^ n23420 ;
  assign n52997 = n41413 ^ n4440 ^ 1'b0 ;
  assign n52998 = n47476 ^ n40526 ^ 1'b0 ;
  assign n52999 = n16764 ^ x215 ^ 1'b0 ;
  assign n53000 = ( ~n3333 & n20144 ) | ( ~n3333 & n24425 ) | ( n20144 & n24425 ) ;
  assign n53001 = ( n1305 & n52999 ) | ( n1305 & n53000 ) | ( n52999 & n53000 ) ;
  assign n53002 = n26569 & ~n53001 ;
  assign n53003 = n53002 ^ n12856 ^ 1'b0 ;
  assign n53004 = n16372 & n48227 ;
  assign n53005 = ~n52746 & n53004 ;
  assign n53006 = n52481 ^ n9596 ^ 1'b0 ;
  assign n53007 = ~n34475 & n53006 ;
  assign n53008 = ~n8017 & n41231 ;
  assign n53009 = n53008 ^ n8619 ^ 1'b0 ;
  assign n53010 = ( n15456 & n30622 ) | ( n15456 & ~n53009 ) | ( n30622 & ~n53009 ) ;
  assign n53011 = ( n2580 & n29353 ) | ( n2580 & ~n41267 ) | ( n29353 & ~n41267 ) ;
  assign n53012 = n52171 ^ n50450 ^ n34033 ;
  assign n53013 = n39891 ^ n27842 ^ n20873 ;
  assign n53014 = n14501 ^ n11861 ^ n722 ;
  assign n53015 = n53014 ^ n31252 ^ n3306 ;
  assign n53016 = n53015 ^ n50389 ^ n26013 ;
  assign n53017 = ~n31392 & n45170 ;
  assign n53018 = n39409 ^ n20061 ^ 1'b0 ;
  assign n53019 = n11238 & ~n16463 ;
  assign n53020 = n53019 ^ n4119 ^ 1'b0 ;
  assign n53021 = n28574 ^ n10453 ^ 1'b0 ;
  assign n53022 = n53020 & ~n53021 ;
  assign n53023 = n22156 | n36473 ;
  assign n53024 = x145 & n16549 ;
  assign n53025 = n53024 ^ n24792 ^ 1'b0 ;
  assign n53026 = n53025 ^ n30273 ^ 1'b0 ;
  assign n53027 = n32703 & n53026 ;
  assign n53028 = n15105 & ~n31692 ;
  assign n53029 = ( n3081 & n11305 ) | ( n3081 & ~n17737 ) | ( n11305 & ~n17737 ) ;
  assign n53030 = ( n1823 & n17013 ) | ( n1823 & ~n35749 ) | ( n17013 & ~n35749 ) ;
  assign n53031 = n20728 ^ n9037 ^ n366 ;
  assign n53033 = n15182 ^ n11494 ^ n2306 ;
  assign n53032 = n11312 & ~n36905 ;
  assign n53034 = n53033 ^ n53032 ^ n21242 ;
  assign n53035 = n53034 ^ n13053 ^ n1935 ;
  assign n53036 = n3094 & n16068 ;
  assign n53037 = ( ~n20495 & n20583 ) | ( ~n20495 & n38986 ) | ( n20583 & n38986 ) ;
  assign n53038 = n53037 ^ n9992 ^ 1'b0 ;
  assign n53039 = n36242 ^ n17574 ^ 1'b0 ;
  assign n53040 = n18141 & ~n28205 ;
  assign n53041 = n53040 ^ n11058 ^ 1'b0 ;
  assign n53042 = ~n6151 & n18281 ;
  assign n53043 = n53042 ^ n51121 ^ 1'b0 ;
  assign n53044 = n51864 ^ n35491 ^ 1'b0 ;
  assign n53045 = ~n53043 & n53044 ;
  assign n53046 = n50281 | n51948 ;
  assign n53047 = n53046 ^ n5271 ^ 1'b0 ;
  assign n53048 = ( n7805 & ~n37490 ) | ( n7805 & n52498 ) | ( ~n37490 & n52498 ) ;
  assign n53049 = ( n14967 & n17858 ) | ( n14967 & n47843 ) | ( n17858 & n47843 ) ;
  assign n53050 = n28398 ^ n14021 ^ n12358 ;
  assign n53051 = n15883 & ~n36279 ;
  assign n53052 = ~n16697 & n53051 ;
  assign n53053 = n53052 ^ n30166 ^ n9444 ;
  assign n53054 = n46526 ^ n24207 ^ 1'b0 ;
  assign n53055 = n27294 ^ n27224 ^ n16360 ;
  assign n53056 = n3263 & n4780 ;
  assign n53057 = n16107 & ~n40592 ;
  assign n53058 = n53057 ^ n49029 ^ 1'b0 ;
  assign n53059 = n12797 & n13670 ;
  assign n53060 = n53059 ^ n16272 ^ 1'b0 ;
  assign n53061 = n2843 & ~n53060 ;
  assign n53062 = n53061 ^ n4681 ^ 1'b0 ;
  assign n53063 = ( n15216 & ~n18031 ) | ( n15216 & n21280 ) | ( ~n18031 & n21280 ) ;
  assign n53064 = n1206 | n1890 ;
  assign n53065 = n53063 | n53064 ;
  assign n53066 = n9140 & n53065 ;
  assign n53067 = n47776 ^ n40412 ^ 1'b0 ;
  assign n53068 = n20305 ^ n12385 ^ n4231 ;
  assign n53069 = ( n14232 & n40695 ) | ( n14232 & n53068 ) | ( n40695 & n53068 ) ;
  assign n53070 = n53069 ^ n20635 ^ n7700 ;
  assign n53071 = n34713 ^ n24656 ^ 1'b0 ;
  assign n53072 = n8117 ^ n2610 ^ 1'b0 ;
  assign n53073 = n19489 | n53072 ;
  assign n53074 = ( n3500 & n4451 ) | ( n3500 & n13508 ) | ( n4451 & n13508 ) ;
  assign n53075 = ( n11231 & n53073 ) | ( n11231 & ~n53074 ) | ( n53073 & ~n53074 ) ;
  assign n53076 = ( n28060 & ~n41060 ) | ( n28060 & n45538 ) | ( ~n41060 & n45538 ) ;
  assign n53077 = n35688 ^ n28989 ^ n19393 ;
  assign n53078 = n2163 | n31526 ;
  assign n53079 = n3837 | n53078 ;
  assign n53080 = ( n8248 & n11466 ) | ( n8248 & n53079 ) | ( n11466 & n53079 ) ;
  assign n53081 = n3462 & ~n8006 ;
  assign n53082 = ~n17330 & n53081 ;
  assign n53083 = n53082 ^ n32978 ^ 1'b0 ;
  assign n53084 = n53080 | n53083 ;
  assign n53085 = n7779 & ~n32980 ;
  assign n53086 = n53085 ^ n35681 ^ 1'b0 ;
  assign n53087 = n43679 | n53086 ;
  assign n53088 = n33239 & ~n53087 ;
  assign n53089 = n50850 ^ n15888 ^ 1'b0 ;
  assign n53090 = n1359 | n9682 ;
  assign n53091 = n23851 & ~n53090 ;
  assign n53092 = ( n12843 & n53015 ) | ( n12843 & n53091 ) | ( n53015 & n53091 ) ;
  assign n53093 = n40815 ^ n19825 ^ n11673 ;
  assign n53094 = n53093 ^ n32410 ^ n20042 ;
  assign n53095 = n46827 ^ n45866 ^ n26585 ;
  assign n53096 = n24289 & ~n41331 ;
  assign n53097 = n30525 ^ n16658 ^ 1'b0 ;
  assign n53098 = ( ~n7330 & n30621 ) | ( ~n7330 & n47326 ) | ( n30621 & n47326 ) ;
  assign n53099 = ~n17667 & n40971 ;
  assign n53100 = ~n35576 & n53099 ;
  assign n53101 = n952 & n33575 ;
  assign n53102 = n17184 & n53101 ;
  assign n53103 = n8117 & ~n35970 ;
  assign n53104 = n53103 ^ n18593 ^ 1'b0 ;
  assign n53105 = n48126 ^ n46537 ^ n358 ;
  assign n53106 = n8324 & ~n9773 ;
  assign n53107 = ~n10342 & n53106 ;
  assign n53108 = ( ~n7870 & n12109 ) | ( ~n7870 & n53107 ) | ( n12109 & n53107 ) ;
  assign n53109 = n21028 | n30017 ;
  assign n53110 = n24293 & ~n53109 ;
  assign n53111 = n53110 ^ n49389 ^ n41589 ;
  assign n53112 = ( n4522 & n11570 ) | ( n4522 & n42827 ) | ( n11570 & n42827 ) ;
  assign n53113 = n1652 & n6972 ;
  assign n53114 = ( n24852 & n28422 ) | ( n24852 & n53113 ) | ( n28422 & n53113 ) ;
  assign n53115 = ( ~n10743 & n36466 ) | ( ~n10743 & n53114 ) | ( n36466 & n53114 ) ;
  assign n53116 = n45305 ^ n16961 ^ 1'b0 ;
  assign n53117 = n46589 | n46963 ;
  assign n53118 = n53116 | n53117 ;
  assign n53119 = n38250 ^ n15188 ^ 1'b0 ;
  assign n53120 = n11480 | n53119 ;
  assign n53121 = n17894 | n46482 ;
  assign n53122 = n53121 ^ n29324 ^ 1'b0 ;
  assign n53123 = n26918 ^ n16419 ^ 1'b0 ;
  assign n53126 = n13132 ^ n10936 ^ n5036 ;
  assign n53124 = ( n4934 & n7737 ) | ( n4934 & ~n33411 ) | ( n7737 & ~n33411 ) ;
  assign n53125 = n53124 ^ n28470 ^ n9350 ;
  assign n53127 = n53126 ^ n53125 ^ n23580 ;
  assign n53128 = n46038 ^ n30364 ^ n5757 ;
  assign n53129 = n12884 ^ n6520 ^ 1'b0 ;
  assign n53130 = ( ~n30313 & n33170 ) | ( ~n30313 & n36027 ) | ( n33170 & n36027 ) ;
  assign n53131 = n7255 & n28342 ;
  assign n53132 = ~n27179 & n33188 ;
  assign n53133 = n5489 | n38042 ;
  assign n53134 = n53133 ^ n26101 ^ 1'b0 ;
  assign n53135 = n28976 & ~n53134 ;
  assign n53136 = ~n29964 & n53135 ;
  assign n53137 = n2851 & ~n21497 ;
  assign n53138 = n53137 ^ n7563 ^ 1'b0 ;
  assign n53139 = ~n27156 & n53138 ;
  assign n53140 = ( ~n16123 & n24044 ) | ( ~n16123 & n53139 ) | ( n24044 & n53139 ) ;
  assign n53141 = ( n15063 & n15813 ) | ( n15063 & ~n26443 ) | ( n15813 & ~n26443 ) ;
  assign n53142 = ~n4960 & n11163 ;
  assign n53143 = n53142 ^ n36795 ^ 1'b0 ;
  assign n53144 = n24514 & ~n53143 ;
  assign n53145 = n53144 ^ n39440 ^ n31820 ;
  assign n53146 = n22218 | n37672 ;
  assign n53147 = ( n6507 & n9140 ) | ( n6507 & ~n53146 ) | ( n9140 & ~n53146 ) ;
  assign n53152 = n6768 ^ n5912 ^ n5376 ;
  assign n53153 = ( ~n2661 & n32093 ) | ( ~n2661 & n53152 ) | ( n32093 & n53152 ) ;
  assign n53148 = n38078 ^ n16133 ^ 1'b0 ;
  assign n53149 = n52390 & n53148 ;
  assign n53150 = ~n33048 & n53149 ;
  assign n53151 = ~n10049 & n53150 ;
  assign n53154 = n53153 ^ n53151 ^ n5004 ;
  assign n53155 = n43846 ^ n20272 ^ 1'b0 ;
  assign n53156 = n23824 & n53155 ;
  assign n53157 = n53156 ^ n42301 ^ 1'b0 ;
  assign n53158 = n53157 ^ n13131 ^ n6077 ;
  assign n53159 = n536 | n53158 ;
  assign n53160 = n1544 & ~n53159 ;
  assign n53161 = n20537 & n42831 ;
  assign n53162 = n18988 & ~n53161 ;
  assign n53163 = n1881 & n53162 ;
  assign n53164 = n53163 ^ n48771 ^ 1'b0 ;
  assign n53165 = n18272 & n37489 ;
  assign n53166 = x221 & n53165 ;
  assign n53167 = ~n8922 & n53166 ;
  assign n53168 = n33198 ^ n19251 ^ n880 ;
  assign n53169 = ~n320 & n43735 ;
  assign n53170 = n53169 ^ n18609 ^ 1'b0 ;
  assign n53171 = n53170 ^ n51432 ^ n49634 ;
  assign n53172 = ( n9742 & n24320 ) | ( n9742 & n33038 ) | ( n24320 & n33038 ) ;
  assign n53173 = ( n1525 & ~n13502 ) | ( n1525 & n22597 ) | ( ~n13502 & n22597 ) ;
  assign n53174 = n35374 & ~n53173 ;
  assign n53175 = n43810 ^ n26256 ^ n15427 ;
  assign n53176 = n47075 ^ n29861 ^ n10827 ;
  assign n53177 = n12013 ^ n3280 ^ n3019 ;
  assign n53178 = ~n40291 & n53177 ;
  assign n53179 = ( n13153 & n13484 ) | ( n13153 & n33543 ) | ( n13484 & n33543 ) ;
  assign n53180 = ~n14245 & n15263 ;
  assign n53181 = n9010 & n53180 ;
  assign n53182 = ( n19760 & n38861 ) | ( n19760 & ~n53181 ) | ( n38861 & ~n53181 ) ;
  assign n53183 = n53182 ^ n40415 ^ 1'b0 ;
  assign n53192 = n2827 & n38832 ;
  assign n53193 = ( n7174 & n21578 ) | ( n7174 & n53192 ) | ( n21578 & n53192 ) ;
  assign n53191 = ~n27501 & n52171 ;
  assign n53194 = n53193 ^ n53191 ^ n1648 ;
  assign n53184 = n4384 & n11677 ;
  assign n53185 = n35095 & n53184 ;
  assign n53186 = ~n29304 & n53185 ;
  assign n53187 = ~n8382 & n20467 ;
  assign n53188 = ~n53186 & n53187 ;
  assign n53189 = n11671 | n53188 ;
  assign n53190 = n53189 ^ n10761 ^ 1'b0 ;
  assign n53195 = n53194 ^ n53190 ^ n7846 ;
  assign n53196 = ( n24941 & n25188 ) | ( n24941 & n33999 ) | ( n25188 & n33999 ) ;
  assign n53197 = ( ~n1910 & n15510 ) | ( ~n1910 & n53196 ) | ( n15510 & n53196 ) ;
  assign n53198 = n32620 ^ n5730 ^ 1'b0 ;
  assign n53199 = ~n15008 & n53198 ;
  assign n53200 = n4175 & ~n15746 ;
  assign n53201 = n31880 & n53200 ;
  assign n53202 = n4115 & ~n10046 ;
  assign n53203 = n53202 ^ n41238 ^ 1'b0 ;
  assign n53204 = ( n25642 & n32302 ) | ( n25642 & ~n43624 ) | ( n32302 & ~n43624 ) ;
  assign n53205 = ~n16757 & n53204 ;
  assign n53206 = n53205 ^ n2605 ^ 1'b0 ;
  assign n53207 = n5131 & n24917 ;
  assign n53208 = n18160 & n53207 ;
  assign n53209 = n13513 | n40451 ;
  assign n53210 = n49500 | n53209 ;
  assign n53211 = n53210 ^ n43525 ^ 1'b0 ;
  assign n53212 = n36581 ^ n14719 ^ n1643 ;
  assign n53213 = ( n14619 & n16472 ) | ( n14619 & ~n45424 ) | ( n16472 & ~n45424 ) ;
  assign n53214 = n30428 & n35638 ;
  assign n53215 = ( ~n20469 & n26252 ) | ( ~n20469 & n41782 ) | ( n26252 & n41782 ) ;
  assign n53216 = n26463 ^ n20427 ^ 1'b0 ;
  assign n53217 = n27904 | n53216 ;
  assign n53218 = ~n13944 & n49750 ;
  assign n53219 = ~n37220 & n50666 ;
  assign n53220 = n37253 & n53219 ;
  assign n53221 = n31543 ^ n14594 ^ 1'b0 ;
  assign n53222 = n22012 | n53221 ;
  assign n53223 = ( n6174 & n30398 ) | ( n6174 & n51858 ) | ( n30398 & n51858 ) ;
  assign n53224 = n34056 ^ n22936 ^ 1'b0 ;
  assign n53226 = ~x83 & n2124 ;
  assign n53227 = n42064 & ~n53226 ;
  assign n53228 = ~n24603 & n53227 ;
  assign n53225 = n31245 ^ n24643 ^ n3307 ;
  assign n53229 = n53228 ^ n53225 ^ n7573 ;
  assign n53230 = n32218 ^ n27180 ^ 1'b0 ;
  assign n53231 = n22066 ^ n21431 ^ n3760 ;
  assign n53232 = n53231 ^ n27816 ^ n17870 ;
  assign n53233 = n30053 ^ n4579 ^ 1'b0 ;
  assign n53234 = n12861 & n53233 ;
  assign n53235 = n35631 ^ n23647 ^ n15849 ;
  assign n53236 = n53235 ^ n50075 ^ n13593 ;
  assign n53237 = ( n11324 & n53234 ) | ( n11324 & n53236 ) | ( n53234 & n53236 ) ;
  assign n53238 = n2145 & n14132 ;
  assign n53239 = n53238 ^ n43588 ^ 1'b0 ;
  assign n53240 = n5981 & n43053 ;
  assign n53241 = n53240 ^ n20385 ^ 1'b0 ;
  assign n53242 = n4937 & n18158 ;
  assign n53243 = n20639 & n53242 ;
  assign n53244 = ( n10132 & n22711 ) | ( n10132 & ~n29647 ) | ( n22711 & ~n29647 ) ;
  assign n53245 = n29436 & ~n53244 ;
  assign n53246 = n53243 & n53245 ;
  assign n53247 = n2670 & ~n13220 ;
  assign n53248 = ~n10446 & n53247 ;
  assign n53249 = n32664 ^ n24855 ^ n16257 ;
  assign n53251 = ( n7956 & n10056 ) | ( n7956 & ~n12258 ) | ( n10056 & ~n12258 ) ;
  assign n53250 = ~n13807 & n24799 ;
  assign n53252 = n53251 ^ n53250 ^ 1'b0 ;
  assign n53253 = n53252 ^ n4495 ^ 1'b0 ;
  assign n53254 = n33657 ^ n20369 ^ 1'b0 ;
  assign n53255 = n17170 & ~n23212 ;
  assign n53256 = ( n12494 & n17982 ) | ( n12494 & n25834 ) | ( n17982 & n25834 ) ;
  assign n53257 = ( n27803 & n33497 ) | ( n27803 & ~n39584 ) | ( n33497 & ~n39584 ) ;
  assign n53258 = n16483 ^ n687 ^ 1'b0 ;
  assign n53259 = ~n53257 & n53258 ;
  assign n53260 = ~n4722 & n29560 ;
  assign n53261 = ~n20538 & n53260 ;
  assign n53262 = n42002 ^ n29044 ^ 1'b0 ;
  assign n53263 = n53261 | n53262 ;
  assign n53264 = n11329 ^ n7417 ^ 1'b0 ;
  assign n53265 = n31941 | n53264 ;
  assign n53266 = n31850 | n53265 ;
  assign n53267 = n52843 | n53266 ;
  assign n53268 = n15670 | n16279 ;
  assign n53269 = ~n26033 & n53268 ;
  assign n53270 = n45838 ^ n37314 ^ 1'b0 ;
  assign n53271 = n42190 ^ n30767 ^ n9075 ;
  assign n53272 = n29171 ^ n28472 ^ n22061 ;
  assign n53273 = ( ~n586 & n1524 ) | ( ~n586 & n12472 ) | ( n1524 & n12472 ) ;
  assign n53274 = ( ~n4580 & n18586 ) | ( ~n4580 & n19189 ) | ( n18586 & n19189 ) ;
  assign n53275 = n14351 ^ n3662 ^ 1'b0 ;
  assign n53276 = n21635 & ~n53275 ;
  assign n53277 = n24707 & n53276 ;
  assign n53278 = n21104 | n52113 ;
  assign n53279 = n4087 & ~n49823 ;
  assign n53280 = n7351 & n53279 ;
  assign n53281 = n51792 ^ n45538 ^ 1'b0 ;
  assign n53282 = n9530 | n53281 ;
  assign n53284 = ( ~n517 & n6092 ) | ( ~n517 & n41173 ) | ( n6092 & n41173 ) ;
  assign n53283 = n26939 | n29461 ;
  assign n53285 = n53284 ^ n53283 ^ 1'b0 ;
  assign n53286 = ( ~n2911 & n9281 ) | ( ~n2911 & n14917 ) | ( n9281 & n14917 ) ;
  assign n53287 = n53286 ^ n45874 ^ n3726 ;
  assign n53288 = n19205 & n53287 ;
  assign n53289 = n39667 ^ n37565 ^ n1131 ;
  assign n53291 = n19316 ^ n2527 ^ 1'b0 ;
  assign n53290 = ( n1626 & n11578 ) | ( n1626 & ~n14840 ) | ( n11578 & ~n14840 ) ;
  assign n53292 = n53291 ^ n53290 ^ n39176 ;
  assign n53293 = n20733 | n51418 ;
  assign n53294 = n53293 ^ n35691 ^ n31483 ;
  assign n53295 = n3615 ^ x189 ^ 1'b0 ;
  assign n53296 = ( ~n13599 & n18575 ) | ( ~n13599 & n53295 ) | ( n18575 & n53295 ) ;
  assign n53297 = n16278 & n47827 ;
  assign n53298 = ( n19945 & n35937 ) | ( n19945 & ~n52058 ) | ( n35937 & ~n52058 ) ;
  assign n53299 = n53297 & n53298 ;
  assign n53300 = n31647 | n44293 ;
  assign n53301 = n9819 | n53300 ;
  assign n53302 = n27898 ^ n13900 ^ 1'b0 ;
  assign n53303 = n53301 & n53302 ;
  assign n53304 = ~n8964 & n53303 ;
  assign n53305 = n15211 ^ n7598 ^ 1'b0 ;
  assign n53306 = n25721 & ~n53305 ;
  assign n53307 = n34745 ^ n30127 ^ 1'b0 ;
  assign n53308 = n53306 & ~n53307 ;
  assign n53309 = ( n3465 & n6951 ) | ( n3465 & ~n13174 ) | ( n6951 & ~n13174 ) ;
  assign n53310 = n4302 & ~n53309 ;
  assign n53311 = n53310 ^ n13157 ^ 1'b0 ;
  assign n53314 = n9907 & ~n20087 ;
  assign n53315 = n53314 ^ n12536 ^ 1'b0 ;
  assign n53312 = ~n3785 & n46144 ;
  assign n53313 = ~n11390 & n53312 ;
  assign n53316 = n53315 ^ n53313 ^ 1'b0 ;
  assign n53317 = ( n1967 & n20928 ) | ( n1967 & n22068 ) | ( n20928 & n22068 ) ;
  assign n53318 = n53317 ^ n49277 ^ 1'b0 ;
  assign n53319 = n3662 | n53318 ;
  assign n53320 = ( n9496 & n19569 ) | ( n9496 & ~n53319 ) | ( n19569 & ~n53319 ) ;
  assign n53321 = ~n3945 & n42071 ;
  assign n53322 = n53321 ^ n46535 ^ n43882 ;
  assign n53323 = n28916 ^ n11408 ^ 1'b0 ;
  assign n53324 = ( n7077 & n34751 ) | ( n7077 & n52061 ) | ( n34751 & n52061 ) ;
  assign n53325 = n27556 ^ n18996 ^ 1'b0 ;
  assign n53326 = n7022 ^ n1370 ^ 1'b0 ;
  assign n53327 = n32914 ^ n15609 ^ 1'b0 ;
  assign n53328 = ~n10905 & n29829 ;
  assign n53329 = n14408 | n27316 ;
  assign n53330 = n53329 ^ n5653 ^ 1'b0 ;
  assign n53331 = ( n5845 & ~n10458 ) | ( n5845 & n53330 ) | ( ~n10458 & n53330 ) ;
  assign n53332 = n53331 ^ n3748 ^ 1'b0 ;
  assign n53333 = ~n53328 & n53332 ;
  assign n53334 = n2173 & n42892 ;
  assign n53335 = n53334 ^ n44862 ^ 1'b0 ;
  assign n53336 = n5265 & ~n23186 ;
  assign n53337 = ~n42719 & n53336 ;
  assign n53338 = ( n16046 & n35005 ) | ( n16046 & ~n42079 ) | ( n35005 & ~n42079 ) ;
  assign n53339 = ~n20928 & n53338 ;
  assign n53340 = n48053 & n53339 ;
  assign n53341 = n2937 & ~n9862 ;
  assign n53342 = n21797 & n53341 ;
  assign n53343 = n53342 ^ n50335 ^ n12719 ;
  assign n53344 = ( n20854 & ~n22055 ) | ( n20854 & n53343 ) | ( ~n22055 & n53343 ) ;
  assign n53345 = ~n7173 & n50771 ;
  assign n53346 = n53345 ^ n20357 ^ 1'b0 ;
  assign n53347 = ( n4759 & n19178 ) | ( n4759 & ~n24085 ) | ( n19178 & ~n24085 ) ;
  assign n53348 = n53347 ^ n2690 ^ n2340 ;
  assign n53349 = n43733 ^ n13453 ^ 1'b0 ;
  assign n53350 = n53348 | n53349 ;
  assign n53351 = ( n51994 & n53346 ) | ( n51994 & n53350 ) | ( n53346 & n53350 ) ;
  assign n53352 = n27599 ^ n25618 ^ 1'b0 ;
  assign n53353 = n53352 ^ n49083 ^ n2360 ;
  assign n53354 = ( n14542 & ~n26684 ) | ( n14542 & n32512 ) | ( ~n26684 & n32512 ) ;
  assign n53355 = n29666 ^ n21271 ^ 1'b0 ;
  assign n53356 = ( n15914 & n22042 ) | ( n15914 & n53355 ) | ( n22042 & n53355 ) ;
  assign n53359 = n28513 ^ n23099 ^ n21287 ;
  assign n53357 = n3906 & n36279 ;
  assign n53358 = n53357 ^ n10208 ^ 1'b0 ;
  assign n53360 = n53359 ^ n53358 ^ 1'b0 ;
  assign n53361 = n37647 ^ n1950 ^ n314 ;
  assign n53362 = n286 | n3111 ;
  assign n53363 = ~n34061 & n53362 ;
  assign n53364 = n53361 & n53363 ;
  assign n53368 = n30483 ^ n12172 ^ 1'b0 ;
  assign n53369 = n49297 & n53368 ;
  assign n53365 = n16957 ^ n7230 ^ 1'b0 ;
  assign n53366 = n15294 | n53365 ;
  assign n53367 = n4070 & ~n53366 ;
  assign n53370 = n53369 ^ n53367 ^ 1'b0 ;
  assign n53371 = n32184 & ~n47447 ;
  assign n53372 = n53371 ^ n35039 ^ 1'b0 ;
  assign n53373 = n1589 | n4743 ;
  assign n53374 = n15551 ^ n15190 ^ 1'b0 ;
  assign n53377 = ~n2865 & n37319 ;
  assign n53375 = n5363 & n32528 ;
  assign n53376 = n53375 ^ n3715 ^ 1'b0 ;
  assign n53378 = n53377 ^ n53376 ^ n20445 ;
  assign n53379 = n24473 | n25997 ;
  assign n53380 = n53379 ^ n37555 ^ n23577 ;
  assign n53381 = n46176 ^ n38338 ^ n35709 ;
  assign n53382 = n24829 ^ n6664 ^ n4493 ;
  assign n53383 = n5997 & n53284 ;
  assign n53384 = n880 & n53383 ;
  assign n53385 = n42713 ^ n36700 ^ 1'b0 ;
  assign n53386 = ~n51579 & n53385 ;
  assign n53387 = n49134 | n52184 ;
  assign n53388 = n34154 | n53387 ;
  assign n53389 = n11314 & ~n38812 ;
  assign n53390 = ~n31846 & n34451 ;
  assign n53391 = n5477 & n53390 ;
  assign n53392 = n13253 & n18119 ;
  assign n53393 = n53391 & n53392 ;
  assign n53394 = n19751 ^ n12303 ^ n6554 ;
  assign n53395 = n14284 ^ n7837 ^ 1'b0 ;
  assign n53396 = ~n4440 & n53395 ;
  assign n53397 = ( n665 & n15931 ) | ( n665 & ~n53396 ) | ( n15931 & ~n53396 ) ;
  assign n53398 = n16002 ^ n10578 ^ n2371 ;
  assign n53399 = ( n1832 & n53146 ) | ( n1832 & ~n53398 ) | ( n53146 & ~n53398 ) ;
  assign n53400 = n53399 ^ n30512 ^ 1'b0 ;
  assign n53401 = n47765 ^ n30763 ^ n20323 ;
  assign n53402 = n53401 ^ n2398 ^ 1'b0 ;
  assign n53403 = n22506 ^ n18052 ^ n7087 ;
  assign n53404 = n24533 | n37256 ;
  assign n53405 = n29060 & ~n37253 ;
  assign n53406 = n53405 ^ n17632 ^ 1'b0 ;
  assign n53407 = n8529 | n23918 ;
  assign n53408 = ~n4068 & n48553 ;
  assign n53409 = ~n38511 & n46095 ;
  assign n53410 = n35091 & ~n53409 ;
  assign n53411 = ~n1455 & n28919 ;
  assign n53412 = ( ~n1418 & n13261 ) | ( ~n1418 & n53411 ) | ( n13261 & n53411 ) ;
  assign n53413 = n53412 ^ n39751 ^ n1783 ;
  assign n53414 = n53413 ^ n22228 ^ n21132 ;
  assign n53415 = n44817 ^ n6612 ^ 1'b0 ;
  assign n53416 = ~n8530 & n19247 ;
  assign n53417 = ~n1308 & n53416 ;
  assign n53418 = ( n4052 & n10163 ) | ( n4052 & ~n53417 ) | ( n10163 & ~n53417 ) ;
  assign n53419 = ~n13078 & n47325 ;
  assign n53420 = ~n53418 & n53419 ;
  assign n53421 = ( n4079 & n16534 ) | ( n4079 & ~n18087 ) | ( n16534 & ~n18087 ) ;
  assign n53422 = n37032 ^ n27175 ^ n21674 ;
  assign n53423 = n1148 & n50052 ;
  assign n53424 = n1431 & n4404 ;
  assign n53425 = n53424 ^ n4020 ^ 1'b0 ;
  assign n53426 = n12247 ^ n9611 ^ 1'b0 ;
  assign n53427 = n21553 & n53426 ;
  assign n53428 = n28490 ^ n11158 ^ n4872 ;
  assign n53429 = n9720 ^ n7475 ^ n6747 ;
  assign n53430 = ( n11974 & n27128 ) | ( n11974 & n40011 ) | ( n27128 & n40011 ) ;
  assign n53431 = ( n38946 & ~n53429 ) | ( n38946 & n53430 ) | ( ~n53429 & n53430 ) ;
  assign n53432 = n13639 ^ n3003 ^ 1'b0 ;
  assign n53433 = ( n701 & ~n2200 ) | ( n701 & n27018 ) | ( ~n2200 & n27018 ) ;
  assign n53434 = n53433 ^ n36431 ^ 1'b0 ;
  assign n53435 = n19137 & n53434 ;
  assign n53436 = n53435 ^ n47354 ^ n3813 ;
  assign n53437 = n6270 & ~n14134 ;
  assign n53438 = n3184 & n53437 ;
  assign n53439 = ( ~n15934 & n40264 ) | ( ~n15934 & n41360 ) | ( n40264 & n41360 ) ;
  assign n53440 = n50121 ^ n26011 ^ n6224 ;
  assign n53441 = n1319 & n53440 ;
  assign n53443 = ( n4402 & n12677 ) | ( n4402 & n18379 ) | ( n12677 & n18379 ) ;
  assign n53442 = n3783 | n14428 ;
  assign n53444 = n53443 ^ n53442 ^ n6334 ;
  assign n53445 = n3834 & ~n14427 ;
  assign n53446 = ~n3005 & n53445 ;
  assign n53447 = n33795 ^ n10334 ^ 1'b0 ;
  assign n53448 = n29196 ^ n12380 ^ 1'b0 ;
  assign n53449 = n53447 & n53448 ;
  assign n53450 = ( n22846 & n53446 ) | ( n22846 & n53449 ) | ( n53446 & n53449 ) ;
  assign n53451 = n53450 ^ n22770 ^ n4495 ;
  assign n53452 = n51990 ^ n25229 ^ n10905 ;
  assign n53453 = n27061 ^ n17451 ^ n1137 ;
  assign n53455 = ( n4046 & ~n15130 ) | ( n4046 & n37018 ) | ( ~n15130 & n37018 ) ;
  assign n53454 = n22437 ^ n14358 ^ n1910 ;
  assign n53456 = n53455 ^ n53454 ^ n27013 ;
  assign n53457 = n40608 ^ n39306 ^ n14055 ;
  assign n53458 = ~n5125 & n19369 ;
  assign n53459 = n25621 & n53458 ;
  assign n53460 = n53459 ^ n34151 ^ 1'b0 ;
  assign n53461 = n53460 ^ n15154 ^ 1'b0 ;
  assign n53462 = n21033 | n53461 ;
  assign n53463 = ~n4268 & n4486 ;
  assign n53464 = n53463 ^ n6567 ^ 1'b0 ;
  assign n53465 = n11299 | n21240 ;
  assign n53466 = n293 & ~n53465 ;
  assign n53467 = ~n21115 & n53466 ;
  assign n53468 = n10036 | n12979 ;
  assign n53469 = n53467 | n53468 ;
  assign n53470 = ( n25450 & ~n28741 ) | ( n25450 & n43051 ) | ( ~n28741 & n43051 ) ;
  assign n53471 = ( n2168 & n11379 ) | ( n2168 & ~n14036 ) | ( n11379 & ~n14036 ) ;
  assign n53472 = n48020 ^ n46165 ^ n874 ;
  assign n53473 = ~n1433 & n13903 ;
  assign n53474 = n53473 ^ n5244 ^ 1'b0 ;
  assign n53475 = n39299 | n53474 ;
  assign n53480 = n21600 & ~n30105 ;
  assign n53481 = n53480 ^ n9537 ^ 1'b0 ;
  assign n53482 = n53481 ^ n353 ^ 1'b0 ;
  assign n53476 = n9543 ^ n3326 ^ 1'b0 ;
  assign n53477 = n24620 & ~n53476 ;
  assign n53478 = n12301 & ~n53477 ;
  assign n53479 = n4227 & ~n53478 ;
  assign n53483 = n53482 ^ n53479 ^ n12552 ;
  assign n53484 = n42117 ^ n31185 ^ n16496 ;
  assign n53485 = ( n12172 & n16441 ) | ( n12172 & n53484 ) | ( n16441 & n53484 ) ;
  assign n53486 = ( x161 & ~x210 ) | ( x161 & n19391 ) | ( ~x210 & n19391 ) ;
  assign n53487 = ( n31580 & ~n34056 ) | ( n31580 & n53486 ) | ( ~n34056 & n53486 ) ;
  assign n53488 = n17611 | n41337 ;
  assign n53489 = n53487 | n53488 ;
  assign n53490 = n26824 & n31817 ;
  assign n53491 = n31299 & n53490 ;
  assign n53492 = n34389 ^ n9505 ^ 1'b0 ;
  assign n53493 = n41845 ^ n11181 ^ 1'b0 ;
  assign n53494 = ( ~n22747 & n36851 ) | ( ~n22747 & n48746 ) | ( n36851 & n48746 ) ;
  assign n53495 = n19489 ^ n17415 ^ n1647 ;
  assign n53496 = n53495 ^ n38033 ^ n26377 ;
  assign n53497 = ~n13437 & n41210 ;
  assign n53498 = ~n1530 & n53497 ;
  assign n53499 = ( n26413 & n41245 ) | ( n26413 & n53498 ) | ( n41245 & n53498 ) ;
  assign n53500 = ~n15491 & n53499 ;
  assign n53501 = n43402 ^ n10306 ^ 1'b0 ;
  assign n53502 = n53501 ^ n49223 ^ n40385 ;
  assign n53503 = n1881 & n31206 ;
  assign n53504 = n53503 ^ n22597 ^ 1'b0 ;
  assign n53505 = n53504 ^ n25573 ^ n14912 ;
  assign n53507 = ~n2881 & n27237 ;
  assign n53508 = n15835 & n53507 ;
  assign n53506 = n15888 ^ n13958 ^ n13453 ;
  assign n53509 = n53508 ^ n53506 ^ n25462 ;
  assign n53510 = n31432 | n53509 ;
  assign n53511 = n10835 & ~n16046 ;
  assign n53512 = n53511 ^ n9040 ^ 1'b0 ;
  assign n53516 = n34121 ^ n29688 ^ n15568 ;
  assign n53513 = ( n1103 & ~n23469 ) | ( n1103 & n27481 ) | ( ~n23469 & n27481 ) ;
  assign n53514 = n53513 ^ n39113 ^ 1'b0 ;
  assign n53515 = n1158 | n53514 ;
  assign n53517 = n53516 ^ n53515 ^ 1'b0 ;
  assign n53518 = n41527 ^ n35250 ^ n10651 ;
  assign n53519 = n20479 & n53518 ;
  assign n53520 = n4659 & n53519 ;
  assign n53522 = n23724 & n26032 ;
  assign n53523 = n53522 ^ n5424 ^ 1'b0 ;
  assign n53521 = n23471 & n34078 ;
  assign n53524 = n53523 ^ n53521 ^ 1'b0 ;
  assign n53525 = n53524 ^ n15548 ^ n7900 ;
  assign n53526 = n44988 ^ n33288 ^ n28692 ;
  assign n53527 = n48097 ^ n40744 ^ n23135 ;
  assign n53528 = n46051 ^ n15918 ^ n8926 ;
  assign n53529 = n53528 ^ n30121 ^ n10592 ;
  assign n53530 = n24051 | n39794 ;
  assign n53531 = n4063 & n47695 ;
  assign n53532 = n53531 ^ n49929 ^ 1'b0 ;
  assign n53533 = n35377 ^ n4580 ^ 1'b0 ;
  assign n53535 = n8566 ^ n6774 ^ 1'b0 ;
  assign n53534 = n42832 ^ n19780 ^ n6113 ;
  assign n53536 = n53535 ^ n53534 ^ n31889 ;
  assign n53537 = ( n36970 & n42852 ) | ( n36970 & n53536 ) | ( n42852 & n53536 ) ;
  assign n53538 = n17929 & ~n42637 ;
  assign n53539 = n53538 ^ n27275 ^ 1'b0 ;
  assign n53540 = ( ~n21957 & n51663 ) | ( ~n21957 & n53539 ) | ( n51663 & n53539 ) ;
  assign n53541 = n450 & ~n53540 ;
  assign n53542 = n25523 ^ n4237 ^ 1'b0 ;
  assign n53543 = n3613 & ~n53542 ;
  assign n53544 = n53543 ^ n12120 ^ 1'b0 ;
  assign n53545 = ~n21137 & n33179 ;
  assign n53546 = ( ~n1010 & n8382 ) | ( ~n1010 & n10500 ) | ( n8382 & n10500 ) ;
  assign n53547 = ( n32625 & n39011 ) | ( n32625 & ~n53546 ) | ( n39011 & ~n53546 ) ;
  assign n53548 = n11431 | n38406 ;
  assign n53549 = n53548 ^ n48654 ^ 1'b0 ;
  assign n53550 = n38660 ^ n25107 ^ 1'b0 ;
  assign n53551 = n47278 ^ n34695 ^ 1'b0 ;
  assign n53552 = n21837 ^ n17054 ^ n12017 ;
  assign n53553 = n13209 | n53552 ;
  assign n53554 = n27356 | n53553 ;
  assign n53555 = ~n18624 & n19009 ;
  assign n53556 = n53555 ^ n3462 ^ 1'b0 ;
  assign n53557 = n53556 ^ n40012 ^ n287 ;
  assign n53558 = n35445 ^ n25808 ^ n22873 ;
  assign n53559 = n53558 ^ n17327 ^ 1'b0 ;
  assign n53560 = n13384 ^ n5638 ^ 1'b0 ;
  assign n53561 = n20449 & n53560 ;
  assign n53562 = n53561 ^ n26720 ^ 1'b0 ;
  assign n53563 = n39204 ^ n6769 ^ 1'b0 ;
  assign n53564 = n15814 ^ n13934 ^ 1'b0 ;
  assign n53565 = n20813 & ~n53564 ;
  assign n53566 = n53565 ^ n26891 ^ 1'b0 ;
  assign n53567 = n38076 & n53566 ;
  assign n53568 = n53567 ^ n11798 ^ 1'b0 ;
  assign n53569 = n14449 & n20126 ;
  assign n53570 = ~x65 & n53569 ;
  assign n53571 = n2935 & n53570 ;
  assign n53572 = n53571 ^ n25700 ^ n14369 ;
  assign n53573 = n53572 ^ n39780 ^ n19229 ;
  assign n53574 = ~n7772 & n19321 ;
  assign n53575 = ~n52117 & n53574 ;
  assign n53578 = ( ~n14542 & n19189 ) | ( ~n14542 & n19859 ) | ( n19189 & n19859 ) ;
  assign n53579 = n53578 ^ n35849 ^ n7005 ;
  assign n53576 = n11795 & ~n22169 ;
  assign n53577 = n11973 & ~n53576 ;
  assign n53580 = n53579 ^ n53577 ^ 1'b0 ;
  assign n53581 = ( n2673 & n7973 ) | ( n2673 & ~n11390 ) | ( n7973 & ~n11390 ) ;
  assign n53582 = n53581 ^ n17667 ^ 1'b0 ;
  assign n53583 = x36 | n5780 ;
  assign n53584 = n14325 & ~n53583 ;
  assign n53585 = n23688 | n32498 ;
  assign n53586 = n48152 ^ n20014 ^ n14472 ;
  assign n53587 = n24415 | n25324 ;
  assign n53588 = n36312 ^ n12352 ^ n12041 ;
  assign n53591 = n36976 ^ n21855 ^ n14797 ;
  assign n53589 = n23218 ^ n14542 ^ n12479 ;
  assign n53590 = n53589 ^ n47018 ^ n2022 ;
  assign n53592 = n53591 ^ n53590 ^ 1'b0 ;
  assign n53593 = n53592 ^ n43469 ^ n39750 ;
  assign n53594 = n18121 ^ n17369 ^ 1'b0 ;
  assign n53595 = n53594 ^ n5335 ^ n5056 ;
  assign n53596 = ~n17935 & n52969 ;
  assign n53597 = ~n43457 & n53596 ;
  assign n53598 = x91 & n4305 ;
  assign n53599 = n53598 ^ n15535 ^ 1'b0 ;
  assign n53600 = n25480 & n48188 ;
  assign n53601 = n53600 ^ n34098 ^ 1'b0 ;
  assign n53602 = ( ~n10969 & n40734 ) | ( ~n10969 & n53601 ) | ( n40734 & n53601 ) ;
  assign n53603 = n39564 ^ n17178 ^ 1'b0 ;
  assign n53604 = ~n2178 & n53603 ;
  assign n53605 = n48635 & n53604 ;
  assign n53606 = ( ~n28395 & n52461 ) | ( ~n28395 & n53605 ) | ( n52461 & n53605 ) ;
  assign n53609 = n34266 ^ n22472 ^ n2183 ;
  assign n53607 = ( n5542 & n26636 ) | ( n5542 & n33469 ) | ( n26636 & n33469 ) ;
  assign n53608 = ( n41356 & n47572 ) | ( n41356 & n53607 ) | ( n47572 & n53607 ) ;
  assign n53610 = n53609 ^ n53608 ^ 1'b0 ;
  assign n53611 = ( n15998 & n31750 ) | ( n15998 & n46368 ) | ( n31750 & n46368 ) ;
  assign n53613 = n7834 ^ n5927 ^ 1'b0 ;
  assign n53612 = n36088 ^ n12811 ^ n12630 ;
  assign n53614 = n53613 ^ n53612 ^ n20354 ;
  assign n53615 = n32211 ^ n9840 ^ n4117 ;
  assign n53616 = n53615 ^ n31835 ^ n19097 ;
  assign n53617 = n28174 ^ n13342 ^ n3732 ;
  assign n53618 = n53617 ^ n14504 ^ n9648 ;
  assign n53619 = ( n26366 & ~n53616 ) | ( n26366 & n53618 ) | ( ~n53616 & n53618 ) ;
  assign n53620 = n13117 ^ n9125 ^ n3075 ;
  assign n53621 = n53620 ^ n53493 ^ 1'b0 ;
  assign n53622 = n8544 & ~n53621 ;
  assign n53623 = ~n2026 & n21287 ;
  assign n53624 = ~n22382 & n53623 ;
  assign n53625 = ( n3381 & n17942 ) | ( n3381 & n37238 ) | ( n17942 & n37238 ) ;
  assign n53626 = ~n24972 & n25725 ;
  assign n53627 = ( ~n7407 & n38992 ) | ( ~n7407 & n53626 ) | ( n38992 & n53626 ) ;
  assign n53628 = n53627 ^ n16058 ^ 1'b0 ;
  assign n53629 = ~n53625 & n53628 ;
  assign n53630 = n20060 ^ n7520 ^ 1'b0 ;
  assign n53631 = n53629 & n53630 ;
  assign n53635 = ( n7224 & ~n8757 ) | ( n7224 & n47127 ) | ( ~n8757 & n47127 ) ;
  assign n53636 = n53635 ^ n11887 ^ n1339 ;
  assign n53633 = n52055 ^ n6999 ^ n6138 ;
  assign n53634 = ~n22357 & n53633 ;
  assign n53637 = n53636 ^ n53634 ^ 1'b0 ;
  assign n53632 = ~n21623 & n49781 ;
  assign n53638 = n53637 ^ n53632 ^ 1'b0 ;
  assign n53639 = n19495 & n19954 ;
  assign n53640 = n53639 ^ n26676 ^ n16501 ;
  assign n53641 = n24955 & n51921 ;
  assign n53642 = n14682 | n30363 ;
  assign n53643 = n27231 ^ n6341 ^ n5269 ;
  assign n53644 = n53643 ^ n6074 ^ 1'b0 ;
  assign n53645 = n11742 | n14987 ;
  assign n53646 = n21231 & ~n53645 ;
  assign n53647 = ( n2319 & n15478 ) | ( n2319 & n53646 ) | ( n15478 & n53646 ) ;
  assign n53648 = ( n18712 & n24465 ) | ( n18712 & n33128 ) | ( n24465 & n33128 ) ;
  assign n53649 = n27046 ^ n22892 ^ n7118 ;
  assign n53650 = n39616 ^ n21075 ^ 1'b0 ;
  assign n53654 = ~n2266 & n4781 ;
  assign n53655 = ~n1896 & n53654 ;
  assign n53651 = ( ~n7650 & n13340 ) | ( ~n7650 & n17914 ) | ( n13340 & n17914 ) ;
  assign n53652 = n53651 ^ n4779 ^ 1'b0 ;
  assign n53653 = n27132 & ~n53652 ;
  assign n53656 = n53655 ^ n53653 ^ 1'b0 ;
  assign n53657 = n12910 ^ n9277 ^ n5609 ;
  assign n53658 = n3773 | n53657 ;
  assign n53659 = n53658 ^ n25512 ^ 1'b0 ;
  assign n53661 = n52835 ^ n43297 ^ n9810 ;
  assign n53660 = n26472 ^ n3662 ^ n2131 ;
  assign n53662 = n53661 ^ n53660 ^ 1'b0 ;
  assign n53663 = n9622 ^ n7466 ^ n6307 ;
  assign n53664 = n40246 ^ n20690 ^ 1'b0 ;
  assign n53665 = ( ~n5270 & n8010 ) | ( ~n5270 & n22988 ) | ( n8010 & n22988 ) ;
  assign n53666 = n43065 ^ n21262 ^ 1'b0 ;
  assign n53667 = n3228 & n32741 ;
  assign n53668 = ~n53666 & n53667 ;
  assign n53669 = n997 & n53668 ;
  assign n53670 = n28464 ^ n25887 ^ n4290 ;
  assign n53671 = n9124 & n53670 ;
  assign n53673 = n50368 ^ n21209 ^ n20433 ;
  assign n53672 = ~n11114 & n11946 ;
  assign n53674 = n53673 ^ n53672 ^ 1'b0 ;
  assign n53675 = n974 | n49049 ;
  assign n53676 = n48065 | n53675 ;
  assign n53678 = ( n12668 & n19398 ) | ( n12668 & n20378 ) | ( n19398 & n20378 ) ;
  assign n53679 = n29370 ^ n11923 ^ n1083 ;
  assign n53680 = n53678 | n53679 ;
  assign n53677 = n5907 & n28842 ;
  assign n53681 = n53680 ^ n53677 ^ n29904 ;
  assign n53682 = n23430 ^ n13623 ^ n1980 ;
  assign n53683 = n48651 ^ n27831 ^ 1'b0 ;
  assign n53684 = ( n725 & n5930 ) | ( n725 & ~n38265 ) | ( n5930 & ~n38265 ) ;
  assign n53685 = n20152 ^ n2927 ^ 1'b0 ;
  assign n53686 = ~n2959 & n20304 ;
  assign n53687 = ( n15973 & n17258 ) | ( n15973 & n53686 ) | ( n17258 & n53686 ) ;
  assign n53688 = ( n33748 & n53685 ) | ( n33748 & ~n53687 ) | ( n53685 & ~n53687 ) ;
  assign n53689 = n52170 & n53433 ;
  assign n53690 = n6481 & ~n38951 ;
  assign n53691 = ~n37540 & n53690 ;
  assign n53692 = n24342 | n26262 ;
  assign n53693 = n53692 ^ n21572 ^ 1'b0 ;
  assign n53694 = ( n10261 & n15824 ) | ( n10261 & n23157 ) | ( n15824 & n23157 ) ;
  assign n53695 = ~n43472 & n53694 ;
  assign n53696 = n47103 ^ n45039 ^ 1'b0 ;
  assign n53697 = ( n11685 & n14493 ) | ( n11685 & ~n37979 ) | ( n14493 & ~n37979 ) ;
  assign n53698 = n34716 ^ n21540 ^ n11095 ;
  assign n53699 = ~n2472 & n38752 ;
  assign n53700 = ~n19264 & n53699 ;
  assign n53701 = n53700 ^ n37771 ^ n10539 ;
  assign n53702 = n44030 ^ n39305 ^ n8992 ;
  assign n53703 = n53702 ^ n1548 ^ 1'b0 ;
  assign n53704 = ( n7497 & ~n42537 ) | ( n7497 & n53703 ) | ( ~n42537 & n53703 ) ;
  assign n53705 = ~n6973 & n11617 ;
  assign n53706 = n53705 ^ n47979 ^ 1'b0 ;
  assign n53707 = n31639 ^ n569 ^ 1'b0 ;
  assign n53708 = n27944 & n37222 ;
  assign n53709 = n47579 ^ n39990 ^ n26498 ;
  assign n53710 = n16964 | n48937 ;
  assign n53711 = n40257 & ~n53710 ;
  assign n53712 = n53711 ^ n19798 ^ 1'b0 ;
  assign n53713 = n17451 ^ n7683 ^ x170 ;
  assign n53714 = n53713 ^ n45273 ^ n4967 ;
  assign n53715 = n32856 ^ n27437 ^ n23726 ;
  assign n53716 = n38651 ^ n11490 ^ 1'b0 ;
  assign n53717 = n19923 ^ n12653 ^ 1'b0 ;
  assign n53718 = n39385 & n53717 ;
  assign n53719 = n53718 ^ n40542 ^ 1'b0 ;
  assign n53720 = n1012 & n53719 ;
  assign n53721 = n35616 ^ n3965 ^ 1'b0 ;
  assign n53722 = ~n6236 & n53721 ;
  assign n53723 = n42687 ^ n33802 ^ 1'b0 ;
  assign n53724 = n13158 ^ n2950 ^ 1'b0 ;
  assign n53725 = ~n8998 & n53724 ;
  assign n53726 = ( ~n12277 & n23209 ) | ( ~n12277 & n53725 ) | ( n23209 & n53725 ) ;
  assign n53727 = n53723 & ~n53726 ;
  assign n53728 = n53727 ^ n36961 ^ n17695 ;
  assign n53729 = n52117 ^ n35886 ^ 1'b0 ;
  assign n53730 = n13949 | n53729 ;
  assign n53731 = ( n3798 & n11830 ) | ( n3798 & ~n53730 ) | ( n11830 & ~n53730 ) ;
  assign n53732 = ( n4384 & ~n28510 ) | ( n4384 & n30248 ) | ( ~n28510 & n30248 ) ;
  assign n53733 = ( n3468 & n32773 ) | ( n3468 & n34691 ) | ( n32773 & n34691 ) ;
  assign n53734 = ( n5900 & n19527 ) | ( n5900 & ~n53733 ) | ( n19527 & ~n53733 ) ;
  assign n53735 = n2766 | n27035 ;
  assign n53736 = ~n12121 & n12843 ;
  assign n53737 = n53736 ^ n15934 ^ 1'b0 ;
  assign n53738 = ( n29928 & ~n52851 ) | ( n29928 & n53737 ) | ( ~n52851 & n53737 ) ;
  assign n53739 = n12290 | n40249 ;
  assign n53740 = n14934 & ~n53739 ;
  assign n53741 = n928 & ~n32856 ;
  assign n53742 = n53740 & n53741 ;
  assign n53743 = n25229 & ~n38271 ;
  assign n53744 = n53743 ^ n2873 ^ 1'b0 ;
  assign n53745 = n53744 ^ n32108 ^ n14960 ;
  assign n53746 = ~n32670 & n53745 ;
  assign n53747 = n53746 ^ n12497 ^ 1'b0 ;
  assign n53748 = ~n33296 & n40115 ;
  assign n53749 = n53748 ^ n43987 ^ 1'b0 ;
  assign n53750 = n35348 ^ n4499 ^ 1'b0 ;
  assign n53751 = n18455 | n53750 ;
  assign n53752 = n29143 ^ n25838 ^ 1'b0 ;
  assign n53753 = n26540 ^ n2824 ^ 1'b0 ;
  assign n53754 = n20959 | n40417 ;
  assign n53755 = n4442 & ~n53754 ;
  assign n53756 = n53755 ^ n48537 ^ n21264 ;
  assign n53757 = ( ~n9691 & n22807 ) | ( ~n9691 & n53756 ) | ( n22807 & n53756 ) ;
  assign n53758 = n24151 ^ n17998 ^ n4203 ;
  assign n53759 = n51903 ^ n45540 ^ n31493 ;
  assign n53760 = n51794 ^ n37093 ^ n1319 ;
  assign n53761 = n7630 ^ n2261 ^ 1'b0 ;
  assign n53762 = n3649 & n53761 ;
  assign n53763 = ( ~n38247 & n53760 ) | ( ~n38247 & n53762 ) | ( n53760 & n53762 ) ;
  assign n53764 = n9291 & ~n20635 ;
  assign n53765 = ~n1288 & n53764 ;
  assign n53766 = n36196 ^ n2365 ^ 1'b0 ;
  assign n53767 = ~n8793 & n53766 ;
  assign n53769 = ( n1564 & n4952 ) | ( n1564 & ~n15813 ) | ( n4952 & ~n15813 ) ;
  assign n53770 = n33757 ^ n24751 ^ n23244 ;
  assign n53771 = ( n14880 & n53769 ) | ( n14880 & ~n53770 ) | ( n53769 & ~n53770 ) ;
  assign n53768 = n6808 & ~n31517 ;
  assign n53772 = n53771 ^ n53768 ^ 1'b0 ;
  assign n53774 = n22362 ^ n19104 ^ n828 ;
  assign n53773 = ( n8336 & n21281 ) | ( n8336 & ~n35467 ) | ( n21281 & ~n35467 ) ;
  assign n53775 = n53774 ^ n53773 ^ n20273 ;
  assign n53776 = n53775 ^ n45084 ^ 1'b0 ;
  assign n53777 = n23586 ^ n15991 ^ 1'b0 ;
  assign n53778 = ~n53776 & n53777 ;
  assign n53779 = n34107 ^ n23666 ^ 1'b0 ;
  assign n53780 = ( n4629 & n51453 ) | ( n4629 & n53779 ) | ( n51453 & n53779 ) ;
  assign n53782 = ~n26571 & n26768 ;
  assign n53783 = n29176 | n53782 ;
  assign n53781 = n7450 & ~n8034 ;
  assign n53784 = n53783 ^ n53781 ^ 1'b0 ;
  assign n53785 = n53784 ^ n46466 ^ n26638 ;
  assign n53786 = n45152 ^ n2301 ^ 1'b0 ;
  assign n53787 = ( n11313 & ~n21099 ) | ( n11313 & n53786 ) | ( ~n21099 & n53786 ) ;
  assign n53788 = ( n30933 & ~n36953 ) | ( n30933 & n53787 ) | ( ~n36953 & n53787 ) ;
  assign n53789 = x85 & n4009 ;
  assign n53790 = n53789 ^ n6659 ^ 1'b0 ;
  assign n53791 = ~n3224 & n53790 ;
  assign n53792 = ( n848 & n6444 ) | ( n848 & n38410 ) | ( n6444 & n38410 ) ;
  assign n53793 = ~n11854 & n53792 ;
  assign n53794 = n53793 ^ n8218 ^ n394 ;
  assign n53795 = ( n5562 & ~n16473 ) | ( n5562 & n40897 ) | ( ~n16473 & n40897 ) ;
  assign n53796 = ( n13413 & n28741 ) | ( n13413 & ~n53795 ) | ( n28741 & ~n53795 ) ;
  assign n53797 = ( n4109 & n19227 ) | ( n4109 & n19566 ) | ( n19227 & n19566 ) ;
  assign n53798 = n53797 ^ n40810 ^ 1'b0 ;
  assign n53799 = n6670 | n53798 ;
  assign n53800 = n28246 ^ n11971 ^ 1'b0 ;
  assign n53801 = n28477 & n53800 ;
  assign n53802 = n13165 ^ n12456 ^ n3221 ;
  assign n53803 = n905 & ~n13165 ;
  assign n53804 = ( n6037 & ~n21733 ) | ( n6037 & n38532 ) | ( ~n21733 & n38532 ) ;
  assign n53805 = n53804 ^ n23767 ^ n3323 ;
  assign n53806 = ( n4087 & n24950 ) | ( n4087 & ~n53805 ) | ( n24950 & ~n53805 ) ;
  assign n53807 = ( n12472 & ~n24602 ) | ( n12472 & n53806 ) | ( ~n24602 & n53806 ) ;
  assign n53808 = n44167 ^ n44029 ^ n25411 ;
  assign n53809 = ( ~n20509 & n32626 ) | ( ~n20509 & n41990 ) | ( n32626 & n41990 ) ;
  assign n53810 = n47002 & n48929 ;
  assign n53811 = n43994 & n53810 ;
  assign n53812 = n13741 & ~n20497 ;
  assign n53813 = n53812 ^ n9325 ^ 1'b0 ;
  assign n53814 = n1610 & n21693 ;
  assign n53815 = n53814 ^ n31357 ^ 1'b0 ;
  assign n53816 = n29066 ^ n14074 ^ n10357 ;
  assign n53817 = n53816 ^ n17774 ^ 1'b0 ;
  assign n53818 = n28330 & n53817 ;
  assign n53819 = n41354 ^ n4989 ^ 1'b0 ;
  assign n53820 = ~n19715 & n53819 ;
  assign n53821 = ~n26975 & n53820 ;
  assign n53822 = n7224 | n11793 ;
  assign n53823 = n11332 ^ n6527 ^ n1388 ;
  assign n53824 = n7425 | n40363 ;
  assign n53825 = n53823 & ~n53824 ;
  assign n53826 = n53825 ^ n12499 ^ n8473 ;
  assign n53827 = n53822 | n53826 ;
  assign n53828 = n6515 & ~n36148 ;
  assign n53829 = n53828 ^ n16410 ^ 1'b0 ;
  assign n53830 = n53829 ^ n39007 ^ 1'b0 ;
  assign n53832 = ( x57 & n1550 ) | ( x57 & n27137 ) | ( n1550 & n27137 ) ;
  assign n53833 = n53832 ^ n37259 ^ n4474 ;
  assign n53831 = n33472 ^ n1823 ^ 1'b0 ;
  assign n53834 = n53833 ^ n53831 ^ 1'b0 ;
  assign n53835 = ~n16625 & n37829 ;
  assign n53836 = n3208 | n5288 ;
  assign n53837 = n53836 ^ n27844 ^ 1'b0 ;
  assign n53838 = n53837 ^ n41496 ^ n13702 ;
  assign n53839 = ( ~n7627 & n25520 ) | ( ~n7627 & n53838 ) | ( n25520 & n53838 ) ;
  assign n53840 = n52802 ^ n44127 ^ n42443 ;
  assign y0 = x8 ;
  assign y1 = x11 ;
  assign y2 = x19 ;
  assign y3 = x28 ;
  assign y4 = x30 ;
  assign y5 = x33 ;
  assign y6 = x37 ;
  assign y7 = x41 ;
  assign y8 = x45 ;
  assign y9 = x50 ;
  assign y10 = x53 ;
  assign y11 = x56 ;
  assign y12 = x60 ;
  assign y13 = x69 ;
  assign y14 = x74 ;
  assign y15 = x77 ;
  assign y16 = x82 ;
  assign y17 = x92 ;
  assign y18 = x95 ;
  assign y19 = x97 ;
  assign y20 = x115 ;
  assign y21 = x116 ;
  assign y22 = x129 ;
  assign y23 = x136 ;
  assign y24 = x143 ;
  assign y25 = x147 ;
  assign y26 = x151 ;
  assign y27 = x153 ;
  assign y28 = x157 ;
  assign y29 = x160 ;
  assign y30 = x163 ;
  assign y31 = x174 ;
  assign y32 = x176 ;
  assign y33 = x189 ;
  assign y34 = x192 ;
  assign y35 = x197 ;
  assign y36 = x198 ;
  assign y37 = x205 ;
  assign y38 = x212 ;
  assign y39 = x221 ;
  assign y40 = x227 ;
  assign y41 = x235 ;
  assign y42 = x237 ;
  assign y43 = x240 ;
  assign y44 = x242 ;
  assign y45 = x250 ;
  assign y46 = x252 ;
  assign y47 = n256 ;
  assign y48 = ~n257 ;
  assign y49 = n258 ;
  assign y50 = n260 ;
  assign y51 = ~1'b0 ;
  assign y52 = n261 ;
  assign y53 = n262 ;
  assign y54 = n264 ;
  assign y55 = n265 ;
  assign y56 = n266 ;
  assign y57 = n271 ;
  assign y58 = ~n273 ;
  assign y59 = ~n276 ;
  assign y60 = ~1'b0 ;
  assign y61 = ~1'b0 ;
  assign y62 = n282 ;
  assign y63 = ~1'b0 ;
  assign y64 = ~n285 ;
  assign y65 = ~n286 ;
  assign y66 = ~1'b0 ;
  assign y67 = ~1'b0 ;
  assign y68 = n289 ;
  assign y69 = ~n290 ;
  assign y70 = n291 ;
  assign y71 = ~n296 ;
  assign y72 = ~n297 ;
  assign y73 = n298 ;
  assign y74 = ~n300 ;
  assign y75 = n301 ;
  assign y76 = ~n257 ;
  assign y77 = ~n303 ;
  assign y78 = ~n309 ;
  assign y79 = ~1'b0 ;
  assign y80 = ~1'b0 ;
  assign y81 = n312 ;
  assign y82 = ~n314 ;
  assign y83 = ~n315 ;
  assign y84 = n318 ;
  assign y85 = n324 ;
  assign y86 = ~n325 ;
  assign y87 = n326 ;
  assign y88 = n333 ;
  assign y89 = ~1'b0 ;
  assign y90 = ~n335 ;
  assign y91 = ~n341 ;
  assign y92 = n345 ;
  assign y93 = n346 ;
  assign y94 = ~n358 ;
  assign y95 = ~1'b0 ;
  assign y96 = ~1'b0 ;
  assign y97 = ~n362 ;
  assign y98 = ~1'b0 ;
  assign y99 = n363 ;
  assign y100 = n372 ;
  assign y101 = ~n376 ;
  assign y102 = ~n391 ;
  assign y103 = n392 ;
  assign y104 = n393 ;
  assign y105 = n400 ;
  assign y106 = ~n401 ;
  assign y107 = n410 ;
  assign y108 = ~n418 ;
  assign y109 = ~n421 ;
  assign y110 = ~n422 ;
  assign y111 = n425 ;
  assign y112 = ~1'b0 ;
  assign y113 = n428 ;
  assign y114 = ~1'b0 ;
  assign y115 = ~n431 ;
  assign y116 = n432 ;
  assign y117 = n433 ;
  assign y118 = ~n437 ;
  assign y119 = n440 ;
  assign y120 = n441 ;
  assign y121 = ~n443 ;
  assign y122 = ~n447 ;
  assign y123 = ~n448 ;
  assign y124 = ~1'b0 ;
  assign y125 = ~n454 ;
  assign y126 = n432 ;
  assign y127 = n462 ;
  assign y128 = n464 ;
  assign y129 = ~n466 ;
  assign y130 = ~n472 ;
  assign y131 = n473 ;
  assign y132 = ~n480 ;
  assign y133 = n485 ;
  assign y134 = ~n492 ;
  assign y135 = n497 ;
  assign y136 = n498 ;
  assign y137 = n500 ;
  assign y138 = ~1'b0 ;
  assign y139 = ~n514 ;
  assign y140 = ~1'b0 ;
  assign y141 = ~n518 ;
  assign y142 = ~n523 ;
  assign y143 = n526 ;
  assign y144 = ~1'b0 ;
  assign y145 = ~n531 ;
  assign y146 = ~n539 ;
  assign y147 = ~n549 ;
  assign y148 = ~n553 ;
  assign y149 = n554 ;
  assign y150 = ~1'b0 ;
  assign y151 = ~n557 ;
  assign y152 = ~1'b0 ;
  assign y153 = ~1'b0 ;
  assign y154 = n558 ;
  assign y155 = ~n560 ;
  assign y156 = ~1'b0 ;
  assign y157 = ~n562 ;
  assign y158 = ~n564 ;
  assign y159 = ~1'b0 ;
  assign y160 = n567 ;
  assign y161 = n570 ;
  assign y162 = ~n575 ;
  assign y163 = n584 ;
  assign y164 = n593 ;
  assign y165 = n595 ;
  assign y166 = ~n604 ;
  assign y167 = ~1'b0 ;
  assign y168 = ~1'b0 ;
  assign y169 = n608 ;
  assign y170 = ~n615 ;
  assign y171 = n623 ;
  assign y172 = ~n627 ;
  assign y173 = n628 ;
  assign y174 = ~1'b0 ;
  assign y175 = n633 ;
  assign y176 = n644 ;
  assign y177 = ~n645 ;
  assign y178 = ~n647 ;
  assign y179 = ~1'b0 ;
  assign y180 = ~n650 ;
  assign y181 = ~n652 ;
  assign y182 = ~n660 ;
  assign y183 = n666 ;
  assign y184 = n670 ;
  assign y185 = n673 ;
  assign y186 = ~1'b0 ;
  assign y187 = ~n681 ;
  assign y188 = ~1'b0 ;
  assign y189 = ~n683 ;
  assign y190 = n688 ;
  assign y191 = n695 ;
  assign y192 = ~1'b0 ;
  assign y193 = ~n702 ;
  assign y194 = ~n712 ;
  assign y195 = n721 ;
  assign y196 = n724 ;
  assign y197 = ~n727 ;
  assign y198 = n741 ;
  assign y199 = ~n742 ;
  assign y200 = ~n744 ;
  assign y201 = ~n746 ;
  assign y202 = n751 ;
  assign y203 = n753 ;
  assign y204 = n766 ;
  assign y205 = n776 ;
  assign y206 = ~n779 ;
  assign y207 = ~n785 ;
  assign y208 = n786 ;
  assign y209 = n801 ;
  assign y210 = n802 ;
  assign y211 = ~n803 ;
  assign y212 = ~n805 ;
  assign y213 = n808 ;
  assign y214 = ~n811 ;
  assign y215 = ~1'b0 ;
  assign y216 = n819 ;
  assign y217 = ~n834 ;
  assign y218 = ~n836 ;
  assign y219 = n841 ;
  assign y220 = n843 ;
  assign y221 = ~n851 ;
  assign y222 = n853 ;
  assign y223 = n862 ;
  assign y224 = ~n864 ;
  assign y225 = n868 ;
  assign y226 = ~n870 ;
  assign y227 = ~n872 ;
  assign y228 = ~1'b0 ;
  assign y229 = ~1'b0 ;
  assign y230 = ~n877 ;
  assign y231 = ~n884 ;
  assign y232 = ~n888 ;
  assign y233 = ~n893 ;
  assign y234 = n894 ;
  assign y235 = n900 ;
  assign y236 = ~1'b0 ;
  assign y237 = n902 ;
  assign y238 = ~n903 ;
  assign y239 = ~1'b0 ;
  assign y240 = n909 ;
  assign y241 = ~n912 ;
  assign y242 = n913 ;
  assign y243 = ~n920 ;
  assign y244 = n925 ;
  assign y245 = ~1'b0 ;
  assign y246 = ~1'b0 ;
  assign y247 = n928 ;
  assign y248 = n929 ;
  assign y249 = n932 ;
  assign y250 = 1'b0 ;
  assign y251 = ~n937 ;
  assign y252 = n938 ;
  assign y253 = ~n945 ;
  assign y254 = ~1'b0 ;
  assign y255 = n948 ;
  assign y256 = ~n949 ;
  assign y257 = n952 ;
  assign y258 = n955 ;
  assign y259 = ~n962 ;
  assign y260 = ~n967 ;
  assign y261 = n972 ;
  assign y262 = ~n975 ;
  assign y263 = n977 ;
  assign y264 = n980 ;
  assign y265 = ~n982 ;
  assign y266 = n984 ;
  assign y267 = n989 ;
  assign y268 = n990 ;
  assign y269 = ~1'b0 ;
  assign y270 = n995 ;
  assign y271 = n999 ;
  assign y272 = ~n1000 ;
  assign y273 = n1002 ;
  assign y274 = n1016 ;
  assign y275 = ~n1023 ;
  assign y276 = ~n1037 ;
  assign y277 = ~n1040 ;
  assign y278 = n1042 ;
  assign y279 = ~n1047 ;
  assign y280 = ~1'b0 ;
  assign y281 = ~1'b0 ;
  assign y282 = ~n1049 ;
  assign y283 = n1052 ;
  assign y284 = n1054 ;
  assign y285 = ~n1058 ;
  assign y286 = ~n1063 ;
  assign y287 = ~n1067 ;
  assign y288 = n1073 ;
  assign y289 = n1077 ;
  assign y290 = n1078 ;
  assign y291 = ~1'b0 ;
  assign y292 = ~n1091 ;
  assign y293 = ~1'b0 ;
  assign y294 = ~n1098 ;
  assign y295 = ~n1100 ;
  assign y296 = n1103 ;
  assign y297 = ~n1114 ;
  assign y298 = n1125 ;
  assign y299 = ~n1133 ;
  assign y300 = ~n1152 ;
  assign y301 = n1152 ;
  assign y302 = ~n1158 ;
  assign y303 = n1162 ;
  assign y304 = ~1'b0 ;
  assign y305 = ~n1166 ;
  assign y306 = n1179 ;
  assign y307 = ~n1180 ;
  assign y308 = ~n1190 ;
  assign y309 = n1191 ;
  assign y310 = n1199 ;
  assign y311 = ~n1203 ;
  assign y312 = ~n1206 ;
  assign y313 = ~n1208 ;
  assign y314 = ~1'b0 ;
  assign y315 = ~n1213 ;
  assign y316 = n1216 ;
  assign y317 = ~n1219 ;
  assign y318 = ~n1226 ;
  assign y319 = ~n1227 ;
  assign y320 = ~n1237 ;
  assign y321 = n1241 ;
  assign y322 = n1243 ;
  assign y323 = n1246 ;
  assign y324 = ~n1274 ;
  assign y325 = n1275 ;
  assign y326 = n1277 ;
  assign y327 = ~1'b0 ;
  assign y328 = ~n1280 ;
  assign y329 = ~n1284 ;
  assign y330 = n1288 ;
  assign y331 = ~n1297 ;
  assign y332 = ~n1300 ;
  assign y333 = ~n1301 ;
  assign y334 = ~n1304 ;
  assign y335 = ~1'b0 ;
  assign y336 = n1308 ;
  assign y337 = ~1'b0 ;
  assign y338 = n1312 ;
  assign y339 = n1317 ;
  assign y340 = ~n1322 ;
  assign y341 = n1325 ;
  assign y342 = ~1'b0 ;
  assign y343 = ~n1330 ;
  assign y344 = ~n1341 ;
  assign y345 = ~n1354 ;
  assign y346 = n1363 ;
  assign y347 = ~1'b0 ;
  assign y348 = n1365 ;
  assign y349 = ~1'b0 ;
  assign y350 = n1368 ;
  assign y351 = ~1'b0 ;
  assign y352 = ~n1373 ;
  assign y353 = n1376 ;
  assign y354 = ~n1385 ;
  assign y355 = ~n1396 ;
  assign y356 = ~n1425 ;
  assign y357 = ~1'b0 ;
  assign y358 = ~n1428 ;
  assign y359 = n1436 ;
  assign y360 = ~n1438 ;
  assign y361 = ~n1448 ;
  assign y362 = ~n1449 ;
  assign y363 = ~n1461 ;
  assign y364 = ~1'b0 ;
  assign y365 = n1468 ;
  assign y366 = ~n1469 ;
  assign y367 = ~n1472 ;
  assign y368 = n1473 ;
  assign y369 = ~1'b0 ;
  assign y370 = ~n1474 ;
  assign y371 = ~n1484 ;
  assign y372 = ~n1491 ;
  assign y373 = ~1'b0 ;
  assign y374 = ~n1492 ;
  assign y375 = n1497 ;
  assign y376 = ~n1507 ;
  assign y377 = ~n1510 ;
  assign y378 = 1'b0 ;
  assign y379 = n1511 ;
  assign y380 = n1513 ;
  assign y381 = n1518 ;
  assign y382 = n1527 ;
  assign y383 = ~1'b0 ;
  assign y384 = ~n1528 ;
  assign y385 = ~n1531 ;
  assign y386 = ~n1534 ;
  assign y387 = n1542 ;
  assign y388 = ~n1546 ;
  assign y389 = ~n1549 ;
  assign y390 = n1553 ;
  assign y391 = n1556 ;
  assign y392 = n1557 ;
  assign y393 = n1562 ;
  assign y394 = n1564 ;
  assign y395 = ~1'b0 ;
  assign y396 = ~n1582 ;
  assign y397 = ~n1583 ;
  assign y398 = ~n1588 ;
  assign y399 = n1590 ;
  assign y400 = ~n1609 ;
  assign y401 = n1610 ;
  assign y402 = n1612 ;
  assign y403 = n1623 ;
  assign y404 = ~n1626 ;
  assign y405 = n1627 ;
  assign y406 = ~n1628 ;
  assign y407 = ~1'b0 ;
  assign y408 = n1631 ;
  assign y409 = ~n1635 ;
  assign y410 = ~n1639 ;
  assign y411 = ~n1643 ;
  assign y412 = ~n1647 ;
  assign y413 = ~1'b0 ;
  assign y414 = ~n1651 ;
  assign y415 = n1656 ;
  assign y416 = n1666 ;
  assign y417 = n1668 ;
  assign y418 = ~n1676 ;
  assign y419 = n1678 ;
  assign y420 = ~1'b0 ;
  assign y421 = ~n1683 ;
  assign y422 = ~n1688 ;
  assign y423 = n1689 ;
  assign y424 = n1690 ;
  assign y425 = ~n1692 ;
  assign y426 = ~n1697 ;
  assign y427 = n1702 ;
  assign y428 = ~n1708 ;
  assign y429 = n1717 ;
  assign y430 = ~n1721 ;
  assign y431 = ~n1724 ;
  assign y432 = n1730 ;
  assign y433 = n1732 ;
  assign y434 = ~n1739 ;
  assign y435 = ~n1747 ;
  assign y436 = n1748 ;
  assign y437 = ~n1754 ;
  assign y438 = ~n1755 ;
  assign y439 = ~n1761 ;
  assign y440 = ~n1763 ;
  assign y441 = ~1'b0 ;
  assign y442 = ~n1768 ;
  assign y443 = ~1'b0 ;
  assign y444 = n1772 ;
  assign y445 = ~n1776 ;
  assign y446 = ~n1779 ;
  assign y447 = n1791 ;
  assign y448 = n1793 ;
  assign y449 = n1798 ;
  assign y450 = n1799 ;
  assign y451 = ~n1800 ;
  assign y452 = n1806 ;
  assign y453 = ~n1818 ;
  assign y454 = n1824 ;
  assign y455 = n1830 ;
  assign y456 = n1840 ;
  assign y457 = ~n1853 ;
  assign y458 = ~n1856 ;
  assign y459 = ~n1862 ;
  assign y460 = n1864 ;
  assign y461 = ~n1869 ;
  assign y462 = ~n1874 ;
  assign y463 = n1881 ;
  assign y464 = ~n1884 ;
  assign y465 = n1886 ;
  assign y466 = n1889 ;
  assign y467 = n1896 ;
  assign y468 = ~1'b0 ;
  assign y469 = ~n1897 ;
  assign y470 = n1906 ;
  assign y471 = ~n1915 ;
  assign y472 = ~n1916 ;
  assign y473 = n1919 ;
  assign y474 = ~n1921 ;
  assign y475 = n1922 ;
  assign y476 = n1932 ;
  assign y477 = n1938 ;
  assign y478 = ~1'b0 ;
  assign y479 = n1945 ;
  assign y480 = ~1'b0 ;
  assign y481 = n1950 ;
  assign y482 = ~1'b0 ;
  assign y483 = ~n536 ;
  assign y484 = ~n1951 ;
  assign y485 = n1952 ;
  assign y486 = ~n1957 ;
  assign y487 = n1968 ;
  assign y488 = n1974 ;
  assign y489 = ~1'b0 ;
  assign y490 = n1975 ;
  assign y491 = n1979 ;
  assign y492 = n1984 ;
  assign y493 = ~n1989 ;
  assign y494 = n1993 ;
  assign y495 = n2003 ;
  assign y496 = ~n2007 ;
  assign y497 = ~n2015 ;
  assign y498 = ~n2022 ;
  assign y499 = ~n2024 ;
  assign y500 = ~1'b0 ;
  assign y501 = ~n2026 ;
  assign y502 = ~n2027 ;
  assign y503 = ~n2031 ;
  assign y504 = ~1'b0 ;
  assign y505 = ~1'b0 ;
  assign y506 = n2043 ;
  assign y507 = n2046 ;
  assign y508 = ~n2049 ;
  assign y509 = ~n2057 ;
  assign y510 = ~n2063 ;
  assign y511 = n2074 ;
  assign y512 = ~n2077 ;
  assign y513 = ~n2087 ;
  assign y514 = n2089 ;
  assign y515 = ~n2091 ;
  assign y516 = n2095 ;
  assign y517 = ~n2099 ;
  assign y518 = ~n2102 ;
  assign y519 = n2106 ;
  assign y520 = ~n2108 ;
  assign y521 = n2110 ;
  assign y522 = ~n2121 ;
  assign y523 = n2123 ;
  assign y524 = n2124 ;
  assign y525 = ~n2127 ;
  assign y526 = ~n2128 ;
  assign y527 = ~n2130 ;
  assign y528 = ~n2132 ;
  assign y529 = ~n2135 ;
  assign y530 = ~n2140 ;
  assign y531 = ~n2143 ;
  assign y532 = ~n2146 ;
  assign y533 = ~n2148 ;
  assign y534 = ~n2150 ;
  assign y535 = n2152 ;
  assign y536 = ~1'b0 ;
  assign y537 = ~n2163 ;
  assign y538 = ~1'b0 ;
  assign y539 = ~n2169 ;
  assign y540 = n2173 ;
  assign y541 = n2174 ;
  assign y542 = n2175 ;
  assign y543 = ~n2178 ;
  assign y544 = n2179 ;
  assign y545 = ~1'b0 ;
  assign y546 = n2182 ;
  assign y547 = ~1'b0 ;
  assign y548 = ~n2185 ;
  assign y549 = ~n2193 ;
  assign y550 = n2195 ;
  assign y551 = n2205 ;
  assign y552 = ~n2207 ;
  assign y553 = ~1'b0 ;
  assign y554 = ~n2208 ;
  assign y555 = n2209 ;
  assign y556 = ~n2213 ;
  assign y557 = ~n2214 ;
  assign y558 = ~n2217 ;
  assign y559 = ~x88 ;
  assign y560 = ~n2218 ;
  assign y561 = ~n2234 ;
  assign y562 = ~n2242 ;
  assign y563 = n2257 ;
  assign y564 = ~1'b0 ;
  assign y565 = ~n2259 ;
  assign y566 = ~n2272 ;
  assign y567 = n2274 ;
  assign y568 = ~n2279 ;
  assign y569 = ~n2288 ;
  assign y570 = n2291 ;
  assign y571 = ~n2298 ;
  assign y572 = ~1'b0 ;
  assign y573 = ~n2304 ;
  assign y574 = ~n2315 ;
  assign y575 = n2320 ;
  assign y576 = n2333 ;
  assign y577 = ~n2348 ;
  assign y578 = ~n2355 ;
  assign y579 = n2370 ;
  assign y580 = ~n2372 ;
  assign y581 = ~n2373 ;
  assign y582 = n2378 ;
  assign y583 = n2386 ;
  assign y584 = n2387 ;
  assign y585 = ~n2393 ;
  assign y586 = n2394 ;
  assign y587 = n2402 ;
  assign y588 = ~1'b0 ;
  assign y589 = ~n2410 ;
  assign y590 = n2411 ;
  assign y591 = n2415 ;
  assign y592 = n2416 ;
  assign y593 = n2419 ;
  assign y594 = n2427 ;
  assign y595 = n2428 ;
  assign y596 = n2429 ;
  assign y597 = ~n2441 ;
  assign y598 = n2444 ;
  assign y599 = n2445 ;
  assign y600 = ~n2446 ;
  assign y601 = ~n2464 ;
  assign y602 = ~n2470 ;
  assign y603 = ~n2472 ;
  assign y604 = n2474 ;
  assign y605 = n1246 ;
  assign y606 = ~n2475 ;
  assign y607 = ~n2476 ;
  assign y608 = ~n2480 ;
  assign y609 = n2494 ;
  assign y610 = ~n2495 ;
  assign y611 = n2501 ;
  assign y612 = n2502 ;
  assign y613 = ~n2511 ;
  assign y614 = ~n1545 ;
  assign y615 = n2514 ;
  assign y616 = ~n2515 ;
  assign y617 = ~n2530 ;
  assign y618 = ~n2535 ;
  assign y619 = ~1'b0 ;
  assign y620 = ~n2536 ;
  assign y621 = n2539 ;
  assign y622 = ~1'b0 ;
  assign y623 = n2543 ;
  assign y624 = ~n2545 ;
  assign y625 = n2552 ;
  assign y626 = ~n2561 ;
  assign y627 = n2569 ;
  assign y628 = ~n2570 ;
  assign y629 = n2571 ;
  assign y630 = ~n2572 ;
  assign y631 = ~1'b0 ;
  assign y632 = n2577 ;
  assign y633 = ~1'b0 ;
  assign y634 = ~1'b0 ;
  assign y635 = ~n2580 ;
  assign y636 = n2582 ;
  assign y637 = ~1'b0 ;
  assign y638 = ~n2583 ;
  assign y639 = ~1'b0 ;
  assign y640 = ~1'b0 ;
  assign y641 = n2584 ;
  assign y642 = ~n2585 ;
  assign y643 = ~n2589 ;
  assign y644 = n2601 ;
  assign y645 = n2603 ;
  assign y646 = ~n2604 ;
  assign y647 = n2606 ;
  assign y648 = ~n2610 ;
  assign y649 = n2627 ;
  assign y650 = ~n2629 ;
  assign y651 = ~1'b0 ;
  assign y652 = n2637 ;
  assign y653 = ~n2643 ;
  assign y654 = n2667 ;
  assign y655 = n2677 ;
  assign y656 = ~n2679 ;
  assign y657 = ~n2684 ;
  assign y658 = n2691 ;
  assign y659 = n2696 ;
  assign y660 = ~1'b0 ;
  assign y661 = ~1'b0 ;
  assign y662 = n2698 ;
  assign y663 = n2704 ;
  assign y664 = n2712 ;
  assign y665 = ~1'b0 ;
  assign y666 = ~n2717 ;
  assign y667 = ~1'b0 ;
  assign y668 = n2724 ;
  assign y669 = ~n2725 ;
  assign y670 = n2733 ;
  assign y671 = ~n2740 ;
  assign y672 = n2744 ;
  assign y673 = n2753 ;
  assign y674 = ~1'b0 ;
  assign y675 = ~1'b0 ;
  assign y676 = n2754 ;
  assign y677 = n2759 ;
  assign y678 = ~1'b0 ;
  assign y679 = n2761 ;
  assign y680 = ~n2771 ;
  assign y681 = ~n2775 ;
  assign y682 = ~n2784 ;
  assign y683 = n2785 ;
  assign y684 = ~n2788 ;
  assign y685 = ~n2793 ;
  assign y686 = n2797 ;
  assign y687 = n2806 ;
  assign y688 = ~n2807 ;
  assign y689 = ~n2809 ;
  assign y690 = n2817 ;
  assign y691 = ~n2826 ;
  assign y692 = ~n2840 ;
  assign y693 = ~n2841 ;
  assign y694 = n2842 ;
  assign y695 = n2843 ;
  assign y696 = ~n2847 ;
  assign y697 = ~1'b0 ;
  assign y698 = n2851 ;
  assign y699 = ~1'b0 ;
  assign y700 = ~n2857 ;
  assign y701 = n2859 ;
  assign y702 = ~1'b0 ;
  assign y703 = ~1'b0 ;
  assign y704 = ~1'b0 ;
  assign y705 = n2864 ;
  assign y706 = n2873 ;
  assign y707 = n2879 ;
  assign y708 = ~n2881 ;
  assign y709 = n2882 ;
  assign y710 = n2891 ;
  assign y711 = n2896 ;
  assign y712 = ~n2906 ;
  assign y713 = ~n2912 ;
  assign y714 = ~1'b0 ;
  assign y715 = n2918 ;
  assign y716 = n2927 ;
  assign y717 = ~1'b0 ;
  assign y718 = ~n2932 ;
  assign y719 = n2934 ;
  assign y720 = n2939 ;
  assign y721 = ~n2947 ;
  assign y722 = ~n2948 ;
  assign y723 = n2951 ;
  assign y724 = n2957 ;
  assign y725 = n2960 ;
  assign y726 = ~n2009 ;
  assign y727 = ~1'b0 ;
  assign y728 = ~n2964 ;
  assign y729 = n2968 ;
  assign y730 = ~n2978 ;
  assign y731 = ~1'b0 ;
  assign y732 = ~n2983 ;
  assign y733 = n2994 ;
  assign y734 = ~1'b0 ;
  assign y735 = ~n2997 ;
  assign y736 = ~n3004 ;
  assign y737 = n3007 ;
  assign y738 = n3008 ;
  assign y739 = ~n3010 ;
  assign y740 = ~1'b0 ;
  assign y741 = n3011 ;
  assign y742 = ~n3015 ;
  assign y743 = n3017 ;
  assign y744 = n3018 ;
  assign y745 = ~n3024 ;
  assign y746 = n3025 ;
  assign y747 = n3026 ;
  assign y748 = ~1'b0 ;
  assign y749 = ~n3033 ;
  assign y750 = ~n3040 ;
  assign y751 = n3043 ;
  assign y752 = n3047 ;
  assign y753 = ~n3055 ;
  assign y754 = ~n3057 ;
  assign y755 = ~n3068 ;
  assign y756 = ~n3080 ;
  assign y757 = ~n3083 ;
  assign y758 = ~n3085 ;
  assign y759 = ~n3087 ;
  assign y760 = ~n3093 ;
  assign y761 = n3105 ;
  assign y762 = n3109 ;
  assign y763 = n3112 ;
  assign y764 = n3123 ;
  assign y765 = ~n3125 ;
  assign y766 = ~n3133 ;
  assign y767 = ~n3136 ;
  assign y768 = n3139 ;
  assign y769 = ~n3141 ;
  assign y770 = n3144 ;
  assign y771 = n3147 ;
  assign y772 = n3149 ;
  assign y773 = n3155 ;
  assign y774 = ~n3156 ;
  assign y775 = ~n3162 ;
  assign y776 = ~n3164 ;
  assign y777 = ~1'b0 ;
  assign y778 = n3171 ;
  assign y779 = ~n3172 ;
  assign y780 = n3173 ;
  assign y781 = ~n3188 ;
  assign y782 = n3189 ;
  assign y783 = ~n3191 ;
  assign y784 = ~1'b0 ;
  assign y785 = n3198 ;
  assign y786 = n3202 ;
  assign y787 = ~n3206 ;
  assign y788 = ~1'b0 ;
  assign y789 = ~n3215 ;
  assign y790 = ~n3219 ;
  assign y791 = n3220 ;
  assign y792 = ~1'b0 ;
  assign y793 = ~1'b0 ;
  assign y794 = ~n3223 ;
  assign y795 = n3228 ;
  assign y796 = ~1'b0 ;
  assign y797 = ~n3229 ;
  assign y798 = n3231 ;
  assign y799 = ~1'b0 ;
  assign y800 = ~n3236 ;
  assign y801 = n3249 ;
  assign y802 = ~1'b0 ;
  assign y803 = ~n3254 ;
  assign y804 = n3255 ;
  assign y805 = n3258 ;
  assign y806 = n3263 ;
  assign y807 = n3266 ;
  assign y808 = ~n3267 ;
  assign y809 = n3272 ;
  assign y810 = ~n3290 ;
  assign y811 = n3294 ;
  assign y812 = ~n3295 ;
  assign y813 = n3300 ;
  assign y814 = ~n3303 ;
  assign y815 = ~n3307 ;
  assign y816 = n3315 ;
  assign y817 = ~n3320 ;
  assign y818 = ~n3325 ;
  assign y819 = n3327 ;
  assign y820 = ~n3330 ;
  assign y821 = ~n3337 ;
  assign y822 = n3342 ;
  assign y823 = n3350 ;
  assign y824 = n3351 ;
  assign y825 = n3359 ;
  assign y826 = ~n3362 ;
  assign y827 = ~n3371 ;
  assign y828 = ~n3375 ;
  assign y829 = ~n3385 ;
  assign y830 = ~n3392 ;
  assign y831 = n3399 ;
  assign y832 = n3401 ;
  assign y833 = ~1'b0 ;
  assign y834 = n3407 ;
  assign y835 = ~n3411 ;
  assign y836 = ~n3413 ;
  assign y837 = ~n3415 ;
  assign y838 = ~n3420 ;
  assign y839 = ~n3421 ;
  assign y840 = ~1'b0 ;
  assign y841 = n3428 ;
  assign y842 = n3430 ;
  assign y843 = ~n3431 ;
  assign y844 = ~n3433 ;
  assign y845 = ~1'b0 ;
  assign y846 = ~n3436 ;
  assign y847 = ~n3444 ;
  assign y848 = ~n3450 ;
  assign y849 = n3452 ;
  assign y850 = ~n3454 ;
  assign y851 = ~n3456 ;
  assign y852 = n3467 ;
  assign y853 = ~n3470 ;
  assign y854 = n3471 ;
  assign y855 = ~n3483 ;
  assign y856 = ~n3500 ;
  assign y857 = ~n3502 ;
  assign y858 = ~n3509 ;
  assign y859 = ~n3510 ;
  assign y860 = ~n3516 ;
  assign y861 = ~n3523 ;
  assign y862 = n3527 ;
  assign y863 = n3529 ;
  assign y864 = n3537 ;
  assign y865 = ~n3542 ;
  assign y866 = ~n3548 ;
  assign y867 = n3549 ;
  assign y868 = ~n3560 ;
  assign y869 = ~1'b0 ;
  assign y870 = ~1'b0 ;
  assign y871 = ~n3562 ;
  assign y872 = ~n3564 ;
  assign y873 = ~n3571 ;
  assign y874 = n3582 ;
  assign y875 = n3583 ;
  assign y876 = ~n3584 ;
  assign y877 = ~n3588 ;
  assign y878 = ~n3589 ;
  assign y879 = n3590 ;
  assign y880 = ~n3591 ;
  assign y881 = n3596 ;
  assign y882 = n3600 ;
  assign y883 = n3603 ;
  assign y884 = n3604 ;
  assign y885 = ~n3608 ;
  assign y886 = ~n3611 ;
  assign y887 = n3613 ;
  assign y888 = ~1'b0 ;
  assign y889 = ~n3620 ;
  assign y890 = n3625 ;
  assign y891 = n3630 ;
  assign y892 = n3637 ;
  assign y893 = ~1'b0 ;
  assign y894 = n3640 ;
  assign y895 = n3642 ;
  assign y896 = n3643 ;
  assign y897 = n3645 ;
  assign y898 = n3647 ;
  assign y899 = n3653 ;
  assign y900 = ~n3658 ;
  assign y901 = n3661 ;
  assign y902 = n3667 ;
  assign y903 = n3671 ;
  assign y904 = ~n3681 ;
  assign y905 = n3692 ;
  assign y906 = n3697 ;
  assign y907 = ~n3703 ;
  assign y908 = n3704 ;
  assign y909 = n3710 ;
  assign y910 = n3722 ;
  assign y911 = ~n3725 ;
  assign y912 = ~n3730 ;
  assign y913 = n3737 ;
  assign y914 = ~n3744 ;
  assign y915 = ~n3746 ;
  assign y916 = ~n3748 ;
  assign y917 = ~n3756 ;
  assign y918 = ~n3774 ;
  assign y919 = ~1'b0 ;
  assign y920 = ~n3780 ;
  assign y921 = n3781 ;
  assign y922 = ~n3785 ;
  assign y923 = ~n3786 ;
  assign y924 = n3793 ;
  assign y925 = ~n3803 ;
  assign y926 = n3809 ;
  assign y927 = n3814 ;
  assign y928 = ~n3819 ;
  assign y929 = ~n3820 ;
  assign y930 = n3824 ;
  assign y931 = ~1'b0 ;
  assign y932 = n3827 ;
  assign y933 = n3200 ;
  assign y934 = n3833 ;
  assign y935 = ~1'b0 ;
  assign y936 = n3843 ;
  assign y937 = n3844 ;
  assign y938 = ~n3846 ;
  assign y939 = n3854 ;
  assign y940 = ~n3857 ;
  assign y941 = n3858 ;
  assign y942 = ~n3871 ;
  assign y943 = n3873 ;
  assign y944 = ~1'b0 ;
  assign y945 = n3874 ;
  assign y946 = ~n3877 ;
  assign y947 = ~1'b0 ;
  assign y948 = n3881 ;
  assign y949 = ~1'b0 ;
  assign y950 = n3895 ;
  assign y951 = ~n3905 ;
  assign y952 = ~1'b0 ;
  assign y953 = n3906 ;
  assign y954 = ~n3909 ;
  assign y955 = ~n3911 ;
  assign y956 = ~n3912 ;
  assign y957 = ~n3920 ;
  assign y958 = ~n3924 ;
  assign y959 = n3931 ;
  assign y960 = n3934 ;
  assign y961 = n3935 ;
  assign y962 = ~1'b0 ;
  assign y963 = ~n3937 ;
  assign y964 = ~1'b0 ;
  assign y965 = ~n3941 ;
  assign y966 = ~n3943 ;
  assign y967 = ~n3958 ;
  assign y968 = n3961 ;
  assign y969 = n3962 ;
  assign y970 = ~n3965 ;
  assign y971 = n3967 ;
  assign y972 = ~n3969 ;
  assign y973 = n3976 ;
  assign y974 = ~n3985 ;
  assign y975 = n3989 ;
  assign y976 = n3996 ;
  assign y977 = ~n4006 ;
  assign y978 = n4009 ;
  assign y979 = ~n4011 ;
  assign y980 = ~n4021 ;
  assign y981 = ~1'b0 ;
  assign y982 = ~n4023 ;
  assign y983 = ~n4025 ;
  assign y984 = ~n4030 ;
  assign y985 = n4032 ;
  assign y986 = ~n4044 ;
  assign y987 = ~n4045 ;
  assign y988 = ~n4049 ;
  assign y989 = ~n4052 ;
  assign y990 = n4056 ;
  assign y991 = n4057 ;
  assign y992 = n4070 ;
  assign y993 = ~n4077 ;
  assign y994 = ~1'b0 ;
  assign y995 = n4093 ;
  assign y996 = ~n4094 ;
  assign y997 = ~n4107 ;
  assign y998 = n4115 ;
  assign y999 = ~1'b0 ;
  assign y1000 = ~n4117 ;
  assign y1001 = ~n4121 ;
  assign y1002 = ~n4123 ;
  assign y1003 = ~n4132 ;
  assign y1004 = ~n4134 ;
  assign y1005 = n4139 ;
  assign y1006 = ~n4151 ;
  assign y1007 = ~n4160 ;
  assign y1008 = n4166 ;
  assign y1009 = n4175 ;
  assign y1010 = n4189 ;
  assign y1011 = n4195 ;
  assign y1012 = ~n4201 ;
  assign y1013 = n4206 ;
  assign y1014 = ~1'b0 ;
  assign y1015 = ~1'b0 ;
  assign y1016 = ~1'b0 ;
  assign y1017 = ~n4210 ;
  assign y1018 = ~n4223 ;
  assign y1019 = ~n4224 ;
  assign y1020 = n4226 ;
  assign y1021 = n4227 ;
  assign y1022 = n4228 ;
  assign y1023 = ~n4231 ;
  assign y1024 = n4232 ;
  assign y1025 = ~n4244 ;
  assign y1026 = ~n4248 ;
  assign y1027 = n4251 ;
  assign y1028 = n4254 ;
  assign y1029 = ~n4262 ;
  assign y1030 = n4263 ;
  assign y1031 = ~n4268 ;
  assign y1032 = ~n4275 ;
  assign y1033 = ~n4280 ;
  assign y1034 = ~n4283 ;
  assign y1035 = ~n4285 ;
  assign y1036 = n4290 ;
  assign y1037 = n4302 ;
  assign y1038 = n4305 ;
  assign y1039 = ~n4309 ;
  assign y1040 = ~n4311 ;
  assign y1041 = ~1'b0 ;
  assign y1042 = n4322 ;
  assign y1043 = n4329 ;
  assign y1044 = ~n4331 ;
  assign y1045 = ~n4338 ;
  assign y1046 = ~n4339 ;
  assign y1047 = ~n4343 ;
  assign y1048 = ~n4345 ;
  assign y1049 = ~n4346 ;
  assign y1050 = n4350 ;
  assign y1051 = ~n4353 ;
  assign y1052 = ~1'b0 ;
  assign y1053 = ~n4356 ;
  assign y1054 = n4357 ;
  assign y1055 = n4365 ;
  assign y1056 = ~n4366 ;
  assign y1057 = n4382 ;
  assign y1058 = ~n4386 ;
  assign y1059 = n4389 ;
  assign y1060 = ~n4390 ;
  assign y1061 = n4394 ;
  assign y1062 = ~n4399 ;
  assign y1063 = n4404 ;
  assign y1064 = n4405 ;
  assign y1065 = ~n4407 ;
  assign y1066 = ~n4415 ;
  assign y1067 = n4424 ;
  assign y1068 = n4425 ;
  assign y1069 = n4434 ;
  assign y1070 = ~1'b0 ;
  assign y1071 = n4438 ;
  assign y1072 = n4443 ;
  assign y1073 = n4449 ;
  assign y1074 = n4452 ;
  assign y1075 = ~n4454 ;
  assign y1076 = n4466 ;
  assign y1077 = n4467 ;
  assign y1078 = ~n4470 ;
  assign y1079 = n4483 ;
  assign y1080 = ~n4487 ;
  assign y1081 = n4488 ;
  assign y1082 = n4492 ;
  assign y1083 = n4494 ;
  assign y1084 = ~1'b0 ;
  assign y1085 = n4498 ;
  assign y1086 = x41 ;
  assign y1087 = n4499 ;
  assign y1088 = n4507 ;
  assign y1089 = n4514 ;
  assign y1090 = ~n4537 ;
  assign y1091 = n4541 ;
  assign y1092 = ~n4546 ;
  assign y1093 = n4547 ;
  assign y1094 = n4555 ;
  assign y1095 = ~1'b0 ;
  assign y1096 = ~n4560 ;
  assign y1097 = ~n4562 ;
  assign y1098 = ~n4574 ;
  assign y1099 = ~1'b0 ;
  assign y1100 = n4579 ;
  assign y1101 = ~n4581 ;
  assign y1102 = 1'b0 ;
  assign y1103 = n4585 ;
  assign y1104 = n4587 ;
  assign y1105 = ~1'b0 ;
  assign y1106 = ~n4589 ;
  assign y1107 = ~n3408 ;
  assign y1108 = ~n4602 ;
  assign y1109 = ~n4605 ;
  assign y1110 = n4617 ;
  assign y1111 = ~n4619 ;
  assign y1112 = ~n4622 ;
  assign y1113 = ~1'b0 ;
  assign y1114 = ~1'b0 ;
  assign y1115 = n4623 ;
  assign y1116 = ~n4624 ;
  assign y1117 = ~n4633 ;
  assign y1118 = n4636 ;
  assign y1119 = ~n4639 ;
  assign y1120 = n4649 ;
  assign y1121 = ~n4656 ;
  assign y1122 = n4661 ;
  assign y1123 = ~n4662 ;
  assign y1124 = ~n4668 ;
  assign y1125 = n4670 ;
  assign y1126 = n4671 ;
  assign y1127 = ~n4673 ;
  assign y1128 = ~n4678 ;
  assign y1129 = n4688 ;
  assign y1130 = ~1'b0 ;
  assign y1131 = ~n4694 ;
  assign y1132 = ~1'b0 ;
  assign y1133 = n4698 ;
  assign y1134 = ~n4700 ;
  assign y1135 = n4703 ;
  assign y1136 = n4717 ;
  assign y1137 = n4726 ;
  assign y1138 = ~n4729 ;
  assign y1139 = ~n4733 ;
  assign y1140 = n4738 ;
  assign y1141 = ~n4748 ;
  assign y1142 = ~n4750 ;
  assign y1143 = ~n4753 ;
  assign y1144 = ~n4755 ;
  assign y1145 = ~n4763 ;
  assign y1146 = n4765 ;
  assign y1147 = ~1'b0 ;
  assign y1148 = n4766 ;
  assign y1149 = ~1'b0 ;
  assign y1150 = n4769 ;
  assign y1151 = n4773 ;
  assign y1152 = n4777 ;
  assign y1153 = n4779 ;
  assign y1154 = n4781 ;
  assign y1155 = n4785 ;
  assign y1156 = ~n4786 ;
  assign y1157 = n4787 ;
  assign y1158 = n4793 ;
  assign y1159 = n4794 ;
  assign y1160 = n4795 ;
  assign y1161 = n4798 ;
  assign y1162 = n4800 ;
  assign y1163 = n4804 ;
  assign y1164 = ~n4811 ;
  assign y1165 = n4815 ;
  assign y1166 = n4816 ;
  assign y1167 = ~n4817 ;
  assign y1168 = n4819 ;
  assign y1169 = n4820 ;
  assign y1170 = n4821 ;
  assign y1171 = n4825 ;
  assign y1172 = n4833 ;
  assign y1173 = n4841 ;
  assign y1174 = ~n4842 ;
  assign y1175 = 1'b0 ;
  assign y1176 = ~n4851 ;
  assign y1177 = ~n4862 ;
  assign y1178 = ~n4871 ;
  assign y1179 = ~n4872 ;
  assign y1180 = n4873 ;
  assign y1181 = ~n4875 ;
  assign y1182 = ~n4883 ;
  assign y1183 = ~n4884 ;
  assign y1184 = n4897 ;
  assign y1185 = n4899 ;
  assign y1186 = ~n4904 ;
  assign y1187 = ~n4913 ;
  assign y1188 = ~n4914 ;
  assign y1189 = n4922 ;
  assign y1190 = n4923 ;
  assign y1191 = n4926 ;
  assign y1192 = ~n4927 ;
  assign y1193 = n4932 ;
  assign y1194 = ~1'b0 ;
  assign y1195 = ~1'b0 ;
  assign y1196 = n4939 ;
  assign y1197 = ~1'b0 ;
  assign y1198 = n959 ;
  assign y1199 = ~n327 ;
  assign y1200 = n4941 ;
  assign y1201 = ~n4945 ;
  assign y1202 = ~n4946 ;
  assign y1203 = ~n4948 ;
  assign y1204 = n4949 ;
  assign y1205 = ~n4951 ;
  assign y1206 = ~n4952 ;
  assign y1207 = n4954 ;
  assign y1208 = ~n4958 ;
  assign y1209 = ~n4963 ;
  assign y1210 = n4969 ;
  assign y1211 = ~1'b0 ;
  assign y1212 = n4971 ;
  assign y1213 = ~1'b0 ;
  assign y1214 = ~n4976 ;
  assign y1215 = ~n4977 ;
  assign y1216 = ~n4981 ;
  assign y1217 = ~1'b0 ;
  assign y1218 = ~n4982 ;
  assign y1219 = ~1'b0 ;
  assign y1220 = ~1'b0 ;
  assign y1221 = ~n4984 ;
  assign y1222 = ~n4990 ;
  assign y1223 = ~n4995 ;
  assign y1224 = ~n4997 ;
  assign y1225 = ~1'b0 ;
  assign y1226 = ~n5002 ;
  assign y1227 = ~n5006 ;
  assign y1228 = ~n5012 ;
  assign y1229 = ~n5013 ;
  assign y1230 = ~n5014 ;
  assign y1231 = ~n5015 ;
  assign y1232 = ~n5022 ;
  assign y1233 = ~1'b0 ;
  assign y1234 = n5025 ;
  assign y1235 = n5027 ;
  assign y1236 = n5033 ;
  assign y1237 = ~n5037 ;
  assign y1238 = ~1'b0 ;
  assign y1239 = ~n5038 ;
  assign y1240 = ~n5040 ;
  assign y1241 = n5046 ;
  assign y1242 = ~n5054 ;
  assign y1243 = ~n5057 ;
  assign y1244 = ~n5059 ;
  assign y1245 = ~n5066 ;
  assign y1246 = n5087 ;
  assign y1247 = ~n5091 ;
  assign y1248 = n5094 ;
  assign y1249 = ~1'b0 ;
  assign y1250 = n5098 ;
  assign y1251 = ~n5101 ;
  assign y1252 = n5108 ;
  assign y1253 = ~n5112 ;
  assign y1254 = ~n5116 ;
  assign y1255 = ~n5118 ;
  assign y1256 = ~n5123 ;
  assign y1257 = ~n5127 ;
  assign y1258 = n5131 ;
  assign y1259 = ~1'b0 ;
  assign y1260 = n5134 ;
  assign y1261 = ~n5135 ;
  assign y1262 = n5137 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = n5139 ;
  assign y1265 = ~n5140 ;
  assign y1266 = ~n5142 ;
  assign y1267 = ~n5158 ;
  assign y1268 = n4662 ;
  assign y1269 = ~n5159 ;
  assign y1270 = ~n5165 ;
  assign y1271 = ~1'b0 ;
  assign y1272 = n5166 ;
  assign y1273 = n5173 ;
  assign y1274 = n326 ;
  assign y1275 = ~n5175 ;
  assign y1276 = ~n5184 ;
  assign y1277 = n5192 ;
  assign y1278 = n5194 ;
  assign y1279 = n5195 ;
  assign y1280 = n5196 ;
  assign y1281 = n5197 ;
  assign y1282 = ~n5202 ;
  assign y1283 = ~1'b0 ;
  assign y1284 = n5206 ;
  assign y1285 = ~n5209 ;
  assign y1286 = n5216 ;
  assign y1287 = ~n5218 ;
  assign y1288 = n5222 ;
  assign y1289 = ~n5225 ;
  assign y1290 = ~n5226 ;
  assign y1291 = ~n5231 ;
  assign y1292 = n5235 ;
  assign y1293 = ~n5239 ;
  assign y1294 = n5264 ;
  assign y1295 = n5272 ;
  assign y1296 = ~n5275 ;
  assign y1297 = n5129 ;
  assign y1298 = n5276 ;
  assign y1299 = n5278 ;
  assign y1300 = ~n5282 ;
  assign y1301 = ~n5283 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = ~n5288 ;
  assign y1304 = ~n5295 ;
  assign y1305 = n5299 ;
  assign y1306 = ~1'b0 ;
  assign y1307 = ~n5301 ;
  assign y1308 = n5303 ;
  assign y1309 = ~n5310 ;
  assign y1310 = ~n5320 ;
  assign y1311 = ~n5323 ;
  assign y1312 = n5326 ;
  assign y1313 = n5327 ;
  assign y1314 = n5339 ;
  assign y1315 = ~n5343 ;
  assign y1316 = ~n5345 ;
  assign y1317 = n5347 ;
  assign y1318 = n5348 ;
  assign y1319 = ~n5359 ;
  assign y1320 = n5362 ;
  assign y1321 = n5367 ;
  assign y1322 = ~n5368 ;
  assign y1323 = n5369 ;
  assign y1324 = ~n5372 ;
  assign y1325 = n5376 ;
  assign y1326 = ~n5377 ;
  assign y1327 = ~n5388 ;
  assign y1328 = ~1'b0 ;
  assign y1329 = n5391 ;
  assign y1330 = ~n5401 ;
  assign y1331 = n5403 ;
  assign y1332 = n5411 ;
  assign y1333 = ~n5414 ;
  assign y1334 = n5416 ;
  assign y1335 = n5417 ;
  assign y1336 = n5421 ;
  assign y1337 = ~n5423 ;
  assign y1338 = ~n5429 ;
  assign y1339 = ~1'b0 ;
  assign y1340 = n5431 ;
  assign y1341 = ~n5435 ;
  assign y1342 = n5439 ;
  assign y1343 = ~1'b0 ;
  assign y1344 = ~n5440 ;
  assign y1345 = n5444 ;
  assign y1346 = ~1'b0 ;
  assign y1347 = n5446 ;
  assign y1348 = ~n5450 ;
  assign y1349 = ~n5452 ;
  assign y1350 = ~n5458 ;
  assign y1351 = ~n5461 ;
  assign y1352 = ~n5465 ;
  assign y1353 = n5474 ;
  assign y1354 = n5478 ;
  assign y1355 = ~n5492 ;
  assign y1356 = n5495 ;
  assign y1357 = n5497 ;
  assign y1358 = n5498 ;
  assign y1359 = ~n5507 ;
  assign y1360 = ~n5514 ;
  assign y1361 = n5521 ;
  assign y1362 = ~n5526 ;
  assign y1363 = ~1'b0 ;
  assign y1364 = ~n5531 ;
  assign y1365 = n5537 ;
  assign y1366 = ~1'b0 ;
  assign y1367 = ~n5548 ;
  assign y1368 = ~n5551 ;
  assign y1369 = ~n5553 ;
  assign y1370 = ~n5555 ;
  assign y1371 = ~n5557 ;
  assign y1372 = n5559 ;
  assign y1373 = ~n5560 ;
  assign y1374 = n5566 ;
  assign y1375 = ~n5573 ;
  assign y1376 = ~n5581 ;
  assign y1377 = ~n5583 ;
  assign y1378 = ~n5585 ;
  assign y1379 = ~1'b0 ;
  assign y1380 = ~1'b0 ;
  assign y1381 = ~n5588 ;
  assign y1382 = n5592 ;
  assign y1383 = n5596 ;
  assign y1384 = ~n5599 ;
  assign y1385 = n5604 ;
  assign y1386 = ~1'b0 ;
  assign y1387 = ~1'b0 ;
  assign y1388 = ~n5606 ;
  assign y1389 = ~n5615 ;
  assign y1390 = ~1'b0 ;
  assign y1391 = ~n5636 ;
  assign y1392 = ~n5642 ;
  assign y1393 = ~n5645 ;
  assign y1394 = n5647 ;
  assign y1395 = ~n5655 ;
  assign y1396 = n5662 ;
  assign y1397 = ~n5663 ;
  assign y1398 = n5676 ;
  assign y1399 = ~n5677 ;
  assign y1400 = ~1'b0 ;
  assign y1401 = ~n5684 ;
  assign y1402 = n5690 ;
  assign y1403 = n5695 ;
  assign y1404 = n5700 ;
  assign y1405 = ~n5705 ;
  assign y1406 = n5712 ;
  assign y1407 = n5721 ;
  assign y1408 = ~n5722 ;
  assign y1409 = ~n5725 ;
  assign y1410 = n5730 ;
  assign y1411 = ~n5731 ;
  assign y1412 = n5734 ;
  assign y1413 = n5735 ;
  assign y1414 = n5752 ;
  assign y1415 = ~n5753 ;
  assign y1416 = ~n5755 ;
  assign y1417 = ~n5756 ;
  assign y1418 = n5758 ;
  assign y1419 = ~n5761 ;
  assign y1420 = ~1'b0 ;
  assign y1421 = ~n5762 ;
  assign y1422 = n4996 ;
  assign y1423 = n5767 ;
  assign y1424 = ~1'b0 ;
  assign y1425 = n5769 ;
  assign y1426 = ~n5771 ;
  assign y1427 = ~n5778 ;
  assign y1428 = ~1'b0 ;
  assign y1429 = ~n5780 ;
  assign y1430 = n5786 ;
  assign y1431 = ~n5788 ;
  assign y1432 = n5789 ;
  assign y1433 = n5793 ;
  assign y1434 = ~n5814 ;
  assign y1435 = ~1'b0 ;
  assign y1436 = ~n5820 ;
  assign y1437 = ~1'b0 ;
  assign y1438 = n5827 ;
  assign y1439 = n5828 ;
  assign y1440 = n5833 ;
  assign y1441 = ~n5836 ;
  assign y1442 = n5838 ;
  assign y1443 = ~1'b0 ;
  assign y1444 = ~n5839 ;
  assign y1445 = n5842 ;
  assign y1446 = n5846 ;
  assign y1447 = n5850 ;
  assign y1448 = ~1'b0 ;
  assign y1449 = n5851 ;
  assign y1450 = n5856 ;
  assign y1451 = n5863 ;
  assign y1452 = ~n5865 ;
  assign y1453 = ~n5867 ;
  assign y1454 = n5868 ;
  assign y1455 = ~1'b0 ;
  assign y1456 = n5871 ;
  assign y1457 = ~n5876 ;
  assign y1458 = ~1'b0 ;
  assign y1459 = ~n5878 ;
  assign y1460 = ~n5880 ;
  assign y1461 = n5884 ;
  assign y1462 = n5897 ;
  assign y1463 = ~1'b0 ;
  assign y1464 = ~1'b0 ;
  assign y1465 = ~n5912 ;
  assign y1466 = ~n5923 ;
  assign y1467 = n5926 ;
  assign y1468 = ~n5927 ;
  assign y1469 = n5928 ;
  assign y1470 = ~n5931 ;
  assign y1471 = ~1'b0 ;
  assign y1472 = ~n5945 ;
  assign y1473 = ~n5947 ;
  assign y1474 = ~n5948 ;
  assign y1475 = n5952 ;
  assign y1476 = n5954 ;
  assign y1477 = n5955 ;
  assign y1478 = n5963 ;
  assign y1479 = ~1'b0 ;
  assign y1480 = n5966 ;
  assign y1481 = ~n5971 ;
  assign y1482 = n5976 ;
  assign y1483 = n5979 ;
  assign y1484 = n5980 ;
  assign y1485 = ~n5984 ;
  assign y1486 = ~1'b0 ;
  assign y1487 = ~1'b0 ;
  assign y1488 = n5994 ;
  assign y1489 = n5997 ;
  assign y1490 = n5998 ;
  assign y1491 = ~n6000 ;
  assign y1492 = n6002 ;
  assign y1493 = n6003 ;
  assign y1494 = ~n6009 ;
  assign y1495 = ~n6012 ;
  assign y1496 = ~n6020 ;
  assign y1497 = n6029 ;
  assign y1498 = ~1'b0 ;
  assign y1499 = n6035 ;
  assign y1500 = n6039 ;
  assign y1501 = n6042 ;
  assign y1502 = ~n6048 ;
  assign y1503 = ~n6053 ;
  assign y1504 = ~n6056 ;
  assign y1505 = ~n6061 ;
  assign y1506 = n6067 ;
  assign y1507 = n6070 ;
  assign y1508 = ~1'b0 ;
  assign y1509 = n6073 ;
  assign y1510 = n6078 ;
  assign y1511 = n6088 ;
  assign y1512 = n6090 ;
  assign y1513 = n6092 ;
  assign y1514 = ~n6103 ;
  assign y1515 = ~n6110 ;
  assign y1516 = n6115 ;
  assign y1517 = n6118 ;
  assign y1518 = ~1'b0 ;
  assign y1519 = n6121 ;
  assign y1520 = ~n6130 ;
  assign y1521 = n6131 ;
  assign y1522 = ~n6134 ;
  assign y1523 = ~n6156 ;
  assign y1524 = ~n6167 ;
  assign y1525 = ~1'b0 ;
  assign y1526 = ~n6168 ;
  assign y1527 = ~n6169 ;
  assign y1528 = ~n6171 ;
  assign y1529 = ~n6173 ;
  assign y1530 = n6176 ;
  assign y1531 = ~n6179 ;
  assign y1532 = ~n6182 ;
  assign y1533 = ~1'b0 ;
  assign y1534 = n6186 ;
  assign y1535 = ~n6189 ;
  assign y1536 = n6192 ;
  assign y1537 = ~n6200 ;
  assign y1538 = ~n6201 ;
  assign y1539 = ~1'b0 ;
  assign y1540 = n5738 ;
  assign y1541 = n6202 ;
  assign y1542 = n6218 ;
  assign y1543 = ~n6219 ;
  assign y1544 = ~n6220 ;
  assign y1545 = ~n6222 ;
  assign y1546 = ~n6224 ;
  assign y1547 = ~n6226 ;
  assign y1548 = ~n6229 ;
  assign y1549 = ~n6230 ;
  assign y1550 = n6233 ;
  assign y1551 = n6234 ;
  assign y1552 = n6238 ;
  assign y1553 = ~n6241 ;
  assign y1554 = n6247 ;
  assign y1555 = ~n6253 ;
  assign y1556 = n6256 ;
  assign y1557 = n6260 ;
  assign y1558 = ~n6261 ;
  assign y1559 = ~n6272 ;
  assign y1560 = ~n6281 ;
  assign y1561 = n6282 ;
  assign y1562 = ~n6283 ;
  assign y1563 = ~1'b0 ;
  assign y1564 = ~n6285 ;
  assign y1565 = ~n6292 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = n6299 ;
  assign y1568 = n6305 ;
  assign y1569 = ~n6308 ;
  assign y1570 = ~n6310 ;
  assign y1571 = ~1'b0 ;
  assign y1572 = n6311 ;
  assign y1573 = ~n5715 ;
  assign y1574 = ~n6312 ;
  assign y1575 = n6313 ;
  assign y1576 = n6315 ;
  assign y1577 = ~n6318 ;
  assign y1578 = ~n6322 ;
  assign y1579 = ~n3625 ;
  assign y1580 = n6325 ;
  assign y1581 = ~n6328 ;
  assign y1582 = ~n6332 ;
  assign y1583 = ~n6336 ;
  assign y1584 = n6339 ;
  assign y1585 = ~1'b0 ;
  assign y1586 = ~n6344 ;
  assign y1587 = ~1'b0 ;
  assign y1588 = ~1'b0 ;
  assign y1589 = n6350 ;
  assign y1590 = n6356 ;
  assign y1591 = n6359 ;
  assign y1592 = ~n6368 ;
  assign y1593 = ~n6372 ;
  assign y1594 = ~n6378 ;
  assign y1595 = ~n6381 ;
  assign y1596 = ~1'b0 ;
  assign y1597 = ~n6387 ;
  assign y1598 = ~n608 ;
  assign y1599 = n6389 ;
  assign y1600 = ~n6392 ;
  assign y1601 = n6396 ;
  assign y1602 = ~n6404 ;
  assign y1603 = ~n6406 ;
  assign y1604 = n6413 ;
  assign y1605 = ~n6417 ;
  assign y1606 = n6418 ;
  assign y1607 = n6420 ;
  assign y1608 = n6424 ;
  assign y1609 = ~n6427 ;
  assign y1610 = n6428 ;
  assign y1611 = ~n6433 ;
  assign y1612 = ~n6439 ;
  assign y1613 = ~1'b0 ;
  assign y1614 = n6440 ;
  assign y1615 = ~n6443 ;
  assign y1616 = ~n6445 ;
  assign y1617 = ~n6456 ;
  assign y1618 = ~n6462 ;
  assign y1619 = n6480 ;
  assign y1620 = n6481 ;
  assign y1621 = n6482 ;
  assign y1622 = n6486 ;
  assign y1623 = ~n6490 ;
  assign y1624 = ~1'b0 ;
  assign y1625 = ~1'b0 ;
  assign y1626 = n6491 ;
  assign y1627 = ~n6498 ;
  assign y1628 = n6499 ;
  assign y1629 = n6502 ;
  assign y1630 = n6504 ;
  assign y1631 = n6516 ;
  assign y1632 = ~n6517 ;
  assign y1633 = n6521 ;
  assign y1634 = n6522 ;
  assign y1635 = ~1'b0 ;
  assign y1636 = ~1'b0 ;
  assign y1637 = n6525 ;
  assign y1638 = n6539 ;
  assign y1639 = n6543 ;
  assign y1640 = n6553 ;
  assign y1641 = ~1'b0 ;
  assign y1642 = ~1'b0 ;
  assign y1643 = ~n6557 ;
  assign y1644 = ~n6561 ;
  assign y1645 = ~n6566 ;
  assign y1646 = ~1'b0 ;
  assign y1647 = ~n6569 ;
  assign y1648 = ~n6578 ;
  assign y1649 = ~n6579 ;
  assign y1650 = n6587 ;
  assign y1651 = n6602 ;
  assign y1652 = 1'b0 ;
  assign y1653 = n6607 ;
  assign y1654 = ~n6609 ;
  assign y1655 = ~n6610 ;
  assign y1656 = n6613 ;
  assign y1657 = n6618 ;
  assign y1658 = n6634 ;
  assign y1659 = n6638 ;
  assign y1660 = ~n6640 ;
  assign y1661 = ~n6643 ;
  assign y1662 = n6647 ;
  assign y1663 = ~n6652 ;
  assign y1664 = ~n6655 ;
  assign y1665 = ~n6658 ;
  assign y1666 = ~n6664 ;
  assign y1667 = ~1'b0 ;
  assign y1668 = ~n6666 ;
  assign y1669 = n6668 ;
  assign y1670 = ~1'b0 ;
  assign y1671 = ~n6674 ;
  assign y1672 = n6676 ;
  assign y1673 = ~n6681 ;
  assign y1674 = n6683 ;
  assign y1675 = n6695 ;
  assign y1676 = n6701 ;
  assign y1677 = ~n6705 ;
  assign y1678 = n6708 ;
  assign y1679 = n6721 ;
  assign y1680 = ~n6728 ;
  assign y1681 = n6729 ;
  assign y1682 = n6730 ;
  assign y1683 = n6735 ;
  assign y1684 = n6740 ;
  assign y1685 = ~n6741 ;
  assign y1686 = n6747 ;
  assign y1687 = n6750 ;
  assign y1688 = ~1'b0 ;
  assign y1689 = ~n6755 ;
  assign y1690 = ~n6756 ;
  assign y1691 = n6765 ;
  assign y1692 = ~1'b0 ;
  assign y1693 = ~n6768 ;
  assign y1694 = ~1'b0 ;
  assign y1695 = ~n6769 ;
  assign y1696 = ~n6771 ;
  assign y1697 = ~n6775 ;
  assign y1698 = n6776 ;
  assign y1699 = ~1'b0 ;
  assign y1700 = ~n6789 ;
  assign y1701 = ~n6791 ;
  assign y1702 = ~n6795 ;
  assign y1703 = ~n6799 ;
  assign y1704 = ~n6802 ;
  assign y1705 = ~n6805 ;
  assign y1706 = n6808 ;
  assign y1707 = ~n6811 ;
  assign y1708 = n6813 ;
  assign y1709 = ~1'b0 ;
  assign y1710 = ~1'b0 ;
  assign y1711 = ~n6825 ;
  assign y1712 = n6827 ;
  assign y1713 = ~1'b0 ;
  assign y1714 = ~1'b0 ;
  assign y1715 = n6828 ;
  assign y1716 = ~n6830 ;
  assign y1717 = ~n6837 ;
  assign y1718 = ~n6838 ;
  assign y1719 = n6842 ;
  assign y1720 = ~n6844 ;
  assign y1721 = n6845 ;
  assign y1722 = n6850 ;
  assign y1723 = ~n6851 ;
  assign y1724 = ~n6857 ;
  assign y1725 = ~1'b0 ;
  assign y1726 = n5176 ;
  assign y1727 = ~1'b0 ;
  assign y1728 = ~1'b0 ;
  assign y1729 = ~n6858 ;
  assign y1730 = ~n6864 ;
  assign y1731 = ~n6868 ;
  assign y1732 = n6871 ;
  assign y1733 = ~n6877 ;
  assign y1734 = n6882 ;
  assign y1735 = ~n6885 ;
  assign y1736 = ~n6896 ;
  assign y1737 = n6898 ;
  assign y1738 = n6903 ;
  assign y1739 = ~1'b0 ;
  assign y1740 = n6904 ;
  assign y1741 = n6908 ;
  assign y1742 = ~n6916 ;
  assign y1743 = n6920 ;
  assign y1744 = n6923 ;
  assign y1745 = ~n6927 ;
  assign y1746 = ~1'b0 ;
  assign y1747 = n6933 ;
  assign y1748 = n6941 ;
  assign y1749 = ~n6946 ;
  assign y1750 = n6947 ;
  assign y1751 = n6949 ;
  assign y1752 = ~1'b0 ;
  assign y1753 = ~n6959 ;
  assign y1754 = ~n6973 ;
  assign y1755 = n6974 ;
  assign y1756 = n6979 ;
  assign y1757 = n6980 ;
  assign y1758 = ~n6982 ;
  assign y1759 = ~n6986 ;
  assign y1760 = ~n7001 ;
  assign y1761 = n7006 ;
  assign y1762 = ~1'b0 ;
  assign y1763 = n7016 ;
  assign y1764 = ~n7025 ;
  assign y1765 = ~n7031 ;
  assign y1766 = ~n7033 ;
  assign y1767 = ~1'b0 ;
  assign y1768 = ~n7035 ;
  assign y1769 = ~n7040 ;
  assign y1770 = n7047 ;
  assign y1771 = ~n7051 ;
  assign y1772 = ~1'b0 ;
  assign y1773 = ~n7056 ;
  assign y1774 = ~n7058 ;
  assign y1775 = n7060 ;
  assign y1776 = n1370 ;
  assign y1777 = ~1'b0 ;
  assign y1778 = ~n7067 ;
  assign y1779 = n7078 ;
  assign y1780 = n7080 ;
  assign y1781 = ~1'b0 ;
  assign y1782 = ~n7081 ;
  assign y1783 = ~n7088 ;
  assign y1784 = ~n7092 ;
  assign y1785 = ~1'b0 ;
  assign y1786 = ~n7094 ;
  assign y1787 = ~n7100 ;
  assign y1788 = ~n7101 ;
  assign y1789 = n7102 ;
  assign y1790 = ~1'b0 ;
  assign y1791 = ~1'b0 ;
  assign y1792 = ~n7104 ;
  assign y1793 = ~n7113 ;
  assign y1794 = n7122 ;
  assign y1795 = n7130 ;
  assign y1796 = 1'b0 ;
  assign y1797 = n7134 ;
  assign y1798 = ~n7137 ;
  assign y1799 = ~n7139 ;
  assign y1800 = n7141 ;
  assign y1801 = ~n7148 ;
  assign y1802 = ~1'b0 ;
  assign y1803 = n7153 ;
  assign y1804 = n7157 ;
  assign y1805 = ~n7160 ;
  assign y1806 = n7168 ;
  assign y1807 = n7179 ;
  assign y1808 = n7181 ;
  assign y1809 = ~n7188 ;
  assign y1810 = n7191 ;
  assign y1811 = n7196 ;
  assign y1812 = n7198 ;
  assign y1813 = n7212 ;
  assign y1814 = n7220 ;
  assign y1815 = ~n7224 ;
  assign y1816 = ~n7229 ;
  assign y1817 = ~n7230 ;
  assign y1818 = ~n7233 ;
  assign y1819 = n7234 ;
  assign y1820 = ~n7246 ;
  assign y1821 = ~n7249 ;
  assign y1822 = ~n7255 ;
  assign y1823 = n7257 ;
  assign y1824 = n7259 ;
  assign y1825 = n7260 ;
  assign y1826 = ~n7261 ;
  assign y1827 = n7262 ;
  assign y1828 = ~1'b0 ;
  assign y1829 = ~n7266 ;
  assign y1830 = ~n7276 ;
  assign y1831 = n7278 ;
  assign y1832 = ~n7282 ;
  assign y1833 = ~n7284 ;
  assign y1834 = n7288 ;
  assign y1835 = ~1'b0 ;
  assign y1836 = ~n7290 ;
  assign y1837 = ~n7292 ;
  assign y1838 = n6667 ;
  assign y1839 = ~n7296 ;
  assign y1840 = ~1'b0 ;
  assign y1841 = ~n7301 ;
  assign y1842 = n7305 ;
  assign y1843 = ~n7312 ;
  assign y1844 = n7313 ;
  assign y1845 = n7316 ;
  assign y1846 = n7323 ;
  assign y1847 = n7332 ;
  assign y1848 = ~1'b0 ;
  assign y1849 = ~n7333 ;
  assign y1850 = ~n7339 ;
  assign y1851 = ~n7356 ;
  assign y1852 = ~n7359 ;
  assign y1853 = n7363 ;
  assign y1854 = n7365 ;
  assign y1855 = ~n7374 ;
  assign y1856 = ~n5548 ;
  assign y1857 = n7378 ;
  assign y1858 = ~1'b0 ;
  assign y1859 = n7385 ;
  assign y1860 = n7388 ;
  assign y1861 = ~n7392 ;
  assign y1862 = ~1'b0 ;
  assign y1863 = ~1'b0 ;
  assign y1864 = ~1'b0 ;
  assign y1865 = ~n7396 ;
  assign y1866 = n7397 ;
  assign y1867 = n7398 ;
  assign y1868 = ~n7400 ;
  assign y1869 = n7401 ;
  assign y1870 = n7402 ;
  assign y1871 = ~n7405 ;
  assign y1872 = ~n7409 ;
  assign y1873 = ~1'b0 ;
  assign y1874 = n7412 ;
  assign y1875 = ~n7413 ;
  assign y1876 = n7418 ;
  assign y1877 = n7419 ;
  assign y1878 = ~1'b0 ;
  assign y1879 = ~n7425 ;
  assign y1880 = ~1'b0 ;
  assign y1881 = n7426 ;
  assign y1882 = n7430 ;
  assign y1883 = ~1'b0 ;
  assign y1884 = n7431 ;
  assign y1885 = ~n7433 ;
  assign y1886 = n7439 ;
  assign y1887 = n7447 ;
  assign y1888 = ~n7462 ;
  assign y1889 = ~1'b0 ;
  assign y1890 = n7468 ;
  assign y1891 = ~n7469 ;
  assign y1892 = ~n7472 ;
  assign y1893 = ~1'b0 ;
  assign y1894 = ~1'b0 ;
  assign y1895 = ~n7473 ;
  assign y1896 = ~n7480 ;
  assign y1897 = ~n7485 ;
  assign y1898 = n7489 ;
  assign y1899 = n7494 ;
  assign y1900 = n7500 ;
  assign y1901 = ~n7502 ;
  assign y1902 = n7504 ;
  assign y1903 = ~n7514 ;
  assign y1904 = ~n7517 ;
  assign y1905 = ~n7520 ;
  assign y1906 = ~n7523 ;
  assign y1907 = ~1'b0 ;
  assign y1908 = n7528 ;
  assign y1909 = n7529 ;
  assign y1910 = n7533 ;
  assign y1911 = n7535 ;
  assign y1912 = n7540 ;
  assign y1913 = ~n7544 ;
  assign y1914 = n7547 ;
  assign y1915 = ~n7549 ;
  assign y1916 = ~1'b0 ;
  assign y1917 = ~n7559 ;
  assign y1918 = n7562 ;
  assign y1919 = n7566 ;
  assign y1920 = ~1'b0 ;
  assign y1921 = ~n7576 ;
  assign y1922 = n7577 ;
  assign y1923 = ~1'b0 ;
  assign y1924 = n7580 ;
  assign y1925 = n7581 ;
  assign y1926 = n7586 ;
  assign y1927 = n7587 ;
  assign y1928 = n7593 ;
  assign y1929 = n7600 ;
  assign y1930 = n7601 ;
  assign y1931 = ~1'b0 ;
  assign y1932 = ~n7604 ;
  assign y1933 = ~1'b0 ;
  assign y1934 = ~n7608 ;
  assign y1935 = n7622 ;
  assign y1936 = n7623 ;
  assign y1937 = n2317 ;
  assign y1938 = ~n7626 ;
  assign y1939 = ~n7629 ;
  assign y1940 = n7632 ;
  assign y1941 = n7639 ;
  assign y1942 = n7648 ;
  assign y1943 = ~1'b0 ;
  assign y1944 = ~1'b0 ;
  assign y1945 = ~n7651 ;
  assign y1946 = ~n7652 ;
  assign y1947 = ~n7654 ;
  assign y1948 = n7662 ;
  assign y1949 = ~1'b0 ;
  assign y1950 = ~1'b0 ;
  assign y1951 = ~n7667 ;
  assign y1952 = ~n7678 ;
  assign y1953 = n7682 ;
  assign y1954 = ~1'b0 ;
  assign y1955 = ~1'b0 ;
  assign y1956 = ~n7684 ;
  assign y1957 = n7686 ;
  assign y1958 = ~n7690 ;
  assign y1959 = n7694 ;
  assign y1960 = ~n1028 ;
  assign y1961 = ~n7703 ;
  assign y1962 = n7712 ;
  assign y1963 = n7715 ;
  assign y1964 = n7716 ;
  assign y1965 = n7735 ;
  assign y1966 = ~1'b0 ;
  assign y1967 = n7738 ;
  assign y1968 = ~n7744 ;
  assign y1969 = ~n7764 ;
  assign y1970 = ~1'b0 ;
  assign y1971 = n7769 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = n7776 ;
  assign y1974 = ~n7786 ;
  assign y1975 = n7792 ;
  assign y1976 = ~n7793 ;
  assign y1977 = n7798 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = ~1'b0 ;
  assign y1980 = ~n7799 ;
  assign y1981 = n7800 ;
  assign y1982 = ~n7801 ;
  assign y1983 = ~n7803 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = n7811 ;
  assign y1986 = n7817 ;
  assign y1987 = ~n7819 ;
  assign y1988 = ~n7830 ;
  assign y1989 = n7833 ;
  assign y1990 = ~n7835 ;
  assign y1991 = ~1'b0 ;
  assign y1992 = ~n7837 ;
  assign y1993 = ~n7840 ;
  assign y1994 = ~1'b0 ;
  assign y1995 = ~n7847 ;
  assign y1996 = ~n7849 ;
  assign y1997 = ~n7850 ;
  assign y1998 = ~n7856 ;
  assign y1999 = ~n7857 ;
  assign y2000 = n7858 ;
  assign y2001 = ~1'b0 ;
  assign y2002 = ~n7863 ;
  assign y2003 = ~n7864 ;
  assign y2004 = ~n7865 ;
  assign y2005 = ~n7874 ;
  assign y2006 = ~1'b0 ;
  assign y2007 = ~n7876 ;
  assign y2008 = ~1'b0 ;
  assign y2009 = n7879 ;
  assign y2010 = ~1'b0 ;
  assign y2011 = ~n7882 ;
  assign y2012 = n7885 ;
  assign y2013 = ~n7886 ;
  assign y2014 = ~n7888 ;
  assign y2015 = n7890 ;
  assign y2016 = ~1'b0 ;
  assign y2017 = ~n7897 ;
  assign y2018 = ~n7904 ;
  assign y2019 = n7907 ;
  assign y2020 = ~n7914 ;
  assign y2021 = ~1'b0 ;
  assign y2022 = n7919 ;
  assign y2023 = n7923 ;
  assign y2024 = ~n7936 ;
  assign y2025 = n7944 ;
  assign y2026 = n7947 ;
  assign y2027 = ~n7950 ;
  assign y2028 = n7952 ;
  assign y2029 = n7953 ;
  assign y2030 = ~n7956 ;
  assign y2031 = n7962 ;
  assign y2032 = ~1'b0 ;
  assign y2033 = ~n7970 ;
  assign y2034 = n7972 ;
  assign y2035 = n7974 ;
  assign y2036 = n7977 ;
  assign y2037 = ~n7978 ;
  assign y2038 = n7985 ;
  assign y2039 = n7987 ;
  assign y2040 = ~n7992 ;
  assign y2041 = ~n7993 ;
  assign y2042 = n7995 ;
  assign y2043 = ~n8006 ;
  assign y2044 = ~n8008 ;
  assign y2045 = n8019 ;
  assign y2046 = ~n8023 ;
  assign y2047 = n8025 ;
  assign y2048 = n8033 ;
  assign y2049 = ~n8034 ;
  assign y2050 = n8035 ;
  assign y2051 = ~1'b0 ;
  assign y2052 = n8036 ;
  assign y2053 = ~n8038 ;
  assign y2054 = ~n8039 ;
  assign y2055 = n8045 ;
  assign y2056 = ~n8049 ;
  assign y2057 = n8056 ;
  assign y2058 = n8057 ;
  assign y2059 = ~1'b0 ;
  assign y2060 = ~n8074 ;
  assign y2061 = n8078 ;
  assign y2062 = ~n8080 ;
  assign y2063 = ~n8083 ;
  assign y2064 = ~n8090 ;
  assign y2065 = n8097 ;
  assign y2066 = ~n8099 ;
  assign y2067 = n8101 ;
  assign y2068 = ~n8104 ;
  assign y2069 = n8106 ;
  assign y2070 = ~n8107 ;
  assign y2071 = n8110 ;
  assign y2072 = n8114 ;
  assign y2073 = ~n8118 ;
  assign y2074 = n8123 ;
  assign y2075 = ~n8127 ;
  assign y2076 = n8133 ;
  assign y2077 = n8134 ;
  assign y2078 = ~n7726 ;
  assign y2079 = n8135 ;
  assign y2080 = ~n8140 ;
  assign y2081 = n8141 ;
  assign y2082 = ~n8150 ;
  assign y2083 = ~n8154 ;
  assign y2084 = ~n8160 ;
  assign y2085 = ~n8171 ;
  assign y2086 = n8183 ;
  assign y2087 = n8184 ;
  assign y2088 = ~n8185 ;
  assign y2089 = ~n8189 ;
  assign y2090 = ~n8196 ;
  assign y2091 = ~n8201 ;
  assign y2092 = n8203 ;
  assign y2093 = n8205 ;
  assign y2094 = ~n8211 ;
  assign y2095 = ~n8214 ;
  assign y2096 = ~n8226 ;
  assign y2097 = n8233 ;
  assign y2098 = ~n8234 ;
  assign y2099 = ~n8237 ;
  assign y2100 = n8243 ;
  assign y2101 = ~n8251 ;
  assign y2102 = n8260 ;
  assign y2103 = ~1'b0 ;
  assign y2104 = n8278 ;
  assign y2105 = n8282 ;
  assign y2106 = ~n8287 ;
  assign y2107 = ~n8293 ;
  assign y2108 = ~1'b0 ;
  assign y2109 = n8301 ;
  assign y2110 = ~n8302 ;
  assign y2111 = n8306 ;
  assign y2112 = n8308 ;
  assign y2113 = n8318 ;
  assign y2114 = n8328 ;
  assign y2115 = 1'b0 ;
  assign y2116 = n8329 ;
  assign y2117 = ~n8332 ;
  assign y2118 = n8345 ;
  assign y2119 = n8346 ;
  assign y2120 = ~1'b0 ;
  assign y2121 = ~1'b0 ;
  assign y2122 = n8347 ;
  assign y2123 = ~n8351 ;
  assign y2124 = ~n8363 ;
  assign y2125 = ~n8368 ;
  assign y2126 = ~n8372 ;
  assign y2127 = ~n8375 ;
  assign y2128 = ~n8380 ;
  assign y2129 = ~n8384 ;
  assign y2130 = n8394 ;
  assign y2131 = n8397 ;
  assign y2132 = ~n8402 ;
  assign y2133 = ~n8406 ;
  assign y2134 = ~n8411 ;
  assign y2135 = ~n8414 ;
  assign y2136 = ~1'b0 ;
  assign y2137 = ~n8418 ;
  assign y2138 = ~n8422 ;
  assign y2139 = ~n8424 ;
  assign y2140 = ~n8427 ;
  assign y2141 = ~n8428 ;
  assign y2142 = ~n8432 ;
  assign y2143 = n8436 ;
  assign y2144 = n8440 ;
  assign y2145 = ~n4373 ;
  assign y2146 = n8443 ;
  assign y2147 = ~1'b0 ;
  assign y2148 = n8449 ;
  assign y2149 = n1239 ;
  assign y2150 = ~n8452 ;
  assign y2151 = n8456 ;
  assign y2152 = ~n8457 ;
  assign y2153 = ~n8460 ;
  assign y2154 = n8462 ;
  assign y2155 = ~1'b0 ;
  assign y2156 = n8470 ;
  assign y2157 = ~n8476 ;
  assign y2158 = ~n8477 ;
  assign y2159 = n8491 ;
  assign y2160 = ~n8493 ;
  assign y2161 = ~n8494 ;
  assign y2162 = ~1'b0 ;
  assign y2163 = ~n8495 ;
  assign y2164 = n8499 ;
  assign y2165 = ~1'b0 ;
  assign y2166 = ~n8506 ;
  assign y2167 = ~n8511 ;
  assign y2168 = n8513 ;
  assign y2169 = ~1'b0 ;
  assign y2170 = ~1'b0 ;
  assign y2171 = ~n8519 ;
  assign y2172 = n8525 ;
  assign y2173 = ~n8529 ;
  assign y2174 = n8531 ;
  assign y2175 = n8534 ;
  assign y2176 = ~1'b0 ;
  assign y2177 = ~n8548 ;
  assign y2178 = n8552 ;
  assign y2179 = n8553 ;
  assign y2180 = n8570 ;
  assign y2181 = n8572 ;
  assign y2182 = ~n8573 ;
  assign y2183 = ~n8575 ;
  assign y2184 = ~n8577 ;
  assign y2185 = ~n8582 ;
  assign y2186 = ~1'b0 ;
  assign y2187 = n8591 ;
  assign y2188 = ~1'b0 ;
  assign y2189 = n8593 ;
  assign y2190 = ~n8599 ;
  assign y2191 = ~n8603 ;
  assign y2192 = n8605 ;
  assign y2193 = n8614 ;
  assign y2194 = ~n8615 ;
  assign y2195 = ~n8625 ;
  assign y2196 = ~1'b0 ;
  assign y2197 = ~n8628 ;
  assign y2198 = n8632 ;
  assign y2199 = ~n8642 ;
  assign y2200 = ~1'b0 ;
  assign y2201 = n8645 ;
  assign y2202 = ~n8648 ;
  assign y2203 = n8653 ;
  assign y2204 = n8654 ;
  assign y2205 = n8656 ;
  assign y2206 = ~1'b0 ;
  assign y2207 = ~n8663 ;
  assign y2208 = ~n8664 ;
  assign y2209 = n8666 ;
  assign y2210 = 1'b0 ;
  assign y2211 = ~1'b0 ;
  assign y2212 = n8671 ;
  assign y2213 = ~n8675 ;
  assign y2214 = n8678 ;
  assign y2215 = ~n8679 ;
  assign y2216 = n8681 ;
  assign y2217 = ~n8684 ;
  assign y2218 = n8688 ;
  assign y2219 = ~n8692 ;
  assign y2220 = n8698 ;
  assign y2221 = n8702 ;
  assign y2222 = n8705 ;
  assign y2223 = n8706 ;
  assign y2224 = n8707 ;
  assign y2225 = ~n8708 ;
  assign y2226 = n8711 ;
  assign y2227 = n8713 ;
  assign y2228 = n8715 ;
  assign y2229 = ~n8716 ;
  assign y2230 = n8720 ;
  assign y2231 = n8725 ;
  assign y2232 = ~n8729 ;
  assign y2233 = ~n8741 ;
  assign y2234 = ~n8747 ;
  assign y2235 = n8753 ;
  assign y2236 = ~n8762 ;
  assign y2237 = ~1'b0 ;
  assign y2238 = ~1'b0 ;
  assign y2239 = ~n8772 ;
  assign y2240 = ~n8774 ;
  assign y2241 = n8777 ;
  assign y2242 = ~1'b0 ;
  assign y2243 = ~n8783 ;
  assign y2244 = ~n8784 ;
  assign y2245 = ~n8787 ;
  assign y2246 = n8794 ;
  assign y2247 = ~1'b0 ;
  assign y2248 = n8795 ;
  assign y2249 = ~n8811 ;
  assign y2250 = n8814 ;
  assign y2251 = n8817 ;
  assign y2252 = n8830 ;
  assign y2253 = ~n8855 ;
  assign y2254 = ~n8856 ;
  assign y2255 = n8863 ;
  assign y2256 = ~1'b0 ;
  assign y2257 = ~n8871 ;
  assign y2258 = ~n8885 ;
  assign y2259 = n8888 ;
  assign y2260 = ~n8890 ;
  assign y2261 = n8892 ;
  assign y2262 = ~n8894 ;
  assign y2263 = ~n8899 ;
  assign y2264 = ~n8902 ;
  assign y2265 = ~n8923 ;
  assign y2266 = n8924 ;
  assign y2267 = ~n8925 ;
  assign y2268 = n8928 ;
  assign y2269 = n8931 ;
  assign y2270 = ~n8932 ;
  assign y2271 = ~1'b0 ;
  assign y2272 = ~n8933 ;
  assign y2273 = ~n8939 ;
  assign y2274 = ~n8941 ;
  assign y2275 = ~1'b0 ;
  assign y2276 = n8946 ;
  assign y2277 = n1708 ;
  assign y2278 = ~n8951 ;
  assign y2279 = n8955 ;
  assign y2280 = ~n8956 ;
  assign y2281 = n8975 ;
  assign y2282 = ~n8991 ;
  assign y2283 = ~n8997 ;
  assign y2284 = ~1'b0 ;
  assign y2285 = ~1'b0 ;
  assign y2286 = ~1'b0 ;
  assign y2287 = ~n8998 ;
  assign y2288 = ~n8999 ;
  assign y2289 = ~n9000 ;
  assign y2290 = ~n3894 ;
  assign y2291 = ~1'b0 ;
  assign y2292 = ~n3177 ;
  assign y2293 = n9001 ;
  assign y2294 = n9002 ;
  assign y2295 = ~n9003 ;
  assign y2296 = n9009 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = ~n9011 ;
  assign y2299 = n9029 ;
  assign y2300 = ~n9033 ;
  assign y2301 = n9036 ;
  assign y2302 = n9044 ;
  assign y2303 = ~1'b0 ;
  assign y2304 = ~n9045 ;
  assign y2305 = n3605 ;
  assign y2306 = ~n9049 ;
  assign y2307 = ~n9050 ;
  assign y2308 = n9051 ;
  assign y2309 = n9052 ;
  assign y2310 = ~1'b0 ;
  assign y2311 = n9062 ;
  assign y2312 = ~n9070 ;
  assign y2313 = ~n9071 ;
  assign y2314 = n9074 ;
  assign y2315 = n9076 ;
  assign y2316 = ~n9080 ;
  assign y2317 = ~n9082 ;
  assign y2318 = n9091 ;
  assign y2319 = n9101 ;
  assign y2320 = ~n9103 ;
  assign y2321 = ~n9104 ;
  assign y2322 = ~n9113 ;
  assign y2323 = n9115 ;
  assign y2324 = ~n9116 ;
  assign y2325 = ~n9118 ;
  assign y2326 = n9120 ;
  assign y2327 = ~1'b0 ;
  assign y2328 = n9122 ;
  assign y2329 = ~n9124 ;
  assign y2330 = ~n9143 ;
  assign y2331 = ~1'b0 ;
  assign y2332 = ~n9146 ;
  assign y2333 = ~1'b0 ;
  assign y2334 = ~n9148 ;
  assign y2335 = ~n2006 ;
  assign y2336 = ~n9149 ;
  assign y2337 = ~n9150 ;
  assign y2338 = ~n9156 ;
  assign y2339 = ~n9164 ;
  assign y2340 = n9166 ;
  assign y2341 = ~n9172 ;
  assign y2342 = n9173 ;
  assign y2343 = n9176 ;
  assign y2344 = ~1'b0 ;
  assign y2345 = ~n9179 ;
  assign y2346 = n9180 ;
  assign y2347 = ~n9194 ;
  assign y2348 = n9203 ;
  assign y2349 = ~n9206 ;
  assign y2350 = n9217 ;
  assign y2351 = ~n9219 ;
  assign y2352 = ~n9221 ;
  assign y2353 = n9225 ;
  assign y2354 = n9226 ;
  assign y2355 = ~n9227 ;
  assign y2356 = ~n9234 ;
  assign y2357 = ~n9244 ;
  assign y2358 = n9246 ;
  assign y2359 = n9252 ;
  assign y2360 = ~n9253 ;
  assign y2361 = n9254 ;
  assign y2362 = n9256 ;
  assign y2363 = ~n9260 ;
  assign y2364 = ~n9263 ;
  assign y2365 = ~n9269 ;
  assign y2366 = n9270 ;
  assign y2367 = n9272 ;
  assign y2368 = n9276 ;
  assign y2369 = n9287 ;
  assign y2370 = n9292 ;
  assign y2371 = ~n9296 ;
  assign y2372 = n9298 ;
  assign y2373 = ~n9303 ;
  assign y2374 = ~n9306 ;
  assign y2375 = n9313 ;
  assign y2376 = n9317 ;
  assign y2377 = ~n9318 ;
  assign y2378 = ~1'b0 ;
  assign y2379 = ~n9322 ;
  assign y2380 = ~n9323 ;
  assign y2381 = ~1'b0 ;
  assign y2382 = n9329 ;
  assign y2383 = n9337 ;
  assign y2384 = ~n9347 ;
  assign y2385 = ~1'b0 ;
  assign y2386 = ~n9354 ;
  assign y2387 = ~1'b0 ;
  assign y2388 = n9358 ;
  assign y2389 = n9362 ;
  assign y2390 = n9370 ;
  assign y2391 = n9371 ;
  assign y2392 = n9374 ;
  assign y2393 = ~n9378 ;
  assign y2394 = ~1'b0 ;
  assign y2395 = n9383 ;
  assign y2396 = ~n9391 ;
  assign y2397 = ~n9392 ;
  assign y2398 = n9397 ;
  assign y2399 = n9401 ;
  assign y2400 = ~n9402 ;
  assign y2401 = ~1'b0 ;
  assign y2402 = n9413 ;
  assign y2403 = ~1'b0 ;
  assign y2404 = n9414 ;
  assign y2405 = ~n9418 ;
  assign y2406 = ~n9420 ;
  assign y2407 = ~n9424 ;
  assign y2408 = ~n9425 ;
  assign y2409 = ~n9426 ;
  assign y2410 = ~n9427 ;
  assign y2411 = ~n9429 ;
  assign y2412 = n9432 ;
  assign y2413 = ~n9449 ;
  assign y2414 = ~1'b0 ;
  assign y2415 = n9450 ;
  assign y2416 = n9456 ;
  assign y2417 = n9459 ;
  assign y2418 = ~1'b0 ;
  assign y2419 = n9463 ;
  assign y2420 = ~n9464 ;
  assign y2421 = ~1'b0 ;
  assign y2422 = n9466 ;
  assign y2423 = n9474 ;
  assign y2424 = ~n9475 ;
  assign y2425 = ~n9481 ;
  assign y2426 = ~n9498 ;
  assign y2427 = ~n9499 ;
  assign y2428 = n9500 ;
  assign y2429 = n9505 ;
  assign y2430 = n9508 ;
  assign y2431 = n9512 ;
  assign y2432 = ~n9515 ;
  assign y2433 = n9518 ;
  assign y2434 = ~n9522 ;
  assign y2435 = ~n9524 ;
  assign y2436 = ~n9525 ;
  assign y2437 = ~n9528 ;
  assign y2438 = ~n9530 ;
  assign y2439 = n4680 ;
  assign y2440 = ~n9533 ;
  assign y2441 = ~n9538 ;
  assign y2442 = ~n9539 ;
  assign y2443 = ~n9549 ;
  assign y2444 = ~1'b0 ;
  assign y2445 = ~n9563 ;
  assign y2446 = ~n9564 ;
  assign y2447 = ~n9568 ;
  assign y2448 = ~1'b0 ;
  assign y2449 = ~n9574 ;
  assign y2450 = n9576 ;
  assign y2451 = ~n9579 ;
  assign y2452 = ~n9587 ;
  assign y2453 = n9596 ;
  assign y2454 = ~1'b0 ;
  assign y2455 = ~n9602 ;
  assign y2456 = ~n9607 ;
  assign y2457 = n9608 ;
  assign y2458 = ~n9609 ;
  assign y2459 = ~n9611 ;
  assign y2460 = ~1'b0 ;
  assign y2461 = n9613 ;
  assign y2462 = n9617 ;
  assign y2463 = ~n9621 ;
  assign y2464 = ~n9624 ;
  assign y2465 = ~n9626 ;
  assign y2466 = n9628 ;
  assign y2467 = n9629 ;
  assign y2468 = ~1'b0 ;
  assign y2469 = ~n9632 ;
  assign y2470 = n9636 ;
  assign y2471 = n9639 ;
  assign y2472 = ~n9642 ;
  assign y2473 = n9652 ;
  assign y2474 = ~n9656 ;
  assign y2475 = ~n9658 ;
  assign y2476 = n9659 ;
  assign y2477 = ~1'b0 ;
  assign y2478 = ~n1666 ;
  assign y2479 = n9667 ;
  assign y2480 = n9669 ;
  assign y2481 = ~n9674 ;
  assign y2482 = ~n9681 ;
  assign y2483 = ~n9682 ;
  assign y2484 = n9689 ;
  assign y2485 = n9693 ;
  assign y2486 = n9706 ;
  assign y2487 = n9708 ;
  assign y2488 = n9725 ;
  assign y2489 = n9734 ;
  assign y2490 = ~n9744 ;
  assign y2491 = n9749 ;
  assign y2492 = ~1'b0 ;
  assign y2493 = n9754 ;
  assign y2494 = ~n9757 ;
  assign y2495 = n9762 ;
  assign y2496 = ~n9777 ;
  assign y2497 = ~n9786 ;
  assign y2498 = n9788 ;
  assign y2499 = ~n9791 ;
  assign y2500 = ~n9794 ;
  assign y2501 = n9795 ;
  assign y2502 = n9799 ;
  assign y2503 = n9801 ;
  assign y2504 = n9805 ;
  assign y2505 = n9807 ;
  assign y2506 = n9809 ;
  assign y2507 = ~n9812 ;
  assign y2508 = ~1'b0 ;
  assign y2509 = ~n9814 ;
  assign y2510 = n9815 ;
  assign y2511 = n9817 ;
  assign y2512 = n9820 ;
  assign y2513 = ~1'b0 ;
  assign y2514 = ~n9824 ;
  assign y2515 = n9830 ;
  assign y2516 = n9833 ;
  assign y2517 = n9852 ;
  assign y2518 = ~n9853 ;
  assign y2519 = ~n9858 ;
  assign y2520 = n9864 ;
  assign y2521 = n9868 ;
  assign y2522 = ~n9876 ;
  assign y2523 = n9877 ;
  assign y2524 = n9901 ;
  assign y2525 = ~n9902 ;
  assign y2526 = n9904 ;
  assign y2527 = n9906 ;
  assign y2528 = ~n9908 ;
  assign y2529 = n9911 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = ~n9917 ;
  assign y2532 = ~1'b0 ;
  assign y2533 = n9925 ;
  assign y2534 = n9927 ;
  assign y2535 = ~n9931 ;
  assign y2536 = n9934 ;
  assign y2537 = ~n9935 ;
  assign y2538 = n9941 ;
  assign y2539 = n9953 ;
  assign y2540 = ~1'b0 ;
  assign y2541 = n9958 ;
  assign y2542 = n9962 ;
  assign y2543 = n9967 ;
  assign y2544 = n9968 ;
  assign y2545 = ~n9982 ;
  assign y2546 = ~n320 ;
  assign y2547 = ~n9986 ;
  assign y2548 = ~1'b0 ;
  assign y2549 = n9993 ;
  assign y2550 = n9998 ;
  assign y2551 = ~n9999 ;
  assign y2552 = n10000 ;
  assign y2553 = ~n10011 ;
  assign y2554 = n10015 ;
  assign y2555 = n10017 ;
  assign y2556 = ~n10027 ;
  assign y2557 = ~n10033 ;
  assign y2558 = ~n10036 ;
  assign y2559 = n10047 ;
  assign y2560 = n10019 ;
  assign y2561 = n10059 ;
  assign y2562 = ~n10060 ;
  assign y2563 = n10061 ;
  assign y2564 = n10076 ;
  assign y2565 = ~n10087 ;
  assign y2566 = ~n10088 ;
  assign y2567 = n10089 ;
  assign y2568 = n10091 ;
  assign y2569 = ~1'b0 ;
  assign y2570 = n10096 ;
  assign y2571 = ~n10098 ;
  assign y2572 = ~n10100 ;
  assign y2573 = n10105 ;
  assign y2574 = ~1'b0 ;
  assign y2575 = n10106 ;
  assign y2576 = ~n10109 ;
  assign y2577 = ~n10111 ;
  assign y2578 = ~n10112 ;
  assign y2579 = ~n10114 ;
  assign y2580 = ~n10120 ;
  assign y2581 = ~n10121 ;
  assign y2582 = n10122 ;
  assign y2583 = ~n10123 ;
  assign y2584 = ~1'b0 ;
  assign y2585 = ~1'b0 ;
  assign y2586 = ~n10125 ;
  assign y2587 = ~n10138 ;
  assign y2588 = ~n10144 ;
  assign y2589 = ~n10150 ;
  assign y2590 = n10154 ;
  assign y2591 = ~n10156 ;
  assign y2592 = ~n10167 ;
  assign y2593 = ~1'b0 ;
  assign y2594 = n10172 ;
  assign y2595 = ~n10174 ;
  assign y2596 = ~n10179 ;
  assign y2597 = ~n10181 ;
  assign y2598 = ~1'b0 ;
  assign y2599 = n10182 ;
  assign y2600 = n10186 ;
  assign y2601 = ~n10190 ;
  assign y2602 = ~n10193 ;
  assign y2603 = ~n10200 ;
  assign y2604 = ~n10202 ;
  assign y2605 = n10210 ;
  assign y2606 = ~n10219 ;
  assign y2607 = n10220 ;
  assign y2608 = n10221 ;
  assign y2609 = n10224 ;
  assign y2610 = ~n10230 ;
  assign y2611 = ~n10233 ;
  assign y2612 = ~n10235 ;
  assign y2613 = ~n10237 ;
  assign y2614 = ~x229 ;
  assign y2615 = n10242 ;
  assign y2616 = ~1'b0 ;
  assign y2617 = n10243 ;
  assign y2618 = ~n10251 ;
  assign y2619 = ~1'b0 ;
  assign y2620 = ~n10269 ;
  assign y2621 = ~1'b0 ;
  assign y2622 = n10275 ;
  assign y2623 = n10280 ;
  assign y2624 = ~n10283 ;
  assign y2625 = n10286 ;
  assign y2626 = ~n5140 ;
  assign y2627 = n10290 ;
  assign y2628 = ~1'b0 ;
  assign y2629 = ~n10301 ;
  assign y2630 = ~1'b0 ;
  assign y2631 = ~1'b0 ;
  assign y2632 = ~n10305 ;
  assign y2633 = n10307 ;
  assign y2634 = n10309 ;
  assign y2635 = n10311 ;
  assign y2636 = n10312 ;
  assign y2637 = n10316 ;
  assign y2638 = n10318 ;
  assign y2639 = n10322 ;
  assign y2640 = n10323 ;
  assign y2641 = ~n10324 ;
  assign y2642 = n10326 ;
  assign y2643 = ~n8561 ;
  assign y2644 = ~n10048 ;
  assign y2645 = n10328 ;
  assign y2646 = ~n10331 ;
  assign y2647 = ~n10332 ;
  assign y2648 = n10333 ;
  assign y2649 = ~n10340 ;
  assign y2650 = n10348 ;
  assign y2651 = ~n10361 ;
  assign y2652 = ~n10366 ;
  assign y2653 = ~n10374 ;
  assign y2654 = ~n10376 ;
  assign y2655 = n10382 ;
  assign y2656 = n10390 ;
  assign y2657 = ~1'b0 ;
  assign y2658 = n10393 ;
  assign y2659 = ~n10397 ;
  assign y2660 = n1462 ;
  assign y2661 = ~n10404 ;
  assign y2662 = n10406 ;
  assign y2663 = ~n10409 ;
  assign y2664 = ~n10420 ;
  assign y2665 = n10421 ;
  assign y2666 = n10429 ;
  assign y2667 = ~n10430 ;
  assign y2668 = n10436 ;
  assign y2669 = n10439 ;
  assign y2670 = ~1'b0 ;
  assign y2671 = ~n10444 ;
  assign y2672 = ~n10451 ;
  assign y2673 = ~1'b0 ;
  assign y2674 = ~n10459 ;
  assign y2675 = n10474 ;
  assign y2676 = ~1'b0 ;
  assign y2677 = ~n10484 ;
  assign y2678 = n10487 ;
  assign y2679 = ~n10492 ;
  assign y2680 = ~n10498 ;
  assign y2681 = ~1'b0 ;
  assign y2682 = ~1'b0 ;
  assign y2683 = n10501 ;
  assign y2684 = n10511 ;
  assign y2685 = n10516 ;
  assign y2686 = n10518 ;
  assign y2687 = n10523 ;
  assign y2688 = n10525 ;
  assign y2689 = n10537 ;
  assign y2690 = ~n10540 ;
  assign y2691 = n10543 ;
  assign y2692 = ~n10545 ;
  assign y2693 = ~1'b0 ;
  assign y2694 = ~n10558 ;
  assign y2695 = n10559 ;
  assign y2696 = n10565 ;
  assign y2697 = n10569 ;
  assign y2698 = n10572 ;
  assign y2699 = ~n10580 ;
  assign y2700 = ~n10590 ;
  assign y2701 = ~n10593 ;
  assign y2702 = ~n10594 ;
  assign y2703 = ~1'b0 ;
  assign y2704 = ~n10598 ;
  assign y2705 = n10600 ;
  assign y2706 = n10602 ;
  assign y2707 = ~n10607 ;
  assign y2708 = ~1'b0 ;
  assign y2709 = ~n10610 ;
  assign y2710 = n10611 ;
  assign y2711 = 1'b0 ;
  assign y2712 = n10620 ;
  assign y2713 = ~n10626 ;
  assign y2714 = n10629 ;
  assign y2715 = n10633 ;
  assign y2716 = n10635 ;
  assign y2717 = n10645 ;
  assign y2718 = n10652 ;
  assign y2719 = ~n10658 ;
  assign y2720 = ~1'b0 ;
  assign y2721 = ~n10659 ;
  assign y2722 = ~n10660 ;
  assign y2723 = ~n10670 ;
  assign y2724 = n10676 ;
  assign y2725 = ~1'b0 ;
  assign y2726 = ~n10682 ;
  assign y2727 = ~n10683 ;
  assign y2728 = ~n10684 ;
  assign y2729 = n10691 ;
  assign y2730 = ~n10693 ;
  assign y2731 = ~n10708 ;
  assign y2732 = ~1'b0 ;
  assign y2733 = 1'b0 ;
  assign y2734 = n10716 ;
  assign y2735 = n10718 ;
  assign y2736 = n10723 ;
  assign y2737 = n10725 ;
  assign y2738 = ~n10728 ;
  assign y2739 = ~1'b0 ;
  assign y2740 = ~1'b0 ;
  assign y2741 = ~n10730 ;
  assign y2742 = ~n10733 ;
  assign y2743 = n10735 ;
  assign y2744 = n10739 ;
  assign y2745 = ~n10763 ;
  assign y2746 = n10768 ;
  assign y2747 = ~n10782 ;
  assign y2748 = ~n10786 ;
  assign y2749 = n10788 ;
  assign y2750 = ~n10794 ;
  assign y2751 = ~n10797 ;
  assign y2752 = n10799 ;
  assign y2753 = n10803 ;
  assign y2754 = n10807 ;
  assign y2755 = ~1'b0 ;
  assign y2756 = ~n10809 ;
  assign y2757 = ~n10810 ;
  assign y2758 = n10811 ;
  assign y2759 = ~n10829 ;
  assign y2760 = n10835 ;
  assign y2761 = ~n10842 ;
  assign y2762 = n304 ;
  assign y2763 = ~n10843 ;
  assign y2764 = ~n10858 ;
  assign y2765 = n10863 ;
  assign y2766 = ~n10864 ;
  assign y2767 = n10867 ;
  assign y2768 = ~n10873 ;
  assign y2769 = n10874 ;
  assign y2770 = n10875 ;
  assign y2771 = ~n10877 ;
  assign y2772 = n10883 ;
  assign y2773 = n10889 ;
  assign y2774 = n10890 ;
  assign y2775 = n10891 ;
  assign y2776 = ~n10892 ;
  assign y2777 = n10893 ;
  assign y2778 = n10895 ;
  assign y2779 = ~1'b0 ;
  assign y2780 = n10903 ;
  assign y2781 = ~1'b0 ;
  assign y2782 = n10906 ;
  assign y2783 = n10908 ;
  assign y2784 = n10909 ;
  assign y2785 = n10916 ;
  assign y2786 = ~n10922 ;
  assign y2787 = ~n10933 ;
  assign y2788 = ~n10937 ;
  assign y2789 = ~n10943 ;
  assign y2790 = n10948 ;
  assign y2791 = n10949 ;
  assign y2792 = n10951 ;
  assign y2793 = ~n10953 ;
  assign y2794 = ~n10957 ;
  assign y2795 = ~1'b0 ;
  assign y2796 = ~1'b0 ;
  assign y2797 = ~n10959 ;
  assign y2798 = ~n10960 ;
  assign y2799 = ~n10963 ;
  assign y2800 = ~1'b0 ;
  assign y2801 = n10966 ;
  assign y2802 = n10971 ;
  assign y2803 = n10975 ;
  assign y2804 = n10988 ;
  assign y2805 = n10990 ;
  assign y2806 = ~1'b0 ;
  assign y2807 = ~n10996 ;
  assign y2808 = ~1'b0 ;
  assign y2809 = n10999 ;
  assign y2810 = ~n11003 ;
  assign y2811 = ~n11004 ;
  assign y2812 = n11006 ;
  assign y2813 = n11013 ;
  assign y2814 = n11015 ;
  assign y2815 = ~n11017 ;
  assign y2816 = n11020 ;
  assign y2817 = ~n11021 ;
  assign y2818 = n11024 ;
  assign y2819 = ~1'b0 ;
  assign y2820 = ~n11025 ;
  assign y2821 = n7772 ;
  assign y2822 = ~n11026 ;
  assign y2823 = n11029 ;
  assign y2824 = n11037 ;
  assign y2825 = ~1'b0 ;
  assign y2826 = ~n11039 ;
  assign y2827 = ~n11040 ;
  assign y2828 = ~1'b0 ;
  assign y2829 = ~1'b0 ;
  assign y2830 = ~n11045 ;
  assign y2831 = n11054 ;
  assign y2832 = n11057 ;
  assign y2833 = ~1'b0 ;
  assign y2834 = ~1'b0 ;
  assign y2835 = ~1'b0 ;
  assign y2836 = ~n11069 ;
  assign y2837 = ~1'b0 ;
  assign y2838 = ~n11075 ;
  assign y2839 = ~1'b0 ;
  assign y2840 = n11080 ;
  assign y2841 = n11084 ;
  assign y2842 = n11092 ;
  assign y2843 = ~n11102 ;
  assign y2844 = ~n11104 ;
  assign y2845 = ~n11109 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = ~n11113 ;
  assign y2848 = ~n11114 ;
  assign y2849 = ~1'b0 ;
  assign y2850 = n11119 ;
  assign y2851 = ~1'b0 ;
  assign y2852 = ~n11125 ;
  assign y2853 = ~1'b0 ;
  assign y2854 = n11127 ;
  assign y2855 = ~n11128 ;
  assign y2856 = ~n11132 ;
  assign y2857 = ~n11134 ;
  assign y2858 = ~n11136 ;
  assign y2859 = n11150 ;
  assign y2860 = n11154 ;
  assign y2861 = ~1'b0 ;
  assign y2862 = n11162 ;
  assign y2863 = ~1'b0 ;
  assign y2864 = ~n11164 ;
  assign y2865 = n11174 ;
  assign y2866 = ~n11177 ;
  assign y2867 = ~1'b0 ;
  assign y2868 = ~n11186 ;
  assign y2869 = n11192 ;
  assign y2870 = ~n11200 ;
  assign y2871 = n11201 ;
  assign y2872 = ~n11203 ;
  assign y2873 = n11208 ;
  assign y2874 = ~n11210 ;
  assign y2875 = ~n11215 ;
  assign y2876 = ~n11225 ;
  assign y2877 = ~1'b0 ;
  assign y2878 = ~n11239 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = ~1'b0 ;
  assign y2881 = n11247 ;
  assign y2882 = n11248 ;
  assign y2883 = ~1'b0 ;
  assign y2884 = n11250 ;
  assign y2885 = ~n11254 ;
  assign y2886 = n11256 ;
  assign y2887 = n9917 ;
  assign y2888 = ~n11265 ;
  assign y2889 = n11268 ;
  assign y2890 = n11270 ;
  assign y2891 = ~n11274 ;
  assign y2892 = n11280 ;
  assign y2893 = n11289 ;
  assign y2894 = n11290 ;
  assign y2895 = ~n11296 ;
  assign y2896 = ~n11299 ;
  assign y2897 = n11304 ;
  assign y2898 = n11306 ;
  assign y2899 = n11314 ;
  assign y2900 = n11319 ;
  assign y2901 = n11321 ;
  assign y2902 = ~1'b0 ;
  assign y2903 = ~n11325 ;
  assign y2904 = ~n11326 ;
  assign y2905 = n11327 ;
  assign y2906 = ~1'b0 ;
  assign y2907 = n11334 ;
  assign y2908 = n11336 ;
  assign y2909 = n11338 ;
  assign y2910 = n11346 ;
  assign y2911 = ~n11347 ;
  assign y2912 = ~1'b0 ;
  assign y2913 = ~n11350 ;
  assign y2914 = ~n11351 ;
  assign y2915 = ~n11352 ;
  assign y2916 = ~1'b0 ;
  assign y2917 = ~n11367 ;
  assign y2918 = ~n11371 ;
  assign y2919 = n4087 ;
  assign y2920 = ~n11372 ;
  assign y2921 = n11373 ;
  assign y2922 = n11380 ;
  assign y2923 = ~n11382 ;
  assign y2924 = n11384 ;
  assign y2925 = ~n11390 ;
  assign y2926 = ~1'b0 ;
  assign y2927 = n11395 ;
  assign y2928 = ~n11404 ;
  assign y2929 = n11411 ;
  assign y2930 = ~n11415 ;
  assign y2931 = n11421 ;
  assign y2932 = ~n11422 ;
  assign y2933 = ~n11423 ;
  assign y2934 = n11424 ;
  assign y2935 = ~n11427 ;
  assign y2936 = n11428 ;
  assign y2937 = n11429 ;
  assign y2938 = ~n11431 ;
  assign y2939 = n11434 ;
  assign y2940 = n11439 ;
  assign y2941 = n11441 ;
  assign y2942 = ~n11445 ;
  assign y2943 = n11448 ;
  assign y2944 = n11451 ;
  assign y2945 = n11465 ;
  assign y2946 = ~n11468 ;
  assign y2947 = ~n11474 ;
  assign y2948 = ~n11476 ;
  assign y2949 = n11479 ;
  assign y2950 = n11487 ;
  assign y2951 = ~n11488 ;
  assign y2952 = n11495 ;
  assign y2953 = ~1'b0 ;
  assign y2954 = ~n11496 ;
  assign y2955 = n11500 ;
  assign y2956 = ~1'b0 ;
  assign y2957 = n11513 ;
  assign y2958 = n11515 ;
  assign y2959 = ~n11518 ;
  assign y2960 = ~n11528 ;
  assign y2961 = ~n11534 ;
  assign y2962 = ~1'b0 ;
  assign y2963 = ~1'b0 ;
  assign y2964 = ~n11537 ;
  assign y2965 = ~n11543 ;
  assign y2966 = n11546 ;
  assign y2967 = n11548 ;
  assign y2968 = n11552 ;
  assign y2969 = n11553 ;
  assign y2970 = ~n11555 ;
  assign y2971 = n11558 ;
  assign y2972 = ~n11564 ;
  assign y2973 = n11566 ;
  assign y2974 = ~n11573 ;
  assign y2975 = n11580 ;
  assign y2976 = ~n11582 ;
  assign y2977 = n11583 ;
  assign y2978 = n11585 ;
  assign y2979 = ~n11599 ;
  assign y2980 = ~n11611 ;
  assign y2981 = n11613 ;
  assign y2982 = ~n11614 ;
  assign y2983 = ~n11620 ;
  assign y2984 = ~1'b0 ;
  assign y2985 = n11624 ;
  assign y2986 = ~1'b0 ;
  assign y2987 = ~1'b0 ;
  assign y2988 = ~n11625 ;
  assign y2989 = ~1'b0 ;
  assign y2990 = n11633 ;
  assign y2991 = ~n11636 ;
  assign y2992 = ~n11637 ;
  assign y2993 = n11644 ;
  assign y2994 = n11645 ;
  assign y2995 = ~n11652 ;
  assign y2996 = ~n11664 ;
  assign y2997 = n11670 ;
  assign y2998 = ~1'b0 ;
  assign y2999 = ~n11671 ;
  assign y3000 = ~n7196 ;
  assign y3001 = n11676 ;
  assign y3002 = ~1'b0 ;
  assign y3003 = n11680 ;
  assign y3004 = n11688 ;
  assign y3005 = ~1'b0 ;
  assign y3006 = n11690 ;
  assign y3007 = n11691 ;
  assign y3008 = ~n11696 ;
  assign y3009 = n11703 ;
  assign y3010 = ~n11714 ;
  assign y3011 = ~1'b0 ;
  assign y3012 = n11724 ;
  assign y3013 = ~n11744 ;
  assign y3014 = n3109 ;
  assign y3015 = ~n11759 ;
  assign y3016 = ~1'b0 ;
  assign y3017 = n11763 ;
  assign y3018 = ~n11764 ;
  assign y3019 = ~1'b0 ;
  assign y3020 = ~n11769 ;
  assign y3021 = ~n11780 ;
  assign y3022 = ~n11786 ;
  assign y3023 = ~n11787 ;
  assign y3024 = n11795 ;
  assign y3025 = ~n11796 ;
  assign y3026 = ~1'b0 ;
  assign y3027 = n11806 ;
  assign y3028 = n11808 ;
  assign y3029 = ~1'b0 ;
  assign y3030 = ~n11814 ;
  assign y3031 = ~n11816 ;
  assign y3032 = n11817 ;
  assign y3033 = ~n11822 ;
  assign y3034 = ~1'b0 ;
  assign y3035 = ~1'b0 ;
  assign y3036 = ~x156 ;
  assign y3037 = ~n11823 ;
  assign y3038 = ~n11839 ;
  assign y3039 = ~n11841 ;
  assign y3040 = ~n11842 ;
  assign y3041 = ~n11843 ;
  assign y3042 = ~n11846 ;
  assign y3043 = n11850 ;
  assign y3044 = ~n11865 ;
  assign y3045 = ~n11871 ;
  assign y3046 = n11874 ;
  assign y3047 = ~n11875 ;
  assign y3048 = ~n11892 ;
  assign y3049 = ~n11897 ;
  assign y3050 = ~n11898 ;
  assign y3051 = ~n11910 ;
  assign y3052 = ~n11919 ;
  assign y3053 = n11920 ;
  assign y3054 = ~n11922 ;
  assign y3055 = ~1'b0 ;
  assign y3056 = n11923 ;
  assign y3057 = ~1'b0 ;
  assign y3058 = ~n11925 ;
  assign y3059 = n11927 ;
  assign y3060 = ~n11935 ;
  assign y3061 = ~1'b0 ;
  assign y3062 = n11937 ;
  assign y3063 = n11943 ;
  assign y3064 = n11952 ;
  assign y3065 = n11957 ;
  assign y3066 = ~1'b0 ;
  assign y3067 = n11958 ;
  assign y3068 = ~n11959 ;
  assign y3069 = ~n11965 ;
  assign y3070 = n11970 ;
  assign y3071 = ~1'b0 ;
  assign y3072 = n11973 ;
  assign y3073 = n11980 ;
  assign y3074 = n11986 ;
  assign y3075 = n11987 ;
  assign y3076 = n11999 ;
  assign y3077 = n12001 ;
  assign y3078 = ~n12006 ;
  assign y3079 = ~n12010 ;
  assign y3080 = ~n12011 ;
  assign y3081 = ~n12014 ;
  assign y3082 = ~n12035 ;
  assign y3083 = ~n12038 ;
  assign y3084 = n12049 ;
  assign y3085 = ~1'b0 ;
  assign y3086 = n12066 ;
  assign y3087 = ~n12068 ;
  assign y3088 = n12071 ;
  assign y3089 = n12076 ;
  assign y3090 = ~1'b0 ;
  assign y3091 = n12078 ;
  assign y3092 = n12084 ;
  assign y3093 = ~1'b0 ;
  assign y3094 = ~n12085 ;
  assign y3095 = ~n12087 ;
  assign y3096 = ~1'b0 ;
  assign y3097 = ~1'b0 ;
  assign y3098 = n12090 ;
  assign y3099 = n12094 ;
  assign y3100 = n12102 ;
  assign y3101 = ~n12105 ;
  assign y3102 = n12106 ;
  assign y3103 = ~1'b0 ;
  assign y3104 = ~1'b0 ;
  assign y3105 = n12108 ;
  assign y3106 = ~n12112 ;
  assign y3107 = ~n12121 ;
  assign y3108 = n12127 ;
  assign y3109 = n12130 ;
  assign y3110 = ~n12134 ;
  assign y3111 = ~n12138 ;
  assign y3112 = n12142 ;
  assign y3113 = n12146 ;
  assign y3114 = ~n12149 ;
  assign y3115 = n12152 ;
  assign y3116 = n12153 ;
  assign y3117 = ~n12155 ;
  assign y3118 = n12157 ;
  assign y3119 = n12158 ;
  assign y3120 = ~n12162 ;
  assign y3121 = n12168 ;
  assign y3122 = n12171 ;
  assign y3123 = ~n12173 ;
  assign y3124 = ~n12182 ;
  assign y3125 = n12187 ;
  assign y3126 = ~n12190 ;
  assign y3127 = n12191 ;
  assign y3128 = n12194 ;
  assign y3129 = ~n12196 ;
  assign y3130 = n12204 ;
  assign y3131 = ~1'b0 ;
  assign y3132 = ~n12208 ;
  assign y3133 = ~n12213 ;
  assign y3134 = n12215 ;
  assign y3135 = n12228 ;
  assign y3136 = ~n12229 ;
  assign y3137 = ~n12232 ;
  assign y3138 = n12236 ;
  assign y3139 = n12237 ;
  assign y3140 = n12242 ;
  assign y3141 = ~n12245 ;
  assign y3142 = x49 ;
  assign y3143 = ~n12248 ;
  assign y3144 = ~n12257 ;
  assign y3145 = n12259 ;
  assign y3146 = n12262 ;
  assign y3147 = n12264 ;
  assign y3148 = ~n12265 ;
  assign y3149 = ~1'b0 ;
  assign y3150 = ~n12270 ;
  assign y3151 = ~n12276 ;
  assign y3152 = ~1'b0 ;
  assign y3153 = n12282 ;
  assign y3154 = ~n12286 ;
  assign y3155 = ~1'b0 ;
  assign y3156 = n12288 ;
  assign y3157 = ~1'b0 ;
  assign y3158 = ~n12290 ;
  assign y3159 = ~n12293 ;
  assign y3160 = ~n12296 ;
  assign y3161 = ~1'b0 ;
  assign y3162 = ~n12298 ;
  assign y3163 = ~n12299 ;
  assign y3164 = n12300 ;
  assign y3165 = n12309 ;
  assign y3166 = ~1'b0 ;
  assign y3167 = n12318 ;
  assign y3168 = n12319 ;
  assign y3169 = ~n12320 ;
  assign y3170 = n12321 ;
  assign y3171 = n12331 ;
  assign y3172 = ~1'b0 ;
  assign y3173 = n12336 ;
  assign y3174 = ~n12342 ;
  assign y3175 = ~n12350 ;
  assign y3176 = ~1'b0 ;
  assign y3177 = n12351 ;
  assign y3178 = n12357 ;
  assign y3179 = ~1'b0 ;
  assign y3180 = ~n3979 ;
  assign y3181 = ~n11429 ;
  assign y3182 = n12359 ;
  assign y3183 = n12361 ;
  assign y3184 = n12366 ;
  assign y3185 = ~n12368 ;
  assign y3186 = ~n12372 ;
  assign y3187 = ~1'b0 ;
  assign y3188 = ~n12378 ;
  assign y3189 = n12382 ;
  assign y3190 = n12386 ;
  assign y3191 = n12396 ;
  assign y3192 = n12401 ;
  assign y3193 = n12402 ;
  assign y3194 = ~n12405 ;
  assign y3195 = n12413 ;
  assign y3196 = n12418 ;
  assign y3197 = ~n12436 ;
  assign y3198 = n12437 ;
  assign y3199 = ~n12439 ;
  assign y3200 = ~n12443 ;
  assign y3201 = ~n12448 ;
  assign y3202 = ~n12449 ;
  assign y3203 = ~n12453 ;
  assign y3204 = n12465 ;
  assign y3205 = n12467 ;
  assign y3206 = ~n12470 ;
  assign y3207 = ~n12473 ;
  assign y3208 = ~n12480 ;
  assign y3209 = ~n12481 ;
  assign y3210 = n12484 ;
  assign y3211 = ~n12485 ;
  assign y3212 = ~n12488 ;
  assign y3213 = n12491 ;
  assign y3214 = ~n12493 ;
  assign y3215 = ~n12501 ;
  assign y3216 = n12502 ;
  assign y3217 = ~n12507 ;
  assign y3218 = ~n12508 ;
  assign y3219 = n12517 ;
  assign y3220 = ~n12518 ;
  assign y3221 = n12522 ;
  assign y3222 = n12525 ;
  assign y3223 = n12530 ;
  assign y3224 = n12534 ;
  assign y3225 = n12535 ;
  assign y3226 = n12536 ;
  assign y3227 = ~1'b0 ;
  assign y3228 = ~n12539 ;
  assign y3229 = ~n12548 ;
  assign y3230 = ~n12550 ;
  assign y3231 = n12555 ;
  assign y3232 = ~1'b0 ;
  assign y3233 = ~n12565 ;
  assign y3234 = ~n12566 ;
  assign y3235 = ~n8947 ;
  assign y3236 = ~n12574 ;
  assign y3237 = ~n12579 ;
  assign y3238 = ~n12580 ;
  assign y3239 = ~n12581 ;
  assign y3240 = n12583 ;
  assign y3241 = ~n12590 ;
  assign y3242 = ~n12593 ;
  assign y3243 = ~n12596 ;
  assign y3244 = ~1'b0 ;
  assign y3245 = ~1'b0 ;
  assign y3246 = n12599 ;
  assign y3247 = n12604 ;
  assign y3248 = ~n12610 ;
  assign y3249 = ~n12614 ;
  assign y3250 = n12620 ;
  assign y3251 = ~n12623 ;
  assign y3252 = ~n12625 ;
  assign y3253 = n12626 ;
  assign y3254 = n12628 ;
  assign y3255 = n12631 ;
  assign y3256 = n12639 ;
  assign y3257 = n4662 ;
  assign y3258 = n12644 ;
  assign y3259 = n12648 ;
  assign y3260 = ~1'b0 ;
  assign y3261 = n12651 ;
  assign y3262 = ~n12665 ;
  assign y3263 = ~n12671 ;
  assign y3264 = n12675 ;
  assign y3265 = ~1'b0 ;
  assign y3266 = ~n12685 ;
  assign y3267 = n12687 ;
  assign y3268 = ~1'b0 ;
  assign y3269 = n12696 ;
  assign y3270 = n12698 ;
  assign y3271 = ~1'b0 ;
  assign y3272 = ~n12704 ;
  assign y3273 = n12705 ;
  assign y3274 = ~n12707 ;
  assign y3275 = ~n12708 ;
  assign y3276 = ~n12717 ;
  assign y3277 = ~n12730 ;
  assign y3278 = ~1'b0 ;
  assign y3279 = n12731 ;
  assign y3280 = ~1'b0 ;
  assign y3281 = n12733 ;
  assign y3282 = ~1'b0 ;
  assign y3283 = ~n12747 ;
  assign y3284 = ~n12752 ;
  assign y3285 = ~n12756 ;
  assign y3286 = n12758 ;
  assign y3287 = n12759 ;
  assign y3288 = n12761 ;
  assign y3289 = ~1'b0 ;
  assign y3290 = ~1'b0 ;
  assign y3291 = ~n12763 ;
  assign y3292 = ~n12770 ;
  assign y3293 = ~n12773 ;
  assign y3294 = n12774 ;
  assign y3295 = n12778 ;
  assign y3296 = ~n12779 ;
  assign y3297 = ~n12781 ;
  assign y3298 = ~n12785 ;
  assign y3299 = ~1'b0 ;
  assign y3300 = n12790 ;
  assign y3301 = n12792 ;
  assign y3302 = ~n12793 ;
  assign y3303 = n12802 ;
  assign y3304 = ~1'b0 ;
  assign y3305 = ~n12809 ;
  assign y3306 = n12813 ;
  assign y3307 = n12820 ;
  assign y3308 = ~1'b0 ;
  assign y3309 = n12828 ;
  assign y3310 = n12831 ;
  assign y3311 = ~n12838 ;
  assign y3312 = ~n12842 ;
  assign y3313 = ~n12845 ;
  assign y3314 = n12851 ;
  assign y3315 = ~n12863 ;
  assign y3316 = n12879 ;
  assign y3317 = ~1'b0 ;
  assign y3318 = n12885 ;
  assign y3319 = ~n12886 ;
  assign y3320 = n12892 ;
  assign y3321 = n12903 ;
  assign y3322 = ~n12904 ;
  assign y3323 = ~n12913 ;
  assign y3324 = ~n12920 ;
  assign y3325 = n12922 ;
  assign y3326 = n12925 ;
  assign y3327 = ~n12928 ;
  assign y3328 = ~n12936 ;
  assign y3329 = ~n12937 ;
  assign y3330 = n12941 ;
  assign y3331 = ~n12942 ;
  assign y3332 = ~n12944 ;
  assign y3333 = ~n12945 ;
  assign y3334 = n12950 ;
  assign y3335 = ~n12952 ;
  assign y3336 = n12954 ;
  assign y3337 = n12958 ;
  assign y3338 = n12961 ;
  assign y3339 = ~n12962 ;
  assign y3340 = n12968 ;
  assign y3341 = ~n12987 ;
  assign y3342 = n12990 ;
  assign y3343 = ~1'b0 ;
  assign y3344 = ~n12994 ;
  assign y3345 = ~1'b0 ;
  assign y3346 = ~1'b0 ;
  assign y3347 = ~n12997 ;
  assign y3348 = n13000 ;
  assign y3349 = ~1'b0 ;
  assign y3350 = ~n13003 ;
  assign y3351 = ~1'b0 ;
  assign y3352 = ~n13007 ;
  assign y3353 = ~n13009 ;
  assign y3354 = n13011 ;
  assign y3355 = n13012 ;
  assign y3356 = n13014 ;
  assign y3357 = ~1'b0 ;
  assign y3358 = ~n13016 ;
  assign y3359 = ~n13017 ;
  assign y3360 = n13018 ;
  assign y3361 = n13019 ;
  assign y3362 = ~n13024 ;
  assign y3363 = ~1'b0 ;
  assign y3364 = ~n13028 ;
  assign y3365 = ~n13029 ;
  assign y3366 = ~n13041 ;
  assign y3367 = ~n13045 ;
  assign y3368 = n13047 ;
  assign y3369 = ~n13051 ;
  assign y3370 = ~n13054 ;
  assign y3371 = n11908 ;
  assign y3372 = n13057 ;
  assign y3373 = ~n13067 ;
  assign y3374 = ~n13078 ;
  assign y3375 = n9312 ;
  assign y3376 = ~n13081 ;
  assign y3377 = ~n13084 ;
  assign y3378 = ~1'b0 ;
  assign y3379 = n13087 ;
  assign y3380 = n13095 ;
  assign y3381 = ~n13101 ;
  assign y3382 = n13102 ;
  assign y3383 = ~n13105 ;
  assign y3384 = n13116 ;
  assign y3385 = n13119 ;
  assign y3386 = ~n13124 ;
  assign y3387 = ~n13125 ;
  assign y3388 = ~1'b0 ;
  assign y3389 = ~n13126 ;
  assign y3390 = n13128 ;
  assign y3391 = ~1'b0 ;
  assign y3392 = ~n13129 ;
  assign y3393 = ~n13130 ;
  assign y3394 = ~n13139 ;
  assign y3395 = n13147 ;
  assign y3396 = ~n13163 ;
  assign y3397 = ~1'b0 ;
  assign y3398 = ~n13169 ;
  assign y3399 = ~n13174 ;
  assign y3400 = n13179 ;
  assign y3401 = n13184 ;
  assign y3402 = n13186 ;
  assign y3403 = ~1'b0 ;
  assign y3404 = n13198 ;
  assign y3405 = ~n13200 ;
  assign y3406 = ~n13203 ;
  assign y3407 = ~n13205 ;
  assign y3408 = ~1'b0 ;
  assign y3409 = ~n13209 ;
  assign y3410 = n13211 ;
  assign y3411 = ~n13217 ;
  assign y3412 = ~n13220 ;
  assign y3413 = ~n13221 ;
  assign y3414 = n13223 ;
  assign y3415 = ~n13235 ;
  assign y3416 = ~n13236 ;
  assign y3417 = n13237 ;
  assign y3418 = n13242 ;
  assign y3419 = ~n13245 ;
  assign y3420 = n13248 ;
  assign y3421 = n13250 ;
  assign y3422 = ~n13251 ;
  assign y3423 = n13256 ;
  assign y3424 = ~n13259 ;
  assign y3425 = ~1'b0 ;
  assign y3426 = n13265 ;
  assign y3427 = n13266 ;
  assign y3428 = ~n13267 ;
  assign y3429 = ~n13268 ;
  assign y3430 = ~n13280 ;
  assign y3431 = n13288 ;
  assign y3432 = n13293 ;
  assign y3433 = ~1'b0 ;
  assign y3434 = n13295 ;
  assign y3435 = n13303 ;
  assign y3436 = ~1'b0 ;
  assign y3437 = ~n13304 ;
  assign y3438 = ~1'b0 ;
  assign y3439 = ~n13308 ;
  assign y3440 = ~n13311 ;
  assign y3441 = n13315 ;
  assign y3442 = ~1'b0 ;
  assign y3443 = n13316 ;
  assign y3444 = ~1'b0 ;
  assign y3445 = ~n13320 ;
  assign y3446 = n13322 ;
  assign y3447 = ~1'b0 ;
  assign y3448 = ~n13323 ;
  assign y3449 = ~1'b0 ;
  assign y3450 = n13325 ;
  assign y3451 = n13334 ;
  assign y3452 = ~1'b0 ;
  assign y3453 = ~1'b0 ;
  assign y3454 = ~n13335 ;
  assign y3455 = ~n13338 ;
  assign y3456 = n13341 ;
  assign y3457 = n13342 ;
  assign y3458 = ~n13343 ;
  assign y3459 = ~n13344 ;
  assign y3460 = n13346 ;
  assign y3461 = ~n13350 ;
  assign y3462 = n13355 ;
  assign y3463 = ~n13361 ;
  assign y3464 = ~1'b0 ;
  assign y3465 = n13370 ;
  assign y3466 = ~n13373 ;
  assign y3467 = ~n13376 ;
  assign y3468 = ~1'b0 ;
  assign y3469 = ~n13380 ;
  assign y3470 = ~n13381 ;
  assign y3471 = ~1'b0 ;
  assign y3472 = ~1'b0 ;
  assign y3473 = ~1'b0 ;
  assign y3474 = ~n13382 ;
  assign y3475 = n13384 ;
  assign y3476 = ~1'b0 ;
  assign y3477 = ~n13391 ;
  assign y3478 = ~n13393 ;
  assign y3479 = ~n13398 ;
  assign y3480 = n13405 ;
  assign y3481 = n13407 ;
  assign y3482 = n13414 ;
  assign y3483 = ~n13415 ;
  assign y3484 = ~n13421 ;
  assign y3485 = ~1'b0 ;
  assign y3486 = n13424 ;
  assign y3487 = ~1'b0 ;
  assign y3488 = n13428 ;
  assign y3489 = ~n13433 ;
  assign y3490 = n13435 ;
  assign y3491 = ~n13437 ;
  assign y3492 = n13438 ;
  assign y3493 = ~n13441 ;
  assign y3494 = n13446 ;
  assign y3495 = n13448 ;
  assign y3496 = n13451 ;
  assign y3497 = n13453 ;
  assign y3498 = ~n13455 ;
  assign y3499 = ~n13460 ;
  assign y3500 = n13470 ;
  assign y3501 = n13473 ;
  assign y3502 = ~n13481 ;
  assign y3503 = ~1'b0 ;
  assign y3504 = ~1'b0 ;
  assign y3505 = ~n13482 ;
  assign y3506 = n13483 ;
  assign y3507 = n13487 ;
  assign y3508 = ~1'b0 ;
  assign y3509 = n13494 ;
  assign y3510 = ~n13496 ;
  assign y3511 = n13510 ;
  assign y3512 = n13517 ;
  assign y3513 = ~n13526 ;
  assign y3514 = ~n13532 ;
  assign y3515 = ~1'b0 ;
  assign y3516 = ~1'b0 ;
  assign y3517 = ~1'b0 ;
  assign y3518 = ~1'b0 ;
  assign y3519 = ~n13540 ;
  assign y3520 = n13541 ;
  assign y3521 = n13545 ;
  assign y3522 = n13547 ;
  assign y3523 = ~n13549 ;
  assign y3524 = ~1'b0 ;
  assign y3525 = ~n13551 ;
  assign y3526 = ~n13554 ;
  assign y3527 = ~1'b0 ;
  assign y3528 = ~n13565 ;
  assign y3529 = n13569 ;
  assign y3530 = ~n13572 ;
  assign y3531 = ~n13577 ;
  assign y3532 = n13595 ;
  assign y3533 = ~n13597 ;
  assign y3534 = n13601 ;
  assign y3535 = n13604 ;
  assign y3536 = n13610 ;
  assign y3537 = n13613 ;
  assign y3538 = n13624 ;
  assign y3539 = n13630 ;
  assign y3540 = n13631 ;
  assign y3541 = ~n13632 ;
  assign y3542 = ~n13637 ;
  assign y3543 = ~n13638 ;
  assign y3544 = n13641 ;
  assign y3545 = ~n3666 ;
  assign y3546 = n13644 ;
  assign y3547 = ~1'b0 ;
  assign y3548 = ~n13645 ;
  assign y3549 = ~n13646 ;
  assign y3550 = n13648 ;
  assign y3551 = ~n13652 ;
  assign y3552 = n13655 ;
  assign y3553 = n13657 ;
  assign y3554 = ~n13660 ;
  assign y3555 = ~n13667 ;
  assign y3556 = n13672 ;
  assign y3557 = n13675 ;
  assign y3558 = n13677 ;
  assign y3559 = ~n13683 ;
  assign y3560 = n10884 ;
  assign y3561 = n13684 ;
  assign y3562 = ~n13685 ;
  assign y3563 = n13687 ;
  assign y3564 = ~n13698 ;
  assign y3565 = n13700 ;
  assign y3566 = ~n13701 ;
  assign y3567 = n13703 ;
  assign y3568 = n13707 ;
  assign y3569 = n13708 ;
  assign y3570 = ~1'b0 ;
  assign y3571 = ~n13719 ;
  assign y3572 = n13723 ;
  assign y3573 = ~1'b0 ;
  assign y3574 = ~n13730 ;
  assign y3575 = n13732 ;
  assign y3576 = n13735 ;
  assign y3577 = ~n4011 ;
  assign y3578 = n13741 ;
  assign y3579 = n13744 ;
  assign y3580 = n13751 ;
  assign y3581 = ~1'b0 ;
  assign y3582 = n13752 ;
  assign y3583 = n13762 ;
  assign y3584 = n13764 ;
  assign y3585 = ~1'b0 ;
  assign y3586 = n13770 ;
  assign y3587 = n13776 ;
  assign y3588 = ~n13777 ;
  assign y3589 = ~n13782 ;
  assign y3590 = n13793 ;
  assign y3591 = ~1'b0 ;
  assign y3592 = n13799 ;
  assign y3593 = ~n13803 ;
  assign y3594 = n13804 ;
  assign y3595 = n13805 ;
  assign y3596 = ~n13808 ;
  assign y3597 = ~n13812 ;
  assign y3598 = n13814 ;
  assign y3599 = ~n13820 ;
  assign y3600 = n13825 ;
  assign y3601 = ~1'b0 ;
  assign y3602 = n13827 ;
  assign y3603 = ~n13828 ;
  assign y3604 = ~n13829 ;
  assign y3605 = n13830 ;
  assign y3606 = ~n13839 ;
  assign y3607 = n13843 ;
  assign y3608 = n13856 ;
  assign y3609 = ~n13866 ;
  assign y3610 = n13867 ;
  assign y3611 = ~n13879 ;
  assign y3612 = ~1'b0 ;
  assign y3613 = ~n13881 ;
  assign y3614 = ~n13882 ;
  assign y3615 = ~1'b0 ;
  assign y3616 = n13883 ;
  assign y3617 = ~1'b0 ;
  assign y3618 = ~n13889 ;
  assign y3619 = ~n13892 ;
  assign y3620 = ~n13893 ;
  assign y3621 = ~n13898 ;
  assign y3622 = ~1'b0 ;
  assign y3623 = n13903 ;
  assign y3624 = n13911 ;
  assign y3625 = n13917 ;
  assign y3626 = n13925 ;
  assign y3627 = ~n13927 ;
  assign y3628 = n13931 ;
  assign y3629 = n13932 ;
  assign y3630 = ~n13936 ;
  assign y3631 = n13939 ;
  assign y3632 = ~1'b0 ;
  assign y3633 = n13951 ;
  assign y3634 = n13954 ;
  assign y3635 = ~n13956 ;
  assign y3636 = n13962 ;
  assign y3637 = n13963 ;
  assign y3638 = ~n13965 ;
  assign y3639 = ~n13967 ;
  assign y3640 = n13968 ;
  assign y3641 = ~n13987 ;
  assign y3642 = ~1'b0 ;
  assign y3643 = n13994 ;
  assign y3644 = ~n6736 ;
  assign y3645 = n13996 ;
  assign y3646 = n14001 ;
  assign y3647 = n14002 ;
  assign y3648 = n14004 ;
  assign y3649 = n14008 ;
  assign y3650 = n14010 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = ~1'b0 ;
  assign y3653 = ~n14011 ;
  assign y3654 = n14024 ;
  assign y3655 = ~1'b0 ;
  assign y3656 = ~n14027 ;
  assign y3657 = n14028 ;
  assign y3658 = ~n14031 ;
  assign y3659 = n14044 ;
  assign y3660 = ~n14045 ;
  assign y3661 = ~n14046 ;
  assign y3662 = n14050 ;
  assign y3663 = ~n14063 ;
  assign y3664 = n14064 ;
  assign y3665 = ~1'b0 ;
  assign y3666 = n14065 ;
  assign y3667 = ~n14068 ;
  assign y3668 = n14077 ;
  assign y3669 = n14080 ;
  assign y3670 = n6797 ;
  assign y3671 = ~n14082 ;
  assign y3672 = n14083 ;
  assign y3673 = ~n14084 ;
  assign y3674 = ~n14090 ;
  assign y3675 = n14091 ;
  assign y3676 = n14093 ;
  assign y3677 = ~n14094 ;
  assign y3678 = ~n14095 ;
  assign y3679 = n14099 ;
  assign y3680 = ~n14104 ;
  assign y3681 = ~n14107 ;
  assign y3682 = n14111 ;
  assign y3683 = ~n14113 ;
  assign y3684 = n1233 ;
  assign y3685 = n14114 ;
  assign y3686 = ~n14122 ;
  assign y3687 = ~n14127 ;
  assign y3688 = n14130 ;
  assign y3689 = ~n14131 ;
  assign y3690 = n14132 ;
  assign y3691 = ~n14135 ;
  assign y3692 = n14137 ;
  assign y3693 = ~n14146 ;
  assign y3694 = ~n14147 ;
  assign y3695 = ~1'b0 ;
  assign y3696 = n14163 ;
  assign y3697 = ~n14173 ;
  assign y3698 = n14174 ;
  assign y3699 = ~1'b0 ;
  assign y3700 = ~n14182 ;
  assign y3701 = n14194 ;
  assign y3702 = n14201 ;
  assign y3703 = n14211 ;
  assign y3704 = n14213 ;
  assign y3705 = ~n14222 ;
  assign y3706 = ~n14224 ;
  assign y3707 = n14230 ;
  assign y3708 = n14237 ;
  assign y3709 = ~n14245 ;
  assign y3710 = ~n14247 ;
  assign y3711 = ~n14253 ;
  assign y3712 = ~n14255 ;
  assign y3713 = n14256 ;
  assign y3714 = ~1'b0 ;
  assign y3715 = n14262 ;
  assign y3716 = n14265 ;
  assign y3717 = n14267 ;
  assign y3718 = ~n14268 ;
  assign y3719 = ~1'b0 ;
  assign y3720 = 1'b0 ;
  assign y3721 = n14269 ;
  assign y3722 = ~n14274 ;
  assign y3723 = ~1'b0 ;
  assign y3724 = n14278 ;
  assign y3725 = n14281 ;
  assign y3726 = n14283 ;
  assign y3727 = ~1'b0 ;
  assign y3728 = n14291 ;
  assign y3729 = n14298 ;
  assign y3730 = ~n14302 ;
  assign y3731 = ~1'b0 ;
  assign y3732 = ~n14306 ;
  assign y3733 = ~n14307 ;
  assign y3734 = ~n14309 ;
  assign y3735 = ~n14312 ;
  assign y3736 = ~n14313 ;
  assign y3737 = ~n14317 ;
  assign y3738 = ~n14318 ;
  assign y3739 = ~n14329 ;
  assign y3740 = ~n14336 ;
  assign y3741 = ~n14338 ;
  assign y3742 = n14340 ;
  assign y3743 = ~n14342 ;
  assign y3744 = n14346 ;
  assign y3745 = ~n14348 ;
  assign y3746 = n14354 ;
  assign y3747 = ~n14363 ;
  assign y3748 = n14364 ;
  assign y3749 = ~n14370 ;
  assign y3750 = n14371 ;
  assign y3751 = n14374 ;
  assign y3752 = ~n10373 ;
  assign y3753 = n14379 ;
  assign y3754 = ~1'b0 ;
  assign y3755 = ~n14383 ;
  assign y3756 = ~n14386 ;
  assign y3757 = ~n14392 ;
  assign y3758 = ~n14397 ;
  assign y3759 = n14402 ;
  assign y3760 = ~n14408 ;
  assign y3761 = ~n14429 ;
  assign y3762 = ~n14436 ;
  assign y3763 = n14438 ;
  assign y3764 = ~1'b0 ;
  assign y3765 = n14440 ;
  assign y3766 = ~n14441 ;
  assign y3767 = ~1'b0 ;
  assign y3768 = n14449 ;
  assign y3769 = ~n14460 ;
  assign y3770 = n14470 ;
  assign y3771 = n14473 ;
  assign y3772 = n14479 ;
  assign y3773 = ~n14483 ;
  assign y3774 = n14484 ;
  assign y3775 = ~n14486 ;
  assign y3776 = n14496 ;
  assign y3777 = n14505 ;
  assign y3778 = ~1'b0 ;
  assign y3779 = ~n14510 ;
  assign y3780 = ~n14512 ;
  assign y3781 = ~1'b0 ;
  assign y3782 = n14522 ;
  assign y3783 = ~1'b0 ;
  assign y3784 = n14524 ;
  assign y3785 = ~n14529 ;
  assign y3786 = n14531 ;
  assign y3787 = ~n14533 ;
  assign y3788 = ~n14537 ;
  assign y3789 = ~n14541 ;
  assign y3790 = n14554 ;
  assign y3791 = ~n14559 ;
  assign y3792 = n14561 ;
  assign y3793 = n14563 ;
  assign y3794 = ~n14568 ;
  assign y3795 = n14581 ;
  assign y3796 = n14589 ;
  assign y3797 = ~1'b0 ;
  assign y3798 = ~1'b0 ;
  assign y3799 = n14592 ;
  assign y3800 = n14594 ;
  assign y3801 = ~n14596 ;
  assign y3802 = ~n14598 ;
  assign y3803 = ~n14610 ;
  assign y3804 = ~n14611 ;
  assign y3805 = n14612 ;
  assign y3806 = ~n14613 ;
  assign y3807 = ~n14618 ;
  assign y3808 = ~n14621 ;
  assign y3809 = n14628 ;
  assign y3810 = n14629 ;
  assign y3811 = ~1'b0 ;
  assign y3812 = ~n14630 ;
  assign y3813 = n14634 ;
  assign y3814 = n14635 ;
  assign y3815 = ~n14642 ;
  assign y3816 = ~1'b0 ;
  assign y3817 = ~1'b0 ;
  assign y3818 = n14651 ;
  assign y3819 = n14657 ;
  assign y3820 = ~n14660 ;
  assign y3821 = n14661 ;
  assign y3822 = ~n14663 ;
  assign y3823 = n14664 ;
  assign y3824 = n14669 ;
  assign y3825 = n14684 ;
  assign y3826 = ~1'b0 ;
  assign y3827 = ~n14686 ;
  assign y3828 = n14692 ;
  assign y3829 = ~n14693 ;
  assign y3830 = ~n14704 ;
  assign y3831 = ~1'b0 ;
  assign y3832 = n14710 ;
  assign y3833 = n14711 ;
  assign y3834 = n14713 ;
  assign y3835 = ~n14714 ;
  assign y3836 = ~n3527 ;
  assign y3837 = ~n14727 ;
  assign y3838 = ~n14729 ;
  assign y3839 = ~n14732 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = n14734 ;
  assign y3842 = n14735 ;
  assign y3843 = n14742 ;
  assign y3844 = ~n14749 ;
  assign y3845 = ~n14752 ;
  assign y3846 = ~1'b0 ;
  assign y3847 = ~n14755 ;
  assign y3848 = ~1'b0 ;
  assign y3849 = ~1'b0 ;
  assign y3850 = n14761 ;
  assign y3851 = n14763 ;
  assign y3852 = ~1'b0 ;
  assign y3853 = n14764 ;
  assign y3854 = ~n14768 ;
  assign y3855 = n14769 ;
  assign y3856 = ~n14785 ;
  assign y3857 = ~1'b0 ;
  assign y3858 = ~n14791 ;
  assign y3859 = ~n14799 ;
  assign y3860 = ~n14804 ;
  assign y3861 = ~n14806 ;
  assign y3862 = ~n14807 ;
  assign y3863 = ~n14812 ;
  assign y3864 = ~n14816 ;
  assign y3865 = n14825 ;
  assign y3866 = ~n14829 ;
  assign y3867 = n14831 ;
  assign y3868 = ~n14838 ;
  assign y3869 = ~n14842 ;
  assign y3870 = ~n14847 ;
  assign y3871 = ~n14849 ;
  assign y3872 = ~n14851 ;
  assign y3873 = n14858 ;
  assign y3874 = ~n14865 ;
  assign y3875 = n14871 ;
  assign y3876 = ~n14881 ;
  assign y3877 = ~n14884 ;
  assign y3878 = n14889 ;
  assign y3879 = ~1'b0 ;
  assign y3880 = ~n14893 ;
  assign y3881 = n14895 ;
  assign y3882 = n14898 ;
  assign y3883 = ~n14906 ;
  assign y3884 = n14909 ;
  assign y3885 = n14916 ;
  assign y3886 = n14920 ;
  assign y3887 = ~1'b0 ;
  assign y3888 = ~n14921 ;
  assign y3889 = ~n14922 ;
  assign y3890 = ~n14923 ;
  assign y3891 = n14924 ;
  assign y3892 = ~1'b0 ;
  assign y3893 = ~n14935 ;
  assign y3894 = ~n14936 ;
  assign y3895 = ~1'b0 ;
  assign y3896 = ~n14937 ;
  assign y3897 = ~n14940 ;
  assign y3898 = ~1'b0 ;
  assign y3899 = ~n14943 ;
  assign y3900 = n14945 ;
  assign y3901 = n14948 ;
  assign y3902 = ~n14956 ;
  assign y3903 = ~n14961 ;
  assign y3904 = ~n14965 ;
  assign y3905 = ~n14971 ;
  assign y3906 = n14986 ;
  assign y3907 = ~1'b0 ;
  assign y3908 = ~n14989 ;
  assign y3909 = ~n14993 ;
  assign y3910 = ~n14995 ;
  assign y3911 = n15002 ;
  assign y3912 = ~1'b0 ;
  assign y3913 = ~n15006 ;
  assign y3914 = n15010 ;
  assign y3915 = ~n15016 ;
  assign y3916 = ~1'b0 ;
  assign y3917 = n15020 ;
  assign y3918 = ~n15027 ;
  assign y3919 = n15032 ;
  assign y3920 = ~n15044 ;
  assign y3921 = n15046 ;
  assign y3922 = ~n15051 ;
  assign y3923 = ~n15054 ;
  assign y3924 = ~1'b0 ;
  assign y3925 = ~n15055 ;
  assign y3926 = n15060 ;
  assign y3927 = ~n15068 ;
  assign y3928 = n15072 ;
  assign y3929 = ~1'b0 ;
  assign y3930 = n10154 ;
  assign y3931 = ~n15081 ;
  assign y3932 = n15088 ;
  assign y3933 = ~n15093 ;
  assign y3934 = n15097 ;
  assign y3935 = ~n15098 ;
  assign y3936 = ~n15099 ;
  assign y3937 = n15102 ;
  assign y3938 = ~n15108 ;
  assign y3939 = n15116 ;
  assign y3940 = ~n15117 ;
  assign y3941 = n15118 ;
  assign y3942 = ~n15122 ;
  assign y3943 = ~1'b0 ;
  assign y3944 = ~n15124 ;
  assign y3945 = ~n15127 ;
  assign y3946 = n15130 ;
  assign y3947 = n15135 ;
  assign y3948 = ~n15136 ;
  assign y3949 = n11494 ;
  assign y3950 = ~1'b0 ;
  assign y3951 = n15138 ;
  assign y3952 = ~n15142 ;
  assign y3953 = n15149 ;
  assign y3954 = n15154 ;
  assign y3955 = n15161 ;
  assign y3956 = n15167 ;
  assign y3957 = n15170 ;
  assign y3958 = ~n15171 ;
  assign y3959 = n15177 ;
  assign y3960 = ~n15179 ;
  assign y3961 = ~n15188 ;
  assign y3962 = ~n15189 ;
  assign y3963 = n15193 ;
  assign y3964 = ~n15198 ;
  assign y3965 = n15206 ;
  assign y3966 = ~n15215 ;
  assign y3967 = n15216 ;
  assign y3968 = n15218 ;
  assign y3969 = ~1'b0 ;
  assign y3970 = ~n15219 ;
  assign y3971 = ~n15220 ;
  assign y3972 = ~n15223 ;
  assign y3973 = ~n15224 ;
  assign y3974 = ~n15230 ;
  assign y3975 = n15232 ;
  assign y3976 = ~n15241 ;
  assign y3977 = n15242 ;
  assign y3978 = n15243 ;
  assign y3979 = ~n15245 ;
  assign y3980 = n15247 ;
  assign y3981 = ~n15253 ;
  assign y3982 = ~n15259 ;
  assign y3983 = ~n15267 ;
  assign y3984 = ~n15275 ;
  assign y3985 = n15279 ;
  assign y3986 = n15281 ;
  assign y3987 = ~n15284 ;
  assign y3988 = ~n15285 ;
  assign y3989 = ~n15287 ;
  assign y3990 = ~n15291 ;
  assign y3991 = ~n15296 ;
  assign y3992 = n15298 ;
  assign y3993 = ~1'b0 ;
  assign y3994 = n15299 ;
  assign y3995 = ~n15311 ;
  assign y3996 = n15312 ;
  assign y3997 = n15317 ;
  assign y3998 = ~n15322 ;
  assign y3999 = ~n15324 ;
  assign y4000 = n15328 ;
  assign y4001 = n15330 ;
  assign y4002 = n15337 ;
  assign y4003 = ~n4409 ;
  assign y4004 = ~n15341 ;
  assign y4005 = n15343 ;
  assign y4006 = ~n15345 ;
  assign y4007 = ~n15350 ;
  assign y4008 = ~n15351 ;
  assign y4009 = ~n15352 ;
  assign y4010 = ~n15356 ;
  assign y4011 = ~n15357 ;
  assign y4012 = n15359 ;
  assign y4013 = n15362 ;
  assign y4014 = ~n15365 ;
  assign y4015 = ~n15372 ;
  assign y4016 = ~1'b0 ;
  assign y4017 = ~n15376 ;
  assign y4018 = ~n15377 ;
  assign y4019 = n15380 ;
  assign y4020 = n15382 ;
  assign y4021 = ~n15384 ;
  assign y4022 = ~n15386 ;
  assign y4023 = ~n15387 ;
  assign y4024 = ~n15405 ;
  assign y4025 = ~1'b0 ;
  assign y4026 = ~n15411 ;
  assign y4027 = ~n15420 ;
  assign y4028 = n15424 ;
  assign y4029 = ~n15438 ;
  assign y4030 = ~n15439 ;
  assign y4031 = ~1'b0 ;
  assign y4032 = ~n15446 ;
  assign y4033 = ~n15448 ;
  assign y4034 = ~n15452 ;
  assign y4035 = n15455 ;
  assign y4036 = ~n15457 ;
  assign y4037 = n15466 ;
  assign y4038 = ~1'b0 ;
  assign y4039 = ~1'b0 ;
  assign y4040 = n15471 ;
  assign y4041 = n15473 ;
  assign y4042 = n15474 ;
  assign y4043 = n15480 ;
  assign y4044 = n15483 ;
  assign y4045 = ~n15485 ;
  assign y4046 = ~1'b0 ;
  assign y4047 = ~n15497 ;
  assign y4048 = ~n15499 ;
  assign y4049 = ~n15501 ;
  assign y4050 = ~n15507 ;
  assign y4051 = n15508 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = ~n15509 ;
  assign y4054 = n15511 ;
  assign y4055 = ~n15514 ;
  assign y4056 = n15523 ;
  assign y4057 = ~n15530 ;
  assign y4058 = n15533 ;
  assign y4059 = ~n15541 ;
  assign y4060 = ~n15544 ;
  assign y4061 = n15554 ;
  assign y4062 = ~n15555 ;
  assign y4063 = ~n15557 ;
  assign y4064 = ~n15559 ;
  assign y4065 = ~n15564 ;
  assign y4066 = n15569 ;
  assign y4067 = n15570 ;
  assign y4068 = n15574 ;
  assign y4069 = n15582 ;
  assign y4070 = ~n15587 ;
  assign y4071 = n15590 ;
  assign y4072 = ~1'b0 ;
  assign y4073 = ~n15593 ;
  assign y4074 = ~n15595 ;
  assign y4075 = n15600 ;
  assign y4076 = n15611 ;
  assign y4077 = ~n15617 ;
  assign y4078 = n15621 ;
  assign y4079 = ~n15626 ;
  assign y4080 = ~1'b0 ;
  assign y4081 = n15628 ;
  assign y4082 = ~n15637 ;
  assign y4083 = n15639 ;
  assign y4084 = ~n15640 ;
  assign y4085 = ~1'b0 ;
  assign y4086 = ~n15644 ;
  assign y4087 = ~1'b0 ;
  assign y4088 = n15645 ;
  assign y4089 = n15649 ;
  assign y4090 = n15655 ;
  assign y4091 = n15664 ;
  assign y4092 = ~n15665 ;
  assign y4093 = ~n15671 ;
  assign y4094 = n15682 ;
  assign y4095 = n15687 ;
  assign y4096 = ~n15691 ;
  assign y4097 = ~1'b0 ;
  assign y4098 = n15693 ;
  assign y4099 = n15696 ;
  assign y4100 = ~1'b0 ;
  assign y4101 = ~n15699 ;
  assign y4102 = ~n15700 ;
  assign y4103 = ~n15701 ;
  assign y4104 = ~n15704 ;
  assign y4105 = ~n15707 ;
  assign y4106 = ~1'b0 ;
  assign y4107 = n15708 ;
  assign y4108 = n15710 ;
  assign y4109 = n15717 ;
  assign y4110 = n15718 ;
  assign y4111 = ~1'b0 ;
  assign y4112 = ~n15721 ;
  assign y4113 = ~n15722 ;
  assign y4114 = ~1'b0 ;
  assign y4115 = ~1'b0 ;
  assign y4116 = ~n15732 ;
  assign y4117 = ~n15733 ;
  assign y4118 = ~n15734 ;
  assign y4119 = n15736 ;
  assign y4120 = ~n15738 ;
  assign y4121 = ~n15748 ;
  assign y4122 = ~n15752 ;
  assign y4123 = n10052 ;
  assign y4124 = ~n15755 ;
  assign y4125 = n15757 ;
  assign y4126 = n15760 ;
  assign y4127 = n15762 ;
  assign y4128 = ~n15768 ;
  assign y4129 = ~n15773 ;
  assign y4130 = n15774 ;
  assign y4131 = n15779 ;
  assign y4132 = n15780 ;
  assign y4133 = n15782 ;
  assign y4134 = n15784 ;
  assign y4135 = ~n15790 ;
  assign y4136 = ~1'b0 ;
  assign y4137 = ~1'b0 ;
  assign y4138 = n15793 ;
  assign y4139 = n15796 ;
  assign y4140 = ~n15797 ;
  assign y4141 = ~n15801 ;
  assign y4142 = n15804 ;
  assign y4143 = ~n15817 ;
  assign y4144 = ~n15819 ;
  assign y4145 = n15820 ;
  assign y4146 = n15824 ;
  assign y4147 = ~n15828 ;
  assign y4148 = n15830 ;
  assign y4149 = n15837 ;
  assign y4150 = ~n3021 ;
  assign y4151 = n15843 ;
  assign y4152 = n15848 ;
  assign y4153 = ~n15857 ;
  assign y4154 = ~n15860 ;
  assign y4155 = n15864 ;
  assign y4156 = ~n15869 ;
  assign y4157 = n15870 ;
  assign y4158 = ~n15872 ;
  assign y4159 = n15874 ;
  assign y4160 = ~1'b0 ;
  assign y4161 = ~n15882 ;
  assign y4162 = ~n15887 ;
  assign y4163 = ~n15893 ;
  assign y4164 = n15897 ;
  assign y4165 = ~n15901 ;
  assign y4166 = n15902 ;
  assign y4167 = n15905 ;
  assign y4168 = n15912 ;
  assign y4169 = ~n15920 ;
  assign y4170 = ~n15922 ;
  assign y4171 = ~n15926 ;
  assign y4172 = n15933 ;
  assign y4173 = n15937 ;
  assign y4174 = ~n15938 ;
  assign y4175 = ~1'b0 ;
  assign y4176 = ~n15947 ;
  assign y4177 = n15948 ;
  assign y4178 = ~n15951 ;
  assign y4179 = n15956 ;
  assign y4180 = n15960 ;
  assign y4181 = n15969 ;
  assign y4182 = n15970 ;
  assign y4183 = ~1'b0 ;
  assign y4184 = ~1'b0 ;
  assign y4185 = ~n15971 ;
  assign y4186 = n15975 ;
  assign y4187 = n15982 ;
  assign y4188 = n15987 ;
  assign y4189 = ~1'b0 ;
  assign y4190 = ~n15990 ;
  assign y4191 = ~n15991 ;
  assign y4192 = n15992 ;
  assign y4193 = ~n16004 ;
  assign y4194 = n16005 ;
  assign y4195 = ~n16008 ;
  assign y4196 = n16010 ;
  assign y4197 = ~n16013 ;
  assign y4198 = n16017 ;
  assign y4199 = n16018 ;
  assign y4200 = ~n16024 ;
  assign y4201 = n16036 ;
  assign y4202 = ~n16037 ;
  assign y4203 = n16053 ;
  assign y4204 = ~n16058 ;
  assign y4205 = ~n16065 ;
  assign y4206 = n16073 ;
  assign y4207 = n13320 ;
  assign y4208 = n16074 ;
  assign y4209 = ~1'b0 ;
  assign y4210 = n16075 ;
  assign y4211 = n16079 ;
  assign y4212 = ~n16081 ;
  assign y4213 = ~n16087 ;
  assign y4214 = ~n16088 ;
  assign y4215 = n16090 ;
  assign y4216 = n16093 ;
  assign y4217 = ~n16097 ;
  assign y4218 = n16099 ;
  assign y4219 = n16100 ;
  assign y4220 = n16101 ;
  assign y4221 = n16104 ;
  assign y4222 = ~1'b0 ;
  assign y4223 = n16112 ;
  assign y4224 = n16115 ;
  assign y4225 = ~1'b0 ;
  assign y4226 = ~n16119 ;
  assign y4227 = ~n16122 ;
  assign y4228 = n16128 ;
  assign y4229 = n16133 ;
  assign y4230 = n16137 ;
  assign y4231 = n16138 ;
  assign y4232 = n16140 ;
  assign y4233 = n16141 ;
  assign y4234 = ~n16142 ;
  assign y4235 = n16146 ;
  assign y4236 = ~n16148 ;
  assign y4237 = n16152 ;
  assign y4238 = ~n16154 ;
  assign y4239 = n16157 ;
  assign y4240 = ~n16166 ;
  assign y4241 = ~1'b0 ;
  assign y4242 = ~n16170 ;
  assign y4243 = ~n16173 ;
  assign y4244 = n16182 ;
  assign y4245 = ~n16183 ;
  assign y4246 = ~n16189 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = n16190 ;
  assign y4249 = ~n16195 ;
  assign y4250 = ~n16201 ;
  assign y4251 = ~n16206 ;
  assign y4252 = ~1'b0 ;
  assign y4253 = ~1'b0 ;
  assign y4254 = ~n16208 ;
  assign y4255 = n16218 ;
  assign y4256 = ~n16229 ;
  assign y4257 = n16233 ;
  assign y4258 = ~1'b0 ;
  assign y4259 = ~1'b0 ;
  assign y4260 = ~n16238 ;
  assign y4261 = ~n16241 ;
  assign y4262 = ~n16260 ;
  assign y4263 = n12296 ;
  assign y4264 = ~n16262 ;
  assign y4265 = n16263 ;
  assign y4266 = n16265 ;
  assign y4267 = ~n16270 ;
  assign y4268 = ~n16277 ;
  assign y4269 = ~n16278 ;
  assign y4270 = n16279 ;
  assign y4271 = n16280 ;
  assign y4272 = n16281 ;
  assign y4273 = n5710 ;
  assign y4274 = ~n16283 ;
  assign y4275 = ~n16285 ;
  assign y4276 = n16286 ;
  assign y4277 = ~n16290 ;
  assign y4278 = ~n16293 ;
  assign y4279 = ~1'b0 ;
  assign y4280 = n16298 ;
  assign y4281 = ~n16300 ;
  assign y4282 = n16301 ;
  assign y4283 = n16303 ;
  assign y4284 = n16305 ;
  assign y4285 = n16306 ;
  assign y4286 = n16309 ;
  assign y4287 = n16312 ;
  assign y4288 = ~1'b0 ;
  assign y4289 = n16320 ;
  assign y4290 = n16322 ;
  assign y4291 = n16323 ;
  assign y4292 = ~n16324 ;
  assign y4293 = ~n16336 ;
  assign y4294 = n16340 ;
  assign y4295 = n16342 ;
  assign y4296 = ~n16358 ;
  assign y4297 = ~n16363 ;
  assign y4298 = n16366 ;
  assign y4299 = n16373 ;
  assign y4300 = ~n16374 ;
  assign y4301 = ~n16377 ;
  assign y4302 = ~n16380 ;
  assign y4303 = ~n16384 ;
  assign y4304 = ~1'b0 ;
  assign y4305 = ~n16385 ;
  assign y4306 = ~n16387 ;
  assign y4307 = ~n16391 ;
  assign y4308 = n16398 ;
  assign y4309 = ~1'b0 ;
  assign y4310 = n16401 ;
  assign y4311 = ~n16409 ;
  assign y4312 = n16416 ;
  assign y4313 = ~n16426 ;
  assign y4314 = n16431 ;
  assign y4315 = ~n16432 ;
  assign y4316 = ~1'b0 ;
  assign y4317 = ~n16438 ;
  assign y4318 = ~n16439 ;
  assign y4319 = 1'b0 ;
  assign y4320 = ~n16443 ;
  assign y4321 = n16447 ;
  assign y4322 = ~n16456 ;
  assign y4323 = ~n16461 ;
  assign y4324 = ~n16465 ;
  assign y4325 = n16467 ;
  assign y4326 = n16468 ;
  assign y4327 = n16470 ;
  assign y4328 = n16474 ;
  assign y4329 = n16477 ;
  assign y4330 = ~n16480 ;
  assign y4331 = ~1'b0 ;
  assign y4332 = ~n16483 ;
  assign y4333 = n16489 ;
  assign y4334 = n16492 ;
  assign y4335 = n16493 ;
  assign y4336 = n16500 ;
  assign y4337 = n16502 ;
  assign y4338 = ~n16511 ;
  assign y4339 = ~1'b0 ;
  assign y4340 = ~1'b0 ;
  assign y4341 = ~n16516 ;
  assign y4342 = ~1'b0 ;
  assign y4343 = ~1'b0 ;
  assign y4344 = n16518 ;
  assign y4345 = ~n6418 ;
  assign y4346 = ~n16519 ;
  assign y4347 = ~n16522 ;
  assign y4348 = ~n16524 ;
  assign y4349 = ~n16529 ;
  assign y4350 = ~n16535 ;
  assign y4351 = ~n16538 ;
  assign y4352 = ~n16539 ;
  assign y4353 = n16545 ;
  assign y4354 = n16549 ;
  assign y4355 = ~n16550 ;
  assign y4356 = n16554 ;
  assign y4357 = ~n16555 ;
  assign y4358 = ~n16557 ;
  assign y4359 = ~n16566 ;
  assign y4360 = ~n16568 ;
  assign y4361 = ~n16569 ;
  assign y4362 = ~n16571 ;
  assign y4363 = ~n16572 ;
  assign y4364 = n16578 ;
  assign y4365 = ~1'b0 ;
  assign y4366 = n16590 ;
  assign y4367 = ~n16592 ;
  assign y4368 = ~n16596 ;
  assign y4369 = ~n16600 ;
  assign y4370 = n16607 ;
  assign y4371 = n16609 ;
  assign y4372 = n16610 ;
  assign y4373 = n16611 ;
  assign y4374 = ~1'b0 ;
  assign y4375 = ~n16619 ;
  assign y4376 = ~n16620 ;
  assign y4377 = ~n16621 ;
  assign y4378 = n16624 ;
  assign y4379 = n16626 ;
  assign y4380 = n16628 ;
  assign y4381 = ~n16629 ;
  assign y4382 = ~n16636 ;
  assign y4383 = n16637 ;
  assign y4384 = n16643 ;
  assign y4385 = ~1'b0 ;
  assign y4386 = ~1'b0 ;
  assign y4387 = ~n16652 ;
  assign y4388 = ~n16657 ;
  assign y4389 = ~n16665 ;
  assign y4390 = n16673 ;
  assign y4391 = ~n16678 ;
  assign y4392 = ~1'b0 ;
  assign y4393 = ~n16682 ;
  assign y4394 = n16693 ;
  assign y4395 = ~n16695 ;
  assign y4396 = n16697 ;
  assign y4397 = ~1'b0 ;
  assign y4398 = n16698 ;
  assign y4399 = ~n16699 ;
  assign y4400 = ~n16708 ;
  assign y4401 = n16710 ;
  assign y4402 = ~n16716 ;
  assign y4403 = n16719 ;
  assign y4404 = n16721 ;
  assign y4405 = n16723 ;
  assign y4406 = ~n16727 ;
  assign y4407 = n16731 ;
  assign y4408 = n16739 ;
  assign y4409 = ~n16748 ;
  assign y4410 = n16749 ;
  assign y4411 = ~n16750 ;
  assign y4412 = ~1'b0 ;
  assign y4413 = ~n16751 ;
  assign y4414 = n16756 ;
  assign y4415 = ~n16757 ;
  assign y4416 = ~n16761 ;
  assign y4417 = ~1'b0 ;
  assign y4418 = ~1'b0 ;
  assign y4419 = n16769 ;
  assign y4420 = n16772 ;
  assign y4421 = n16777 ;
  assign y4422 = ~n16778 ;
  assign y4423 = ~n16779 ;
  assign y4424 = ~n16793 ;
  assign y4425 = ~n16794 ;
  assign y4426 = ~n16797 ;
  assign y4427 = ~n16799 ;
  assign y4428 = ~n16800 ;
  assign y4429 = ~n16802 ;
  assign y4430 = ~n16803 ;
  assign y4431 = ~n16804 ;
  assign y4432 = ~n16805 ;
  assign y4433 = ~n16806 ;
  assign y4434 = ~n16807 ;
  assign y4435 = n16808 ;
  assign y4436 = n16809 ;
  assign y4437 = ~n16810 ;
  assign y4438 = ~n16812 ;
  assign y4439 = n16816 ;
  assign y4440 = n16817 ;
  assign y4441 = n16819 ;
  assign y4442 = n16821 ;
  assign y4443 = n16823 ;
  assign y4444 = ~n16825 ;
  assign y4445 = n16826 ;
  assign y4446 = n16828 ;
  assign y4447 = n16834 ;
  assign y4448 = n16836 ;
  assign y4449 = n2282 ;
  assign y4450 = ~n16848 ;
  assign y4451 = ~n16850 ;
  assign y4452 = ~n16852 ;
  assign y4453 = ~n16854 ;
  assign y4454 = ~n16855 ;
  assign y4455 = ~n7732 ;
  assign y4456 = ~n16860 ;
  assign y4457 = ~n16861 ;
  assign y4458 = n16862 ;
  assign y4459 = ~n16865 ;
  assign y4460 = n16872 ;
  assign y4461 = ~n16878 ;
  assign y4462 = ~n16880 ;
  assign y4463 = ~n16884 ;
  assign y4464 = ~1'b0 ;
  assign y4465 = n16889 ;
  assign y4466 = n16893 ;
  assign y4467 = n16902 ;
  assign y4468 = n16915 ;
  assign y4469 = n16919 ;
  assign y4470 = ~n16933 ;
  assign y4471 = ~n16939 ;
  assign y4472 = ~n16940 ;
  assign y4473 = ~n16953 ;
  assign y4474 = n16960 ;
  assign y4475 = n16965 ;
  assign y4476 = n16973 ;
  assign y4477 = n16975 ;
  assign y4478 = ~n16982 ;
  assign y4479 = ~1'b0 ;
  assign y4480 = n16987 ;
  assign y4481 = ~n16990 ;
  assign y4482 = ~n16996 ;
  assign y4483 = n16998 ;
  assign y4484 = ~n17001 ;
  assign y4485 = n17003 ;
  assign y4486 = n17005 ;
  assign y4487 = n17009 ;
  assign y4488 = ~1'b0 ;
  assign y4489 = n17014 ;
  assign y4490 = n17028 ;
  assign y4491 = ~n17032 ;
  assign y4492 = n17034 ;
  assign y4493 = ~n17035 ;
  assign y4494 = ~n17040 ;
  assign y4495 = ~1'b0 ;
  assign y4496 = ~n17050 ;
  assign y4497 = ~1'b0 ;
  assign y4498 = ~1'b0 ;
  assign y4499 = ~1'b0 ;
  assign y4500 = ~n17052 ;
  assign y4501 = ~n17056 ;
  assign y4502 = ~n17060 ;
  assign y4503 = ~n17063 ;
  assign y4504 = ~1'b0 ;
  assign y4505 = n17068 ;
  assign y4506 = ~n17071 ;
  assign y4507 = n17074 ;
  assign y4508 = n17083 ;
  assign y4509 = ~n17085 ;
  assign y4510 = ~1'b0 ;
  assign y4511 = ~1'b0 ;
  assign y4512 = ~n17089 ;
  assign y4513 = ~n17092 ;
  assign y4514 = ~n17094 ;
  assign y4515 = ~n5818 ;
  assign y4516 = ~1'b0 ;
  assign y4517 = ~n17095 ;
  assign y4518 = n17096 ;
  assign y4519 = ~n17099 ;
  assign y4520 = n17101 ;
  assign y4521 = n17102 ;
  assign y4522 = n17105 ;
  assign y4523 = ~n17107 ;
  assign y4524 = n17108 ;
  assign y4525 = n17109 ;
  assign y4526 = ~n17111 ;
  assign y4527 = ~1'b0 ;
  assign y4528 = n17113 ;
  assign y4529 = ~n17130 ;
  assign y4530 = ~n17133 ;
  assign y4531 = ~n17138 ;
  assign y4532 = ~n17142 ;
  assign y4533 = n17143 ;
  assign y4534 = n17149 ;
  assign y4535 = n17153 ;
  assign y4536 = n17158 ;
  assign y4537 = ~n17161 ;
  assign y4538 = n17167 ;
  assign y4539 = ~n17173 ;
  assign y4540 = ~n17175 ;
  assign y4541 = n17176 ;
  assign y4542 = n17182 ;
  assign y4543 = ~1'b0 ;
  assign y4544 = n17187 ;
  assign y4545 = ~n17192 ;
  assign y4546 = n17200 ;
  assign y4547 = n17209 ;
  assign y4548 = n17210 ;
  assign y4549 = n17215 ;
  assign y4550 = n17217 ;
  assign y4551 = n17220 ;
  assign y4552 = n17221 ;
  assign y4553 = ~n17231 ;
  assign y4554 = n17234 ;
  assign y4555 = ~n17241 ;
  assign y4556 = ~n17247 ;
  assign y4557 = ~n17250 ;
  assign y4558 = ~n17254 ;
  assign y4559 = n17256 ;
  assign y4560 = ~n17261 ;
  assign y4561 = n17269 ;
  assign y4562 = ~n17271 ;
  assign y4563 = ~n8548 ;
  assign y4564 = n17276 ;
  assign y4565 = n17281 ;
  assign y4566 = n17282 ;
  assign y4567 = ~n17290 ;
  assign y4568 = ~n17296 ;
  assign y4569 = ~n17300 ;
  assign y4570 = n17302 ;
  assign y4571 = ~n17304 ;
  assign y4572 = n17310 ;
  assign y4573 = n17312 ;
  assign y4574 = n17317 ;
  assign y4575 = ~n17328 ;
  assign y4576 = n17332 ;
  assign y4577 = ~n17334 ;
  assign y4578 = ~1'b0 ;
  assign y4579 = n17341 ;
  assign y4580 = ~n17347 ;
  assign y4581 = ~n17348 ;
  assign y4582 = n17357 ;
  assign y4583 = n17362 ;
  assign y4584 = ~n17365 ;
  assign y4585 = ~n17366 ;
  assign y4586 = ~n17375 ;
  assign y4587 = ~n17378 ;
  assign y4588 = n17380 ;
  assign y4589 = ~n17383 ;
  assign y4590 = n17388 ;
  assign y4591 = n17390 ;
  assign y4592 = ~n17392 ;
  assign y4593 = ~1'b0 ;
  assign y4594 = n17399 ;
  assign y4595 = ~n17401 ;
  assign y4596 = ~n17407 ;
  assign y4597 = n17409 ;
  assign y4598 = ~n17417 ;
  assign y4599 = ~n17418 ;
  assign y4600 = ~n17420 ;
  assign y4601 = n17428 ;
  assign y4602 = n17429 ;
  assign y4603 = ~1'b0 ;
  assign y4604 = ~n17437 ;
  assign y4605 = n17441 ;
  assign y4606 = n17452 ;
  assign y4607 = ~n17458 ;
  assign y4608 = n17459 ;
  assign y4609 = ~n17464 ;
  assign y4610 = ~1'b0 ;
  assign y4611 = n17467 ;
  assign y4612 = n17484 ;
  assign y4613 = ~n17491 ;
  assign y4614 = n17495 ;
  assign y4615 = ~1'b0 ;
  assign y4616 = n17501 ;
  assign y4617 = n17504 ;
  assign y4618 = ~1'b0 ;
  assign y4619 = ~n17505 ;
  assign y4620 = ~n17508 ;
  assign y4621 = n17517 ;
  assign y4622 = n17521 ;
  assign y4623 = n17524 ;
  assign y4624 = ~n17527 ;
  assign y4625 = ~n17533 ;
  assign y4626 = n17536 ;
  assign y4627 = ~1'b0 ;
  assign y4628 = ~n17537 ;
  assign y4629 = ~n17550 ;
  assign y4630 = ~n17551 ;
  assign y4631 = n17559 ;
  assign y4632 = n17560 ;
  assign y4633 = ~n17563 ;
  assign y4634 = n17565 ;
  assign y4635 = ~n17567 ;
  assign y4636 = n17575 ;
  assign y4637 = ~n17580 ;
  assign y4638 = n17587 ;
  assign y4639 = ~n17588 ;
  assign y4640 = n17589 ;
  assign y4641 = n17591 ;
  assign y4642 = ~n17597 ;
  assign y4643 = ~n17602 ;
  assign y4644 = ~1'b0 ;
  assign y4645 = ~n17603 ;
  assign y4646 = ~n17605 ;
  assign y4647 = ~n17606 ;
  assign y4648 = n17620 ;
  assign y4649 = n17623 ;
  assign y4650 = ~1'b0 ;
  assign y4651 = n17625 ;
  assign y4652 = ~n17630 ;
  assign y4653 = n17633 ;
  assign y4654 = ~n17643 ;
  assign y4655 = ~n17646 ;
  assign y4656 = ~n17647 ;
  assign y4657 = n17648 ;
  assign y4658 = ~n17649 ;
  assign y4659 = ~n17651 ;
  assign y4660 = ~1'b0 ;
  assign y4661 = ~1'b0 ;
  assign y4662 = ~n17654 ;
  assign y4663 = ~n17660 ;
  assign y4664 = n17664 ;
  assign y4665 = ~1'b0 ;
  assign y4666 = ~n17667 ;
  assign y4667 = n17672 ;
  assign y4668 = n17676 ;
  assign y4669 = n17677 ;
  assign y4670 = ~n17683 ;
  assign y4671 = ~n17684 ;
  assign y4672 = ~1'b0 ;
  assign y4673 = n17685 ;
  assign y4674 = ~n17689 ;
  assign y4675 = n17690 ;
  assign y4676 = n17691 ;
  assign y4677 = n17694 ;
  assign y4678 = n17702 ;
  assign y4679 = ~n17704 ;
  assign y4680 = n17708 ;
  assign y4681 = ~n17711 ;
  assign y4682 = ~n17715 ;
  assign y4683 = ~n17716 ;
  assign y4684 = ~1'b0 ;
  assign y4685 = ~n17717 ;
  assign y4686 = n17718 ;
  assign y4687 = ~n17721 ;
  assign y4688 = n17729 ;
  assign y4689 = n17734 ;
  assign y4690 = n17736 ;
  assign y4691 = n17741 ;
  assign y4692 = ~n17745 ;
  assign y4693 = ~n17747 ;
  assign y4694 = n17754 ;
  assign y4695 = n17758 ;
  assign y4696 = n17759 ;
  assign y4697 = ~n17764 ;
  assign y4698 = n17766 ;
  assign y4699 = n17772 ;
  assign y4700 = n17774 ;
  assign y4701 = n17776 ;
  assign y4702 = n17777 ;
  assign y4703 = n17780 ;
  assign y4704 = ~1'b0 ;
  assign y4705 = n17785 ;
  assign y4706 = n17792 ;
  assign y4707 = n17794 ;
  assign y4708 = n17802 ;
  assign y4709 = ~n10621 ;
  assign y4710 = n17806 ;
  assign y4711 = ~n3546 ;
  assign y4712 = ~1'b0 ;
  assign y4713 = ~n17809 ;
  assign y4714 = ~n17810 ;
  assign y4715 = ~n17818 ;
  assign y4716 = n17823 ;
  assign y4717 = ~n17827 ;
  assign y4718 = ~n17835 ;
  assign y4719 = n17839 ;
  assign y4720 = ~1'b0 ;
  assign y4721 = n17841 ;
  assign y4722 = ~1'b0 ;
  assign y4723 = n17845 ;
  assign y4724 = ~n17846 ;
  assign y4725 = ~1'b0 ;
  assign y4726 = ~n17849 ;
  assign y4727 = n17854 ;
  assign y4728 = n17857 ;
  assign y4729 = ~1'b0 ;
  assign y4730 = n17864 ;
  assign y4731 = ~n17865 ;
  assign y4732 = ~1'b0 ;
  assign y4733 = n17868 ;
  assign y4734 = ~n1988 ;
  assign y4735 = n17869 ;
  assign y4736 = ~n17871 ;
  assign y4737 = ~n17873 ;
  assign y4738 = n17875 ;
  assign y4739 = n17877 ;
  assign y4740 = ~n17886 ;
  assign y4741 = ~n17894 ;
  assign y4742 = ~n17896 ;
  assign y4743 = n17901 ;
  assign y4744 = ~n17903 ;
  assign y4745 = n17917 ;
  assign y4746 = ~n17920 ;
  assign y4747 = n17929 ;
  assign y4748 = n17930 ;
  assign y4749 = ~n17933 ;
  assign y4750 = ~n17934 ;
  assign y4751 = ~n17935 ;
  assign y4752 = ~n17942 ;
  assign y4753 = n17953 ;
  assign y4754 = n17961 ;
  assign y4755 = n17964 ;
  assign y4756 = n17970 ;
  assign y4757 = n17981 ;
  assign y4758 = ~n17984 ;
  assign y4759 = n17989 ;
  assign y4760 = n17992 ;
  assign y4761 = ~n17995 ;
  assign y4762 = ~n17997 ;
  assign y4763 = ~n18002 ;
  assign y4764 = ~n18016 ;
  assign y4765 = ~n18024 ;
  assign y4766 = ~n18027 ;
  assign y4767 = ~1'b0 ;
  assign y4768 = ~n18028 ;
  assign y4769 = n18032 ;
  assign y4770 = ~1'b0 ;
  assign y4771 = ~n18034 ;
  assign y4772 = ~n18045 ;
  assign y4773 = n18048 ;
  assign y4774 = n18049 ;
  assign y4775 = n18051 ;
  assign y4776 = ~n18054 ;
  assign y4777 = n18060 ;
  assign y4778 = n18063 ;
  assign y4779 = ~n18068 ;
  assign y4780 = n18078 ;
  assign y4781 = ~n18094 ;
  assign y4782 = ~1'b0 ;
  assign y4783 = ~n18098 ;
  assign y4784 = ~n18102 ;
  assign y4785 = ~n18103 ;
  assign y4786 = ~n18107 ;
  assign y4787 = n18109 ;
  assign y4788 = ~n18113 ;
  assign y4789 = ~n18114 ;
  assign y4790 = n18119 ;
  assign y4791 = n18121 ;
  assign y4792 = n18127 ;
  assign y4793 = n5927 ;
  assign y4794 = ~n18128 ;
  assign y4795 = n18135 ;
  assign y4796 = ~1'b0 ;
  assign y4797 = ~1'b0 ;
  assign y4798 = ~n18139 ;
  assign y4799 = ~1'b0 ;
  assign y4800 = ~1'b0 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = n18141 ;
  assign y4803 = ~n18145 ;
  assign y4804 = n18148 ;
  assign y4805 = ~1'b0 ;
  assign y4806 = n18155 ;
  assign y4807 = n18158 ;
  assign y4808 = ~1'b0 ;
  assign y4809 = ~n18162 ;
  assign y4810 = ~n18164 ;
  assign y4811 = n18171 ;
  assign y4812 = ~n18178 ;
  assign y4813 = ~n18181 ;
  assign y4814 = ~n18185 ;
  assign y4815 = ~n18189 ;
  assign y4816 = ~n18196 ;
  assign y4817 = ~n3615 ;
  assign y4818 = ~n17110 ;
  assign y4819 = ~1'b0 ;
  assign y4820 = n18202 ;
  assign y4821 = n18203 ;
  assign y4822 = n18208 ;
  assign y4823 = ~n18210 ;
  assign y4824 = ~n18212 ;
  assign y4825 = ~n18214 ;
  assign y4826 = n18219 ;
  assign y4827 = ~1'b0 ;
  assign y4828 = ~n18220 ;
  assign y4829 = ~n18222 ;
  assign y4830 = n18224 ;
  assign y4831 = n18234 ;
  assign y4832 = ~n18238 ;
  assign y4833 = n18244 ;
  assign y4834 = ~n18247 ;
  assign y4835 = ~n18251 ;
  assign y4836 = ~n18252 ;
  assign y4837 = n18261 ;
  assign y4838 = 1'b0 ;
  assign y4839 = ~n18263 ;
  assign y4840 = n18270 ;
  assign y4841 = ~n18271 ;
  assign y4842 = ~1'b0 ;
  assign y4843 = n18273 ;
  assign y4844 = ~1'b0 ;
  assign y4845 = n18283 ;
  assign y4846 = n18286 ;
  assign y4847 = ~n18289 ;
  assign y4848 = ~n18291 ;
  assign y4849 = ~n18292 ;
  assign y4850 = n18296 ;
  assign y4851 = n18303 ;
  assign y4852 = ~n18305 ;
  assign y4853 = ~n18316 ;
  assign y4854 = ~1'b0 ;
  assign y4855 = ~1'b0 ;
  assign y4856 = ~1'b0 ;
  assign y4857 = ~1'b0 ;
  assign y4858 = ~n18317 ;
  assign y4859 = n18319 ;
  assign y4860 = n18324 ;
  assign y4861 = n18331 ;
  assign y4862 = ~n18336 ;
  assign y4863 = n18338 ;
  assign y4864 = ~n18339 ;
  assign y4865 = ~1'b0 ;
  assign y4866 = ~n18340 ;
  assign y4867 = 1'b0 ;
  assign y4868 = ~n18344 ;
  assign y4869 = ~1'b0 ;
  assign y4870 = n18347 ;
  assign y4871 = n18351 ;
  assign y4872 = ~1'b0 ;
  assign y4873 = ~n18357 ;
  assign y4874 = n18360 ;
  assign y4875 = ~1'b0 ;
  assign y4876 = ~1'b0 ;
  assign y4877 = ~n18362 ;
  assign y4878 = n18364 ;
  assign y4879 = ~n18365 ;
  assign y4880 = 1'b0 ;
  assign y4881 = n18369 ;
  assign y4882 = ~n18373 ;
  assign y4883 = n18377 ;
  assign y4884 = ~n18387 ;
  assign y4885 = ~n1396 ;
  assign y4886 = n18390 ;
  assign y4887 = n18395 ;
  assign y4888 = n18396 ;
  assign y4889 = n18397 ;
  assign y4890 = ~1'b0 ;
  assign y4891 = ~1'b0 ;
  assign y4892 = ~n18399 ;
  assign y4893 = ~n18400 ;
  assign y4894 = ~n18406 ;
  assign y4895 = ~1'b0 ;
  assign y4896 = ~n18408 ;
  assign y4897 = n18409 ;
  assign y4898 = ~n18411 ;
  assign y4899 = ~n18415 ;
  assign y4900 = ~n18417 ;
  assign y4901 = n18419 ;
  assign y4902 = n18420 ;
  assign y4903 = n18426 ;
  assign y4904 = ~n18431 ;
  assign y4905 = n18433 ;
  assign y4906 = n18437 ;
  assign y4907 = n18438 ;
  assign y4908 = ~n18444 ;
  assign y4909 = n18446 ;
  assign y4910 = n18448 ;
  assign y4911 = n18449 ;
  assign y4912 = n18451 ;
  assign y4913 = ~1'b0 ;
  assign y4914 = ~1'b0 ;
  assign y4915 = n18459 ;
  assign y4916 = ~n18462 ;
  assign y4917 = n18480 ;
  assign y4918 = ~1'b0 ;
  assign y4919 = ~n18482 ;
  assign y4920 = ~n18489 ;
  assign y4921 = ~n18492 ;
  assign y4922 = ~n18497 ;
  assign y4923 = n18503 ;
  assign y4924 = n18507 ;
  assign y4925 = ~1'b0 ;
  assign y4926 = ~n18511 ;
  assign y4927 = n18512 ;
  assign y4928 = ~1'b0 ;
  assign y4929 = 1'b0 ;
  assign y4930 = n18522 ;
  assign y4931 = n18526 ;
  assign y4932 = ~1'b0 ;
  assign y4933 = n18529 ;
  assign y4934 = ~1'b0 ;
  assign y4935 = ~1'b0 ;
  assign y4936 = n18531 ;
  assign y4937 = ~n18535 ;
  assign y4938 = ~n18538 ;
  assign y4939 = n18539 ;
  assign y4940 = n18546 ;
  assign y4941 = n18548 ;
  assign y4942 = ~1'b0 ;
  assign y4943 = n18551 ;
  assign y4944 = ~1'b0 ;
  assign y4945 = ~n18554 ;
  assign y4946 = ~n18556 ;
  assign y4947 = n18557 ;
  assign y4948 = n18562 ;
  assign y4949 = n18566 ;
  assign y4950 = ~1'b0 ;
  assign y4951 = ~n18572 ;
  assign y4952 = ~n18583 ;
  assign y4953 = ~n18585 ;
  assign y4954 = n18595 ;
  assign y4955 = ~n18596 ;
  assign y4956 = n18599 ;
  assign y4957 = 1'b0 ;
  assign y4958 = n18602 ;
  assign y4959 = ~n18607 ;
  assign y4960 = ~n18614 ;
  assign y4961 = n18618 ;
  assign y4962 = ~1'b0 ;
  assign y4963 = ~n18621 ;
  assign y4964 = n18625 ;
  assign y4965 = ~n18636 ;
  assign y4966 = ~1'b0 ;
  assign y4967 = n18640 ;
  assign y4968 = ~n18642 ;
  assign y4969 = ~n18647 ;
  assign y4970 = ~n18649 ;
  assign y4971 = n18652 ;
  assign y4972 = ~n18656 ;
  assign y4973 = ~n18657 ;
  assign y4974 = n18660 ;
  assign y4975 = n18664 ;
  assign y4976 = n18668 ;
  assign y4977 = ~n18669 ;
  assign y4978 = n18673 ;
  assign y4979 = n18683 ;
  assign y4980 = ~n18689 ;
  assign y4981 = ~n18691 ;
  assign y4982 = n18692 ;
  assign y4983 = n18700 ;
  assign y4984 = ~n18701 ;
  assign y4985 = n18705 ;
  assign y4986 = ~1'b0 ;
  assign y4987 = ~n18706 ;
  assign y4988 = ~n18708 ;
  assign y4989 = n18709 ;
  assign y4990 = n18714 ;
  assign y4991 = ~n18717 ;
  assign y4992 = n18719 ;
  assign y4993 = ~n18723 ;
  assign y4994 = n18725 ;
  assign y4995 = n18735 ;
  assign y4996 = ~n18738 ;
  assign y4997 = ~n18739 ;
  assign y4998 = n18741 ;
  assign y4999 = ~n18742 ;
  assign y5000 = n18743 ;
  assign y5001 = ~n18748 ;
  assign y5002 = ~n18749 ;
  assign y5003 = n18750 ;
  assign y5004 = ~1'b0 ;
  assign y5005 = n18758 ;
  assign y5006 = n18759 ;
  assign y5007 = ~n18761 ;
  assign y5008 = ~n18763 ;
  assign y5009 = ~n18764 ;
  assign y5010 = n18770 ;
  assign y5011 = n18781 ;
  assign y5012 = n18787 ;
  assign y5013 = n18788 ;
  assign y5014 = ~n18791 ;
  assign y5015 = n18793 ;
  assign y5016 = n18796 ;
  assign y5017 = n18798 ;
  assign y5018 = n18806 ;
  assign y5019 = ~n18814 ;
  assign y5020 = n18816 ;
  assign y5021 = ~n18817 ;
  assign y5022 = n18820 ;
  assign y5023 = n18822 ;
  assign y5024 = n18824 ;
  assign y5025 = n18825 ;
  assign y5026 = ~1'b0 ;
  assign y5027 = ~1'b0 ;
  assign y5028 = n18828 ;
  assign y5029 = ~n18834 ;
  assign y5030 = ~n18840 ;
  assign y5031 = ~1'b0 ;
  assign y5032 = ~1'b0 ;
  assign y5033 = ~1'b0 ;
  assign y5034 = ~n18848 ;
  assign y5035 = n18864 ;
  assign y5036 = ~n18869 ;
  assign y5037 = n18876 ;
  assign y5038 = ~n18882 ;
  assign y5039 = ~n18886 ;
  assign y5040 = n18888 ;
  assign y5041 = ~n18897 ;
  assign y5042 = n18898 ;
  assign y5043 = ~n18901 ;
  assign y5044 = ~n18904 ;
  assign y5045 = ~1'b0 ;
  assign y5046 = n18906 ;
  assign y5047 = ~n18910 ;
  assign y5048 = n18917 ;
  assign y5049 = n18919 ;
  assign y5050 = n18920 ;
  assign y5051 = ~n18926 ;
  assign y5052 = ~1'b0 ;
  assign y5053 = n18927 ;
  assign y5054 = ~1'b0 ;
  assign y5055 = n18931 ;
  assign y5056 = ~1'b0 ;
  assign y5057 = n18940 ;
  assign y5058 = n18943 ;
  assign y5059 = n18946 ;
  assign y5060 = n18947 ;
  assign y5061 = ~n18954 ;
  assign y5062 = n18955 ;
  assign y5063 = n18957 ;
  assign y5064 = ~n18960 ;
  assign y5065 = n18963 ;
  assign y5066 = n18966 ;
  assign y5067 = ~n18968 ;
  assign y5068 = n18983 ;
  assign y5069 = ~n18984 ;
  assign y5070 = ~1'b0 ;
  assign y5071 = n18987 ;
  assign y5072 = ~n18988 ;
  assign y5073 = n18989 ;
  assign y5074 = ~n18993 ;
  assign y5075 = ~n18994 ;
  assign y5076 = ~n18995 ;
  assign y5077 = n18999 ;
  assign y5078 = n19002 ;
  assign y5079 = ~n19007 ;
  assign y5080 = ~n19013 ;
  assign y5081 = ~1'b0 ;
  assign y5082 = ~n19018 ;
  assign y5083 = n19025 ;
  assign y5084 = ~n19027 ;
  assign y5085 = ~n19031 ;
  assign y5086 = n19032 ;
  assign y5087 = ~n19040 ;
  assign y5088 = ~n19047 ;
  assign y5089 = n19048 ;
  assign y5090 = ~1'b0 ;
  assign y5091 = ~n19054 ;
  assign y5092 = ~1'b0 ;
  assign y5093 = n19059 ;
  assign y5094 = ~n19060 ;
  assign y5095 = n19063 ;
  assign y5096 = ~n19075 ;
  assign y5097 = n19078 ;
  assign y5098 = n19082 ;
  assign y5099 = n19085 ;
  assign y5100 = ~1'b0 ;
  assign y5101 = n19089 ;
  assign y5102 = ~n19090 ;
  assign y5103 = ~n19093 ;
  assign y5104 = n19099 ;
  assign y5105 = ~n19104 ;
  assign y5106 = ~n19105 ;
  assign y5107 = n19109 ;
  assign y5108 = ~1'b0 ;
  assign y5109 = ~n19110 ;
  assign y5110 = ~n19115 ;
  assign y5111 = ~1'b0 ;
  assign y5112 = ~1'b0 ;
  assign y5113 = n19120 ;
  assign y5114 = ~n19126 ;
  assign y5115 = ~1'b0 ;
  assign y5116 = ~n19132 ;
  assign y5117 = n19138 ;
  assign y5118 = ~n19147 ;
  assign y5119 = ~n19150 ;
  assign y5120 = ~n19162 ;
  assign y5121 = n19169 ;
  assign y5122 = n19172 ;
  assign y5123 = ~n19176 ;
  assign y5124 = ~n19179 ;
  assign y5125 = ~n19181 ;
  assign y5126 = n19182 ;
  assign y5127 = ~1'b0 ;
  assign y5128 = n19185 ;
  assign y5129 = ~n19194 ;
  assign y5130 = ~n19198 ;
  assign y5131 = ~1'b0 ;
  assign y5132 = n19204 ;
  assign y5133 = n19206 ;
  assign y5134 = n19207 ;
  assign y5135 = ~n19218 ;
  assign y5136 = ~n19225 ;
  assign y5137 = ~n19226 ;
  assign y5138 = ~n19228 ;
  assign y5139 = ~1'b0 ;
  assign y5140 = ~n19230 ;
  assign y5141 = n19232 ;
  assign y5142 = n19241 ;
  assign y5143 = ~n19249 ;
  assign y5144 = n19256 ;
  assign y5145 = ~1'b0 ;
  assign y5146 = n19261 ;
  assign y5147 = ~n19262 ;
  assign y5148 = n19263 ;
  assign y5149 = ~n19267 ;
  assign y5150 = ~1'b0 ;
  assign y5151 = n19278 ;
  assign y5152 = n19283 ;
  assign y5153 = ~n19286 ;
  assign y5154 = ~n19287 ;
  assign y5155 = n19288 ;
  assign y5156 = ~1'b0 ;
  assign y5157 = ~n19292 ;
  assign y5158 = ~n19293 ;
  assign y5159 = ~n19294 ;
  assign y5160 = n19301 ;
  assign y5161 = n19305 ;
  assign y5162 = n19307 ;
  assign y5163 = ~n19313 ;
  assign y5164 = n19318 ;
  assign y5165 = ~1'b0 ;
  assign y5166 = ~n19320 ;
  assign y5167 = n19321 ;
  assign y5168 = ~n19326 ;
  assign y5169 = ~n19334 ;
  assign y5170 = ~n19335 ;
  assign y5171 = ~n19338 ;
  assign y5172 = ~1'b0 ;
  assign y5173 = n19356 ;
  assign y5174 = n19362 ;
  assign y5175 = ~n19365 ;
  assign y5176 = ~n19366 ;
  assign y5177 = ~n19367 ;
  assign y5178 = ~n19372 ;
  assign y5179 = ~n19375 ;
  assign y5180 = n19380 ;
  assign y5181 = n19385 ;
  assign y5182 = n19387 ;
  assign y5183 = n19390 ;
  assign y5184 = n19394 ;
  assign y5185 = n19396 ;
  assign y5186 = ~n19407 ;
  assign y5187 = ~n19414 ;
  assign y5188 = n5305 ;
  assign y5189 = n19416 ;
  assign y5190 = n19418 ;
  assign y5191 = ~n19421 ;
  assign y5192 = ~1'b0 ;
  assign y5193 = n19429 ;
  assign y5194 = ~n19431 ;
  assign y5195 = n19437 ;
  assign y5196 = n19440 ;
  assign y5197 = ~n19441 ;
  assign y5198 = n19444 ;
  assign y5199 = ~n19447 ;
  assign y5200 = ~n19449 ;
  assign y5201 = n19450 ;
  assign y5202 = ~n19452 ;
  assign y5203 = ~n19457 ;
  assign y5204 = ~1'b0 ;
  assign y5205 = n19462 ;
  assign y5206 = n19468 ;
  assign y5207 = n19473 ;
  assign y5208 = n19475 ;
  assign y5209 = ~1'b0 ;
  assign y5210 = ~1'b0 ;
  assign y5211 = ~n19476 ;
  assign y5212 = ~n19481 ;
  assign y5213 = n19482 ;
  assign y5214 = ~n19483 ;
  assign y5215 = ~n19484 ;
  assign y5216 = ~1'b0 ;
  assign y5217 = n19488 ;
  assign y5218 = ~n19490 ;
  assign y5219 = n19494 ;
  assign y5220 = n19495 ;
  assign y5221 = ~n19504 ;
  assign y5222 = ~1'b0 ;
  assign y5223 = ~n19506 ;
  assign y5224 = ~n19509 ;
  assign y5225 = ~1'b0 ;
  assign y5226 = n19512 ;
  assign y5227 = ~n19513 ;
  assign y5228 = ~n19522 ;
  assign y5229 = n19531 ;
  assign y5230 = n19534 ;
  assign y5231 = n19537 ;
  assign y5232 = ~n19548 ;
  assign y5233 = ~n19549 ;
  assign y5234 = n19550 ;
  assign y5235 = n19553 ;
  assign y5236 = ~n19555 ;
  assign y5237 = ~n19562 ;
  assign y5238 = n19572 ;
  assign y5239 = ~n2208 ;
  assign y5240 = ~n19574 ;
  assign y5241 = n19576 ;
  assign y5242 = n19578 ;
  assign y5243 = n19587 ;
  assign y5244 = ~n15104 ;
  assign y5245 = ~n19591 ;
  assign y5246 = ~n19594 ;
  assign y5247 = n19597 ;
  assign y5248 = ~1'b0 ;
  assign y5249 = n19598 ;
  assign y5250 = ~n19600 ;
  assign y5251 = ~n19608 ;
  assign y5252 = n19609 ;
  assign y5253 = ~1'b0 ;
  assign y5254 = n19618 ;
  assign y5255 = ~n19622 ;
  assign y5256 = n19623 ;
  assign y5257 = ~1'b0 ;
  assign y5258 = ~n19627 ;
  assign y5259 = ~n19644 ;
  assign y5260 = ~n19650 ;
  assign y5261 = ~1'b0 ;
  assign y5262 = ~1'b0 ;
  assign y5263 = n19651 ;
  assign y5264 = ~n19654 ;
  assign y5265 = ~1'b0 ;
  assign y5266 = n19657 ;
  assign y5267 = n19662 ;
  assign y5268 = ~n19668 ;
  assign y5269 = n19673 ;
  assign y5270 = ~n19676 ;
  assign y5271 = ~n19677 ;
  assign y5272 = n19681 ;
  assign y5273 = n19683 ;
  assign y5274 = ~n19684 ;
  assign y5275 = n19686 ;
  assign y5276 = ~1'b0 ;
  assign y5277 = n19690 ;
  assign y5278 = n19694 ;
  assign y5279 = n19696 ;
  assign y5280 = ~n19699 ;
  assign y5281 = n19700 ;
  assign y5282 = ~1'b0 ;
  assign y5283 = n19704 ;
  assign y5284 = ~n19708 ;
  assign y5285 = ~n19715 ;
  assign y5286 = n19718 ;
  assign y5287 = ~n19720 ;
  assign y5288 = ~1'b0 ;
  assign y5289 = n19724 ;
  assign y5290 = n19725 ;
  assign y5291 = n19726 ;
  assign y5292 = ~n19729 ;
  assign y5293 = n19743 ;
  assign y5294 = n19745 ;
  assign y5295 = ~n19747 ;
  assign y5296 = ~n19756 ;
  assign y5297 = ~1'b0 ;
  assign y5298 = n19758 ;
  assign y5299 = ~n19759 ;
  assign y5300 = n19765 ;
  assign y5301 = ~1'b0 ;
  assign y5302 = ~n19770 ;
  assign y5303 = ~1'b0 ;
  assign y5304 = ~n19771 ;
  assign y5305 = n19773 ;
  assign y5306 = ~n19778 ;
  assign y5307 = ~n19781 ;
  assign y5308 = 1'b0 ;
  assign y5309 = n19783 ;
  assign y5310 = n19785 ;
  assign y5311 = ~1'b0 ;
  assign y5312 = ~n19789 ;
  assign y5313 = ~n19790 ;
  assign y5314 = n19793 ;
  assign y5315 = ~n19797 ;
  assign y5316 = n19800 ;
  assign y5317 = n19810 ;
  assign y5318 = n19813 ;
  assign y5319 = n19816 ;
  assign y5320 = ~1'b0 ;
  assign y5321 = ~n19822 ;
  assign y5322 = n19827 ;
  assign y5323 = ~n19836 ;
  assign y5324 = n19843 ;
  assign y5325 = ~n19845 ;
  assign y5326 = n19850 ;
  assign y5327 = ~n19857 ;
  assign y5328 = n19858 ;
  assign y5329 = ~n19860 ;
  assign y5330 = ~n19861 ;
  assign y5331 = ~n7024 ;
  assign y5332 = ~n19863 ;
  assign y5333 = ~n19864 ;
  assign y5334 = n19871 ;
  assign y5335 = ~n19872 ;
  assign y5336 = ~n19876 ;
  assign y5337 = ~n19878 ;
  assign y5338 = ~n19880 ;
  assign y5339 = ~n19883 ;
  assign y5340 = n19887 ;
  assign y5341 = ~n19889 ;
  assign y5342 = ~n19897 ;
  assign y5343 = ~1'b0 ;
  assign y5344 = n19898 ;
  assign y5345 = ~n19899 ;
  assign y5346 = n19902 ;
  assign y5347 = n19903 ;
  assign y5348 = n19912 ;
  assign y5349 = n19914 ;
  assign y5350 = n19916 ;
  assign y5351 = 1'b0 ;
  assign y5352 = n19919 ;
  assign y5353 = ~n19924 ;
  assign y5354 = ~n19927 ;
  assign y5355 = ~n19930 ;
  assign y5356 = ~n19935 ;
  assign y5357 = n19936 ;
  assign y5358 = ~n19940 ;
  assign y5359 = n19942 ;
  assign y5360 = ~1'b0 ;
  assign y5361 = ~n19950 ;
  assign y5362 = ~n19956 ;
  assign y5363 = ~n19957 ;
  assign y5364 = ~n19958 ;
  assign y5365 = ~n19960 ;
  assign y5366 = ~n19962 ;
  assign y5367 = ~n19967 ;
  assign y5368 = n19971 ;
  assign y5369 = ~n19975 ;
  assign y5370 = ~n19978 ;
  assign y5371 = ~n19979 ;
  assign y5372 = n19983 ;
  assign y5373 = ~n19987 ;
  assign y5374 = ~n19990 ;
  assign y5375 = 1'b0 ;
  assign y5376 = n19997 ;
  assign y5377 = ~1'b0 ;
  assign y5378 = n20002 ;
  assign y5379 = ~n20004 ;
  assign y5380 = n20005 ;
  assign y5381 = ~n20007 ;
  assign y5382 = ~n20022 ;
  assign y5383 = n20023 ;
  assign y5384 = ~1'b0 ;
  assign y5385 = n20028 ;
  assign y5386 = ~1'b0 ;
  assign y5387 = n20036 ;
  assign y5388 = n20046 ;
  assign y5389 = ~n20049 ;
  assign y5390 = n18188 ;
  assign y5391 = ~n20050 ;
  assign y5392 = ~n20059 ;
  assign y5393 = n20060 ;
  assign y5394 = ~n20064 ;
  assign y5395 = n20071 ;
  assign y5396 = n20072 ;
  assign y5397 = ~1'b0 ;
  assign y5398 = n20074 ;
  assign y5399 = n20078 ;
  assign y5400 = ~n20083 ;
  assign y5401 = ~n20090 ;
  assign y5402 = ~n20094 ;
  assign y5403 = n20099 ;
  assign y5404 = n20100 ;
  assign y5405 = n20104 ;
  assign y5406 = n20107 ;
  assign y5407 = ~n20109 ;
  assign y5408 = ~n20110 ;
  assign y5409 = ~n20114 ;
  assign y5410 = ~n20116 ;
  assign y5411 = ~1'b0 ;
  assign y5412 = ~n20117 ;
  assign y5413 = n20120 ;
  assign y5414 = n20122 ;
  assign y5415 = n20125 ;
  assign y5416 = n20131 ;
  assign y5417 = ~n20132 ;
  assign y5418 = ~n20137 ;
  assign y5419 = ~n20150 ;
  assign y5420 = n20155 ;
  assign y5421 = n20160 ;
  assign y5422 = ~1'b0 ;
  assign y5423 = n20161 ;
  assign y5424 = n20171 ;
  assign y5425 = ~n20173 ;
  assign y5426 = n20179 ;
  assign y5427 = ~n20182 ;
  assign y5428 = n20183 ;
  assign y5429 = ~n20184 ;
  assign y5430 = ~n20187 ;
  assign y5431 = ~n20192 ;
  assign y5432 = ~n20193 ;
  assign y5433 = n20194 ;
  assign y5434 = n20196 ;
  assign y5435 = ~n20197 ;
  assign y5436 = ~n20198 ;
  assign y5437 = ~n20200 ;
  assign y5438 = ~n20202 ;
  assign y5439 = ~n20211 ;
  assign y5440 = ~n20212 ;
  assign y5441 = ~n20217 ;
  assign y5442 = n20218 ;
  assign y5443 = n20228 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = n20231 ;
  assign y5446 = ~n20242 ;
  assign y5447 = ~n20250 ;
  assign y5448 = n20251 ;
  assign y5449 = n20262 ;
  assign y5450 = ~n20276 ;
  assign y5451 = n20280 ;
  assign y5452 = n20285 ;
  assign y5453 = n20286 ;
  assign y5454 = n20290 ;
  assign y5455 = n20291 ;
  assign y5456 = ~n20292 ;
  assign y5457 = n20298 ;
  assign y5458 = ~n20303 ;
  assign y5459 = ~n20307 ;
  assign y5460 = ~1'b0 ;
  assign y5461 = ~n20326 ;
  assign y5462 = ~n20333 ;
  assign y5463 = ~n20342 ;
  assign y5464 = n20345 ;
  assign y5465 = ~n20351 ;
  assign y5466 = ~n20353 ;
  assign y5467 = n20358 ;
  assign y5468 = ~n20361 ;
  assign y5469 = ~n20362 ;
  assign y5470 = ~n20365 ;
  assign y5471 = ~n20368 ;
  assign y5472 = ~n20372 ;
  assign y5473 = ~1'b0 ;
  assign y5474 = ~1'b0 ;
  assign y5475 = ~1'b0 ;
  assign y5476 = n20377 ;
  assign y5477 = ~1'b0 ;
  assign y5478 = n20380 ;
  assign y5479 = n20381 ;
  assign y5480 = ~n20388 ;
  assign y5481 = n20390 ;
  assign y5482 = n20392 ;
  assign y5483 = ~n20397 ;
  assign y5484 = ~n20400 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = n20406 ;
  assign y5487 = n20407 ;
  assign y5488 = ~n20411 ;
  assign y5489 = ~n20412 ;
  assign y5490 = ~1'b0 ;
  assign y5491 = n20413 ;
  assign y5492 = n20416 ;
  assign y5493 = n20424 ;
  assign y5494 = n20425 ;
  assign y5495 = ~1'b0 ;
  assign y5496 = ~n20427 ;
  assign y5497 = n20429 ;
  assign y5498 = ~n20435 ;
  assign y5499 = n20436 ;
  assign y5500 = ~1'b0 ;
  assign y5501 = ~1'b0 ;
  assign y5502 = ~1'b0 ;
  assign y5503 = ~n20438 ;
  assign y5504 = ~n20439 ;
  assign y5505 = n20440 ;
  assign y5506 = ~n20443 ;
  assign y5507 = ~n20451 ;
  assign y5508 = n20453 ;
  assign y5509 = n20459 ;
  assign y5510 = ~1'b0 ;
  assign y5511 = ~n20461 ;
  assign y5512 = ~n20462 ;
  assign y5513 = n20470 ;
  assign y5514 = n20475 ;
  assign y5515 = n20477 ;
  assign y5516 = n20478 ;
  assign y5517 = n20479 ;
  assign y5518 = n20480 ;
  assign y5519 = ~n20481 ;
  assign y5520 = n20485 ;
  assign y5521 = n20488 ;
  assign y5522 = ~n20489 ;
  assign y5523 = ~n7485 ;
  assign y5524 = n20492 ;
  assign y5525 = ~1'b0 ;
  assign y5526 = ~n20502 ;
  assign y5527 = n20503 ;
  assign y5528 = ~n20507 ;
  assign y5529 = ~n20514 ;
  assign y5530 = ~n20517 ;
  assign y5531 = ~n20518 ;
  assign y5532 = n20519 ;
  assign y5533 = 1'b0 ;
  assign y5534 = ~n20521 ;
  assign y5535 = n20524 ;
  assign y5536 = n20526 ;
  assign y5537 = ~n20530 ;
  assign y5538 = ~n20539 ;
  assign y5539 = n20543 ;
  assign y5540 = n20544 ;
  assign y5541 = n20545 ;
  assign y5542 = ~n20548 ;
  assign y5543 = ~n20554 ;
  assign y5544 = ~1'b0 ;
  assign y5545 = n20557 ;
  assign y5546 = n20560 ;
  assign y5547 = n20563 ;
  assign y5548 = ~n20569 ;
  assign y5549 = ~1'b0 ;
  assign y5550 = n20570 ;
  assign y5551 = ~n20575 ;
  assign y5552 = ~1'b0 ;
  assign y5553 = n20577 ;
  assign y5554 = ~n20578 ;
  assign y5555 = ~n20580 ;
  assign y5556 = n20584 ;
  assign y5557 = ~n20590 ;
  assign y5558 = ~1'b0 ;
  assign y5559 = ~1'b0 ;
  assign y5560 = ~n20593 ;
  assign y5561 = ~n20603 ;
  assign y5562 = ~n20606 ;
  assign y5563 = n20608 ;
  assign y5564 = n20612 ;
  assign y5565 = n20614 ;
  assign y5566 = n20615 ;
  assign y5567 = ~1'b0 ;
  assign y5568 = n20618 ;
  assign y5569 = ~n20628 ;
  assign y5570 = ~1'b0 ;
  assign y5571 = n20629 ;
  assign y5572 = ~n20635 ;
  assign y5573 = ~n20637 ;
  assign y5574 = ~1'b0 ;
  assign y5575 = ~1'b0 ;
  assign y5576 = n20640 ;
  assign y5577 = ~n20644 ;
  assign y5578 = ~n20646 ;
  assign y5579 = n20647 ;
  assign y5580 = n20651 ;
  assign y5581 = ~n20658 ;
  assign y5582 = n20661 ;
  assign y5583 = n20666 ;
  assign y5584 = ~n20667 ;
  assign y5585 = n20675 ;
  assign y5586 = ~n20676 ;
  assign y5587 = n20681 ;
  assign y5588 = ~n20682 ;
  assign y5589 = ~n20693 ;
  assign y5590 = ~1'b0 ;
  assign y5591 = ~n20702 ;
  assign y5592 = ~1'b0 ;
  assign y5593 = ~n20706 ;
  assign y5594 = ~n20708 ;
  assign y5595 = ~1'b0 ;
  assign y5596 = ~n20714 ;
  assign y5597 = ~n20718 ;
  assign y5598 = ~n20725 ;
  assign y5599 = n20730 ;
  assign y5600 = n20735 ;
  assign y5601 = ~n20745 ;
  assign y5602 = n20748 ;
  assign y5603 = 1'b0 ;
  assign y5604 = ~n20750 ;
  assign y5605 = ~1'b0 ;
  assign y5606 = ~n20754 ;
  assign y5607 = n20756 ;
  assign y5608 = ~n20757 ;
  assign y5609 = n20758 ;
  assign y5610 = n20770 ;
  assign y5611 = ~n20771 ;
  assign y5612 = n20777 ;
  assign y5613 = ~n20785 ;
  assign y5614 = ~n20787 ;
  assign y5615 = n20789 ;
  assign y5616 = ~n20791 ;
  assign y5617 = ~n20795 ;
  assign y5618 = ~n20796 ;
  assign y5619 = ~1'b0 ;
  assign y5620 = n20798 ;
  assign y5621 = ~n20800 ;
  assign y5622 = ~1'b0 ;
  assign y5623 = ~n20803 ;
  assign y5624 = ~n20805 ;
  assign y5625 = n20810 ;
  assign y5626 = n20812 ;
  assign y5627 = n20817 ;
  assign y5628 = n20819 ;
  assign y5629 = n20822 ;
  assign y5630 = n20827 ;
  assign y5631 = ~1'b0 ;
  assign y5632 = ~n20831 ;
  assign y5633 = ~1'b0 ;
  assign y5634 = ~n20832 ;
  assign y5635 = ~n20833 ;
  assign y5636 = n20835 ;
  assign y5637 = ~n20838 ;
  assign y5638 = n20843 ;
  assign y5639 = ~n20844 ;
  assign y5640 = ~1'b0 ;
  assign y5641 = ~n20848 ;
  assign y5642 = ~n20850 ;
  assign y5643 = n20852 ;
  assign y5644 = n20857 ;
  assign y5645 = ~n20859 ;
  assign y5646 = n20861 ;
  assign y5647 = ~n20864 ;
  assign y5648 = n20869 ;
  assign y5649 = n20874 ;
  assign y5650 = n20876 ;
  assign y5651 = n20883 ;
  assign y5652 = n20894 ;
  assign y5653 = ~1'b0 ;
  assign y5654 = n20903 ;
  assign y5655 = ~n20906 ;
  assign y5656 = n20916 ;
  assign y5657 = ~n20917 ;
  assign y5658 = n9835 ;
  assign y5659 = ~n20924 ;
  assign y5660 = ~n20928 ;
  assign y5661 = ~1'b0 ;
  assign y5662 = ~n20933 ;
  assign y5663 = ~n20936 ;
  assign y5664 = n20940 ;
  assign y5665 = ~n20946 ;
  assign y5666 = n20949 ;
  assign y5667 = ~n20951 ;
  assign y5668 = n20955 ;
  assign y5669 = ~1'b0 ;
  assign y5670 = n20958 ;
  assign y5671 = ~n20959 ;
  assign y5672 = ~n20961 ;
  assign y5673 = ~n20964 ;
  assign y5674 = n20970 ;
  assign y5675 = n20973 ;
  assign y5676 = n20975 ;
  assign y5677 = ~n20980 ;
  assign y5678 = ~1'b0 ;
  assign y5679 = n20982 ;
  assign y5680 = ~1'b0 ;
  assign y5681 = n20983 ;
  assign y5682 = ~1'b0 ;
  assign y5683 = ~n13807 ;
  assign y5684 = n20992 ;
  assign y5685 = n20993 ;
  assign y5686 = n20997 ;
  assign y5687 = ~n21001 ;
  assign y5688 = n6181 ;
  assign y5689 = ~n21007 ;
  assign y5690 = n21010 ;
  assign y5691 = ~n21011 ;
  assign y5692 = n21022 ;
  assign y5693 = ~n21028 ;
  assign y5694 = n21030 ;
  assign y5695 = ~n4263 ;
  assign y5696 = n21035 ;
  assign y5697 = n21043 ;
  assign y5698 = ~n21044 ;
  assign y5699 = ~n21053 ;
  assign y5700 = ~n21055 ;
  assign y5701 = n21056 ;
  assign y5702 = ~n21057 ;
  assign y5703 = ~n21060 ;
  assign y5704 = ~n21065 ;
  assign y5705 = n21068 ;
  assign y5706 = n21069 ;
  assign y5707 = ~n21072 ;
  assign y5708 = n21073 ;
  assign y5709 = ~1'b0 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = ~n21075 ;
  assign y5712 = n21083 ;
  assign y5713 = ~n21084 ;
  assign y5714 = n21091 ;
  assign y5715 = n21102 ;
  assign y5716 = ~n21104 ;
  assign y5717 = ~n21105 ;
  assign y5718 = n21109 ;
  assign y5719 = ~n21111 ;
  assign y5720 = n21118 ;
  assign y5721 = ~n21124 ;
  assign y5722 = ~n21125 ;
  assign y5723 = ~n21128 ;
  assign y5724 = n21134 ;
  assign y5725 = n21138 ;
  assign y5726 = ~n21139 ;
  assign y5727 = n21144 ;
  assign y5728 = n21145 ;
  assign y5729 = n21159 ;
  assign y5730 = ~n21162 ;
  assign y5731 = n21164 ;
  assign y5732 = ~n21168 ;
  assign y5733 = n21173 ;
  assign y5734 = n21179 ;
  assign y5735 = n21183 ;
  assign y5736 = ~n21185 ;
  assign y5737 = ~1'b0 ;
  assign y5738 = ~n21189 ;
  assign y5739 = ~n21192 ;
  assign y5740 = n21193 ;
  assign y5741 = n21194 ;
  assign y5742 = n21195 ;
  assign y5743 = ~n21198 ;
  assign y5744 = ~n12818 ;
  assign y5745 = n21202 ;
  assign y5746 = ~n21208 ;
  assign y5747 = ~n21210 ;
  assign y5748 = ~n21211 ;
  assign y5749 = ~n21212 ;
  assign y5750 = ~1'b0 ;
  assign y5751 = n21213 ;
  assign y5752 = n21217 ;
  assign y5753 = ~n21220 ;
  assign y5754 = ~1'b0 ;
  assign y5755 = ~n21225 ;
  assign y5756 = ~n21226 ;
  assign y5757 = ~n21229 ;
  assign y5758 = ~n21231 ;
  assign y5759 = ~n21236 ;
  assign y5760 = ~n21244 ;
  assign y5761 = n21245 ;
  assign y5762 = n21247 ;
  assign y5763 = ~n21248 ;
  assign y5764 = ~1'b0 ;
  assign y5765 = n21252 ;
  assign y5766 = ~n21260 ;
  assign y5767 = n21262 ;
  assign y5768 = n21265 ;
  assign y5769 = ~n21267 ;
  assign y5770 = ~n21268 ;
  assign y5771 = ~n21274 ;
  assign y5772 = ~n21277 ;
  assign y5773 = ~1'b0 ;
  assign y5774 = ~n21282 ;
  assign y5775 = ~n21284 ;
  assign y5776 = ~1'b0 ;
  assign y5777 = n21286 ;
  assign y5778 = n21296 ;
  assign y5779 = ~n21297 ;
  assign y5780 = ~n21301 ;
  assign y5781 = n21305 ;
  assign y5782 = n21308 ;
  assign y5783 = n21312 ;
  assign y5784 = ~n21314 ;
  assign y5785 = ~1'b0 ;
  assign y5786 = n21317 ;
  assign y5787 = ~n21320 ;
  assign y5788 = ~1'b0 ;
  assign y5789 = n21323 ;
  assign y5790 = ~n21324 ;
  assign y5791 = ~n21325 ;
  assign y5792 = n21329 ;
  assign y5793 = ~1'b0 ;
  assign y5794 = n21331 ;
  assign y5795 = n21338 ;
  assign y5796 = ~n21339 ;
  assign y5797 = n21349 ;
  assign y5798 = ~n21350 ;
  assign y5799 = n21354 ;
  assign y5800 = ~1'b0 ;
  assign y5801 = ~n21357 ;
  assign y5802 = n21365 ;
  assign y5803 = ~n21371 ;
  assign y5804 = n21374 ;
  assign y5805 = n21382 ;
  assign y5806 = ~n21384 ;
  assign y5807 = n21386 ;
  assign y5808 = ~n21394 ;
  assign y5809 = n21396 ;
  assign y5810 = ~n21397 ;
  assign y5811 = ~n21407 ;
  assign y5812 = ~n21411 ;
  assign y5813 = n21413 ;
  assign y5814 = n21418 ;
  assign y5815 = ~1'b0 ;
  assign y5816 = ~n21423 ;
  assign y5817 = n21424 ;
  assign y5818 = n21425 ;
  assign y5819 = ~n21427 ;
  assign y5820 = n21434 ;
  assign y5821 = n21438 ;
  assign y5822 = n21444 ;
  assign y5823 = n21450 ;
  assign y5824 = n21451 ;
  assign y5825 = n21464 ;
  assign y5826 = ~n21465 ;
  assign y5827 = ~n21467 ;
  assign y5828 = n21469 ;
  assign y5829 = n21474 ;
  assign y5830 = ~n21478 ;
  assign y5831 = n21483 ;
  assign y5832 = ~n21484 ;
  assign y5833 = ~1'b0 ;
  assign y5834 = ~n21486 ;
  assign y5835 = ~1'b0 ;
  assign y5836 = n21493 ;
  assign y5837 = ~n21494 ;
  assign y5838 = ~n21496 ;
  assign y5839 = ~n21499 ;
  assign y5840 = ~n21500 ;
  assign y5841 = ~n21501 ;
  assign y5842 = ~n21504 ;
  assign y5843 = n21507 ;
  assign y5844 = n21514 ;
  assign y5845 = n21516 ;
  assign y5846 = ~x49 ;
  assign y5847 = ~1'b0 ;
  assign y5848 = ~1'b0 ;
  assign y5849 = n21519 ;
  assign y5850 = ~n21523 ;
  assign y5851 = n21529 ;
  assign y5852 = ~1'b0 ;
  assign y5853 = ~n21530 ;
  assign y5854 = n21531 ;
  assign y5855 = ~n21535 ;
  assign y5856 = n21543 ;
  assign y5857 = n21544 ;
  assign y5858 = ~n21545 ;
  assign y5859 = ~1'b0 ;
  assign y5860 = ~n21548 ;
  assign y5861 = ~1'b0 ;
  assign y5862 = n21550 ;
  assign y5863 = n21551 ;
  assign y5864 = n21555 ;
  assign y5865 = ~n21558 ;
  assign y5866 = ~n21559 ;
  assign y5867 = ~1'b0 ;
  assign y5868 = ~1'b0 ;
  assign y5869 = ~1'b0 ;
  assign y5870 = n21564 ;
  assign y5871 = ~1'b0 ;
  assign y5872 = ~n21568 ;
  assign y5873 = ~n21569 ;
  assign y5874 = n21571 ;
  assign y5875 = ~1'b0 ;
  assign y5876 = ~n21583 ;
  assign y5877 = ~n21584 ;
  assign y5878 = n21590 ;
  assign y5879 = ~n21593 ;
  assign y5880 = ~n21596 ;
  assign y5881 = ~1'b0 ;
  assign y5882 = ~1'b0 ;
  assign y5883 = ~1'b0 ;
  assign y5884 = ~n21597 ;
  assign y5885 = ~1'b0 ;
  assign y5886 = ~1'b0 ;
  assign y5887 = ~1'b0 ;
  assign y5888 = n21601 ;
  assign y5889 = n21602 ;
  assign y5890 = n21604 ;
  assign y5891 = ~n21608 ;
  assign y5892 = ~n21612 ;
  assign y5893 = n21613 ;
  assign y5894 = ~n21617 ;
  assign y5895 = ~n21619 ;
  assign y5896 = ~n21621 ;
  assign y5897 = ~n21623 ;
  assign y5898 = n21631 ;
  assign y5899 = n21632 ;
  assign y5900 = ~n21633 ;
  assign y5901 = n21635 ;
  assign y5902 = ~n21637 ;
  assign y5903 = n21641 ;
  assign y5904 = n21645 ;
  assign y5905 = n21656 ;
  assign y5906 = n21659 ;
  assign y5907 = ~n21664 ;
  assign y5908 = n21666 ;
  assign y5909 = n21667 ;
  assign y5910 = ~n21672 ;
  assign y5911 = n21675 ;
  assign y5912 = ~1'b0 ;
  assign y5913 = ~n21679 ;
  assign y5914 = ~n21680 ;
  assign y5915 = n21686 ;
  assign y5916 = ~n21688 ;
  assign y5917 = n21689 ;
  assign y5918 = n21692 ;
  assign y5919 = ~1'b0 ;
  assign y5920 = n21700 ;
  assign y5921 = n21704 ;
  assign y5922 = ~n21718 ;
  assign y5923 = n21725 ;
  assign y5924 = n21726 ;
  assign y5925 = ~n21727 ;
  assign y5926 = ~1'b0 ;
  assign y5927 = ~n21729 ;
  assign y5928 = n21730 ;
  assign y5929 = ~n21735 ;
  assign y5930 = ~n21744 ;
  assign y5931 = n21746 ;
  assign y5932 = ~n21747 ;
  assign y5933 = n21751 ;
  assign y5934 = n21752 ;
  assign y5935 = n21757 ;
  assign y5936 = n21759 ;
  assign y5937 = ~n21765 ;
  assign y5938 = ~n21767 ;
  assign y5939 = ~n21773 ;
  assign y5940 = n21776 ;
  assign y5941 = ~n21782 ;
  assign y5942 = ~n21784 ;
  assign y5943 = ~n21786 ;
  assign y5944 = ~n21787 ;
  assign y5945 = ~n21797 ;
  assign y5946 = n21798 ;
  assign y5947 = n21800 ;
  assign y5948 = ~n21802 ;
  assign y5949 = ~n21805 ;
  assign y5950 = n21807 ;
  assign y5951 = ~n21812 ;
  assign y5952 = ~n14087 ;
  assign y5953 = ~n21815 ;
  assign y5954 = n21824 ;
  assign y5955 = ~n21826 ;
  assign y5956 = n21827 ;
  assign y5957 = n21830 ;
  assign y5958 = ~n21836 ;
  assign y5959 = ~n21838 ;
  assign y5960 = n21844 ;
  assign y5961 = ~n21854 ;
  assign y5962 = ~1'b0 ;
  assign y5963 = ~n21856 ;
  assign y5964 = ~n21863 ;
  assign y5965 = ~n21868 ;
  assign y5966 = ~1'b0 ;
  assign y5967 = ~n2504 ;
  assign y5968 = ~1'b0 ;
  assign y5969 = 1'b0 ;
  assign y5970 = ~n21874 ;
  assign y5971 = ~n21875 ;
  assign y5972 = ~n21877 ;
  assign y5973 = ~n21878 ;
  assign y5974 = ~n21880 ;
  assign y5975 = ~n21883 ;
  assign y5976 = n21886 ;
  assign y5977 = n21892 ;
  assign y5978 = ~n21895 ;
  assign y5979 = n21898 ;
  assign y5980 = ~n21902 ;
  assign y5981 = n21909 ;
  assign y5982 = n21912 ;
  assign y5983 = ~n21920 ;
  assign y5984 = ~1'b0 ;
  assign y5985 = ~n21928 ;
  assign y5986 = n21933 ;
  assign y5987 = n21937 ;
  assign y5988 = n21943 ;
  assign y5989 = ~n21944 ;
  assign y5990 = n21946 ;
  assign y5991 = ~1'b0 ;
  assign y5992 = n21947 ;
  assign y5993 = ~n21951 ;
  assign y5994 = ~n21957 ;
  assign y5995 = n21958 ;
  assign y5996 = n21962 ;
  assign y5997 = n21963 ;
  assign y5998 = n21967 ;
  assign y5999 = ~n21968 ;
  assign y6000 = ~n21969 ;
  assign y6001 = ~n21971 ;
  assign y6002 = ~n21972 ;
  assign y6003 = ~n21977 ;
  assign y6004 = ~x65 ;
  assign y6005 = n21978 ;
  assign y6006 = ~1'b0 ;
  assign y6007 = n21984 ;
  assign y6008 = n21986 ;
  assign y6009 = ~n21996 ;
  assign y6010 = ~1'b0 ;
  assign y6011 = n22000 ;
  assign y6012 = n22001 ;
  assign y6013 = n22006 ;
  assign y6014 = n22009 ;
  assign y6015 = n22013 ;
  assign y6016 = n22016 ;
  assign y6017 = n22018 ;
  assign y6018 = n22021 ;
  assign y6019 = ~n22023 ;
  assign y6020 = ~n22025 ;
  assign y6021 = ~n22027 ;
  assign y6022 = ~n22030 ;
  assign y6023 = n22033 ;
  assign y6024 = ~n22052 ;
  assign y6025 = n22056 ;
  assign y6026 = n22063 ;
  assign y6027 = n22065 ;
  assign y6028 = n22071 ;
  assign y6029 = n22074 ;
  assign y6030 = n22082 ;
  assign y6031 = ~n22083 ;
  assign y6032 = ~1'b0 ;
  assign y6033 = ~n22085 ;
  assign y6034 = n22088 ;
  assign y6035 = n22092 ;
  assign y6036 = ~n22095 ;
  assign y6037 = n22097 ;
  assign y6038 = n22099 ;
  assign y6039 = n22107 ;
  assign y6040 = n22115 ;
  assign y6041 = ~1'b0 ;
  assign y6042 = n22116 ;
  assign y6043 = ~n5086 ;
  assign y6044 = n22117 ;
  assign y6045 = n22120 ;
  assign y6046 = ~n22124 ;
  assign y6047 = ~1'b0 ;
  assign y6048 = n22127 ;
  assign y6049 = ~n22128 ;
  assign y6050 = ~n22132 ;
  assign y6051 = n22141 ;
  assign y6052 = n22154 ;
  assign y6053 = ~n22157 ;
  assign y6054 = n22160 ;
  assign y6055 = n22161 ;
  assign y6056 = n22167 ;
  assign y6057 = ~1'b0 ;
  assign y6058 = n22168 ;
  assign y6059 = ~n22176 ;
  assign y6060 = n22177 ;
  assign y6061 = ~n22178 ;
  assign y6062 = n22181 ;
  assign y6063 = n22185 ;
  assign y6064 = n22187 ;
  assign y6065 = n22190 ;
  assign y6066 = ~1'b0 ;
  assign y6067 = ~1'b0 ;
  assign y6068 = n22195 ;
  assign y6069 = ~n22196 ;
  assign y6070 = n22199 ;
  assign y6071 = ~n22205 ;
  assign y6072 = n22206 ;
  assign y6073 = ~n22211 ;
  assign y6074 = ~n22215 ;
  assign y6075 = ~1'b0 ;
  assign y6076 = ~n22216 ;
  assign y6077 = n22224 ;
  assign y6078 = n22226 ;
  assign y6079 = n22233 ;
  assign y6080 = ~n22240 ;
  assign y6081 = ~n22248 ;
  assign y6082 = ~n22251 ;
  assign y6083 = ~n22259 ;
  assign y6084 = ~n22263 ;
  assign y6085 = n22264 ;
  assign y6086 = n22271 ;
  assign y6087 = ~n22273 ;
  assign y6088 = ~1'b0 ;
  assign y6089 = ~n22277 ;
  assign y6090 = n22279 ;
  assign y6091 = n22281 ;
  assign y6092 = n22284 ;
  assign y6093 = n22289 ;
  assign y6094 = ~n22290 ;
  assign y6095 = ~n22291 ;
  assign y6096 = n22292 ;
  assign y6097 = ~n22300 ;
  assign y6098 = ~n22302 ;
  assign y6099 = n22303 ;
  assign y6100 = ~n22311 ;
  assign y6101 = n22314 ;
  assign y6102 = ~n22315 ;
  assign y6103 = ~1'b0 ;
  assign y6104 = ~1'b0 ;
  assign y6105 = ~n22317 ;
  assign y6106 = ~n22319 ;
  assign y6107 = ~n22320 ;
  assign y6108 = n22328 ;
  assign y6109 = ~1'b0 ;
  assign y6110 = ~n22334 ;
  assign y6111 = ~n22335 ;
  assign y6112 = n22344 ;
  assign y6113 = n22345 ;
  assign y6114 = n22348 ;
  assign y6115 = ~n22357 ;
  assign y6116 = n22364 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = ~n22367 ;
  assign y6119 = n22371 ;
  assign y6120 = ~n22373 ;
  assign y6121 = n22376 ;
  assign y6122 = ~n22380 ;
  assign y6123 = n22383 ;
  assign y6124 = ~n22385 ;
  assign y6125 = ~n22387 ;
  assign y6126 = n22388 ;
  assign y6127 = n22394 ;
  assign y6128 = ~n22398 ;
  assign y6129 = ~n22403 ;
  assign y6130 = n22407 ;
  assign y6131 = ~n22411 ;
  assign y6132 = n22412 ;
  assign y6133 = ~n22420 ;
  assign y6134 = n22426 ;
  assign y6135 = n22428 ;
  assign y6136 = n22430 ;
  assign y6137 = ~1'b0 ;
  assign y6138 = ~n22438 ;
  assign y6139 = n22440 ;
  assign y6140 = ~n22441 ;
  assign y6141 = ~1'b0 ;
  assign y6142 = ~n22444 ;
  assign y6143 = n22446 ;
  assign y6144 = n22450 ;
  assign y6145 = ~n22452 ;
  assign y6146 = n22453 ;
  assign y6147 = ~n22457 ;
  assign y6148 = ~n22459 ;
  assign y6149 = ~n22463 ;
  assign y6150 = ~1'b0 ;
  assign y6151 = n22467 ;
  assign y6152 = ~n22468 ;
  assign y6153 = ~n22481 ;
  assign y6154 = n22489 ;
  assign y6155 = n22492 ;
  assign y6156 = n22500 ;
  assign y6157 = ~1'b0 ;
  assign y6158 = ~n22504 ;
  assign y6159 = ~n22507 ;
  assign y6160 = ~n22513 ;
  assign y6161 = n22515 ;
  assign y6162 = n22518 ;
  assign y6163 = n22519 ;
  assign y6164 = ~n22523 ;
  assign y6165 = ~n22525 ;
  assign y6166 = ~n22526 ;
  assign y6167 = n22528 ;
  assign y6168 = ~n20135 ;
  assign y6169 = n22529 ;
  assign y6170 = n22531 ;
  assign y6171 = n22534 ;
  assign y6172 = n22540 ;
  assign y6173 = ~n22542 ;
  assign y6174 = n22544 ;
  assign y6175 = ~n22549 ;
  assign y6176 = n22552 ;
  assign y6177 = n22553 ;
  assign y6178 = ~n22556 ;
  assign y6179 = n22559 ;
  assign y6180 = n22562 ;
  assign y6181 = ~n18467 ;
  assign y6182 = n22563 ;
  assign y6183 = n22564 ;
  assign y6184 = ~1'b0 ;
  assign y6185 = n22568 ;
  assign y6186 = n22569 ;
  assign y6187 = n22575 ;
  assign y6188 = n22579 ;
  assign y6189 = n22580 ;
  assign y6190 = ~n22585 ;
  assign y6191 = n22589 ;
  assign y6192 = ~n22590 ;
  assign y6193 = n22598 ;
  assign y6194 = ~n22599 ;
  assign y6195 = ~n22602 ;
  assign y6196 = ~n22603 ;
  assign y6197 = ~1'b0 ;
  assign y6198 = ~n22605 ;
  assign y6199 = n22606 ;
  assign y6200 = n22624 ;
  assign y6201 = ~1'b0 ;
  assign y6202 = n22625 ;
  assign y6203 = ~n22626 ;
  assign y6204 = ~n22628 ;
  assign y6205 = ~n22637 ;
  assign y6206 = ~n22639 ;
  assign y6207 = ~n22645 ;
  assign y6208 = ~1'b0 ;
  assign y6209 = ~n22649 ;
  assign y6210 = n22650 ;
  assign y6211 = ~1'b0 ;
  assign y6212 = n22654 ;
  assign y6213 = n22655 ;
  assign y6214 = n22661 ;
  assign y6215 = ~n22665 ;
  assign y6216 = n22668 ;
  assign y6217 = ~n22671 ;
  assign y6218 = n22672 ;
  assign y6219 = ~n22675 ;
  assign y6220 = ~n22679 ;
  assign y6221 = ~n22681 ;
  assign y6222 = ~n22684 ;
  assign y6223 = ~n22688 ;
  assign y6224 = ~1'b0 ;
  assign y6225 = n22694 ;
  assign y6226 = n22699 ;
  assign y6227 = ~n22700 ;
  assign y6228 = n22701 ;
  assign y6229 = n22705 ;
  assign y6230 = ~n22706 ;
  assign y6231 = n22707 ;
  assign y6232 = n22714 ;
  assign y6233 = ~n22716 ;
  assign y6234 = n22719 ;
  assign y6235 = n22721 ;
  assign y6236 = ~n22723 ;
  assign y6237 = ~n22724 ;
  assign y6238 = ~n22725 ;
  assign y6239 = ~n22726 ;
  assign y6240 = ~1'b0 ;
  assign y6241 = ~n22727 ;
  assign y6242 = n22728 ;
  assign y6243 = ~1'b0 ;
  assign y6244 = n22733 ;
  assign y6245 = ~n22738 ;
  assign y6246 = ~n22740 ;
  assign y6247 = ~n22742 ;
  assign y6248 = ~n22751 ;
  assign y6249 = ~n22754 ;
  assign y6250 = n22759 ;
  assign y6251 = n22762 ;
  assign y6252 = n22763 ;
  assign y6253 = n22767 ;
  assign y6254 = n22772 ;
  assign y6255 = ~n22775 ;
  assign y6256 = ~n22782 ;
  assign y6257 = ~n22783 ;
  assign y6258 = ~n22785 ;
  assign y6259 = ~1'b0 ;
  assign y6260 = ~n22789 ;
  assign y6261 = n22793 ;
  assign y6262 = n22794 ;
  assign y6263 = n22797 ;
  assign y6264 = ~n22804 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = ~n22806 ;
  assign y6267 = n22813 ;
  assign y6268 = n22814 ;
  assign y6269 = ~n22816 ;
  assign y6270 = n22817 ;
  assign y6271 = ~n22818 ;
  assign y6272 = n22823 ;
  assign y6273 = ~n22828 ;
  assign y6274 = ~n22831 ;
  assign y6275 = n22833 ;
  assign y6276 = ~1'b0 ;
  assign y6277 = n22837 ;
  assign y6278 = n22848 ;
  assign y6279 = n22855 ;
  assign y6280 = ~n22857 ;
  assign y6281 = ~n22858 ;
  assign y6282 = n22865 ;
  assign y6283 = n22873 ;
  assign y6284 = n22878 ;
  assign y6285 = ~n22881 ;
  assign y6286 = ~1'b0 ;
  assign y6287 = ~n22885 ;
  assign y6288 = ~1'b0 ;
  assign y6289 = ~n22887 ;
  assign y6290 = n22894 ;
  assign y6291 = ~1'b0 ;
  assign y6292 = n22898 ;
  assign y6293 = ~n22900 ;
  assign y6294 = n22905 ;
  assign y6295 = n22906 ;
  assign y6296 = ~n22908 ;
  assign y6297 = n22912 ;
  assign y6298 = n22913 ;
  assign y6299 = n22915 ;
  assign y6300 = n22916 ;
  assign y6301 = ~n22918 ;
  assign y6302 = ~n22919 ;
  assign y6303 = n22926 ;
  assign y6304 = ~n22929 ;
  assign y6305 = ~n22932 ;
  assign y6306 = n22934 ;
  assign y6307 = n22940 ;
  assign y6308 = ~n22947 ;
  assign y6309 = ~n22948 ;
  assign y6310 = n22950 ;
  assign y6311 = n22966 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = n22967 ;
  assign y6314 = ~1'b0 ;
  assign y6315 = ~1'b0 ;
  assign y6316 = n22968 ;
  assign y6317 = ~1'b0 ;
  assign y6318 = n22971 ;
  assign y6319 = ~n22973 ;
  assign y6320 = ~n22978 ;
  assign y6321 = n22982 ;
  assign y6322 = ~1'b0 ;
  assign y6323 = n22986 ;
  assign y6324 = ~n22989 ;
  assign y6325 = ~n22992 ;
  assign y6326 = ~n22993 ;
  assign y6327 = ~n22994 ;
  assign y6328 = n22995 ;
  assign y6329 = n22999 ;
  assign y6330 = n23005 ;
  assign y6331 = ~n23006 ;
  assign y6332 = ~n23010 ;
  assign y6333 = ~n23016 ;
  assign y6334 = n23017 ;
  assign y6335 = n23018 ;
  assign y6336 = ~n23021 ;
  assign y6337 = n23028 ;
  assign y6338 = n23030 ;
  assign y6339 = ~n23035 ;
  assign y6340 = ~n23040 ;
  assign y6341 = n23041 ;
  assign y6342 = ~n23044 ;
  assign y6343 = n23045 ;
  assign y6344 = ~1'b0 ;
  assign y6345 = ~1'b0 ;
  assign y6346 = n23048 ;
  assign y6347 = ~n23053 ;
  assign y6348 = ~n23057 ;
  assign y6349 = n23061 ;
  assign y6350 = n23063 ;
  assign y6351 = n23064 ;
  assign y6352 = ~n23065 ;
  assign y6353 = n23069 ;
  assign y6354 = n23073 ;
  assign y6355 = ~n23075 ;
  assign y6356 = ~n23078 ;
  assign y6357 = n23083 ;
  assign y6358 = n23085 ;
  assign y6359 = n23089 ;
  assign y6360 = n23096 ;
  assign y6361 = ~1'b0 ;
  assign y6362 = n23098 ;
  assign y6363 = ~n23107 ;
  assign y6364 = ~1'b0 ;
  assign y6365 = ~n23114 ;
  assign y6366 = ~n23115 ;
  assign y6367 = n23117 ;
  assign y6368 = n23118 ;
  assign y6369 = ~n23124 ;
  assign y6370 = ~n23126 ;
  assign y6371 = n23127 ;
  assign y6372 = n23131 ;
  assign y6373 = ~n23134 ;
  assign y6374 = n23139 ;
  assign y6375 = ~1'b0 ;
  assign y6376 = ~1'b0 ;
  assign y6377 = ~n23143 ;
  assign y6378 = ~1'b0 ;
  assign y6379 = n23148 ;
  assign y6380 = ~n23153 ;
  assign y6381 = ~n23155 ;
  assign y6382 = n23159 ;
  assign y6383 = n23161 ;
  assign y6384 = n23162 ;
  assign y6385 = ~n23163 ;
  assign y6386 = ~n23165 ;
  assign y6387 = n23181 ;
  assign y6388 = ~n23184 ;
  assign y6389 = ~n23186 ;
  assign y6390 = ~1'b0 ;
  assign y6391 = ~n23188 ;
  assign y6392 = ~n23191 ;
  assign y6393 = ~n23200 ;
  assign y6394 = ~n23205 ;
  assign y6395 = ~1'b0 ;
  assign y6396 = n23208 ;
  assign y6397 = n23213 ;
  assign y6398 = n23217 ;
  assign y6399 = n23219 ;
  assign y6400 = ~n23221 ;
  assign y6401 = n23222 ;
  assign y6402 = ~n23225 ;
  assign y6403 = n23229 ;
  assign y6404 = ~n23230 ;
  assign y6405 = n23235 ;
  assign y6406 = ~1'b0 ;
  assign y6407 = ~1'b0 ;
  assign y6408 = n23236 ;
  assign y6409 = ~n23237 ;
  assign y6410 = 1'b0 ;
  assign y6411 = ~1'b0 ;
  assign y6412 = n23244 ;
  assign y6413 = n23247 ;
  assign y6414 = ~n23249 ;
  assign y6415 = ~n23255 ;
  assign y6416 = n23263 ;
  assign y6417 = ~n23267 ;
  assign y6418 = ~1'b0 ;
  assign y6419 = ~n23273 ;
  assign y6420 = ~n23275 ;
  assign y6421 = ~n23277 ;
  assign y6422 = n23282 ;
  assign y6423 = n23283 ;
  assign y6424 = ~n23290 ;
  assign y6425 = n23295 ;
  assign y6426 = ~n23298 ;
  assign y6427 = ~1'b0 ;
  assign y6428 = n23306 ;
  assign y6429 = n23312 ;
  assign y6430 = ~n23323 ;
  assign y6431 = ~n23329 ;
  assign y6432 = ~1'b0 ;
  assign y6433 = ~n23335 ;
  assign y6434 = ~n10068 ;
  assign y6435 = ~n23337 ;
  assign y6436 = n23341 ;
  assign y6437 = ~1'b0 ;
  assign y6438 = ~n23350 ;
  assign y6439 = ~n23351 ;
  assign y6440 = ~n23352 ;
  assign y6441 = ~n23354 ;
  assign y6442 = ~n23360 ;
  assign y6443 = ~1'b0 ;
  assign y6444 = ~n23361 ;
  assign y6445 = ~1'b0 ;
  assign y6446 = n6226 ;
  assign y6447 = n23365 ;
  assign y6448 = n23366 ;
  assign y6449 = ~1'b0 ;
  assign y6450 = ~1'b0 ;
  assign y6451 = ~n23368 ;
  assign y6452 = ~n23369 ;
  assign y6453 = n23370 ;
  assign y6454 = ~n23375 ;
  assign y6455 = ~1'b0 ;
  assign y6456 = ~1'b0 ;
  assign y6457 = ~n23377 ;
  assign y6458 = ~n23378 ;
  assign y6459 = ~n23379 ;
  assign y6460 = n23380 ;
  assign y6461 = n23381 ;
  assign y6462 = ~n23383 ;
  assign y6463 = n9214 ;
  assign y6464 = ~n23393 ;
  assign y6465 = n23394 ;
  assign y6466 = ~n23396 ;
  assign y6467 = n23399 ;
  assign y6468 = n23400 ;
  assign y6469 = n23404 ;
  assign y6470 = ~1'b0 ;
  assign y6471 = n23407 ;
  assign y6472 = ~n23415 ;
  assign y6473 = ~n23418 ;
  assign y6474 = ~1'b0 ;
  assign y6475 = n23419 ;
  assign y6476 = ~n23422 ;
  assign y6477 = ~1'b0 ;
  assign y6478 = n23426 ;
  assign y6479 = ~1'b0 ;
  assign y6480 = n23427 ;
  assign y6481 = ~n23430 ;
  assign y6482 = n23435 ;
  assign y6483 = n2937 ;
  assign y6484 = n23445 ;
  assign y6485 = ~n23449 ;
  assign y6486 = ~n23453 ;
  assign y6487 = ~n23468 ;
  assign y6488 = n23471 ;
  assign y6489 = ~1'b0 ;
  assign y6490 = n23475 ;
  assign y6491 = n23476 ;
  assign y6492 = n23479 ;
  assign y6493 = ~1'b0 ;
  assign y6494 = n23485 ;
  assign y6495 = n23491 ;
  assign y6496 = ~n23494 ;
  assign y6497 = ~n23499 ;
  assign y6498 = n23506 ;
  assign y6499 = n23513 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = n23515 ;
  assign y6502 = n23522 ;
  assign y6503 = ~n23527 ;
  assign y6504 = 1'b0 ;
  assign y6505 = n23531 ;
  assign y6506 = ~n23532 ;
  assign y6507 = ~n23537 ;
  assign y6508 = ~n23539 ;
  assign y6509 = n23542 ;
  assign y6510 = ~n23546 ;
  assign y6511 = n23547 ;
  assign y6512 = ~1'b0 ;
  assign y6513 = ~n23554 ;
  assign y6514 = ~n23555 ;
  assign y6515 = ~n23559 ;
  assign y6516 = ~n23560 ;
  assign y6517 = ~n23562 ;
  assign y6518 = ~1'b0 ;
  assign y6519 = n23565 ;
  assign y6520 = n23566 ;
  assign y6521 = ~n23568 ;
  assign y6522 = n23571 ;
  assign y6523 = n6536 ;
  assign y6524 = ~n23572 ;
  assign y6525 = n23573 ;
  assign y6526 = ~n23581 ;
  assign y6527 = ~1'b0 ;
  assign y6528 = ~1'b0 ;
  assign y6529 = n23584 ;
  assign y6530 = n23592 ;
  assign y6531 = ~n23596 ;
  assign y6532 = n23597 ;
  assign y6533 = ~n23602 ;
  assign y6534 = ~n23606 ;
  assign y6535 = n23613 ;
  assign y6536 = n23618 ;
  assign y6537 = ~1'b0 ;
  assign y6538 = ~1'b0 ;
  assign y6539 = ~n23619 ;
  assign y6540 = ~n23621 ;
  assign y6541 = n23623 ;
  assign y6542 = n23625 ;
  assign y6543 = ~n23629 ;
  assign y6544 = n23634 ;
  assign y6545 = n23635 ;
  assign y6546 = n23639 ;
  assign y6547 = ~n23640 ;
  assign y6548 = n23643 ;
  assign y6549 = ~n23645 ;
  assign y6550 = ~n23646 ;
  assign y6551 = ~n23648 ;
  assign y6552 = n23652 ;
  assign y6553 = n23655 ;
  assign y6554 = n23658 ;
  assign y6555 = n6476 ;
  assign y6556 = n23659 ;
  assign y6557 = n23661 ;
  assign y6558 = ~n23662 ;
  assign y6559 = ~n23664 ;
  assign y6560 = n23667 ;
  assign y6561 = n23670 ;
  assign y6562 = n23672 ;
  assign y6563 = n23674 ;
  assign y6564 = ~n23684 ;
  assign y6565 = ~n23695 ;
  assign y6566 = n23698 ;
  assign y6567 = n23699 ;
  assign y6568 = ~1'b0 ;
  assign y6569 = ~1'b0 ;
  assign y6570 = ~n23703 ;
  assign y6571 = ~n23707 ;
  assign y6572 = n23710 ;
  assign y6573 = n23713 ;
  assign y6574 = ~1'b0 ;
  assign y6575 = ~n23717 ;
  assign y6576 = n23718 ;
  assign y6577 = n23727 ;
  assign y6578 = n23731 ;
  assign y6579 = ~n23734 ;
  assign y6580 = ~1'b0 ;
  assign y6581 = ~n23739 ;
  assign y6582 = n23740 ;
  assign y6583 = n23745 ;
  assign y6584 = ~n23749 ;
  assign y6585 = ~n23752 ;
  assign y6586 = ~n23753 ;
  assign y6587 = ~n23756 ;
  assign y6588 = n23762 ;
  assign y6589 = ~1'b0 ;
  assign y6590 = ~n23764 ;
  assign y6591 = ~n23769 ;
  assign y6592 = ~n23771 ;
  assign y6593 = ~1'b0 ;
  assign y6594 = ~n23776 ;
  assign y6595 = n23778 ;
  assign y6596 = n23780 ;
  assign y6597 = n23782 ;
  assign y6598 = n23785 ;
  assign y6599 = ~n23786 ;
  assign y6600 = n23787 ;
  assign y6601 = ~1'b0 ;
  assign y6602 = n23788 ;
  assign y6603 = n23789 ;
  assign y6604 = n23794 ;
  assign y6605 = ~n23795 ;
  assign y6606 = n23800 ;
  assign y6607 = ~n23801 ;
  assign y6608 = n23803 ;
  assign y6609 = n23806 ;
  assign y6610 = ~1'b0 ;
  assign y6611 = ~n23814 ;
  assign y6612 = n23817 ;
  assign y6613 = n23820 ;
  assign y6614 = ~1'b0 ;
  assign y6615 = ~n23830 ;
  assign y6616 = n23831 ;
  assign y6617 = ~n23832 ;
  assign y6618 = n23835 ;
  assign y6619 = n23837 ;
  assign y6620 = ~n23838 ;
  assign y6621 = ~n23840 ;
  assign y6622 = ~n23845 ;
  assign y6623 = n23846 ;
  assign y6624 = ~n23851 ;
  assign y6625 = ~n23859 ;
  assign y6626 = n23860 ;
  assign y6627 = ~n23864 ;
  assign y6628 = ~n23865 ;
  assign y6629 = n23877 ;
  assign y6630 = n23879 ;
  assign y6631 = ~n23880 ;
  assign y6632 = n23887 ;
  assign y6633 = n23895 ;
  assign y6634 = ~1'b0 ;
  assign y6635 = ~n23898 ;
  assign y6636 = n23900 ;
  assign y6637 = ~n23901 ;
  assign y6638 = ~n23902 ;
  assign y6639 = n23905 ;
  assign y6640 = ~1'b0 ;
  assign y6641 = ~n3248 ;
  assign y6642 = ~n23913 ;
  assign y6643 = ~1'b0 ;
  assign y6644 = ~n23915 ;
  assign y6645 = n23924 ;
  assign y6646 = n23927 ;
  assign y6647 = n23931 ;
  assign y6648 = ~n23934 ;
  assign y6649 = n23936 ;
  assign y6650 = ~n23937 ;
  assign y6651 = n23939 ;
  assign y6652 = ~n23940 ;
  assign y6653 = ~n23942 ;
  assign y6654 = ~n23944 ;
  assign y6655 = n23952 ;
  assign y6656 = ~n23954 ;
  assign y6657 = ~1'b0 ;
  assign y6658 = n23964 ;
  assign y6659 = n23965 ;
  assign y6660 = n23968 ;
  assign y6661 = n7759 ;
  assign y6662 = ~1'b0 ;
  assign y6663 = ~n23970 ;
  assign y6664 = n23974 ;
  assign y6665 = ~n23977 ;
  assign y6666 = ~n23983 ;
  assign y6667 = ~n23985 ;
  assign y6668 = n23988 ;
  assign y6669 = ~n23991 ;
  assign y6670 = n19073 ;
  assign y6671 = n23996 ;
  assign y6672 = ~1'b0 ;
  assign y6673 = ~n23998 ;
  assign y6674 = ~n24007 ;
  assign y6675 = ~n24015 ;
  assign y6676 = n24019 ;
  assign y6677 = n24020 ;
  assign y6678 = n24023 ;
  assign y6679 = ~n24024 ;
  assign y6680 = ~n24028 ;
  assign y6681 = n24030 ;
  assign y6682 = ~1'b0 ;
  assign y6683 = n24035 ;
  assign y6684 = ~1'b0 ;
  assign y6685 = ~1'b0 ;
  assign y6686 = n24039 ;
  assign y6687 = ~n24042 ;
  assign y6688 = n24045 ;
  assign y6689 = n24048 ;
  assign y6690 = ~n24053 ;
  assign y6691 = ~n24055 ;
  assign y6692 = ~1'b0 ;
  assign y6693 = ~n24058 ;
  assign y6694 = ~n24061 ;
  assign y6695 = ~n24062 ;
  assign y6696 = n24068 ;
  assign y6697 = n24069 ;
  assign y6698 = ~n24073 ;
  assign y6699 = ~1'b0 ;
  assign y6700 = n24074 ;
  assign y6701 = ~n24077 ;
  assign y6702 = ~1'b0 ;
  assign y6703 = n24079 ;
  assign y6704 = ~n24083 ;
  assign y6705 = ~n24091 ;
  assign y6706 = ~n24098 ;
  assign y6707 = ~n24099 ;
  assign y6708 = ~n24100 ;
  assign y6709 = ~n24102 ;
  assign y6710 = ~1'b0 ;
  assign y6711 = ~n24110 ;
  assign y6712 = n24113 ;
  assign y6713 = ~n24114 ;
  assign y6714 = ~n24117 ;
  assign y6715 = ~n24118 ;
  assign y6716 = n24121 ;
  assign y6717 = n24125 ;
  assign y6718 = ~n24131 ;
  assign y6719 = n24134 ;
  assign y6720 = ~n24141 ;
  assign y6721 = n24143 ;
  assign y6722 = ~1'b0 ;
  assign y6723 = ~1'b0 ;
  assign y6724 = n24146 ;
  assign y6725 = ~n24148 ;
  assign y6726 = ~1'b0 ;
  assign y6727 = ~1'b0 ;
  assign y6728 = ~1'b0 ;
  assign y6729 = ~n24152 ;
  assign y6730 = ~1'b0 ;
  assign y6731 = n24159 ;
  assign y6732 = ~n24165 ;
  assign y6733 = n24170 ;
  assign y6734 = n24171 ;
  assign y6735 = n24172 ;
  assign y6736 = ~1'b0 ;
  assign y6737 = ~1'b0 ;
  assign y6738 = ~n24173 ;
  assign y6739 = ~n24175 ;
  assign y6740 = ~1'b0 ;
  assign y6741 = n24178 ;
  assign y6742 = n24183 ;
  assign y6743 = ~n24184 ;
  assign y6744 = ~n24187 ;
  assign y6745 = ~1'b0 ;
  assign y6746 = ~1'b0 ;
  assign y6747 = n24190 ;
  assign y6748 = n24198 ;
  assign y6749 = ~n24202 ;
  assign y6750 = n24203 ;
  assign y6751 = ~n24204 ;
  assign y6752 = n13723 ;
  assign y6753 = ~n24209 ;
  assign y6754 = ~n24211 ;
  assign y6755 = n24212 ;
  assign y6756 = n24214 ;
  assign y6757 = n24216 ;
  assign y6758 = n24218 ;
  assign y6759 = n24222 ;
  assign y6760 = n24223 ;
  assign y6761 = n24224 ;
  assign y6762 = n24228 ;
  assign y6763 = n24230 ;
  assign y6764 = ~n24236 ;
  assign y6765 = ~n24244 ;
  assign y6766 = n24247 ;
  assign y6767 = ~n24248 ;
  assign y6768 = n24250 ;
  assign y6769 = ~n24255 ;
  assign y6770 = ~n24261 ;
  assign y6771 = ~n24263 ;
  assign y6772 = ~n24265 ;
  assign y6773 = n24267 ;
  assign y6774 = ~1'b0 ;
  assign y6775 = ~1'b0 ;
  assign y6776 = ~n24271 ;
  assign y6777 = n24273 ;
  assign y6778 = ~n24274 ;
  assign y6779 = n24276 ;
  assign y6780 = ~n24279 ;
  assign y6781 = n24284 ;
  assign y6782 = ~n24294 ;
  assign y6783 = ~1'b0 ;
  assign y6784 = n24296 ;
  assign y6785 = n24298 ;
  assign y6786 = ~1'b0 ;
  assign y6787 = ~n24301 ;
  assign y6788 = ~n24302 ;
  assign y6789 = n24303 ;
  assign y6790 = n24305 ;
  assign y6791 = ~1'b0 ;
  assign y6792 = ~1'b0 ;
  assign y6793 = n24307 ;
  assign y6794 = n24308 ;
  assign y6795 = n24313 ;
  assign y6796 = ~1'b0 ;
  assign y6797 = ~n24314 ;
  assign y6798 = ~n24316 ;
  assign y6799 = n24321 ;
  assign y6800 = n24325 ;
  assign y6801 = ~n24326 ;
  assign y6802 = n24328 ;
  assign y6803 = n24329 ;
  assign y6804 = n24331 ;
  assign y6805 = n24339 ;
  assign y6806 = ~n20494 ;
  assign y6807 = n24340 ;
  assign y6808 = ~1'b0 ;
  assign y6809 = ~n24345 ;
  assign y6810 = ~n24347 ;
  assign y6811 = n24348 ;
  assign y6812 = n24354 ;
  assign y6813 = n24355 ;
  assign y6814 = ~n24359 ;
  assign y6815 = ~n24360 ;
  assign y6816 = ~n24361 ;
  assign y6817 = ~n24362 ;
  assign y6818 = ~1'b0 ;
  assign y6819 = ~n24363 ;
  assign y6820 = ~1'b0 ;
  assign y6821 = n24365 ;
  assign y6822 = ~n24367 ;
  assign y6823 = n24369 ;
  assign y6824 = ~n24372 ;
  assign y6825 = ~n24377 ;
  assign y6826 = ~1'b0 ;
  assign y6827 = ~n24380 ;
  assign y6828 = ~n24387 ;
  assign y6829 = n24389 ;
  assign y6830 = ~n24392 ;
  assign y6831 = ~n24393 ;
  assign y6832 = ~1'b0 ;
  assign y6833 = ~n24396 ;
  assign y6834 = ~n24398 ;
  assign y6835 = ~n24402 ;
  assign y6836 = ~n24403 ;
  assign y6837 = ~1'b0 ;
  assign y6838 = ~1'b0 ;
  assign y6839 = n24405 ;
  assign y6840 = ~n24406 ;
  assign y6841 = ~1'b0 ;
  assign y6842 = ~n24412 ;
  assign y6843 = n24417 ;
  assign y6844 = n24419 ;
  assign y6845 = ~n24420 ;
  assign y6846 = n24424 ;
  assign y6847 = ~1'b0 ;
  assign y6848 = n24430 ;
  assign y6849 = n24432 ;
  assign y6850 = ~1'b0 ;
  assign y6851 = ~n24434 ;
  assign y6852 = n24439 ;
  assign y6853 = ~n24444 ;
  assign y6854 = n24451 ;
  assign y6855 = ~1'b0 ;
  assign y6856 = ~n24460 ;
  assign y6857 = ~n24462 ;
  assign y6858 = n24463 ;
  assign y6859 = ~1'b0 ;
  assign y6860 = ~n24467 ;
  assign y6861 = ~n24474 ;
  assign y6862 = ~n24478 ;
  assign y6863 = ~n24483 ;
  assign y6864 = ~n24485 ;
  assign y6865 = n24487 ;
  assign y6866 = n24489 ;
  assign y6867 = ~1'b0 ;
  assign y6868 = ~n24491 ;
  assign y6869 = n24494 ;
  assign y6870 = ~n24495 ;
  assign y6871 = ~n24498 ;
  assign y6872 = ~n24500 ;
  assign y6873 = ~n24513 ;
  assign y6874 = ~n24524 ;
  assign y6875 = n24527 ;
  assign y6876 = n24528 ;
  assign y6877 = ~n24534 ;
  assign y6878 = n24536 ;
  assign y6879 = ~n24541 ;
  assign y6880 = ~n24544 ;
  assign y6881 = ~n24545 ;
  assign y6882 = ~n24547 ;
  assign y6883 = n24550 ;
  assign y6884 = ~1'b0 ;
  assign y6885 = n24551 ;
  assign y6886 = n24554 ;
  assign y6887 = n24557 ;
  assign y6888 = n24561 ;
  assign y6889 = ~1'b0 ;
  assign y6890 = n24575 ;
  assign y6891 = ~n24589 ;
  assign y6892 = n24590 ;
  assign y6893 = n24592 ;
  assign y6894 = ~1'b0 ;
  assign y6895 = n24594 ;
  assign y6896 = n24595 ;
  assign y6897 = n24599 ;
  assign y6898 = ~n24601 ;
  assign y6899 = ~n24607 ;
  assign y6900 = ~n24610 ;
  assign y6901 = n24611 ;
  assign y6902 = n24613 ;
  assign y6903 = ~n24615 ;
  assign y6904 = ~n24616 ;
  assign y6905 = n24623 ;
  assign y6906 = n24626 ;
  assign y6907 = ~n24629 ;
  assign y6908 = n4975 ;
  assign y6909 = n24632 ;
  assign y6910 = ~n24633 ;
  assign y6911 = ~1'b0 ;
  assign y6912 = ~n24635 ;
  assign y6913 = ~n24637 ;
  assign y6914 = ~n24639 ;
  assign y6915 = ~n24646 ;
  assign y6916 = ~n24652 ;
  assign y6917 = n24660 ;
  assign y6918 = ~1'b0 ;
  assign y6919 = ~n24663 ;
  assign y6920 = ~1'b0 ;
  assign y6921 = n24664 ;
  assign y6922 = n24673 ;
  assign y6923 = ~n24674 ;
  assign y6924 = ~n24677 ;
  assign y6925 = n24681 ;
  assign y6926 = ~n24684 ;
  assign y6927 = n24685 ;
  assign y6928 = ~n24686 ;
  assign y6929 = n21888 ;
  assign y6930 = ~n24690 ;
  assign y6931 = ~n24694 ;
  assign y6932 = ~n24697 ;
  assign y6933 = ~n24701 ;
  assign y6934 = n24706 ;
  assign y6935 = n24710 ;
  assign y6936 = ~n24713 ;
  assign y6937 = n24714 ;
  assign y6938 = n24726 ;
  assign y6939 = ~1'b0 ;
  assign y6940 = n24728 ;
  assign y6941 = ~n24731 ;
  assign y6942 = ~n24732 ;
  assign y6943 = n24733 ;
  assign y6944 = ~n24736 ;
  assign y6945 = n24737 ;
  assign y6946 = n24740 ;
  assign y6947 = ~n24741 ;
  assign y6948 = ~n24743 ;
  assign y6949 = n24749 ;
  assign y6950 = ~1'b0 ;
  assign y6951 = ~n24751 ;
  assign y6952 = ~1'b0 ;
  assign y6953 = ~n24752 ;
  assign y6954 = ~n24757 ;
  assign y6955 = n24758 ;
  assign y6956 = ~n24760 ;
  assign y6957 = ~1'b0 ;
  assign y6958 = n24761 ;
  assign y6959 = ~n24762 ;
  assign y6960 = n24764 ;
  assign y6961 = n24765 ;
  assign y6962 = ~n24773 ;
  assign y6963 = n24778 ;
  assign y6964 = ~n24781 ;
  assign y6965 = n24787 ;
  assign y6966 = ~n24788 ;
  assign y6967 = ~n24791 ;
  assign y6968 = ~n24795 ;
  assign y6969 = n24796 ;
  assign y6970 = n24797 ;
  assign y6971 = n24799 ;
  assign y6972 = n24804 ;
  assign y6973 = n24808 ;
  assign y6974 = ~n24815 ;
  assign y6975 = n24825 ;
  assign y6976 = ~n24827 ;
  assign y6977 = ~n24839 ;
  assign y6978 = n24840 ;
  assign y6979 = n24844 ;
  assign y6980 = ~n24849 ;
  assign y6981 = n24852 ;
  assign y6982 = n24858 ;
  assign y6983 = n24866 ;
  assign y6984 = ~1'b0 ;
  assign y6985 = ~1'b0 ;
  assign y6986 = ~n24867 ;
  assign y6987 = ~1'b0 ;
  assign y6988 = ~n24870 ;
  assign y6989 = ~n24877 ;
  assign y6990 = n24881 ;
  assign y6991 = n24883 ;
  assign y6992 = n24885 ;
  assign y6993 = ~n24888 ;
  assign y6994 = n24889 ;
  assign y6995 = n2130 ;
  assign y6996 = ~n24891 ;
  assign y6997 = n24900 ;
  assign y6998 = n24902 ;
  assign y6999 = n24903 ;
  assign y7000 = ~n24907 ;
  assign y7001 = n24912 ;
  assign y7002 = ~n24916 ;
  assign y7003 = ~n24920 ;
  assign y7004 = ~1'b0 ;
  assign y7005 = n24921 ;
  assign y7006 = n24922 ;
  assign y7007 = ~n24923 ;
  assign y7008 = n24930 ;
  assign y7009 = n24931 ;
  assign y7010 = n24936 ;
  assign y7011 = n24938 ;
  assign y7012 = n24939 ;
  assign y7013 = n24947 ;
  assign y7014 = ~1'b0 ;
  assign y7015 = n24954 ;
  assign y7016 = n24956 ;
  assign y7017 = n24958 ;
  assign y7018 = ~n10987 ;
  assign y7019 = ~1'b0 ;
  assign y7020 = ~n24963 ;
  assign y7021 = n24969 ;
  assign y7022 = n24973 ;
  assign y7023 = ~n24975 ;
  assign y7024 = ~1'b0 ;
  assign y7025 = ~n24977 ;
  assign y7026 = ~n24982 ;
  assign y7027 = ~n24983 ;
  assign y7028 = n24987 ;
  assign y7029 = n24990 ;
  assign y7030 = ~n24993 ;
  assign y7031 = ~1'b0 ;
  assign y7032 = n24995 ;
  assign y7033 = n25000 ;
  assign y7034 = n25002 ;
  assign y7035 = ~n25005 ;
  assign y7036 = ~n25006 ;
  assign y7037 = ~1'b0 ;
  assign y7038 = n25007 ;
  assign y7039 = ~n25009 ;
  assign y7040 = ~n25010 ;
  assign y7041 = n25011 ;
  assign y7042 = n25015 ;
  assign y7043 = ~1'b0 ;
  assign y7044 = n25020 ;
  assign y7045 = n25022 ;
  assign y7046 = ~n25024 ;
  assign y7047 = ~1'b0 ;
  assign y7048 = ~n25026 ;
  assign y7049 = n25029 ;
  assign y7050 = n25034 ;
  assign y7051 = ~1'b0 ;
  assign y7052 = n25040 ;
  assign y7053 = ~n25045 ;
  assign y7054 = n25049 ;
  assign y7055 = ~n25055 ;
  assign y7056 = ~n25065 ;
  assign y7057 = ~1'b0 ;
  assign y7058 = n25070 ;
  assign y7059 = n25071 ;
  assign y7060 = ~n25076 ;
  assign y7061 = ~1'b0 ;
  assign y7062 = ~n25078 ;
  assign y7063 = ~n25082 ;
  assign y7064 = n25083 ;
  assign y7065 = n25086 ;
  assign y7066 = ~n25090 ;
  assign y7067 = n25091 ;
  assign y7068 = ~n25092 ;
  assign y7069 = n25098 ;
  assign y7070 = ~n25100 ;
  assign y7071 = ~n25101 ;
  assign y7072 = n25105 ;
  assign y7073 = ~n25106 ;
  assign y7074 = n25110 ;
  assign y7075 = n25112 ;
  assign y7076 = ~n25115 ;
  assign y7077 = ~n25116 ;
  assign y7078 = ~n25118 ;
  assign y7079 = ~n25120 ;
  assign y7080 = n25121 ;
  assign y7081 = ~1'b0 ;
  assign y7082 = ~1'b0 ;
  assign y7083 = ~1'b0 ;
  assign y7084 = n25124 ;
  assign y7085 = n6671 ;
  assign y7086 = ~n25130 ;
  assign y7087 = ~1'b0 ;
  assign y7088 = ~n25138 ;
  assign y7089 = n25139 ;
  assign y7090 = ~n25142 ;
  assign y7091 = ~n25148 ;
  assign y7092 = ~n25152 ;
  assign y7093 = ~1'b0 ;
  assign y7094 = ~n25154 ;
  assign y7095 = ~n25155 ;
  assign y7096 = n25159 ;
  assign y7097 = ~1'b0 ;
  assign y7098 = ~1'b0 ;
  assign y7099 = ~n25167 ;
  assign y7100 = n25168 ;
  assign y7101 = 1'b0 ;
  assign y7102 = ~n25169 ;
  assign y7103 = ~n25171 ;
  assign y7104 = ~n25178 ;
  assign y7105 = ~n25180 ;
  assign y7106 = ~n25182 ;
  assign y7107 = ~1'b0 ;
  assign y7108 = n25184 ;
  assign y7109 = ~1'b0 ;
  assign y7110 = n25189 ;
  assign y7111 = n25191 ;
  assign y7112 = ~n25195 ;
  assign y7113 = ~n25201 ;
  assign y7114 = n25202 ;
  assign y7115 = ~n25213 ;
  assign y7116 = n25216 ;
  assign y7117 = n25217 ;
  assign y7118 = n25220 ;
  assign y7119 = n25222 ;
  assign y7120 = n25223 ;
  assign y7121 = ~n25226 ;
  assign y7122 = ~1'b0 ;
  assign y7123 = ~1'b0 ;
  assign y7124 = 1'b0 ;
  assign y7125 = n25233 ;
  assign y7126 = n25235 ;
  assign y7127 = n25236 ;
  assign y7128 = ~n25240 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = ~1'b0 ;
  assign y7131 = n25243 ;
  assign y7132 = n25244 ;
  assign y7133 = n25247 ;
  assign y7134 = ~n25252 ;
  assign y7135 = n25254 ;
  assign y7136 = ~1'b0 ;
  assign y7137 = n25255 ;
  assign y7138 = ~1'b0 ;
  assign y7139 = n25259 ;
  assign y7140 = n25260 ;
  assign y7141 = ~n25265 ;
  assign y7142 = ~n25268 ;
  assign y7143 = ~n25274 ;
  assign y7144 = n25278 ;
  assign y7145 = ~n25282 ;
  assign y7146 = ~n25283 ;
  assign y7147 = ~n25284 ;
  assign y7148 = n25285 ;
  assign y7149 = ~n25287 ;
  assign y7150 = ~1'b0 ;
  assign y7151 = n25288 ;
  assign y7152 = ~n25292 ;
  assign y7153 = n25295 ;
  assign y7154 = ~n25297 ;
  assign y7155 = ~n25301 ;
  assign y7156 = ~n25302 ;
  assign y7157 = ~n25308 ;
  assign y7158 = n25309 ;
  assign y7159 = n25311 ;
  assign y7160 = ~n25317 ;
  assign y7161 = n25320 ;
  assign y7162 = ~n25327 ;
  assign y7163 = n25333 ;
  assign y7164 = ~n25340 ;
  assign y7165 = ~n25344 ;
  assign y7166 = n25347 ;
  assign y7167 = n25355 ;
  assign y7168 = n25367 ;
  assign y7169 = n25372 ;
  assign y7170 = n25374 ;
  assign y7171 = ~n25383 ;
  assign y7172 = ~n25387 ;
  assign y7173 = ~n25389 ;
  assign y7174 = ~1'b0 ;
  assign y7175 = n25393 ;
  assign y7176 = ~n25395 ;
  assign y7177 = n25398 ;
  assign y7178 = ~n25400 ;
  assign y7179 = ~n25402 ;
  assign y7180 = ~n23320 ;
  assign y7181 = ~n25403 ;
  assign y7182 = n25405 ;
  assign y7183 = ~n25406 ;
  assign y7184 = n25407 ;
  assign y7185 = ~n25409 ;
  assign y7186 = ~n25410 ;
  assign y7187 = ~n25413 ;
  assign y7188 = n25415 ;
  assign y7189 = ~n25418 ;
  assign y7190 = n25426 ;
  assign y7191 = n25429 ;
  assign y7192 = ~n25435 ;
  assign y7193 = n25441 ;
  assign y7194 = n25445 ;
  assign y7195 = n25447 ;
  assign y7196 = ~n25453 ;
  assign y7197 = ~n25455 ;
  assign y7198 = ~1'b0 ;
  assign y7199 = ~n25457 ;
  assign y7200 = ~n25462 ;
  assign y7201 = ~n25463 ;
  assign y7202 = ~n25464 ;
  assign y7203 = ~n25465 ;
  assign y7204 = ~1'b0 ;
  assign y7205 = ~n25466 ;
  assign y7206 = n25468 ;
  assign y7207 = ~n25469 ;
  assign y7208 = ~n25470 ;
  assign y7209 = ~n25472 ;
  assign y7210 = n25475 ;
  assign y7211 = n25477 ;
  assign y7212 = n25480 ;
  assign y7213 = ~n25482 ;
  assign y7214 = n25485 ;
  assign y7215 = ~n25489 ;
  assign y7216 = ~1'b0 ;
  assign y7217 = ~n25493 ;
  assign y7218 = ~n25502 ;
  assign y7219 = ~n25504 ;
  assign y7220 = n25507 ;
  assign y7221 = n25508 ;
  assign y7222 = ~n25509 ;
  assign y7223 = n25510 ;
  assign y7224 = n25513 ;
  assign y7225 = n25526 ;
  assign y7226 = ~n25530 ;
  assign y7227 = ~n25531 ;
  assign y7228 = ~n25532 ;
  assign y7229 = n25538 ;
  assign y7230 = ~n25544 ;
  assign y7231 = ~n25545 ;
  assign y7232 = n25547 ;
  assign y7233 = n25551 ;
  assign y7234 = n25552 ;
  assign y7235 = n25556 ;
  assign y7236 = n25558 ;
  assign y7237 = ~1'b0 ;
  assign y7238 = ~1'b0 ;
  assign y7239 = ~n25559 ;
  assign y7240 = n25566 ;
  assign y7241 = 1'b0 ;
  assign y7242 = n25571 ;
  assign y7243 = n25572 ;
  assign y7244 = n25577 ;
  assign y7245 = ~n25582 ;
  assign y7246 = ~n25583 ;
  assign y7247 = ~n25590 ;
  assign y7248 = n25592 ;
  assign y7249 = ~1'b0 ;
  assign y7250 = ~n25593 ;
  assign y7251 = n25595 ;
  assign y7252 = n25598 ;
  assign y7253 = ~n25602 ;
  assign y7254 = ~1'b0 ;
  assign y7255 = n25606 ;
  assign y7256 = ~n25615 ;
  assign y7257 = n22046 ;
  assign y7258 = n25620 ;
  assign y7259 = ~n25624 ;
  assign y7260 = n25625 ;
  assign y7261 = ~1'b0 ;
  assign y7262 = n25637 ;
  assign y7263 = ~1'b0 ;
  assign y7264 = ~n25646 ;
  assign y7265 = ~n25647 ;
  assign y7266 = ~n25649 ;
  assign y7267 = ~n25185 ;
  assign y7268 = ~n25652 ;
  assign y7269 = n25655 ;
  assign y7270 = ~n25659 ;
  assign y7271 = n25662 ;
  assign y7272 = ~n25665 ;
  assign y7273 = ~1'b0 ;
  assign y7274 = ~n25669 ;
  assign y7275 = n25673 ;
  assign y7276 = n25675 ;
  assign y7277 = n25679 ;
  assign y7278 = n25683 ;
  assign y7279 = ~n25688 ;
  assign y7280 = ~n25695 ;
  assign y7281 = n25696 ;
  assign y7282 = ~n25701 ;
  assign y7283 = ~n25704 ;
  assign y7284 = n25714 ;
  assign y7285 = ~n25719 ;
  assign y7286 = n25720 ;
  assign y7287 = ~n25722 ;
  assign y7288 = 1'b0 ;
  assign y7289 = ~n25728 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = ~n25729 ;
  assign y7292 = ~n25730 ;
  assign y7293 = ~1'b0 ;
  assign y7294 = n25731 ;
  assign y7295 = ~n25733 ;
  assign y7296 = ~n25736 ;
  assign y7297 = ~1'b0 ;
  assign y7298 = ~n25745 ;
  assign y7299 = ~1'b0 ;
  assign y7300 = n25750 ;
  assign y7301 = ~n25755 ;
  assign y7302 = ~n25756 ;
  assign y7303 = ~n25757 ;
  assign y7304 = ~1'b0 ;
  assign y7305 = ~n25758 ;
  assign y7306 = ~n25765 ;
  assign y7307 = ~1'b0 ;
  assign y7308 = ~n25776 ;
  assign y7309 = ~n25778 ;
  assign y7310 = ~n25784 ;
  assign y7311 = ~n25787 ;
  assign y7312 = ~n25788 ;
  assign y7313 = ~n25793 ;
  assign y7314 = n25798 ;
  assign y7315 = n25801 ;
  assign y7316 = ~n25802 ;
  assign y7317 = ~n25810 ;
  assign y7318 = ~n25812 ;
  assign y7319 = n25813 ;
  assign y7320 = ~n25815 ;
  assign y7321 = ~n25817 ;
  assign y7322 = ~n25821 ;
  assign y7323 = n25825 ;
  assign y7324 = ~n25826 ;
  assign y7325 = n25828 ;
  assign y7326 = ~1'b0 ;
  assign y7327 = n25830 ;
  assign y7328 = ~n25831 ;
  assign y7329 = ~n25832 ;
  assign y7330 = n25835 ;
  assign y7331 = n25837 ;
  assign y7332 = ~n25846 ;
  assign y7333 = ~1'b0 ;
  assign y7334 = n25847 ;
  assign y7335 = ~n25854 ;
  assign y7336 = n25857 ;
  assign y7337 = ~n25865 ;
  assign y7338 = n25868 ;
  assign y7339 = ~n25871 ;
  assign y7340 = n25873 ;
  assign y7341 = n25874 ;
  assign y7342 = ~n25878 ;
  assign y7343 = ~n25879 ;
  assign y7344 = n25880 ;
  assign y7345 = ~n25883 ;
  assign y7346 = ~1'b0 ;
  assign y7347 = n22878 ;
  assign y7348 = n25885 ;
  assign y7349 = n25886 ;
  assign y7350 = n25902 ;
  assign y7351 = n25904 ;
  assign y7352 = n25906 ;
  assign y7353 = n25911 ;
  assign y7354 = n25917 ;
  assign y7355 = ~n25920 ;
  assign y7356 = n25921 ;
  assign y7357 = ~n25922 ;
  assign y7358 = n25925 ;
  assign y7359 = ~n25927 ;
  assign y7360 = n25930 ;
  assign y7361 = ~n25936 ;
  assign y7362 = ~n25944 ;
  assign y7363 = n25945 ;
  assign y7364 = ~1'b0 ;
  assign y7365 = ~n25953 ;
  assign y7366 = n25955 ;
  assign y7367 = ~n25958 ;
  assign y7368 = n25964 ;
  assign y7369 = ~n25968 ;
  assign y7370 = ~n25969 ;
  assign y7371 = ~n25976 ;
  assign y7372 = n25983 ;
  assign y7373 = ~n10210 ;
  assign y7374 = n25990 ;
  assign y7375 = ~1'b0 ;
  assign y7376 = n25993 ;
  assign y7377 = ~n26001 ;
  assign y7378 = ~n26004 ;
  assign y7379 = ~1'b0 ;
  assign y7380 = n26006 ;
  assign y7381 = n26022 ;
  assign y7382 = ~n26027 ;
  assign y7383 = n26028 ;
  assign y7384 = ~n26035 ;
  assign y7385 = ~n26037 ;
  assign y7386 = ~1'b0 ;
  assign y7387 = ~n26039 ;
  assign y7388 = n26040 ;
  assign y7389 = ~n26043 ;
  assign y7390 = ~n26049 ;
  assign y7391 = ~n26050 ;
  assign y7392 = ~n26051 ;
  assign y7393 = ~n26052 ;
  assign y7394 = ~n26059 ;
  assign y7395 = ~n26061 ;
  assign y7396 = ~1'b0 ;
  assign y7397 = ~n26065 ;
  assign y7398 = n26066 ;
  assign y7399 = n26067 ;
  assign y7400 = ~n26072 ;
  assign y7401 = n26085 ;
  assign y7402 = n26087 ;
  assign y7403 = ~1'b0 ;
  assign y7404 = n26088 ;
  assign y7405 = ~n26091 ;
  assign y7406 = n26092 ;
  assign y7407 = ~n26094 ;
  assign y7408 = ~n26099 ;
  assign y7409 = ~n26104 ;
  assign y7410 = n26108 ;
  assign y7411 = ~n26109 ;
  assign y7412 = ~n26110 ;
  assign y7413 = n26122 ;
  assign y7414 = ~1'b0 ;
  assign y7415 = ~1'b0 ;
  assign y7416 = ~n26125 ;
  assign y7417 = ~n26128 ;
  assign y7418 = ~n26130 ;
  assign y7419 = ~1'b0 ;
  assign y7420 = ~n26133 ;
  assign y7421 = ~n26136 ;
  assign y7422 = n26137 ;
  assign y7423 = ~1'b0 ;
  assign y7424 = ~n26147 ;
  assign y7425 = ~n26148 ;
  assign y7426 = ~n26149 ;
  assign y7427 = ~1'b0 ;
  assign y7428 = ~n26153 ;
  assign y7429 = ~n26160 ;
  assign y7430 = ~n26167 ;
  assign y7431 = n26170 ;
  assign y7432 = ~n26172 ;
  assign y7433 = ~n26173 ;
  assign y7434 = n26175 ;
  assign y7435 = n26177 ;
  assign y7436 = ~n26178 ;
  assign y7437 = ~n26180 ;
  assign y7438 = n26182 ;
  assign y7439 = n26191 ;
  assign y7440 = n26197 ;
  assign y7441 = n26200 ;
  assign y7442 = ~1'b0 ;
  assign y7443 = ~n26203 ;
  assign y7444 = ~n26207 ;
  assign y7445 = n26209 ;
  assign y7446 = n26212 ;
  assign y7447 = ~n26215 ;
  assign y7448 = n26219 ;
  assign y7449 = ~n26222 ;
  assign y7450 = n26223 ;
  assign y7451 = n26224 ;
  assign y7452 = ~n26230 ;
  assign y7453 = ~n26231 ;
  assign y7454 = n26234 ;
  assign y7455 = ~1'b0 ;
  assign y7456 = n26235 ;
  assign y7457 = ~n26236 ;
  assign y7458 = n26238 ;
  assign y7459 = ~n26242 ;
  assign y7460 = ~n26245 ;
  assign y7461 = ~n26246 ;
  assign y7462 = n26247 ;
  assign y7463 = ~n26248 ;
  assign y7464 = n26250 ;
  assign y7465 = n26253 ;
  assign y7466 = n26254 ;
  assign y7467 = ~1'b0 ;
  assign y7468 = ~1'b0 ;
  assign y7469 = ~n26262 ;
  assign y7470 = n26266 ;
  assign y7471 = ~n26270 ;
  assign y7472 = ~1'b0 ;
  assign y7473 = ~n26279 ;
  assign y7474 = ~n26281 ;
  assign y7475 = n26282 ;
  assign y7476 = ~n26286 ;
  assign y7477 = n26288 ;
  assign y7478 = ~n26291 ;
  assign y7479 = n7124 ;
  assign y7480 = n26294 ;
  assign y7481 = n26298 ;
  assign y7482 = n26300 ;
  assign y7483 = ~n26302 ;
  assign y7484 = n26303 ;
  assign y7485 = ~n26305 ;
  assign y7486 = n26307 ;
  assign y7487 = ~n26308 ;
  assign y7488 = n26311 ;
  assign y7489 = ~n26313 ;
  assign y7490 = n3228 ;
  assign y7491 = n26316 ;
  assign y7492 = n26317 ;
  assign y7493 = n26320 ;
  assign y7494 = ~n26325 ;
  assign y7495 = n26326 ;
  assign y7496 = ~n26331 ;
  assign y7497 = n26332 ;
  assign y7498 = n26333 ;
  assign y7499 = ~n26337 ;
  assign y7500 = n26340 ;
  assign y7501 = ~n26348 ;
  assign y7502 = ~1'b0 ;
  assign y7503 = ~n26350 ;
  assign y7504 = n26353 ;
  assign y7505 = n26354 ;
  assign y7506 = n26359 ;
  assign y7507 = n26373 ;
  assign y7508 = ~n17391 ;
  assign y7509 = ~n26382 ;
  assign y7510 = n26388 ;
  assign y7511 = ~n26397 ;
  assign y7512 = ~n26401 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = n26403 ;
  assign y7515 = ~1'b0 ;
  assign y7516 = ~1'b0 ;
  assign y7517 = ~n26404 ;
  assign y7518 = n26406 ;
  assign y7519 = n26407 ;
  assign y7520 = ~n26419 ;
  assign y7521 = n26421 ;
  assign y7522 = n26426 ;
  assign y7523 = ~n26428 ;
  assign y7524 = n26434 ;
  assign y7525 = ~n26437 ;
  assign y7526 = n26438 ;
  assign y7527 = ~1'b0 ;
  assign y7528 = ~n26445 ;
  assign y7529 = ~n26449 ;
  assign y7530 = n26451 ;
  assign y7531 = n26456 ;
  assign y7532 = n26458 ;
  assign y7533 = n26459 ;
  assign y7534 = n26469 ;
  assign y7535 = n26470 ;
  assign y7536 = ~n26471 ;
  assign y7537 = ~n26479 ;
  assign y7538 = ~n26480 ;
  assign y7539 = n26483 ;
  assign y7540 = ~1'b0 ;
  assign y7541 = ~n26484 ;
  assign y7542 = ~n26490 ;
  assign y7543 = ~n26491 ;
  assign y7544 = n26494 ;
  assign y7545 = n26496 ;
  assign y7546 = ~1'b0 ;
  assign y7547 = ~1'b0 ;
  assign y7548 = ~n26498 ;
  assign y7549 = ~n26503 ;
  assign y7550 = ~n26509 ;
  assign y7551 = ~n26511 ;
  assign y7552 = ~n26514 ;
  assign y7553 = ~n26519 ;
  assign y7554 = ~n26521 ;
  assign y7555 = n26522 ;
  assign y7556 = n26524 ;
  assign y7557 = ~1'b0 ;
  assign y7558 = n26528 ;
  assign y7559 = n26533 ;
  assign y7560 = ~1'b0 ;
  assign y7561 = ~n26537 ;
  assign y7562 = ~n26542 ;
  assign y7563 = ~n26543 ;
  assign y7564 = ~n26544 ;
  assign y7565 = n26546 ;
  assign y7566 = ~1'b0 ;
  assign y7567 = ~1'b0 ;
  assign y7568 = n26547 ;
  assign y7569 = ~n26552 ;
  assign y7570 = n26553 ;
  assign y7571 = ~n26554 ;
  assign y7572 = ~n10238 ;
  assign y7573 = ~n26556 ;
  assign y7574 = n26560 ;
  assign y7575 = n26564 ;
  assign y7576 = n26569 ;
  assign y7577 = n26574 ;
  assign y7578 = ~n26576 ;
  assign y7579 = n26581 ;
  assign y7580 = n26582 ;
  assign y7581 = ~n26586 ;
  assign y7582 = n26593 ;
  assign y7583 = n26594 ;
  assign y7584 = ~1'b0 ;
  assign y7585 = ~1'b0 ;
  assign y7586 = ~n26595 ;
  assign y7587 = n26596 ;
  assign y7588 = n26598 ;
  assign y7589 = ~n26601 ;
  assign y7590 = n26604 ;
  assign y7591 = n26609 ;
  assign y7592 = n26612 ;
  assign y7593 = ~n26614 ;
  assign y7594 = ~n26616 ;
  assign y7595 = ~n26619 ;
  assign y7596 = n26620 ;
  assign y7597 = ~n26622 ;
  assign y7598 = ~n26625 ;
  assign y7599 = ~n26629 ;
  assign y7600 = ~n26632 ;
  assign y7601 = ~n26633 ;
  assign y7602 = ~n26634 ;
  assign y7603 = n26641 ;
  assign y7604 = n26643 ;
  assign y7605 = ~1'b0 ;
  assign y7606 = ~1'b0 ;
  assign y7607 = ~n26646 ;
  assign y7608 = ~n26651 ;
  assign y7609 = n26656 ;
  assign y7610 = ~1'b0 ;
  assign y7611 = ~1'b0 ;
  assign y7612 = ~n26663 ;
  assign y7613 = ~n26666 ;
  assign y7614 = ~n26667 ;
  assign y7615 = ~n26668 ;
  assign y7616 = n26669 ;
  assign y7617 = n26670 ;
  assign y7618 = n26675 ;
  assign y7619 = n26692 ;
  assign y7620 = ~1'b0 ;
  assign y7621 = n26696 ;
  assign y7622 = ~n26698 ;
  assign y7623 = ~n26709 ;
  assign y7624 = n26711 ;
  assign y7625 = n26712 ;
  assign y7626 = n26718 ;
  assign y7627 = n26724 ;
  assign y7628 = n26726 ;
  assign y7629 = ~n26731 ;
  assign y7630 = n26732 ;
  assign y7631 = n18522 ;
  assign y7632 = ~n26734 ;
  assign y7633 = n26740 ;
  assign y7634 = ~n26744 ;
  assign y7635 = n26746 ;
  assign y7636 = n26751 ;
  assign y7637 = ~n26756 ;
  assign y7638 = n26762 ;
  assign y7639 = n26765 ;
  assign y7640 = n26768 ;
  assign y7641 = ~n26773 ;
  assign y7642 = ~n26775 ;
  assign y7643 = ~n26777 ;
  assign y7644 = n26783 ;
  assign y7645 = n26787 ;
  assign y7646 = ~n26794 ;
  assign y7647 = n26795 ;
  assign y7648 = ~n26804 ;
  assign y7649 = ~n26806 ;
  assign y7650 = n26810 ;
  assign y7651 = n26814 ;
  assign y7652 = ~n26817 ;
  assign y7653 = n26818 ;
  assign y7654 = n26820 ;
  assign y7655 = n26822 ;
  assign y7656 = ~n26828 ;
  assign y7657 = ~n26829 ;
  assign y7658 = n26835 ;
  assign y7659 = ~n26839 ;
  assign y7660 = ~1'b0 ;
  assign y7661 = ~n26850 ;
  assign y7662 = ~n26853 ;
  assign y7663 = n26855 ;
  assign y7664 = ~n26860 ;
  assign y7665 = n26862 ;
  assign y7666 = ~1'b0 ;
  assign y7667 = n26864 ;
  assign y7668 = ~n26865 ;
  assign y7669 = n26870 ;
  assign y7670 = ~n26872 ;
  assign y7671 = n26873 ;
  assign y7672 = ~1'b0 ;
  assign y7673 = ~1'b0 ;
  assign y7674 = ~1'b0 ;
  assign y7675 = n26876 ;
  assign y7676 = ~1'b0 ;
  assign y7677 = ~n26877 ;
  assign y7678 = ~n26879 ;
  assign y7679 = ~n26881 ;
  assign y7680 = n26884 ;
  assign y7681 = n26889 ;
  assign y7682 = ~n26890 ;
  assign y7683 = n26891 ;
  assign y7684 = ~n26898 ;
  assign y7685 = ~n26900 ;
  assign y7686 = n26664 ;
  assign y7687 = n26902 ;
  assign y7688 = n26903 ;
  assign y7689 = ~n26905 ;
  assign y7690 = n26909 ;
  assign y7691 = ~n26917 ;
  assign y7692 = ~1'b0 ;
  assign y7693 = ~1'b0 ;
  assign y7694 = n26923 ;
  assign y7695 = ~n26926 ;
  assign y7696 = ~n26928 ;
  assign y7697 = ~n26930 ;
  assign y7698 = ~n26931 ;
  assign y7699 = n26934 ;
  assign y7700 = ~1'b0 ;
  assign y7701 = n26937 ;
  assign y7702 = ~n26941 ;
  assign y7703 = n26942 ;
  assign y7704 = ~n26946 ;
  assign y7705 = n26947 ;
  assign y7706 = ~n26954 ;
  assign y7707 = ~1'b0 ;
  assign y7708 = ~1'b0 ;
  assign y7709 = ~n26965 ;
  assign y7710 = ~n26966 ;
  assign y7711 = n26968 ;
  assign y7712 = ~n4263 ;
  assign y7713 = n26969 ;
  assign y7714 = ~n26971 ;
  assign y7715 = ~1'b0 ;
  assign y7716 = n26973 ;
  assign y7717 = n26984 ;
  assign y7718 = n26985 ;
  assign y7719 = ~1'b0 ;
  assign y7720 = ~1'b0 ;
  assign y7721 = ~n26997 ;
  assign y7722 = ~n26998 ;
  assign y7723 = n27002 ;
  assign y7724 = ~1'b0 ;
  assign y7725 = n27003 ;
  assign y7726 = ~n27009 ;
  assign y7727 = n27011 ;
  assign y7728 = ~1'b0 ;
  assign y7729 = n24928 ;
  assign y7730 = ~n27016 ;
  assign y7731 = n27019 ;
  assign y7732 = ~n27021 ;
  assign y7733 = n27024 ;
  assign y7734 = ~n27025 ;
  assign y7735 = n27028 ;
  assign y7736 = n27036 ;
  assign y7737 = ~n27038 ;
  assign y7738 = n27039 ;
  assign y7739 = n27042 ;
  assign y7740 = ~n27043 ;
  assign y7741 = n27045 ;
  assign y7742 = ~n27053 ;
  assign y7743 = n27060 ;
  assign y7744 = ~n27064 ;
  assign y7745 = ~1'b0 ;
  assign y7746 = n27067 ;
  assign y7747 = ~n27068 ;
  assign y7748 = ~n27070 ;
  assign y7749 = n27082 ;
  assign y7750 = ~n27083 ;
  assign y7751 = ~n27085 ;
  assign y7752 = ~n27087 ;
  assign y7753 = n27089 ;
  assign y7754 = ~n27095 ;
  assign y7755 = n27097 ;
  assign y7756 = ~n27102 ;
  assign y7757 = n27106 ;
  assign y7758 = ~n27110 ;
  assign y7759 = n27113 ;
  assign y7760 = ~1'b0 ;
  assign y7761 = n27115 ;
  assign y7762 = ~1'b0 ;
  assign y7763 = n27118 ;
  assign y7764 = ~1'b0 ;
  assign y7765 = n27120 ;
  assign y7766 = ~1'b0 ;
  assign y7767 = ~1'b0 ;
  assign y7768 = ~1'b0 ;
  assign y7769 = ~n27124 ;
  assign y7770 = ~n27126 ;
  assign y7771 = ~n27129 ;
  assign y7772 = n27132 ;
  assign y7773 = ~1'b0 ;
  assign y7774 = ~1'b0 ;
  assign y7775 = ~n27134 ;
  assign y7776 = n27142 ;
  assign y7777 = ~n27149 ;
  assign y7778 = ~n27151 ;
  assign y7779 = ~1'b0 ;
  assign y7780 = ~n27157 ;
  assign y7781 = ~n27164 ;
  assign y7782 = n27167 ;
  assign y7783 = n27172 ;
  assign y7784 = n27174 ;
  assign y7785 = ~n27175 ;
  assign y7786 = n27177 ;
  assign y7787 = ~n27179 ;
  assign y7788 = n27184 ;
  assign y7789 = ~n27186 ;
  assign y7790 = ~n27189 ;
  assign y7791 = ~n27190 ;
  assign y7792 = n27198 ;
  assign y7793 = ~1'b0 ;
  assign y7794 = n27215 ;
  assign y7795 = n27216 ;
  assign y7796 = n27217 ;
  assign y7797 = ~1'b0 ;
  assign y7798 = ~n27221 ;
  assign y7799 = ~1'b0 ;
  assign y7800 = n26484 ;
  assign y7801 = ~n27228 ;
  assign y7802 = n27230 ;
  assign y7803 = n27235 ;
  assign y7804 = ~n27236 ;
  assign y7805 = n27241 ;
  assign y7806 = ~n27242 ;
  assign y7807 = ~1'b0 ;
  assign y7808 = ~n27251 ;
  assign y7809 = n27252 ;
  assign y7810 = n27253 ;
  assign y7811 = ~n27260 ;
  assign y7812 = n27261 ;
  assign y7813 = ~n27262 ;
  assign y7814 = ~1'b0 ;
  assign y7815 = ~n27264 ;
  assign y7816 = n27268 ;
  assign y7817 = ~n25737 ;
  assign y7818 = n27271 ;
  assign y7819 = n27272 ;
  assign y7820 = ~n27274 ;
  assign y7821 = ~n27279 ;
  assign y7822 = ~n27283 ;
  assign y7823 = ~n27284 ;
  assign y7824 = n27286 ;
  assign y7825 = n27290 ;
  assign y7826 = ~n27296 ;
  assign y7827 = ~n27298 ;
  assign y7828 = ~n27300 ;
  assign y7829 = ~1'b0 ;
  assign y7830 = ~1'b0 ;
  assign y7831 = ~n27301 ;
  assign y7832 = ~n27308 ;
  assign y7833 = ~n27311 ;
  assign y7834 = ~1'b0 ;
  assign y7835 = ~n27313 ;
  assign y7836 = ~n27318 ;
  assign y7837 = ~n27320 ;
  assign y7838 = n27325 ;
  assign y7839 = ~n27326 ;
  assign y7840 = n27329 ;
  assign y7841 = n27332 ;
  assign y7842 = ~n27342 ;
  assign y7843 = ~n27347 ;
  assign y7844 = ~n27349 ;
  assign y7845 = n27358 ;
  assign y7846 = ~n27362 ;
  assign y7847 = n27367 ;
  assign y7848 = n27368 ;
  assign y7849 = ~n27369 ;
  assign y7850 = n27373 ;
  assign y7851 = ~1'b0 ;
  assign y7852 = ~n27377 ;
  assign y7853 = n27382 ;
  assign y7854 = ~n27385 ;
  assign y7855 = ~n27387 ;
  assign y7856 = ~1'b0 ;
  assign y7857 = ~n27388 ;
  assign y7858 = n27391 ;
  assign y7859 = n27394 ;
  assign y7860 = ~1'b0 ;
  assign y7861 = ~n27396 ;
  assign y7862 = ~1'b0 ;
  assign y7863 = ~n27397 ;
  assign y7864 = ~1'b0 ;
  assign y7865 = ~n27402 ;
  assign y7866 = n27403 ;
  assign y7867 = ~n27407 ;
  assign y7868 = ~1'b0 ;
  assign y7869 = n27411 ;
  assign y7870 = n27412 ;
  assign y7871 = ~n27413 ;
  assign y7872 = n27414 ;
  assign y7873 = ~n27416 ;
  assign y7874 = n27422 ;
  assign y7875 = n27428 ;
  assign y7876 = n27429 ;
  assign y7877 = ~1'b0 ;
  assign y7878 = n27432 ;
  assign y7879 = n27433 ;
  assign y7880 = n25337 ;
  assign y7881 = n27435 ;
  assign y7882 = n27445 ;
  assign y7883 = ~1'b0 ;
  assign y7884 = ~1'b0 ;
  assign y7885 = ~n27446 ;
  assign y7886 = n27447 ;
  assign y7887 = n27450 ;
  assign y7888 = ~n7544 ;
  assign y7889 = ~n27451 ;
  assign y7890 = ~n27455 ;
  assign y7891 = ~n27460 ;
  assign y7892 = ~n27463 ;
  assign y7893 = ~n27467 ;
  assign y7894 = n27470 ;
  assign y7895 = ~1'b0 ;
  assign y7896 = n27479 ;
  assign y7897 = ~n27484 ;
  assign y7898 = n27490 ;
  assign y7899 = ~n27492 ;
  assign y7900 = n27493 ;
  assign y7901 = ~1'b0 ;
  assign y7902 = ~n27507 ;
  assign y7903 = ~1'b0 ;
  assign y7904 = ~n25160 ;
  assign y7905 = ~n27509 ;
  assign y7906 = ~1'b0 ;
  assign y7907 = n27511 ;
  assign y7908 = n27518 ;
  assign y7909 = n27524 ;
  assign y7910 = n27526 ;
  assign y7911 = n27527 ;
  assign y7912 = n27531 ;
  assign y7913 = ~n27532 ;
  assign y7914 = ~n27533 ;
  assign y7915 = ~1'b0 ;
  assign y7916 = ~1'b0 ;
  assign y7917 = n27534 ;
  assign y7918 = ~n27535 ;
  assign y7919 = ~n27538 ;
  assign y7920 = n27541 ;
  assign y7921 = ~n27554 ;
  assign y7922 = ~1'b0 ;
  assign y7923 = n27557 ;
  assign y7924 = ~1'b0 ;
  assign y7925 = ~1'b0 ;
  assign y7926 = ~n27558 ;
  assign y7927 = ~n22801 ;
  assign y7928 = n27560 ;
  assign y7929 = ~n27563 ;
  assign y7930 = n27565 ;
  assign y7931 = ~n27568 ;
  assign y7932 = n27570 ;
  assign y7933 = n27576 ;
  assign y7934 = n27581 ;
  assign y7935 = ~n27582 ;
  assign y7936 = ~1'b0 ;
  assign y7937 = n27585 ;
  assign y7938 = ~1'b0 ;
  assign y7939 = n27586 ;
  assign y7940 = n27589 ;
  assign y7941 = n27591 ;
  assign y7942 = ~n27593 ;
  assign y7943 = ~n27595 ;
  assign y7944 = n27596 ;
  assign y7945 = ~n27600 ;
  assign y7946 = n27609 ;
  assign y7947 = ~1'b0 ;
  assign y7948 = ~n27612 ;
  assign y7949 = n27613 ;
  assign y7950 = n27616 ;
  assign y7951 = n27619 ;
  assign y7952 = ~n27625 ;
  assign y7953 = n27626 ;
  assign y7954 = ~n27633 ;
  assign y7955 = n27638 ;
  assign y7956 = ~n27641 ;
  assign y7957 = ~n27646 ;
  assign y7958 = n27650 ;
  assign y7959 = n27651 ;
  assign y7960 = n27656 ;
  assign y7961 = n27657 ;
  assign y7962 = ~1'b0 ;
  assign y7963 = ~n27662 ;
  assign y7964 = n27665 ;
  assign y7965 = ~1'b0 ;
  assign y7966 = ~1'b0 ;
  assign y7967 = ~n27666 ;
  assign y7968 = ~n27669 ;
  assign y7969 = ~n27672 ;
  assign y7970 = ~n27674 ;
  assign y7971 = ~1'b0 ;
  assign y7972 = ~1'b0 ;
  assign y7973 = ~n27678 ;
  assign y7974 = n27684 ;
  assign y7975 = ~n27691 ;
  assign y7976 = ~n27695 ;
  assign y7977 = ~n27702 ;
  assign y7978 = n27703 ;
  assign y7979 = n27707 ;
  assign y7980 = n27708 ;
  assign y7981 = ~n27710 ;
  assign y7982 = ~n27711 ;
  assign y7983 = ~n27712 ;
  assign y7984 = ~1'b0 ;
  assign y7985 = ~1'b0 ;
  assign y7986 = n27714 ;
  assign y7987 = n27717 ;
  assign y7988 = ~n27722 ;
  assign y7989 = ~n27724 ;
  assign y7990 = n27729 ;
  assign y7991 = ~n27735 ;
  assign y7992 = ~1'b0 ;
  assign y7993 = n27748 ;
  assign y7994 = ~n27753 ;
  assign y7995 = ~n27756 ;
  assign y7996 = ~n27758 ;
  assign y7997 = ~n27761 ;
  assign y7998 = ~n27764 ;
  assign y7999 = ~n27767 ;
  assign y8000 = n27773 ;
  assign y8001 = ~1'b0 ;
  assign y8002 = n27777 ;
  assign y8003 = ~n27782 ;
  assign y8004 = n27785 ;
  assign y8005 = ~1'b0 ;
  assign y8006 = ~n27787 ;
  assign y8007 = ~n27791 ;
  assign y8008 = n27799 ;
  assign y8009 = n27800 ;
  assign y8010 = ~n27804 ;
  assign y8011 = ~n27811 ;
  assign y8012 = ~n27812 ;
  assign y8013 = ~n27818 ;
  assign y8014 = ~1'b0 ;
  assign y8015 = n27820 ;
  assign y8016 = ~n27823 ;
  assign y8017 = ~1'b0 ;
  assign y8018 = n27824 ;
  assign y8019 = ~n27829 ;
  assign y8020 = n27832 ;
  assign y8021 = ~n27841 ;
  assign y8022 = ~n27846 ;
  assign y8023 = n27847 ;
  assign y8024 = n27848 ;
  assign y8025 = ~n27852 ;
  assign y8026 = ~1'b0 ;
  assign y8027 = n27855 ;
  assign y8028 = ~n27856 ;
  assign y8029 = n27858 ;
  assign y8030 = n27861 ;
  assign y8031 = n27864 ;
  assign y8032 = ~n27868 ;
  assign y8033 = ~n15314 ;
  assign y8034 = ~n27873 ;
  assign y8035 = ~n27879 ;
  assign y8036 = n27882 ;
  assign y8037 = ~n27898 ;
  assign y8038 = n27903 ;
  assign y8039 = ~n27905 ;
  assign y8040 = n27906 ;
  assign y8041 = ~n27908 ;
  assign y8042 = n27909 ;
  assign y8043 = ~n27910 ;
  assign y8044 = ~n27914 ;
  assign y8045 = n27916 ;
  assign y8046 = ~n27920 ;
  assign y8047 = ~1'b0 ;
  assign y8048 = n27924 ;
  assign y8049 = ~n27925 ;
  assign y8050 = n27928 ;
  assign y8051 = ~1'b0 ;
  assign y8052 = n27930 ;
  assign y8053 = n27931 ;
  assign y8054 = ~n27936 ;
  assign y8055 = ~n27948 ;
  assign y8056 = ~1'b0 ;
  assign y8057 = ~n27952 ;
  assign y8058 = ~1'b0 ;
  assign y8059 = n27958 ;
  assign y8060 = ~n27959 ;
  assign y8061 = ~1'b0 ;
  assign y8062 = ~1'b0 ;
  assign y8063 = n27961 ;
  assign y8064 = n27967 ;
  assign y8065 = ~n27971 ;
  assign y8066 = ~n27978 ;
  assign y8067 = ~1'b0 ;
  assign y8068 = n27979 ;
  assign y8069 = ~1'b0 ;
  assign y8070 = ~n27981 ;
  assign y8071 = n27984 ;
  assign y8072 = ~n27986 ;
  assign y8073 = ~n27997 ;
  assign y8074 = ~1'b0 ;
  assign y8075 = n28003 ;
  assign y8076 = ~n28006 ;
  assign y8077 = n28009 ;
  assign y8078 = n28012 ;
  assign y8079 = ~n28014 ;
  assign y8080 = n28017 ;
  assign y8081 = n28018 ;
  assign y8082 = ~1'b0 ;
  assign y8083 = ~1'b0 ;
  assign y8084 = ~1'b0 ;
  assign y8085 = ~n28025 ;
  assign y8086 = n28028 ;
  assign y8087 = ~n28030 ;
  assign y8088 = ~n28034 ;
  assign y8089 = n28037 ;
  assign y8090 = ~n28039 ;
  assign y8091 = n28041 ;
  assign y8092 = ~1'b0 ;
  assign y8093 = ~n28043 ;
  assign y8094 = ~n5937 ;
  assign y8095 = n28045 ;
  assign y8096 = ~n28048 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = ~1'b0 ;
  assign y8099 = ~1'b0 ;
  assign y8100 = ~1'b0 ;
  assign y8101 = ~n28049 ;
  assign y8102 = n28052 ;
  assign y8103 = ~n28053 ;
  assign y8104 = ~1'b0 ;
  assign y8105 = ~n28054 ;
  assign y8106 = ~n28058 ;
  assign y8107 = n28064 ;
  assign y8108 = ~n28069 ;
  assign y8109 = ~n28070 ;
  assign y8110 = n28071 ;
  assign y8111 = n28072 ;
  assign y8112 = ~n28073 ;
  assign y8113 = ~1'b0 ;
  assign y8114 = n28075 ;
  assign y8115 = ~1'b0 ;
  assign y8116 = n28079 ;
  assign y8117 = ~n28083 ;
  assign y8118 = n28090 ;
  assign y8119 = n28091 ;
  assign y8120 = ~1'b0 ;
  assign y8121 = n28092 ;
  assign y8122 = n28100 ;
  assign y8123 = ~n28107 ;
  assign y8124 = ~1'b0 ;
  assign y8125 = n28109 ;
  assign y8126 = ~1'b0 ;
  assign y8127 = n28112 ;
  assign y8128 = n28113 ;
  assign y8129 = ~n28114 ;
  assign y8130 = n28116 ;
  assign y8131 = ~1'b0 ;
  assign y8132 = n28118 ;
  assign y8133 = n28119 ;
  assign y8134 = ~n28120 ;
  assign y8135 = ~n28122 ;
  assign y8136 = ~1'b0 ;
  assign y8137 = ~1'b0 ;
  assign y8138 = n28124 ;
  assign y8139 = ~n28127 ;
  assign y8140 = ~n28131 ;
  assign y8141 = ~n3254 ;
  assign y8142 = ~n28133 ;
  assign y8143 = ~1'b0 ;
  assign y8144 = ~1'b0 ;
  assign y8145 = ~n28138 ;
  assign y8146 = n28142 ;
  assign y8147 = n28143 ;
  assign y8148 = n28146 ;
  assign y8149 = n28147 ;
  assign y8150 = n28156 ;
  assign y8151 = ~1'b0 ;
  assign y8152 = ~1'b0 ;
  assign y8153 = ~n21014 ;
  assign y8154 = ~n28158 ;
  assign y8155 = ~n28159 ;
  assign y8156 = ~n28163 ;
  assign y8157 = n28165 ;
  assign y8158 = ~1'b0 ;
  assign y8159 = n28166 ;
  assign y8160 = n28168 ;
  assign y8161 = n28169 ;
  assign y8162 = n28171 ;
  assign y8163 = ~n7271 ;
  assign y8164 = ~1'b0 ;
  assign y8165 = ~n28183 ;
  assign y8166 = n28187 ;
  assign y8167 = n28194 ;
  assign y8168 = n28195 ;
  assign y8169 = ~1'b0 ;
  assign y8170 = ~1'b0 ;
  assign y8171 = ~1'b0 ;
  assign y8172 = ~n28197 ;
  assign y8173 = n28200 ;
  assign y8174 = ~n28204 ;
  assign y8175 = ~n28206 ;
  assign y8176 = ~n28208 ;
  assign y8177 = ~n28209 ;
  assign y8178 = n28210 ;
  assign y8179 = ~n28215 ;
  assign y8180 = ~n28217 ;
  assign y8181 = n28218 ;
  assign y8182 = ~1'b0 ;
  assign y8183 = ~n28221 ;
  assign y8184 = ~n28222 ;
  assign y8185 = n28223 ;
  assign y8186 = n28226 ;
  assign y8187 = n28227 ;
  assign y8188 = ~n28229 ;
  assign y8189 = n28235 ;
  assign y8190 = n28236 ;
  assign y8191 = ~n28240 ;
  assign y8192 = ~1'b0 ;
  assign y8193 = ~n28243 ;
  assign y8194 = n28244 ;
  assign y8195 = ~1'b0 ;
  assign y8196 = ~n28246 ;
  assign y8197 = ~n28248 ;
  assign y8198 = ~1'b0 ;
  assign y8199 = n28251 ;
  assign y8200 = ~n28257 ;
  assign y8201 = ~n28263 ;
  assign y8202 = ~n28265 ;
  assign y8203 = ~n28269 ;
  assign y8204 = ~1'b0 ;
  assign y8205 = n28270 ;
  assign y8206 = ~n28274 ;
  assign y8207 = n28276 ;
  assign y8208 = ~n28277 ;
  assign y8209 = n28279 ;
  assign y8210 = ~n28287 ;
  assign y8211 = ~n28297 ;
  assign y8212 = n28298 ;
  assign y8213 = ~n28300 ;
  assign y8214 = ~1'b0 ;
  assign y8215 = ~n28306 ;
  assign y8216 = n28308 ;
  assign y8217 = ~n28309 ;
  assign y8218 = ~n28312 ;
  assign y8219 = n28314 ;
  assign y8220 = n28316 ;
  assign y8221 = n28317 ;
  assign y8222 = ~n28319 ;
  assign y8223 = ~n28325 ;
  assign y8224 = n28326 ;
  assign y8225 = 1'b0 ;
  assign y8226 = n28332 ;
  assign y8227 = ~1'b0 ;
  assign y8228 = ~n28335 ;
  assign y8229 = n28338 ;
  assign y8230 = ~n28339 ;
  assign y8231 = ~n28347 ;
  assign y8232 = n28354 ;
  assign y8233 = ~n28361 ;
  assign y8234 = ~1'b0 ;
  assign y8235 = n28363 ;
  assign y8236 = ~1'b0 ;
  assign y8237 = n28376 ;
  assign y8238 = n28379 ;
  assign y8239 = n12488 ;
  assign y8240 = ~1'b0 ;
  assign y8241 = ~n28380 ;
  assign y8242 = n28381 ;
  assign y8243 = n28386 ;
  assign y8244 = n28392 ;
  assign y8245 = n28393 ;
  assign y8246 = n28394 ;
  assign y8247 = ~n28400 ;
  assign y8248 = ~n1989 ;
  assign y8249 = n28405 ;
  assign y8250 = ~1'b0 ;
  assign y8251 = ~n28407 ;
  assign y8252 = n28412 ;
  assign y8253 = ~n28419 ;
  assign y8254 = n28420 ;
  assign y8255 = ~n28421 ;
  assign y8256 = n28425 ;
  assign y8257 = n28432 ;
  assign y8258 = ~n28433 ;
  assign y8259 = ~n28435 ;
  assign y8260 = n28436 ;
  assign y8261 = ~n28443 ;
  assign y8262 = ~n28448 ;
  assign y8263 = n28449 ;
  assign y8264 = ~1'b0 ;
  assign y8265 = ~n28454 ;
  assign y8266 = n28458 ;
  assign y8267 = ~n28467 ;
  assign y8268 = n28468 ;
  assign y8269 = ~n28471 ;
  assign y8270 = ~n28474 ;
  assign y8271 = n28476 ;
  assign y8272 = n28482 ;
  assign y8273 = ~n28485 ;
  assign y8274 = n28486 ;
  assign y8275 = n28491 ;
  assign y8276 = ~n28497 ;
  assign y8277 = ~n28505 ;
  assign y8278 = n28508 ;
  assign y8279 = n28511 ;
  assign y8280 = ~n28515 ;
  assign y8281 = n28519 ;
  assign y8282 = ~1'b0 ;
  assign y8283 = ~n28520 ;
  assign y8284 = ~n28524 ;
  assign y8285 = n28525 ;
  assign y8286 = n28526 ;
  assign y8287 = n28528 ;
  assign y8288 = ~n28529 ;
  assign y8289 = ~n28530 ;
  assign y8290 = n28533 ;
  assign y8291 = ~n28538 ;
  assign y8292 = ~n28539 ;
  assign y8293 = n28540 ;
  assign y8294 = n28542 ;
  assign y8295 = ~n28544 ;
  assign y8296 = ~n28546 ;
  assign y8297 = n28548 ;
  assign y8298 = n28550 ;
  assign y8299 = n28554 ;
  assign y8300 = n28560 ;
  assign y8301 = n28565 ;
  assign y8302 = ~1'b0 ;
  assign y8303 = n28566 ;
  assign y8304 = n28571 ;
  assign y8305 = ~1'b0 ;
  assign y8306 = n28574 ;
  assign y8307 = ~n28577 ;
  assign y8308 = ~n5392 ;
  assign y8309 = ~n28585 ;
  assign y8310 = n28601 ;
  assign y8311 = ~1'b0 ;
  assign y8312 = ~n28603 ;
  assign y8313 = n28604 ;
  assign y8314 = ~n28613 ;
  assign y8315 = ~1'b0 ;
  assign y8316 = ~1'b0 ;
  assign y8317 = ~n28615 ;
  assign y8318 = ~n28619 ;
  assign y8319 = ~n28622 ;
  assign y8320 = n28624 ;
  assign y8321 = ~1'b0 ;
  assign y8322 = n28626 ;
  assign y8323 = ~n28630 ;
  assign y8324 = ~1'b0 ;
  assign y8325 = n28636 ;
  assign y8326 = n28638 ;
  assign y8327 = ~n28639 ;
  assign y8328 = ~n28641 ;
  assign y8329 = n28643 ;
  assign y8330 = ~1'b0 ;
  assign y8331 = n28647 ;
  assign y8332 = ~1'b0 ;
  assign y8333 = ~n28649 ;
  assign y8334 = ~n28652 ;
  assign y8335 = ~n28654 ;
  assign y8336 = n28656 ;
  assign y8337 = n28662 ;
  assign y8338 = ~n28670 ;
  assign y8339 = n28671 ;
  assign y8340 = n28672 ;
  assign y8341 = n28675 ;
  assign y8342 = ~n28680 ;
  assign y8343 = n28688 ;
  assign y8344 = ~n28697 ;
  assign y8345 = n28698 ;
  assign y8346 = ~n28699 ;
  assign y8347 = ~1'b0 ;
  assign y8348 = ~n28700 ;
  assign y8349 = n28701 ;
  assign y8350 = n28703 ;
  assign y8351 = ~n28715 ;
  assign y8352 = ~1'b0 ;
  assign y8353 = n28716 ;
  assign y8354 = n28723 ;
  assign y8355 = n28725 ;
  assign y8356 = n28726 ;
  assign y8357 = ~1'b0 ;
  assign y8358 = ~n28727 ;
  assign y8359 = ~n28734 ;
  assign y8360 = n28736 ;
  assign y8361 = n28747 ;
  assign y8362 = ~1'b0 ;
  assign y8363 = ~1'b0 ;
  assign y8364 = n28751 ;
  assign y8365 = ~n28754 ;
  assign y8366 = n28756 ;
  assign y8367 = ~n28757 ;
  assign y8368 = n28762 ;
  assign y8369 = ~n28769 ;
  assign y8370 = ~n28772 ;
  assign y8371 = ~n28776 ;
  assign y8372 = n28779 ;
  assign y8373 = n28781 ;
  assign y8374 = ~1'b0 ;
  assign y8375 = ~n28783 ;
  assign y8376 = ~1'b0 ;
  assign y8377 = n28786 ;
  assign y8378 = n28789 ;
  assign y8379 = n28796 ;
  assign y8380 = ~1'b0 ;
  assign y8381 = ~n28799 ;
  assign y8382 = n28805 ;
  assign y8383 = n28806 ;
  assign y8384 = ~n28807 ;
  assign y8385 = ~n28808 ;
  assign y8386 = n28809 ;
  assign y8387 = n28810 ;
  assign y8388 = ~n28818 ;
  assign y8389 = n28820 ;
  assign y8390 = ~n28822 ;
  assign y8391 = ~n28829 ;
  assign y8392 = n28835 ;
  assign y8393 = ~1'b0 ;
  assign y8394 = n28837 ;
  assign y8395 = ~n28841 ;
  assign y8396 = ~1'b0 ;
  assign y8397 = n28847 ;
  assign y8398 = ~1'b0 ;
  assign y8399 = n28849 ;
  assign y8400 = n28850 ;
  assign y8401 = ~n28852 ;
  assign y8402 = n28858 ;
  assign y8403 = ~n28861 ;
  assign y8404 = n28862 ;
  assign y8405 = n28868 ;
  assign y8406 = n28871 ;
  assign y8407 = ~n28877 ;
  assign y8408 = n28878 ;
  assign y8409 = ~n28882 ;
  assign y8410 = n28884 ;
  assign y8411 = ~n28888 ;
  assign y8412 = ~1'b0 ;
  assign y8413 = n28889 ;
  assign y8414 = ~n28891 ;
  assign y8415 = ~1'b0 ;
  assign y8416 = ~n28895 ;
  assign y8417 = n28898 ;
  assign y8418 = n28905 ;
  assign y8419 = ~1'b0 ;
  assign y8420 = ~1'b0 ;
  assign y8421 = ~1'b0 ;
  assign y8422 = n28906 ;
  assign y8423 = n28909 ;
  assign y8424 = n28910 ;
  assign y8425 = n28913 ;
  assign y8426 = ~1'b0 ;
  assign y8427 = ~1'b0 ;
  assign y8428 = ~n28914 ;
  assign y8429 = ~1'b0 ;
  assign y8430 = ~n28918 ;
  assign y8431 = n28923 ;
  assign y8432 = ~n28924 ;
  assign y8433 = n28925 ;
  assign y8434 = ~1'b0 ;
  assign y8435 = n28928 ;
  assign y8436 = n28929 ;
  assign y8437 = ~n28933 ;
  assign y8438 = ~1'b0 ;
  assign y8439 = ~n28938 ;
  assign y8440 = n28939 ;
  assign y8441 = n28945 ;
  assign y8442 = ~n28947 ;
  assign y8443 = ~n28949 ;
  assign y8444 = ~1'b0 ;
  assign y8445 = ~1'b0 ;
  assign y8446 = ~1'b0 ;
  assign y8447 = ~n28951 ;
  assign y8448 = n28955 ;
  assign y8449 = ~n28962 ;
  assign y8450 = ~n28969 ;
  assign y8451 = ~n28972 ;
  assign y8452 = ~n28973 ;
  assign y8453 = ~1'b0 ;
  assign y8454 = n28976 ;
  assign y8455 = ~n28977 ;
  assign y8456 = ~n28980 ;
  assign y8457 = ~1'b0 ;
  assign y8458 = ~1'b0 ;
  assign y8459 = ~n28981 ;
  assign y8460 = n28982 ;
  assign y8461 = n28995 ;
  assign y8462 = n4483 ;
  assign y8463 = ~1'b0 ;
  assign y8464 = ~1'b0 ;
  assign y8465 = ~n28998 ;
  assign y8466 = ~n28999 ;
  assign y8467 = ~n29000 ;
  assign y8468 = ~1'b0 ;
  assign y8469 = n29006 ;
  assign y8470 = ~1'b0 ;
  assign y8471 = n29008 ;
  assign y8472 = n29010 ;
  assign y8473 = ~n29012 ;
  assign y8474 = n29013 ;
  assign y8475 = ~n29016 ;
  assign y8476 = ~1'b0 ;
  assign y8477 = n29018 ;
  assign y8478 = n29025 ;
  assign y8479 = ~n29028 ;
  assign y8480 = n29029 ;
  assign y8481 = ~1'b0 ;
  assign y8482 = n29030 ;
  assign y8483 = ~n29032 ;
  assign y8484 = n29033 ;
  assign y8485 = ~1'b0 ;
  assign y8486 = ~n29041 ;
  assign y8487 = n29044 ;
  assign y8488 = ~n29046 ;
  assign y8489 = n29047 ;
  assign y8490 = ~n29051 ;
  assign y8491 = ~1'b0 ;
  assign y8492 = ~1'b0 ;
  assign y8493 = n29057 ;
  assign y8494 = n29060 ;
  assign y8495 = ~n29064 ;
  assign y8496 = n29065 ;
  assign y8497 = n29070 ;
  assign y8498 = ~n29075 ;
  assign y8499 = ~n29078 ;
  assign y8500 = n29083 ;
  assign y8501 = n29097 ;
  assign y8502 = ~n29102 ;
  assign y8503 = n29105 ;
  assign y8504 = n29116 ;
  assign y8505 = n29117 ;
  assign y8506 = ~n29120 ;
  assign y8507 = n28228 ;
  assign y8508 = n29121 ;
  assign y8509 = ~n29123 ;
  assign y8510 = n29124 ;
  assign y8511 = ~n29129 ;
  assign y8512 = ~n29131 ;
  assign y8513 = n29132 ;
  assign y8514 = ~n29134 ;
  assign y8515 = ~n29137 ;
  assign y8516 = ~n29139 ;
  assign y8517 = n29140 ;
  assign y8518 = ~n29141 ;
  assign y8519 = n29142 ;
  assign y8520 = n29150 ;
  assign y8521 = ~n29151 ;
  assign y8522 = ~n29153 ;
  assign y8523 = n29158 ;
  assign y8524 = n29161 ;
  assign y8525 = n29162 ;
  assign y8526 = ~n29165 ;
  assign y8527 = ~1'b0 ;
  assign y8528 = ~n29167 ;
  assign y8529 = ~n29174 ;
  assign y8530 = ~n29179 ;
  assign y8531 = ~n29184 ;
  assign y8532 = ~n29187 ;
  assign y8533 = n29193 ;
  assign y8534 = ~n29194 ;
  assign y8535 = ~n29202 ;
  assign y8536 = n29206 ;
  assign y8537 = n29207 ;
  assign y8538 = n29209 ;
  assign y8539 = n29211 ;
  assign y8540 = ~n29219 ;
  assign y8541 = n29222 ;
  assign y8542 = n29223 ;
  assign y8543 = ~n29225 ;
  assign y8544 = n29229 ;
  assign y8545 = ~n29235 ;
  assign y8546 = ~n13257 ;
  assign y8547 = ~n29237 ;
  assign y8548 = ~n29242 ;
  assign y8549 = ~n29246 ;
  assign y8550 = n29248 ;
  assign y8551 = ~n29250 ;
  assign y8552 = n29253 ;
  assign y8553 = ~n29255 ;
  assign y8554 = 1'b0 ;
  assign y8555 = n29258 ;
  assign y8556 = ~n29265 ;
  assign y8557 = ~n29271 ;
  assign y8558 = ~n29277 ;
  assign y8559 = ~n29279 ;
  assign y8560 = ~1'b0 ;
  assign y8561 = ~1'b0 ;
  assign y8562 = ~n29282 ;
  assign y8563 = n29286 ;
  assign y8564 = ~n29291 ;
  assign y8565 = ~1'b0 ;
  assign y8566 = ~n29293 ;
  assign y8567 = n29294 ;
  assign y8568 = n29295 ;
  assign y8569 = ~n29296 ;
  assign y8570 = ~n29297 ;
  assign y8571 = ~1'b0 ;
  assign y8572 = n29299 ;
  assign y8573 = n29303 ;
  assign y8574 = ~n29312 ;
  assign y8575 = ~n29315 ;
  assign y8576 = ~1'b0 ;
  assign y8577 = ~1'b0 ;
  assign y8578 = n29318 ;
  assign y8579 = ~1'b0 ;
  assign y8580 = n29325 ;
  assign y8581 = ~n29326 ;
  assign y8582 = ~n29328 ;
  assign y8583 = ~n29330 ;
  assign y8584 = ~n29338 ;
  assign y8585 = ~n29339 ;
  assign y8586 = ~n29343 ;
  assign y8587 = ~n29347 ;
  assign y8588 = ~n29352 ;
  assign y8589 = n29357 ;
  assign y8590 = 1'b0 ;
  assign y8591 = n29358 ;
  assign y8592 = n29360 ;
  assign y8593 = ~n29367 ;
  assign y8594 = ~n29370 ;
  assign y8595 = n29372 ;
  assign y8596 = ~1'b0 ;
  assign y8597 = ~n29375 ;
  assign y8598 = n29377 ;
  assign y8599 = n29383 ;
  assign y8600 = n29384 ;
  assign y8601 = ~n29386 ;
  assign y8602 = ~1'b0 ;
  assign y8603 = ~n29387 ;
  assign y8604 = n29388 ;
  assign y8605 = n29395 ;
  assign y8606 = ~n29397 ;
  assign y8607 = n29400 ;
  assign y8608 = ~n29401 ;
  assign y8609 = ~n29402 ;
  assign y8610 = ~n29403 ;
  assign y8611 = ~n29404 ;
  assign y8612 = ~n29405 ;
  assign y8613 = n29408 ;
  assign y8614 = ~n29412 ;
  assign y8615 = ~n29413 ;
  assign y8616 = n29414 ;
  assign y8617 = n29415 ;
  assign y8618 = ~n29418 ;
  assign y8619 = n29425 ;
  assign y8620 = ~n24873 ;
  assign y8621 = ~1'b0 ;
  assign y8622 = ~1'b0 ;
  assign y8623 = ~n29426 ;
  assign y8624 = ~n5978 ;
  assign y8625 = ~n29428 ;
  assign y8626 = ~1'b0 ;
  assign y8627 = n29436 ;
  assign y8628 = n29437 ;
  assign y8629 = ~n29443 ;
  assign y8630 = ~1'b0 ;
  assign y8631 = n29445 ;
  assign y8632 = ~1'b0 ;
  assign y8633 = n29448 ;
  assign y8634 = n29451 ;
  assign y8635 = n29452 ;
  assign y8636 = ~n29453 ;
  assign y8637 = ~n29456 ;
  assign y8638 = ~n29459 ;
  assign y8639 = ~n29461 ;
  assign y8640 = n29462 ;
  assign y8641 = n29464 ;
  assign y8642 = ~n29465 ;
  assign y8643 = ~n29467 ;
  assign y8644 = n29470 ;
  assign y8645 = n29476 ;
  assign y8646 = n29481 ;
  assign y8647 = ~n29482 ;
  assign y8648 = ~1'b0 ;
  assign y8649 = ~n29484 ;
  assign y8650 = ~n29490 ;
  assign y8651 = n29491 ;
  assign y8652 = n29496 ;
  assign y8653 = n29497 ;
  assign y8654 = ~n29498 ;
  assign y8655 = ~n29501 ;
  assign y8656 = ~1'b0 ;
  assign y8657 = ~n29504 ;
  assign y8658 = n29508 ;
  assign y8659 = n29512 ;
  assign y8660 = ~n29513 ;
  assign y8661 = ~1'b0 ;
  assign y8662 = n29517 ;
  assign y8663 = ~1'b0 ;
  assign y8664 = ~n29525 ;
  assign y8665 = ~n29531 ;
  assign y8666 = n29532 ;
  assign y8667 = ~n29534 ;
  assign y8668 = 1'b0 ;
  assign y8669 = n29535 ;
  assign y8670 = ~n29537 ;
  assign y8671 = ~n29538 ;
  assign y8672 = n29540 ;
  assign y8673 = n29543 ;
  assign y8674 = n29551 ;
  assign y8675 = n29556 ;
  assign y8676 = n29560 ;
  assign y8677 = n29565 ;
  assign y8678 = ~n29567 ;
  assign y8679 = ~n29568 ;
  assign y8680 = ~n29573 ;
  assign y8681 = ~n29577 ;
  assign y8682 = ~n29579 ;
  assign y8683 = n29583 ;
  assign y8684 = ~n29585 ;
  assign y8685 = ~n29588 ;
  assign y8686 = n29590 ;
  assign y8687 = ~1'b0 ;
  assign y8688 = ~n29596 ;
  assign y8689 = n29597 ;
  assign y8690 = n29601 ;
  assign y8691 = ~n29603 ;
  assign y8692 = n29606 ;
  assign y8693 = n29609 ;
  assign y8694 = n29615 ;
  assign y8695 = n29619 ;
  assign y8696 = n29622 ;
  assign y8697 = ~n29624 ;
  assign y8698 = n29626 ;
  assign y8699 = ~1'b0 ;
  assign y8700 = n19852 ;
  assign y8701 = n29631 ;
  assign y8702 = n29633 ;
  assign y8703 = ~n29637 ;
  assign y8704 = ~n565 ;
  assign y8705 = n29641 ;
  assign y8706 = n29645 ;
  assign y8707 = n29658 ;
  assign y8708 = ~n29660 ;
  assign y8709 = n29661 ;
  assign y8710 = n29665 ;
  assign y8711 = n29667 ;
  assign y8712 = ~n15779 ;
  assign y8713 = ~1'b0 ;
  assign y8714 = ~n29683 ;
  assign y8715 = n29684 ;
  assign y8716 = n29685 ;
  assign y8717 = ~n29689 ;
  assign y8718 = n29693 ;
  assign y8719 = n29695 ;
  assign y8720 = ~n29697 ;
  assign y8721 = ~n29702 ;
  assign y8722 = n29705 ;
  assign y8723 = ~n29706 ;
  assign y8724 = ~n29713 ;
  assign y8725 = n29716 ;
  assign y8726 = ~n29717 ;
  assign y8727 = ~n29721 ;
  assign y8728 = n29723 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = n29724 ;
  assign y8731 = n29726 ;
  assign y8732 = n29730 ;
  assign y8733 = n29731 ;
  assign y8734 = n29732 ;
  assign y8735 = n29734 ;
  assign y8736 = ~n29736 ;
  assign y8737 = ~n29738 ;
  assign y8738 = n29748 ;
  assign y8739 = ~n29749 ;
  assign y8740 = ~n29753 ;
  assign y8741 = n29754 ;
  assign y8742 = ~n29756 ;
  assign y8743 = ~1'b0 ;
  assign y8744 = ~n29760 ;
  assign y8745 = ~n29766 ;
  assign y8746 = n29768 ;
  assign y8747 = ~n29773 ;
  assign y8748 = n29778 ;
  assign y8749 = ~n29779 ;
  assign y8750 = n29780 ;
  assign y8751 = ~n29785 ;
  assign y8752 = ~1'b0 ;
  assign y8753 = ~1'b0 ;
  assign y8754 = n17405 ;
  assign y8755 = ~n29788 ;
  assign y8756 = n29789 ;
  assign y8757 = ~n29793 ;
  assign y8758 = ~n29795 ;
  assign y8759 = n29798 ;
  assign y8760 = n29801 ;
  assign y8761 = ~n29806 ;
  assign y8762 = ~n29810 ;
  assign y8763 = n29818 ;
  assign y8764 = ~n29824 ;
  assign y8765 = ~1'b0 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = n29828 ;
  assign y8768 = n29831 ;
  assign y8769 = ~n29832 ;
  assign y8770 = ~n29836 ;
  assign y8771 = ~n29837 ;
  assign y8772 = n29840 ;
  assign y8773 = n29849 ;
  assign y8774 = ~n29851 ;
  assign y8775 = n29853 ;
  assign y8776 = n29857 ;
  assign y8777 = ~n29860 ;
  assign y8778 = ~n29867 ;
  assign y8779 = n29868 ;
  assign y8780 = ~n29875 ;
  assign y8781 = ~n29882 ;
  assign y8782 = ~1'b0 ;
  assign y8783 = n29887 ;
  assign y8784 = ~1'b0 ;
  assign y8785 = n29888 ;
  assign y8786 = ~n29889 ;
  assign y8787 = ~n29895 ;
  assign y8788 = n29901 ;
  assign y8789 = ~n29905 ;
  assign y8790 = n29907 ;
  assign y8791 = ~n29910 ;
  assign y8792 = n29911 ;
  assign y8793 = n29915 ;
  assign y8794 = ~n29917 ;
  assign y8795 = n29918 ;
  assign y8796 = ~n29925 ;
  assign y8797 = n29926 ;
  assign y8798 = ~n29927 ;
  assign y8799 = ~1'b0 ;
  assign y8800 = ~1'b0 ;
  assign y8801 = n29929 ;
  assign y8802 = n29933 ;
  assign y8803 = ~n29934 ;
  assign y8804 = ~n29937 ;
  assign y8805 = n29938 ;
  assign y8806 = ~n29939 ;
  assign y8807 = ~n29940 ;
  assign y8808 = ~1'b0 ;
  assign y8809 = n29945 ;
  assign y8810 = n29949 ;
  assign y8811 = ~n29950 ;
  assign y8812 = ~1'b0 ;
  assign y8813 = ~n29959 ;
  assign y8814 = ~1'b0 ;
  assign y8815 = n29962 ;
  assign y8816 = n29971 ;
  assign y8817 = ~n29973 ;
  assign y8818 = n29975 ;
  assign y8819 = n29978 ;
  assign y8820 = n29979 ;
  assign y8821 = n29981 ;
  assign y8822 = n29982 ;
  assign y8823 = ~n29984 ;
  assign y8824 = ~n29992 ;
  assign y8825 = n29993 ;
  assign y8826 = ~n29994 ;
  assign y8827 = ~n29998 ;
  assign y8828 = ~n30000 ;
  assign y8829 = 1'b0 ;
  assign y8830 = n30002 ;
  assign y8831 = ~n30009 ;
  assign y8832 = n30012 ;
  assign y8833 = ~n30013 ;
  assign y8834 = n30023 ;
  assign y8835 = ~n30027 ;
  assign y8836 = ~n30035 ;
  assign y8837 = ~n30038 ;
  assign y8838 = ~n30042 ;
  assign y8839 = n30046 ;
  assign y8840 = ~1'b0 ;
  assign y8841 = ~n30049 ;
  assign y8842 = n30050 ;
  assign y8843 = n30054 ;
  assign y8844 = n30056 ;
  assign y8845 = n30061 ;
  assign y8846 = ~n30063 ;
  assign y8847 = n30065 ;
  assign y8848 = ~n30066 ;
  assign y8849 = ~1'b0 ;
  assign y8850 = ~n30069 ;
  assign y8851 = n30071 ;
  assign y8852 = ~n30073 ;
  assign y8853 = ~n30075 ;
  assign y8854 = ~1'b0 ;
  assign y8855 = ~1'b0 ;
  assign y8856 = ~n30080 ;
  assign y8857 = n30081 ;
  assign y8858 = n30083 ;
  assign y8859 = ~n30084 ;
  assign y8860 = n30086 ;
  assign y8861 = n30090 ;
  assign y8862 = ~n30095 ;
  assign y8863 = ~n30099 ;
  assign y8864 = ~n30100 ;
  assign y8865 = ~n30104 ;
  assign y8866 = n30108 ;
  assign y8867 = ~1'b0 ;
  assign y8868 = ~n30110 ;
  assign y8869 = ~n30113 ;
  assign y8870 = ~n30115 ;
  assign y8871 = ~n30119 ;
  assign y8872 = n30122 ;
  assign y8873 = ~n30125 ;
  assign y8874 = n4671 ;
  assign y8875 = ~n30127 ;
  assign y8876 = n30132 ;
  assign y8877 = n30135 ;
  assign y8878 = n30138 ;
  assign y8879 = n30140 ;
  assign y8880 = ~n30144 ;
  assign y8881 = ~n30151 ;
  assign y8882 = n30156 ;
  assign y8883 = n30157 ;
  assign y8884 = ~1'b0 ;
  assign y8885 = ~n28398 ;
  assign y8886 = ~n30160 ;
  assign y8887 = ~n21014 ;
  assign y8888 = n30165 ;
  assign y8889 = ~n30168 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = n30172 ;
  assign y8892 = n30174 ;
  assign y8893 = ~n30181 ;
  assign y8894 = n30185 ;
  assign y8895 = ~1'b0 ;
  assign y8896 = ~1'b0 ;
  assign y8897 = n30186 ;
  assign y8898 = n30192 ;
  assign y8899 = n30193 ;
  assign y8900 = n30209 ;
  assign y8901 = n30210 ;
  assign y8902 = ~1'b0 ;
  assign y8903 = n30215 ;
  assign y8904 = n30217 ;
  assign y8905 = ~1'b0 ;
  assign y8906 = n30219 ;
  assign y8907 = n30220 ;
  assign y8908 = n30222 ;
  assign y8909 = ~n30225 ;
  assign y8910 = n30229 ;
  assign y8911 = n30230 ;
  assign y8912 = ~n30233 ;
  assign y8913 = ~n30236 ;
  assign y8914 = n30237 ;
  assign y8915 = ~n30241 ;
  assign y8916 = n30246 ;
  assign y8917 = ~1'b0 ;
  assign y8918 = ~n30249 ;
  assign y8919 = n30250 ;
  assign y8920 = ~n30252 ;
  assign y8921 = n30253 ;
  assign y8922 = ~n30259 ;
  assign y8923 = ~n30263 ;
  assign y8924 = n30264 ;
  assign y8925 = ~n30265 ;
  assign y8926 = ~n30267 ;
  assign y8927 = n30273 ;
  assign y8928 = ~1'b0 ;
  assign y8929 = ~n30277 ;
  assign y8930 = ~n30278 ;
  assign y8931 = ~1'b0 ;
  assign y8932 = ~1'b0 ;
  assign y8933 = n30279 ;
  assign y8934 = n30280 ;
  assign y8935 = ~1'b0 ;
  assign y8936 = ~n30281 ;
  assign y8937 = ~n28439 ;
  assign y8938 = ~n30283 ;
  assign y8939 = ~n30284 ;
  assign y8940 = ~1'b0 ;
  assign y8941 = ~n30288 ;
  assign y8942 = n30294 ;
  assign y8943 = ~n30302 ;
  assign y8944 = n30306 ;
  assign y8945 = ~n30310 ;
  assign y8946 = ~1'b0 ;
  assign y8947 = n30316 ;
  assign y8948 = n30322 ;
  assign y8949 = ~n30324 ;
  assign y8950 = ~n30332 ;
  assign y8951 = n30337 ;
  assign y8952 = ~1'b0 ;
  assign y8953 = ~n30339 ;
  assign y8954 = ~n30344 ;
  assign y8955 = n30346 ;
  assign y8956 = ~n30348 ;
  assign y8957 = ~1'b0 ;
  assign y8958 = ~n30349 ;
  assign y8959 = ~n30356 ;
  assign y8960 = ~n30359 ;
  assign y8961 = ~n30360 ;
  assign y8962 = n30361 ;
  assign y8963 = n30366 ;
  assign y8964 = n30369 ;
  assign y8965 = ~n30376 ;
  assign y8966 = n30382 ;
  assign y8967 = ~n30383 ;
  assign y8968 = ~n30386 ;
  assign y8969 = ~1'b0 ;
  assign y8970 = ~1'b0 ;
  assign y8971 = n30399 ;
  assign y8972 = n30404 ;
  assign y8973 = ~n30407 ;
  assign y8974 = ~n30410 ;
  assign y8975 = n30411 ;
  assign y8976 = n30414 ;
  assign y8977 = n30420 ;
  assign y8978 = n30427 ;
  assign y8979 = ~n30432 ;
  assign y8980 = ~n30435 ;
  assign y8981 = ~n30437 ;
  assign y8982 = ~n30439 ;
  assign y8983 = ~n30440 ;
  assign y8984 = n30441 ;
  assign y8985 = n30442 ;
  assign y8986 = ~n30446 ;
  assign y8987 = ~1'b0 ;
  assign y8988 = n30451 ;
  assign y8989 = n30453 ;
  assign y8990 = ~n30462 ;
  assign y8991 = ~n30467 ;
  assign y8992 = ~n30469 ;
  assign y8993 = n30471 ;
  assign y8994 = ~n30482 ;
  assign y8995 = n30484 ;
  assign y8996 = ~n30486 ;
  assign y8997 = ~1'b0 ;
  assign y8998 = n30487 ;
  assign y8999 = n30490 ;
  assign y9000 = n30492 ;
  assign y9001 = n30493 ;
  assign y9002 = n30496 ;
  assign y9003 = ~n30497 ;
  assign y9004 = ~1'b0 ;
  assign y9005 = n30498 ;
  assign y9006 = n30499 ;
  assign y9007 = ~n30502 ;
  assign y9008 = n30505 ;
  assign y9009 = ~1'b0 ;
  assign y9010 = ~1'b0 ;
  assign y9011 = ~1'b0 ;
  assign y9012 = n30507 ;
  assign y9013 = ~n30511 ;
  assign y9014 = n30513 ;
  assign y9015 = n30515 ;
  assign y9016 = n30518 ;
  assign y9017 = n30520 ;
  assign y9018 = n30523 ;
  assign y9019 = n30524 ;
  assign y9020 = ~n30531 ;
  assign y9021 = ~1'b0 ;
  assign y9022 = ~n30533 ;
  assign y9023 = ~1'b0 ;
  assign y9024 = n30534 ;
  assign y9025 = ~n30538 ;
  assign y9026 = ~n30543 ;
  assign y9027 = ~1'b0 ;
  assign y9028 = n30552 ;
  assign y9029 = n30554 ;
  assign y9030 = ~n30555 ;
  assign y9031 = ~n30557 ;
  assign y9032 = ~n30559 ;
  assign y9033 = n30561 ;
  assign y9034 = ~n30563 ;
  assign y9035 = ~n30567 ;
  assign y9036 = ~n30571 ;
  assign y9037 = ~n20146 ;
  assign y9038 = ~1'b0 ;
  assign y9039 = ~n30573 ;
  assign y9040 = ~n30575 ;
  assign y9041 = ~n30578 ;
  assign y9042 = n30579 ;
  assign y9043 = ~n30581 ;
  assign y9044 = ~n30584 ;
  assign y9045 = ~n30585 ;
  assign y9046 = n30587 ;
  assign y9047 = n30588 ;
  assign y9048 = n30589 ;
  assign y9049 = n30591 ;
  assign y9050 = n30593 ;
  assign y9051 = ~n30601 ;
  assign y9052 = ~n30602 ;
  assign y9053 = n30605 ;
  assign y9054 = ~n30611 ;
  assign y9055 = n30614 ;
  assign y9056 = n30618 ;
  assign y9057 = n30619 ;
  assign y9058 = ~n30627 ;
  assign y9059 = ~n30630 ;
  assign y9060 = ~n30637 ;
  assign y9061 = n30641 ;
  assign y9062 = ~1'b0 ;
  assign y9063 = n30648 ;
  assign y9064 = n30653 ;
  assign y9065 = ~n30655 ;
  assign y9066 = ~n30656 ;
  assign y9067 = ~n30657 ;
  assign y9068 = n30658 ;
  assign y9069 = ~n30660 ;
  assign y9070 = n30664 ;
  assign y9071 = ~n30673 ;
  assign y9072 = n30675 ;
  assign y9073 = ~n30677 ;
  assign y9074 = ~n30678 ;
  assign y9075 = ~n30680 ;
  assign y9076 = n30681 ;
  assign y9077 = n30684 ;
  assign y9078 = ~n30686 ;
  assign y9079 = ~n30688 ;
  assign y9080 = n30691 ;
  assign y9081 = ~1'b0 ;
  assign y9082 = n30696 ;
  assign y9083 = n30698 ;
  assign y9084 = ~n30701 ;
  assign y9085 = n30705 ;
  assign y9086 = ~1'b0 ;
  assign y9087 = n30708 ;
  assign y9088 = n30712 ;
  assign y9089 = ~n30716 ;
  assign y9090 = n30718 ;
  assign y9091 = n30720 ;
  assign y9092 = ~n7301 ;
  assign y9093 = ~n30722 ;
  assign y9094 = n30723 ;
  assign y9095 = ~n30729 ;
  assign y9096 = ~1'b0 ;
  assign y9097 = ~n30732 ;
  assign y9098 = n30735 ;
  assign y9099 = n17637 ;
  assign y9100 = ~n30737 ;
  assign y9101 = n30738 ;
  assign y9102 = ~n30741 ;
  assign y9103 = n30742 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = n30747 ;
  assign y9106 = ~n30748 ;
  assign y9107 = ~n30751 ;
  assign y9108 = ~n30752 ;
  assign y9109 = n30755 ;
  assign y9110 = n30759 ;
  assign y9111 = ~n30762 ;
  assign y9112 = n30773 ;
  assign y9113 = ~n30774 ;
  assign y9114 = ~n30775 ;
  assign y9115 = ~n30779 ;
  assign y9116 = n30793 ;
  assign y9117 = n30803 ;
  assign y9118 = n30811 ;
  assign y9119 = ~n30815 ;
  assign y9120 = ~n30816 ;
  assign y9121 = ~1'b0 ;
  assign y9122 = ~1'b0 ;
  assign y9123 = n30818 ;
  assign y9124 = ~n30819 ;
  assign y9125 = n30823 ;
  assign y9126 = ~n2375 ;
  assign y9127 = ~n30826 ;
  assign y9128 = ~n30828 ;
  assign y9129 = n30829 ;
  assign y9130 = ~1'b0 ;
  assign y9131 = ~n30833 ;
  assign y9132 = n30839 ;
  assign y9133 = n30841 ;
  assign y9134 = ~1'b0 ;
  assign y9135 = ~n30842 ;
  assign y9136 = ~n30856 ;
  assign y9137 = ~n30857 ;
  assign y9138 = n30865 ;
  assign y9139 = ~n30868 ;
  assign y9140 = ~n30870 ;
  assign y9141 = ~n30873 ;
  assign y9142 = ~1'b0 ;
  assign y9143 = ~1'b0 ;
  assign y9144 = ~n30879 ;
  assign y9145 = n30887 ;
  assign y9146 = n30888 ;
  assign y9147 = n30889 ;
  assign y9148 = ~n30891 ;
  assign y9149 = n30893 ;
  assign y9150 = n30895 ;
  assign y9151 = ~n30896 ;
  assign y9152 = ~n30897 ;
  assign y9153 = n30898 ;
  assign y9154 = ~n30901 ;
  assign y9155 = ~n30903 ;
  assign y9156 = ~n30905 ;
  assign y9157 = n30906 ;
  assign y9158 = ~n30907 ;
  assign y9159 = n30909 ;
  assign y9160 = ~n30912 ;
  assign y9161 = ~n30914 ;
  assign y9162 = n30915 ;
  assign y9163 = ~1'b0 ;
  assign y9164 = n30918 ;
  assign y9165 = n30923 ;
  assign y9166 = n30924 ;
  assign y9167 = n30926 ;
  assign y9168 = n30928 ;
  assign y9169 = ~n30930 ;
  assign y9170 = n30931 ;
  assign y9171 = n30934 ;
  assign y9172 = n30942 ;
  assign y9173 = n30944 ;
  assign y9174 = ~1'b0 ;
  assign y9175 = ~n30945 ;
  assign y9176 = n30948 ;
  assign y9177 = n30957 ;
  assign y9178 = n30958 ;
  assign y9179 = ~1'b0 ;
  assign y9180 = n30960 ;
  assign y9181 = n30961 ;
  assign y9182 = n30965 ;
  assign y9183 = ~n30966 ;
  assign y9184 = ~n30970 ;
  assign y9185 = ~n30973 ;
  assign y9186 = ~n30974 ;
  assign y9187 = ~n30977 ;
  assign y9188 = n30978 ;
  assign y9189 = ~n30979 ;
  assign y9190 = ~n30980 ;
  assign y9191 = ~1'b0 ;
  assign y9192 = ~n30985 ;
  assign y9193 = n30996 ;
  assign y9194 = ~n30999 ;
  assign y9195 = ~n31002 ;
  assign y9196 = n4141 ;
  assign y9197 = ~1'b0 ;
  assign y9198 = ~1'b0 ;
  assign y9199 = n31004 ;
  assign y9200 = ~n31006 ;
  assign y9201 = n31009 ;
  assign y9202 = ~n31012 ;
  assign y9203 = n31015 ;
  assign y9204 = n31016 ;
  assign y9205 = ~n31018 ;
  assign y9206 = ~1'b0 ;
  assign y9207 = ~1'b0 ;
  assign y9208 = ~n27033 ;
  assign y9209 = n31023 ;
  assign y9210 = ~n31024 ;
  assign y9211 = n31025 ;
  assign y9212 = ~n31027 ;
  assign y9213 = ~n31029 ;
  assign y9214 = n31031 ;
  assign y9215 = ~n31032 ;
  assign y9216 = n31038 ;
  assign y9217 = ~n31039 ;
  assign y9218 = ~n31043 ;
  assign y9219 = n31045 ;
  assign y9220 = n31050 ;
  assign y9221 = ~n31053 ;
  assign y9222 = ~n31056 ;
  assign y9223 = ~n31059 ;
  assign y9224 = ~n31063 ;
  assign y9225 = ~n31065 ;
  assign y9226 = n31067 ;
  assign y9227 = ~n31070 ;
  assign y9228 = 1'b0 ;
  assign y9229 = n31080 ;
  assign y9230 = ~n31081 ;
  assign y9231 = ~n31083 ;
  assign y9232 = n31085 ;
  assign y9233 = n31086 ;
  assign y9234 = n31087 ;
  assign y9235 = ~n31093 ;
  assign y9236 = ~n31097 ;
  assign y9237 = ~n31100 ;
  assign y9238 = ~n31106 ;
  assign y9239 = ~n31107 ;
  assign y9240 = n31110 ;
  assign y9241 = ~n31111 ;
  assign y9242 = n31114 ;
  assign y9243 = n31122 ;
  assign y9244 = ~n31126 ;
  assign y9245 = ~n31127 ;
  assign y9246 = n31128 ;
  assign y9247 = ~n31131 ;
  assign y9248 = ~n31134 ;
  assign y9249 = ~n31136 ;
  assign y9250 = n31137 ;
  assign y9251 = ~n31138 ;
  assign y9252 = ~n31139 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = n31141 ;
  assign y9255 = ~n31148 ;
  assign y9256 = ~n31152 ;
  assign y9257 = ~n31155 ;
  assign y9258 = ~n31159 ;
  assign y9259 = ~n31163 ;
  assign y9260 = ~n31164 ;
  assign y9261 = n31169 ;
  assign y9262 = 1'b0 ;
  assign y9263 = ~1'b0 ;
  assign y9264 = n31174 ;
  assign y9265 = ~n31176 ;
  assign y9266 = ~n31178 ;
  assign y9267 = n31179 ;
  assign y9268 = ~1'b0 ;
  assign y9269 = ~1'b0 ;
  assign y9270 = ~n31181 ;
  assign y9271 = ~n31184 ;
  assign y9272 = ~n31190 ;
  assign y9273 = ~1'b0 ;
  assign y9274 = n31191 ;
  assign y9275 = n31194 ;
  assign y9276 = n31197 ;
  assign y9277 = n31199 ;
  assign y9278 = 1'b0 ;
  assign y9279 = n31202 ;
  assign y9280 = n31204 ;
  assign y9281 = ~n31209 ;
  assign y9282 = n31211 ;
  assign y9283 = n31213 ;
  assign y9284 = n31215 ;
  assign y9285 = n31216 ;
  assign y9286 = ~n31220 ;
  assign y9287 = ~1'b0 ;
  assign y9288 = ~n31221 ;
  assign y9289 = n31226 ;
  assign y9290 = ~n31230 ;
  assign y9291 = n31233 ;
  assign y9292 = ~n31235 ;
  assign y9293 = n31237 ;
  assign y9294 = ~n31242 ;
  assign y9295 = ~1'b0 ;
  assign y9296 = ~1'b0 ;
  assign y9297 = n31244 ;
  assign y9298 = ~n31246 ;
  assign y9299 = n31250 ;
  assign y9300 = ~n31254 ;
  assign y9301 = n31257 ;
  assign y9302 = n31259 ;
  assign y9303 = ~n31261 ;
  assign y9304 = ~n31262 ;
  assign y9305 = n31265 ;
  assign y9306 = n31270 ;
  assign y9307 = ~1'b0 ;
  assign y9308 = ~1'b0 ;
  assign y9309 = ~n31278 ;
  assign y9310 = n31279 ;
  assign y9311 = n31280 ;
  assign y9312 = ~n31283 ;
  assign y9313 = ~1'b0 ;
  assign y9314 = ~n31289 ;
  assign y9315 = n31291 ;
  assign y9316 = n31296 ;
  assign y9317 = ~n31297 ;
  assign y9318 = ~n31300 ;
  assign y9319 = n31302 ;
  assign y9320 = n31304 ;
  assign y9321 = ~n31309 ;
  assign y9322 = ~n31311 ;
  assign y9323 = ~n31312 ;
  assign y9324 = n31315 ;
  assign y9325 = n31321 ;
  assign y9326 = ~n31322 ;
  assign y9327 = ~n31325 ;
  assign y9328 = ~n31326 ;
  assign y9329 = ~n31327 ;
  assign y9330 = n31331 ;
  assign y9331 = ~n31332 ;
  assign y9332 = ~n31333 ;
  assign y9333 = ~1'b0 ;
  assign y9334 = ~1'b0 ;
  assign y9335 = n31334 ;
  assign y9336 = ~n31337 ;
  assign y9337 = n31341 ;
  assign y9338 = ~n31348 ;
  assign y9339 = ~1'b0 ;
  assign y9340 = n31351 ;
  assign y9341 = ~1'b0 ;
  assign y9342 = ~n31359 ;
  assign y9343 = n31364 ;
  assign y9344 = ~n31367 ;
  assign y9345 = ~n31368 ;
  assign y9346 = n31374 ;
  assign y9347 = ~n31379 ;
  assign y9348 = n31381 ;
  assign y9349 = n31384 ;
  assign y9350 = ~1'b0 ;
  assign y9351 = ~n31386 ;
  assign y9352 = ~n31388 ;
  assign y9353 = ~n31389 ;
  assign y9354 = n31391 ;
  assign y9355 = n31396 ;
  assign y9356 = n31399 ;
  assign y9357 = ~n31401 ;
  assign y9358 = ~n31403 ;
  assign y9359 = n31413 ;
  assign y9360 = n31414 ;
  assign y9361 = ~n31416 ;
  assign y9362 = n31419 ;
  assign y9363 = n31423 ;
  assign y9364 = ~n31426 ;
  assign y9365 = n31427 ;
  assign y9366 = ~n31431 ;
  assign y9367 = ~n31441 ;
  assign y9368 = ~n31445 ;
  assign y9369 = ~n31447 ;
  assign y9370 = n31453 ;
  assign y9371 = n31458 ;
  assign y9372 = n31463 ;
  assign y9373 = ~1'b0 ;
  assign y9374 = ~n31466 ;
  assign y9375 = n31467 ;
  assign y9376 = ~n31468 ;
  assign y9377 = n31471 ;
  assign y9378 = n31476 ;
  assign y9379 = ~n31479 ;
  assign y9380 = ~n31481 ;
  assign y9381 = ~n31486 ;
  assign y9382 = ~n31488 ;
  assign y9383 = ~1'b0 ;
  assign y9384 = n31489 ;
  assign y9385 = ~n31491 ;
  assign y9386 = ~n31498 ;
  assign y9387 = ~n31501 ;
  assign y9388 = n31503 ;
  assign y9389 = n31505 ;
  assign y9390 = ~n31507 ;
  assign y9391 = ~n31513 ;
  assign y9392 = ~n31514 ;
  assign y9393 = ~n31518 ;
  assign y9394 = ~n31520 ;
  assign y9395 = ~1'b0 ;
  assign y9396 = ~n31522 ;
  assign y9397 = ~n31523 ;
  assign y9398 = ~n31524 ;
  assign y9399 = n31530 ;
  assign y9400 = n31535 ;
  assign y9401 = n31536 ;
  assign y9402 = ~1'b0 ;
  assign y9403 = ~n31538 ;
  assign y9404 = ~n31541 ;
  assign y9405 = n31542 ;
  assign y9406 = ~1'b0 ;
  assign y9407 = n31544 ;
  assign y9408 = n31546 ;
  assign y9409 = n31547 ;
  assign y9410 = ~n31550 ;
  assign y9411 = n31556 ;
  assign y9412 = ~n31558 ;
  assign y9413 = ~1'b0 ;
  assign y9414 = ~1'b0 ;
  assign y9415 = ~n24188 ;
  assign y9416 = ~n31559 ;
  assign y9417 = n31560 ;
  assign y9418 = n31567 ;
  assign y9419 = n31569 ;
  assign y9420 = n31570 ;
  assign y9421 = ~n31573 ;
  assign y9422 = ~n31574 ;
  assign y9423 = ~n31582 ;
  assign y9424 = ~n31585 ;
  assign y9425 = n31588 ;
  assign y9426 = ~n31590 ;
  assign y9427 = ~n31592 ;
  assign y9428 = ~n31601 ;
  assign y9429 = n31606 ;
  assign y9430 = ~n31607 ;
  assign y9431 = ~n31609 ;
  assign y9432 = n31611 ;
  assign y9433 = n31612 ;
  assign y9434 = ~n31616 ;
  assign y9435 = ~n31617 ;
  assign y9436 = ~n31621 ;
  assign y9437 = ~n31627 ;
  assign y9438 = n31628 ;
  assign y9439 = n31631 ;
  assign y9440 = ~1'b0 ;
  assign y9441 = ~n31633 ;
  assign y9442 = ~n31636 ;
  assign y9443 = ~n31639 ;
  assign y9444 = ~n31641 ;
  assign y9445 = ~n31646 ;
  assign y9446 = ~n31648 ;
  assign y9447 = n31652 ;
  assign y9448 = n31653 ;
  assign y9449 = n31659 ;
  assign y9450 = ~n31660 ;
  assign y9451 = n31664 ;
  assign y9452 = ~n31666 ;
  assign y9453 = ~n31671 ;
  assign y9454 = n31672 ;
  assign y9455 = ~n31673 ;
  assign y9456 = n31676 ;
  assign y9457 = n31677 ;
  assign y9458 = n31678 ;
  assign y9459 = ~n31681 ;
  assign y9460 = ~n31685 ;
  assign y9461 = n31686 ;
  assign y9462 = n31689 ;
  assign y9463 = ~n31692 ;
  assign y9464 = ~n31694 ;
  assign y9465 = n31696 ;
  assign y9466 = n31702 ;
  assign y9467 = ~n31706 ;
  assign y9468 = n31708 ;
  assign y9469 = ~n31711 ;
  assign y9470 = ~n31713 ;
  assign y9471 = ~n31715 ;
  assign y9472 = n31717 ;
  assign y9473 = n31719 ;
  assign y9474 = n31720 ;
  assign y9475 = ~n31721 ;
  assign y9476 = n31722 ;
  assign y9477 = ~1'b0 ;
  assign y9478 = ~n31723 ;
  assign y9479 = n31727 ;
  assign y9480 = ~n31732 ;
  assign y9481 = ~n31736 ;
  assign y9482 = n31738 ;
  assign y9483 = n31743 ;
  assign y9484 = ~n31744 ;
  assign y9485 = ~n31745 ;
  assign y9486 = ~n31746 ;
  assign y9487 = n31752 ;
  assign y9488 = n31754 ;
  assign y9489 = ~n31759 ;
  assign y9490 = ~1'b0 ;
  assign y9491 = ~n31762 ;
  assign y9492 = ~1'b0 ;
  assign y9493 = n31763 ;
  assign y9494 = n31770 ;
  assign y9495 = ~n31771 ;
  assign y9496 = n31773 ;
  assign y9497 = n31775 ;
  assign y9498 = n31783 ;
  assign y9499 = ~n31789 ;
  assign y9500 = n31791 ;
  assign y9501 = n31794 ;
  assign y9502 = n31795 ;
  assign y9503 = n31797 ;
  assign y9504 = ~n31798 ;
  assign y9505 = ~n31804 ;
  assign y9506 = n14697 ;
  assign y9507 = n31805 ;
  assign y9508 = n31808 ;
  assign y9509 = ~n31809 ;
  assign y9510 = ~n31814 ;
  assign y9511 = ~1'b0 ;
  assign y9512 = n31817 ;
  assign y9513 = n31819 ;
  assign y9514 = n31825 ;
  assign y9515 = ~1'b0 ;
  assign y9516 = ~n31829 ;
  assign y9517 = n31833 ;
  assign y9518 = ~n31836 ;
  assign y9519 = ~n31837 ;
  assign y9520 = n31838 ;
  assign y9521 = ~n31840 ;
  assign y9522 = n31842 ;
  assign y9523 = ~n31850 ;
  assign y9524 = n31851 ;
  assign y9525 = n31854 ;
  assign y9526 = ~n9045 ;
  assign y9527 = n31856 ;
  assign y9528 = ~n31859 ;
  assign y9529 = n31862 ;
  assign y9530 = ~n31868 ;
  assign y9531 = n31875 ;
  assign y9532 = ~n31877 ;
  assign y9533 = n31881 ;
  assign y9534 = ~n31882 ;
  assign y9535 = ~1'b0 ;
  assign y9536 = ~1'b0 ;
  assign y9537 = ~n31886 ;
  assign y9538 = n31893 ;
  assign y9539 = n31894 ;
  assign y9540 = ~1'b0 ;
  assign y9541 = n31897 ;
  assign y9542 = n31901 ;
  assign y9543 = ~n31905 ;
  assign y9544 = ~n31909 ;
  assign y9545 = 1'b0 ;
  assign y9546 = ~n31910 ;
  assign y9547 = ~n31911 ;
  assign y9548 = n22725 ;
  assign y9549 = n31914 ;
  assign y9550 = ~1'b0 ;
  assign y9551 = n31915 ;
  assign y9552 = ~n31920 ;
  assign y9553 = n31925 ;
  assign y9554 = ~n31926 ;
  assign y9555 = ~n31931 ;
  assign y9556 = ~1'b0 ;
  assign y9557 = ~n31933 ;
  assign y9558 = n31939 ;
  assign y9559 = n31940 ;
  assign y9560 = n31943 ;
  assign y9561 = n31948 ;
  assign y9562 = ~1'b0 ;
  assign y9563 = ~n31949 ;
  assign y9564 = n31953 ;
  assign y9565 = ~n31954 ;
  assign y9566 = ~n31955 ;
  assign y9567 = n31964 ;
  assign y9568 = n31968 ;
  assign y9569 = ~n31969 ;
  assign y9570 = n31971 ;
  assign y9571 = n31973 ;
  assign y9572 = n31979 ;
  assign y9573 = ~n31981 ;
  assign y9574 = n31986 ;
  assign y9575 = ~n31988 ;
  assign y9576 = ~n31989 ;
  assign y9577 = n31997 ;
  assign y9578 = n32000 ;
  assign y9579 = ~n32003 ;
  assign y9580 = ~n32009 ;
  assign y9581 = ~1'b0 ;
  assign y9582 = ~n32010 ;
  assign y9583 = n32021 ;
  assign y9584 = n32023 ;
  assign y9585 = ~1'b0 ;
  assign y9586 = n32026 ;
  assign y9587 = n32031 ;
  assign y9588 = ~n32033 ;
  assign y9589 = n10530 ;
  assign y9590 = ~n32034 ;
  assign y9591 = ~n32039 ;
  assign y9592 = ~1'b0 ;
  assign y9593 = n32041 ;
  assign y9594 = ~n32045 ;
  assign y9595 = ~n32050 ;
  assign y9596 = ~n32056 ;
  assign y9597 = ~n32062 ;
  assign y9598 = ~n32063 ;
  assign y9599 = n32064 ;
  assign y9600 = ~n32068 ;
  assign y9601 = ~1'b0 ;
  assign y9602 = ~1'b0 ;
  assign y9603 = ~n32074 ;
  assign y9604 = n32075 ;
  assign y9605 = ~n32076 ;
  assign y9606 = ~1'b0 ;
  assign y9607 = ~1'b0 ;
  assign y9608 = ~n32077 ;
  assign y9609 = ~n32080 ;
  assign y9610 = ~n7817 ;
  assign y9611 = ~n32083 ;
  assign y9612 = ~1'b0 ;
  assign y9613 = n32085 ;
  assign y9614 = n32096 ;
  assign y9615 = ~n32097 ;
  assign y9616 = n32100 ;
  assign y9617 = n32102 ;
  assign y9618 = ~n32106 ;
  assign y9619 = ~n32112 ;
  assign y9620 = ~1'b0 ;
  assign y9621 = n32113 ;
  assign y9622 = ~n32115 ;
  assign y9623 = n32116 ;
  assign y9624 = n32117 ;
  assign y9625 = ~1'b0 ;
  assign y9626 = ~n32118 ;
  assign y9627 = ~n32119 ;
  assign y9628 = ~n32120 ;
  assign y9629 = ~1'b0 ;
  assign y9630 = n32123 ;
  assign y9631 = n32125 ;
  assign y9632 = ~n32127 ;
  assign y9633 = ~n32131 ;
  assign y9634 = n32132 ;
  assign y9635 = ~n32140 ;
  assign y9636 = ~n32150 ;
  assign y9637 = n32151 ;
  assign y9638 = ~n32154 ;
  assign y9639 = n32157 ;
  assign y9640 = ~1'b0 ;
  assign y9641 = ~1'b0 ;
  assign y9642 = ~n32158 ;
  assign y9643 = ~n32159 ;
  assign y9644 = n32161 ;
  assign y9645 = ~n32164 ;
  assign y9646 = ~1'b0 ;
  assign y9647 = ~n32166 ;
  assign y9648 = n32173 ;
  assign y9649 = n32174 ;
  assign y9650 = n32175 ;
  assign y9651 = n32178 ;
  assign y9652 = ~n32186 ;
  assign y9653 = ~n32187 ;
  assign y9654 = n27285 ;
  assign y9655 = ~n32188 ;
  assign y9656 = ~n32190 ;
  assign y9657 = n18623 ;
  assign y9658 = n32191 ;
  assign y9659 = n32195 ;
  assign y9660 = n32196 ;
  assign y9661 = ~n32198 ;
  assign y9662 = ~n32203 ;
  assign y9663 = n32204 ;
  assign y9664 = ~n32206 ;
  assign y9665 = n32208 ;
  assign y9666 = ~n32212 ;
  assign y9667 = ~n32214 ;
  assign y9668 = ~1'b0 ;
  assign y9669 = ~n32215 ;
  assign y9670 = n32216 ;
  assign y9671 = ~1'b0 ;
  assign y9672 = ~1'b0 ;
  assign y9673 = ~n32219 ;
  assign y9674 = n32225 ;
  assign y9675 = ~n32233 ;
  assign y9676 = ~n32234 ;
  assign y9677 = ~n32235 ;
  assign y9678 = ~n32236 ;
  assign y9679 = ~n32239 ;
  assign y9680 = ~n32241 ;
  assign y9681 = ~1'b0 ;
  assign y9682 = n32245 ;
  assign y9683 = ~1'b0 ;
  assign y9684 = n32246 ;
  assign y9685 = ~n32248 ;
  assign y9686 = ~n32249 ;
  assign y9687 = ~n32252 ;
  assign y9688 = n32255 ;
  assign y9689 = n32259 ;
  assign y9690 = n32260 ;
  assign y9691 = n32261 ;
  assign y9692 = n32266 ;
  assign y9693 = ~n32269 ;
  assign y9694 = n32270 ;
  assign y9695 = n32274 ;
  assign y9696 = ~1'b0 ;
  assign y9697 = n32278 ;
  assign y9698 = ~n32286 ;
  assign y9699 = ~n32289 ;
  assign y9700 = n32291 ;
  assign y9701 = n32292 ;
  assign y9702 = ~n32298 ;
  assign y9703 = ~1'b0 ;
  assign y9704 = n32300 ;
  assign y9705 = n32301 ;
  assign y9706 = n32306 ;
  assign y9707 = ~n32307 ;
  assign y9708 = ~n32310 ;
  assign y9709 = ~n32316 ;
  assign y9710 = n32317 ;
  assign y9711 = ~n32321 ;
  assign y9712 = ~n32323 ;
  assign y9713 = n32324 ;
  assign y9714 = ~n32328 ;
  assign y9715 = ~n32331 ;
  assign y9716 = ~n32336 ;
  assign y9717 = ~1'b0 ;
  assign y9718 = ~n32340 ;
  assign y9719 = ~1'b0 ;
  assign y9720 = ~n32342 ;
  assign y9721 = n32346 ;
  assign y9722 = n32349 ;
  assign y9723 = ~1'b0 ;
  assign y9724 = n32355 ;
  assign y9725 = ~n32356 ;
  assign y9726 = ~n32357 ;
  assign y9727 = ~1'b0 ;
  assign y9728 = ~1'b0 ;
  assign y9729 = ~1'b0 ;
  assign y9730 = n32359 ;
  assign y9731 = n32361 ;
  assign y9732 = ~n32363 ;
  assign y9733 = ~n32366 ;
  assign y9734 = ~n32367 ;
  assign y9735 = ~n32368 ;
  assign y9736 = ~n32369 ;
  assign y9737 = ~n32377 ;
  assign y9738 = ~n32378 ;
  assign y9739 = n32379 ;
  assign y9740 = ~n32381 ;
  assign y9741 = ~1'b0 ;
  assign y9742 = ~n32384 ;
  assign y9743 = n32386 ;
  assign y9744 = n32387 ;
  assign y9745 = n32390 ;
  assign y9746 = ~n32396 ;
  assign y9747 = ~n32397 ;
  assign y9748 = ~n32399 ;
  assign y9749 = n32402 ;
  assign y9750 = n32404 ;
  assign y9751 = n32412 ;
  assign y9752 = n32414 ;
  assign y9753 = ~n32415 ;
  assign y9754 = n32416 ;
  assign y9755 = n32418 ;
  assign y9756 = n32419 ;
  assign y9757 = ~n32420 ;
  assign y9758 = ~1'b0 ;
  assign y9759 = n32422 ;
  assign y9760 = ~n32424 ;
  assign y9761 = ~n32428 ;
  assign y9762 = ~n32434 ;
  assign y9763 = ~n32438 ;
  assign y9764 = ~n32440 ;
  assign y9765 = n32441 ;
  assign y9766 = n32442 ;
  assign y9767 = ~n32450 ;
  assign y9768 = ~n32454 ;
  assign y9769 = ~n32462 ;
  assign y9770 = n32464 ;
  assign y9771 = ~n32467 ;
  assign y9772 = n32468 ;
  assign y9773 = ~n32470 ;
  assign y9774 = ~1'b0 ;
  assign y9775 = ~1'b0 ;
  assign y9776 = n32473 ;
  assign y9777 = n32481 ;
  assign y9778 = ~n32484 ;
  assign y9779 = ~n32485 ;
  assign y9780 = ~1'b0 ;
  assign y9781 = ~n32487 ;
  assign y9782 = ~n32489 ;
  assign y9783 = n32491 ;
  assign y9784 = n32494 ;
  assign y9785 = ~n32500 ;
  assign y9786 = ~n32501 ;
  assign y9787 = ~n32507 ;
  assign y9788 = ~n32508 ;
  assign y9789 = n32518 ;
  assign y9790 = n21973 ;
  assign y9791 = ~1'b0 ;
  assign y9792 = ~n32519 ;
  assign y9793 = n32522 ;
  assign y9794 = n32529 ;
  assign y9795 = ~n32536 ;
  assign y9796 = ~n32537 ;
  assign y9797 = ~1'b0 ;
  assign y9798 = ~n32542 ;
  assign y9799 = ~n32544 ;
  assign y9800 = n32549 ;
  assign y9801 = ~n32551 ;
  assign y9802 = n32552 ;
  assign y9803 = ~1'b0 ;
  assign y9804 = ~1'b0 ;
  assign y9805 = n32554 ;
  assign y9806 = ~n32564 ;
  assign y9807 = ~n32566 ;
  assign y9808 = n32568 ;
  assign y9809 = ~n32577 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = ~1'b0 ;
  assign y9812 = n32579 ;
  assign y9813 = ~n32582 ;
  assign y9814 = n32587 ;
  assign y9815 = ~1'b0 ;
  assign y9816 = n32590 ;
  assign y9817 = ~n32593 ;
  assign y9818 = ~1'b0 ;
  assign y9819 = ~n32596 ;
  assign y9820 = ~n32597 ;
  assign y9821 = ~n32601 ;
  assign y9822 = ~n32604 ;
  assign y9823 = n32606 ;
  assign y9824 = ~n32615 ;
  assign y9825 = ~n32616 ;
  assign y9826 = ~n32617 ;
  assign y9827 = n32623 ;
  assign y9828 = ~n32627 ;
  assign y9829 = ~n32629 ;
  assign y9830 = n32631 ;
  assign y9831 = ~n32633 ;
  assign y9832 = n32634 ;
  assign y9833 = n32636 ;
  assign y9834 = ~n32637 ;
  assign y9835 = n32640 ;
  assign y9836 = n32644 ;
  assign y9837 = ~n32651 ;
  assign y9838 = ~n32654 ;
  assign y9839 = ~n32655 ;
  assign y9840 = ~n32657 ;
  assign y9841 = ~n32658 ;
  assign y9842 = n32660 ;
  assign y9843 = ~n32667 ;
  assign y9844 = ~n32669 ;
  assign y9845 = ~n32670 ;
  assign y9846 = ~1'b0 ;
  assign y9847 = ~n32674 ;
  assign y9848 = n32675 ;
  assign y9849 = n32676 ;
  assign y9850 = ~n32681 ;
  assign y9851 = ~n32683 ;
  assign y9852 = n32686 ;
  assign y9853 = n32688 ;
  assign y9854 = n32690 ;
  assign y9855 = ~n32693 ;
  assign y9856 = ~1'b0 ;
  assign y9857 = ~1'b0 ;
  assign y9858 = ~n32699 ;
  assign y9859 = ~n32700 ;
  assign y9860 = n32701 ;
  assign y9861 = ~1'b0 ;
  assign y9862 = ~1'b0 ;
  assign y9863 = n32706 ;
  assign y9864 = ~1'b0 ;
  assign y9865 = ~n32708 ;
  assign y9866 = ~n32711 ;
  assign y9867 = ~n32712 ;
  assign y9868 = ~n32713 ;
  assign y9869 = ~1'b0 ;
  assign y9870 = n32716 ;
  assign y9871 = n32717 ;
  assign y9872 = n32722 ;
  assign y9873 = ~n32723 ;
  assign y9874 = n32727 ;
  assign y9875 = ~1'b0 ;
  assign y9876 = ~1'b0 ;
  assign y9877 = ~n7494 ;
  assign y9878 = n32730 ;
  assign y9879 = n32741 ;
  assign y9880 = ~n32744 ;
  assign y9881 = ~n32747 ;
  assign y9882 = n32761 ;
  assign y9883 = n32764 ;
  assign y9884 = ~n32770 ;
  assign y9885 = n32778 ;
  assign y9886 = ~1'b0 ;
  assign y9887 = ~1'b0 ;
  assign y9888 = ~n32784 ;
  assign y9889 = n32785 ;
  assign y9890 = ~n32786 ;
  assign y9891 = ~n32788 ;
  assign y9892 = ~1'b0 ;
  assign y9893 = n32789 ;
  assign y9894 = ~n32791 ;
  assign y9895 = n32792 ;
  assign y9896 = n32794 ;
  assign y9897 = n32799 ;
  assign y9898 = n32808 ;
  assign y9899 = ~n32812 ;
  assign y9900 = ~n32814 ;
  assign y9901 = ~n32828 ;
  assign y9902 = ~n32830 ;
  assign y9903 = n32835 ;
  assign y9904 = n32836 ;
  assign y9905 = ~n32837 ;
  assign y9906 = n32838 ;
  assign y9907 = n32839 ;
  assign y9908 = ~n32843 ;
  assign y9909 = n32844 ;
  assign y9910 = n4627 ;
  assign y9911 = n32845 ;
  assign y9912 = n32848 ;
  assign y9913 = n32850 ;
  assign y9914 = n32858 ;
  assign y9915 = ~n32860 ;
  assign y9916 = n32861 ;
  assign y9917 = ~1'b0 ;
  assign y9918 = ~n32862 ;
  assign y9919 = ~n32865 ;
  assign y9920 = ~n32869 ;
  assign y9921 = ~n32870 ;
  assign y9922 = n32874 ;
  assign y9923 = ~1'b0 ;
  assign y9924 = ~n32875 ;
  assign y9925 = ~1'b0 ;
  assign y9926 = ~1'b0 ;
  assign y9927 = n32882 ;
  assign y9928 = n32885 ;
  assign y9929 = n32889 ;
  assign y9930 = n32893 ;
  assign y9931 = n32904 ;
  assign y9932 = n32907 ;
  assign y9933 = ~1'b0 ;
  assign y9934 = ~1'b0 ;
  assign y9935 = ~1'b0 ;
  assign y9936 = ~n32910 ;
  assign y9937 = n32915 ;
  assign y9938 = ~n32916 ;
  assign y9939 = ~n32918 ;
  assign y9940 = ~n32921 ;
  assign y9941 = ~n32926 ;
  assign y9942 = ~1'b0 ;
  assign y9943 = ~n32927 ;
  assign y9944 = ~n32937 ;
  assign y9945 = ~n32938 ;
  assign y9946 = ~1'b0 ;
  assign y9947 = ~n32940 ;
  assign y9948 = n32941 ;
  assign y9949 = n32945 ;
  assign y9950 = ~n32947 ;
  assign y9951 = ~n32951 ;
  assign y9952 = ~n32953 ;
  assign y9953 = ~n32955 ;
  assign y9954 = ~1'b0 ;
  assign y9955 = n32958 ;
  assign y9956 = ~n32959 ;
  assign y9957 = ~n32960 ;
  assign y9958 = ~n32962 ;
  assign y9959 = n32965 ;
  assign y9960 = n32968 ;
  assign y9961 = ~n32969 ;
  assign y9962 = ~n32976 ;
  assign y9963 = ~n32977 ;
  assign y9964 = n32978 ;
  assign y9965 = ~n32987 ;
  assign y9966 = n1544 ;
  assign y9967 = ~n32991 ;
  assign y9968 = ~n32992 ;
  assign y9969 = n32995 ;
  assign y9970 = ~n33001 ;
  assign y9971 = n33007 ;
  assign y9972 = ~1'b0 ;
  assign y9973 = ~n33012 ;
  assign y9974 = ~n33017 ;
  assign y9975 = ~n33022 ;
  assign y9976 = n33027 ;
  assign y9977 = n33028 ;
  assign y9978 = ~n33031 ;
  assign y9979 = n33035 ;
  assign y9980 = n33040 ;
  assign y9981 = n33042 ;
  assign y9982 = ~1'b0 ;
  assign y9983 = ~n33048 ;
  assign y9984 = ~n33050 ;
  assign y9985 = n33051 ;
  assign y9986 = ~n33059 ;
  assign y9987 = ~1'b0 ;
  assign y9988 = n33064 ;
  assign y9989 = ~n33065 ;
  assign y9990 = n33068 ;
  assign y9991 = n33069 ;
  assign y9992 = ~n33072 ;
  assign y9993 = ~1'b0 ;
  assign y9994 = n33076 ;
  assign y9995 = n33077 ;
  assign y9996 = n33080 ;
  assign y9997 = ~n33081 ;
  assign y9998 = ~1'b0 ;
  assign y9999 = ~n33085 ;
  assign y10000 = ~n33087 ;
  assign y10001 = 1'b0 ;
  assign y10002 = n33090 ;
  assign y10003 = ~n33091 ;
  assign y10004 = ~n33101 ;
  assign y10005 = n33102 ;
  assign y10006 = ~n33105 ;
  assign y10007 = n33107 ;
  assign y10008 = n33108 ;
  assign y10009 = n22612 ;
  assign y10010 = n33118 ;
  assign y10011 = 1'b0 ;
  assign y10012 = ~n33120 ;
  assign y10013 = ~1'b0 ;
  assign y10014 = ~1'b0 ;
  assign y10015 = ~1'b0 ;
  assign y10016 = n33126 ;
  assign y10017 = n33131 ;
  assign y10018 = ~n33133 ;
  assign y10019 = ~n33134 ;
  assign y10020 = n33136 ;
  assign y10021 = ~1'b0 ;
  assign y10022 = ~1'b0 ;
  assign y10023 = n33142 ;
  assign y10024 = ~1'b0 ;
  assign y10025 = ~n33145 ;
  assign y10026 = n33148 ;
  assign y10027 = n33150 ;
  assign y10028 = n21724 ;
  assign y10029 = ~1'b0 ;
  assign y10030 = n33151 ;
  assign y10031 = ~1'b0 ;
  assign y10032 = ~n33156 ;
  assign y10033 = n33158 ;
  assign y10034 = n33159 ;
  assign y10035 = n33160 ;
  assign y10036 = n33163 ;
  assign y10037 = n33165 ;
  assign y10038 = ~n33169 ;
  assign y10039 = ~1'b0 ;
  assign y10040 = ~n33172 ;
  assign y10041 = n33175 ;
  assign y10042 = ~n33178 ;
  assign y10043 = n33180 ;
  assign y10044 = ~n33181 ;
  assign y10045 = ~1'b0 ;
  assign y10046 = ~1'b0 ;
  assign y10047 = n33182 ;
  assign y10048 = ~n33186 ;
  assign y10049 = ~1'b0 ;
  assign y10050 = n33190 ;
  assign y10051 = ~n33191 ;
  assign y10052 = ~n33192 ;
  assign y10053 = ~n33193 ;
  assign y10054 = n6584 ;
  assign y10055 = n33197 ;
  assign y10056 = n33200 ;
  assign y10057 = ~n33202 ;
  assign y10058 = ~n33203 ;
  assign y10059 = n33204 ;
  assign y10060 = ~n33209 ;
  assign y10061 = ~n33216 ;
  assign y10062 = n33220 ;
  assign y10063 = ~n33224 ;
  assign y10064 = n33225 ;
  assign y10065 = n33227 ;
  assign y10066 = n33230 ;
  assign y10067 = ~n33234 ;
  assign y10068 = ~1'b0 ;
  assign y10069 = ~n33241 ;
  assign y10070 = n33243 ;
  assign y10071 = n33245 ;
  assign y10072 = ~n33247 ;
  assign y10073 = ~n33248 ;
  assign y10074 = ~n33250 ;
  assign y10075 = ~n33253 ;
  assign y10076 = ~1'b0 ;
  assign y10077 = ~1'b0 ;
  assign y10078 = ~1'b0 ;
  assign y10079 = n33257 ;
  assign y10080 = n33258 ;
  assign y10081 = n33260 ;
  assign y10082 = ~n33263 ;
  assign y10083 = n33264 ;
  assign y10084 = ~1'b0 ;
  assign y10085 = ~n33266 ;
  assign y10086 = ~1'b0 ;
  assign y10087 = ~n33267 ;
  assign y10088 = n13983 ;
  assign y10089 = ~n33273 ;
  assign y10090 = n33278 ;
  assign y10091 = n33280 ;
  assign y10092 = ~1'b0 ;
  assign y10093 = ~n33282 ;
  assign y10094 = ~1'b0 ;
  assign y10095 = ~n33289 ;
  assign y10096 = n33293 ;
  assign y10097 = ~n33297 ;
  assign y10098 = ~n33298 ;
  assign y10099 = ~n33299 ;
  assign y10100 = ~1'b0 ;
  assign y10101 = ~n33306 ;
  assign y10102 = ~1'b0 ;
  assign y10103 = ~n33307 ;
  assign y10104 = ~n33309 ;
  assign y10105 = n33310 ;
  assign y10106 = n33311 ;
  assign y10107 = ~1'b0 ;
  assign y10108 = ~1'b0 ;
  assign y10109 = ~n33318 ;
  assign y10110 = n5809 ;
  assign y10111 = ~n33320 ;
  assign y10112 = n33321 ;
  assign y10113 = ~n33325 ;
  assign y10114 = ~n33327 ;
  assign y10115 = ~n33329 ;
  assign y10116 = n33331 ;
  assign y10117 = ~n33332 ;
  assign y10118 = ~n33336 ;
  assign y10119 = n33342 ;
  assign y10120 = ~n33343 ;
  assign y10121 = ~n33347 ;
  assign y10122 = n33348 ;
  assign y10123 = n33355 ;
  assign y10124 = n33359 ;
  assign y10125 = n33366 ;
  assign y10126 = ~n33369 ;
  assign y10127 = ~1'b0 ;
  assign y10128 = n33374 ;
  assign y10129 = n33375 ;
  assign y10130 = n33376 ;
  assign y10131 = n33378 ;
  assign y10132 = n33393 ;
  assign y10133 = n33397 ;
  assign y10134 = ~1'b0 ;
  assign y10135 = n33399 ;
  assign y10136 = ~n33402 ;
  assign y10137 = ~n33405 ;
  assign y10138 = n33406 ;
  assign y10139 = ~n33418 ;
  assign y10140 = n33419 ;
  assign y10141 = n33422 ;
  assign y10142 = 1'b0 ;
  assign y10143 = n33429 ;
  assign y10144 = n33430 ;
  assign y10145 = n33435 ;
  assign y10146 = ~1'b0 ;
  assign y10147 = ~n33440 ;
  assign y10148 = ~n33443 ;
  assign y10149 = ~n33444 ;
  assign y10150 = ~n33445 ;
  assign y10151 = n33446 ;
  assign y10152 = n33447 ;
  assign y10153 = ~n33453 ;
  assign y10154 = n33455 ;
  assign y10155 = ~n33460 ;
  assign y10156 = n33461 ;
  assign y10157 = n33465 ;
  assign y10158 = ~1'b0 ;
  assign y10159 = n33466 ;
  assign y10160 = ~n33467 ;
  assign y10161 = ~n33468 ;
  assign y10162 = ~n33471 ;
  assign y10163 = ~1'b0 ;
  assign y10164 = ~1'b0 ;
  assign y10165 = ~n33476 ;
  assign y10166 = ~n33477 ;
  assign y10167 = n33478 ;
  assign y10168 = n33484 ;
  assign y10169 = ~1'b0 ;
  assign y10170 = ~1'b0 ;
  assign y10171 = n33493 ;
  assign y10172 = ~n33494 ;
  assign y10173 = n33495 ;
  assign y10174 = ~n33499 ;
  assign y10175 = ~n33501 ;
  assign y10176 = n33502 ;
  assign y10177 = ~n32805 ;
  assign y10178 = ~1'b0 ;
  assign y10179 = ~1'b0 ;
  assign y10180 = n33504 ;
  assign y10181 = ~1'b0 ;
  assign y10182 = n33512 ;
  assign y10183 = n9736 ;
  assign y10184 = ~n31748 ;
  assign y10185 = n33516 ;
  assign y10186 = n33517 ;
  assign y10187 = ~1'b0 ;
  assign y10188 = n33518 ;
  assign y10189 = ~n33521 ;
  assign y10190 = ~n33523 ;
  assign y10191 = n33526 ;
  assign y10192 = ~n33528 ;
  assign y10193 = ~n33530 ;
  assign y10194 = ~n33531 ;
  assign y10195 = n33536 ;
  assign y10196 = n33538 ;
  assign y10197 = ~n33542 ;
  assign y10198 = n33545 ;
  assign y10199 = ~n33548 ;
  assign y10200 = n33549 ;
  assign y10201 = n33554 ;
  assign y10202 = n33556 ;
  assign y10203 = ~n33557 ;
  assign y10204 = ~1'b0 ;
  assign y10205 = ~1'b0 ;
  assign y10206 = n33559 ;
  assign y10207 = ~1'b0 ;
  assign y10208 = ~n33562 ;
  assign y10209 = n33563 ;
  assign y10210 = ~n3070 ;
  assign y10211 = ~n33565 ;
  assign y10212 = ~1'b0 ;
  assign y10213 = n33568 ;
  assign y10214 = ~n33571 ;
  assign y10215 = n33574 ;
  assign y10216 = n33577 ;
  assign y10217 = ~1'b0 ;
  assign y10218 = ~n33579 ;
  assign y10219 = ~n33583 ;
  assign y10220 = ~n33586 ;
  assign y10221 = n33592 ;
  assign y10222 = n33594 ;
  assign y10223 = ~n33596 ;
  assign y10224 = ~1'b0 ;
  assign y10225 = n33599 ;
  assign y10226 = n33601 ;
  assign y10227 = ~n33602 ;
  assign y10228 = ~n33603 ;
  assign y10229 = ~1'b0 ;
  assign y10230 = ~1'b0 ;
  assign y10231 = ~1'b0 ;
  assign y10232 = ~n33605 ;
  assign y10233 = n33607 ;
  assign y10234 = n33612 ;
  assign y10235 = ~n33616 ;
  assign y10236 = ~n33617 ;
  assign y10237 = ~n33618 ;
  assign y10238 = ~n33622 ;
  assign y10239 = ~n33626 ;
  assign y10240 = ~n33628 ;
  assign y10241 = n33630 ;
  assign y10242 = n33631 ;
  assign y10243 = ~n33632 ;
  assign y10244 = n33633 ;
  assign y10245 = ~n33639 ;
  assign y10246 = n33641 ;
  assign y10247 = n33648 ;
  assign y10248 = ~n33649 ;
  assign y10249 = n33652 ;
  assign y10250 = n33654 ;
  assign y10251 = n33659 ;
  assign y10252 = ~n33661 ;
  assign y10253 = ~n33662 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = n33666 ;
  assign y10256 = ~n33667 ;
  assign y10257 = n33672 ;
  assign y10258 = ~n33676 ;
  assign y10259 = n33679 ;
  assign y10260 = ~n33684 ;
  assign y10261 = ~n33690 ;
  assign y10262 = ~n33693 ;
  assign y10263 = ~n33699 ;
  assign y10264 = ~n33701 ;
  assign y10265 = n33705 ;
  assign y10266 = ~n33706 ;
  assign y10267 = n33708 ;
  assign y10268 = n33709 ;
  assign y10269 = n33712 ;
  assign y10270 = ~n33713 ;
  assign y10271 = n33714 ;
  assign y10272 = ~n33717 ;
  assign y10273 = n33718 ;
  assign y10274 = ~n33719 ;
  assign y10275 = n33720 ;
  assign y10276 = n33723 ;
  assign y10277 = ~n33724 ;
  assign y10278 = n33725 ;
  assign y10279 = ~1'b0 ;
  assign y10280 = ~n33727 ;
  assign y10281 = ~1'b0 ;
  assign y10282 = n33731 ;
  assign y10283 = ~n33732 ;
  assign y10284 = ~n33734 ;
  assign y10285 = ~n33739 ;
  assign y10286 = ~n33742 ;
  assign y10287 = ~n33745 ;
  assign y10288 = ~n33752 ;
  assign y10289 = n33756 ;
  assign y10290 = ~n33759 ;
  assign y10291 = ~n33762 ;
  assign y10292 = ~n33764 ;
  assign y10293 = ~n33768 ;
  assign y10294 = n33770 ;
  assign y10295 = ~1'b0 ;
  assign y10296 = n33774 ;
  assign y10297 = ~1'b0 ;
  assign y10298 = ~n33776 ;
  assign y10299 = ~n33778 ;
  assign y10300 = ~n33779 ;
  assign y10301 = n33780 ;
  assign y10302 = ~1'b0 ;
  assign y10303 = n17877 ;
  assign y10304 = ~n33781 ;
  assign y10305 = ~n33784 ;
  assign y10306 = n33789 ;
  assign y10307 = n33796 ;
  assign y10308 = ~n33798 ;
  assign y10309 = ~n33799 ;
  assign y10310 = ~n33803 ;
  assign y10311 = n33805 ;
  assign y10312 = ~n33807 ;
  assign y10313 = n33808 ;
  assign y10314 = n33814 ;
  assign y10315 = ~n33817 ;
  assign y10316 = ~n33821 ;
  assign y10317 = 1'b0 ;
  assign y10318 = ~1'b0 ;
  assign y10319 = n33827 ;
  assign y10320 = n33829 ;
  assign y10321 = ~n33830 ;
  assign y10322 = n33832 ;
  assign y10323 = n33833 ;
  assign y10324 = ~n33834 ;
  assign y10325 = ~n33839 ;
  assign y10326 = ~n33841 ;
  assign y10327 = n33845 ;
  assign y10328 = ~n33855 ;
  assign y10329 = n33860 ;
  assign y10330 = n5617 ;
  assign y10331 = ~n33861 ;
  assign y10332 = ~1'b0 ;
  assign y10333 = ~n33864 ;
  assign y10334 = ~n33869 ;
  assign y10335 = n33872 ;
  assign y10336 = ~n33875 ;
  assign y10337 = n33876 ;
  assign y10338 = ~n33879 ;
  assign y10339 = n33882 ;
  assign y10340 = n33890 ;
  assign y10341 = ~n33891 ;
  assign y10342 = ~n33893 ;
  assign y10343 = ~n33894 ;
  assign y10344 = n33897 ;
  assign y10345 = ~1'b0 ;
  assign y10346 = n33902 ;
  assign y10347 = ~1'b0 ;
  assign y10348 = n33904 ;
  assign y10349 = n33905 ;
  assign y10350 = ~n33906 ;
  assign y10351 = n33909 ;
  assign y10352 = ~n33910 ;
  assign y10353 = ~n33912 ;
  assign y10354 = ~n33917 ;
  assign y10355 = ~n33918 ;
  assign y10356 = n33922 ;
  assign y10357 = ~n33923 ;
  assign y10358 = n33925 ;
  assign y10359 = n5949 ;
  assign y10360 = ~1'b0 ;
  assign y10361 = n33927 ;
  assign y10362 = ~n33931 ;
  assign y10363 = ~n33934 ;
  assign y10364 = n33935 ;
  assign y10365 = ~n33943 ;
  assign y10366 = ~1'b0 ;
  assign y10367 = n33944 ;
  assign y10368 = n33947 ;
  assign y10369 = ~n33948 ;
  assign y10370 = n33951 ;
  assign y10371 = ~n33956 ;
  assign y10372 = ~n33961 ;
  assign y10373 = ~n33962 ;
  assign y10374 = ~1'b0 ;
  assign y10375 = ~n33964 ;
  assign y10376 = n33968 ;
  assign y10377 = ~n33972 ;
  assign y10378 = ~1'b0 ;
  assign y10379 = n33976 ;
  assign y10380 = n33979 ;
  assign y10381 = n33982 ;
  assign y10382 = ~n33989 ;
  assign y10383 = n33991 ;
  assign y10384 = ~n33997 ;
  assign y10385 = n33998 ;
  assign y10386 = n34001 ;
  assign y10387 = ~1'b0 ;
  assign y10388 = n34003 ;
  assign y10389 = ~n34005 ;
  assign y10390 = n34016 ;
  assign y10391 = n34019 ;
  assign y10392 = n34020 ;
  assign y10393 = n34021 ;
  assign y10394 = n34022 ;
  assign y10395 = ~n34024 ;
  assign y10396 = n34031 ;
  assign y10397 = ~n34036 ;
  assign y10398 = ~n34039 ;
  assign y10399 = n34040 ;
  assign y10400 = ~n34047 ;
  assign y10401 = n34049 ;
  assign y10402 = ~1'b0 ;
  assign y10403 = ~n34051 ;
  assign y10404 = ~n34052 ;
  assign y10405 = ~n34054 ;
  assign y10406 = ~n34057 ;
  assign y10407 = n34059 ;
  assign y10408 = ~n34061 ;
  assign y10409 = ~n34063 ;
  assign y10410 = ~n34065 ;
  assign y10411 = n34070 ;
  assign y10412 = n34073 ;
  assign y10413 = ~n34076 ;
  assign y10414 = ~n34082 ;
  assign y10415 = ~n34083 ;
  assign y10416 = ~n34084 ;
  assign y10417 = ~n34090 ;
  assign y10418 = n34094 ;
  assign y10419 = ~1'b0 ;
  assign y10420 = ~n34095 ;
  assign y10421 = ~n34100 ;
  assign y10422 = n34102 ;
  assign y10423 = ~n34105 ;
  assign y10424 = ~n34108 ;
  assign y10425 = ~n34109 ;
  assign y10426 = n34113 ;
  assign y10427 = n34117 ;
  assign y10428 = ~n34118 ;
  assign y10429 = n34119 ;
  assign y10430 = ~n34127 ;
  assign y10431 = ~n34132 ;
  assign y10432 = ~1'b0 ;
  assign y10433 = n34137 ;
  assign y10434 = ~n34138 ;
  assign y10435 = ~n34139 ;
  assign y10436 = n34140 ;
  assign y10437 = n34142 ;
  assign y10438 = n34147 ;
  assign y10439 = ~1'b0 ;
  assign y10440 = ~1'b0 ;
  assign y10441 = n34153 ;
  assign y10442 = n34155 ;
  assign y10443 = ~n34160 ;
  assign y10444 = ~n34162 ;
  assign y10445 = ~1'b0 ;
  assign y10446 = ~1'b0 ;
  assign y10447 = ~n34169 ;
  assign y10448 = n34170 ;
  assign y10449 = ~n5754 ;
  assign y10450 = ~n34171 ;
  assign y10451 = ~1'b0 ;
  assign y10452 = n34174 ;
  assign y10453 = n34183 ;
  assign y10454 = n34185 ;
  assign y10455 = n34190 ;
  assign y10456 = ~1'b0 ;
  assign y10457 = n34191 ;
  assign y10458 = ~n34196 ;
  assign y10459 = n34198 ;
  assign y10460 = n34201 ;
  assign y10461 = n34202 ;
  assign y10462 = ~1'b0 ;
  assign y10463 = n34204 ;
  assign y10464 = n26440 ;
  assign y10465 = ~n13811 ;
  assign y10466 = n34206 ;
  assign y10467 = ~1'b0 ;
  assign y10468 = ~1'b0 ;
  assign y10469 = ~n34210 ;
  assign y10470 = n34211 ;
  assign y10471 = n34212 ;
  assign y10472 = ~1'b0 ;
  assign y10473 = ~1'b0 ;
  assign y10474 = ~n34213 ;
  assign y10475 = ~n34214 ;
  assign y10476 = n34219 ;
  assign y10477 = n34222 ;
  assign y10478 = ~n34223 ;
  assign y10479 = ~n34224 ;
  assign y10480 = n34225 ;
  assign y10481 = ~n34228 ;
  assign y10482 = n34240 ;
  assign y10483 = ~n34248 ;
  assign y10484 = ~n34249 ;
  assign y10485 = n34251 ;
  assign y10486 = ~1'b0 ;
  assign y10487 = ~1'b0 ;
  assign y10488 = n34252 ;
  assign y10489 = n34253 ;
  assign y10490 = n34254 ;
  assign y10491 = n34259 ;
  assign y10492 = n34261 ;
  assign y10493 = ~1'b0 ;
  assign y10494 = ~n34264 ;
  assign y10495 = ~1'b0 ;
  assign y10496 = ~n34269 ;
  assign y10497 = n34273 ;
  assign y10498 = n34277 ;
  assign y10499 = ~n34280 ;
  assign y10500 = ~n34282 ;
  assign y10501 = n12596 ;
  assign y10502 = ~n34284 ;
  assign y10503 = ~n34286 ;
  assign y10504 = ~n34288 ;
  assign y10505 = ~n34291 ;
  assign y10506 = ~n21573 ;
  assign y10507 = ~n34292 ;
  assign y10508 = n34294 ;
  assign y10509 = ~1'b0 ;
  assign y10510 = ~1'b0 ;
  assign y10511 = ~n34299 ;
  assign y10512 = n34301 ;
  assign y10513 = n34305 ;
  assign y10514 = n34307 ;
  assign y10515 = n34314 ;
  assign y10516 = ~1'b0 ;
  assign y10517 = n34316 ;
  assign y10518 = ~n34319 ;
  assign y10519 = n34320 ;
  assign y10520 = ~n34324 ;
  assign y10521 = n34327 ;
  assign y10522 = ~1'b0 ;
  assign y10523 = ~n34328 ;
  assign y10524 = ~n34331 ;
  assign y10525 = ~n34337 ;
  assign y10526 = n34339 ;
  assign y10527 = ~n34341 ;
  assign y10528 = ~n34342 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = ~1'b0 ;
  assign y10531 = ~1'b0 ;
  assign y10532 = ~1'b0 ;
  assign y10533 = ~n34344 ;
  assign y10534 = n34347 ;
  assign y10535 = ~n34348 ;
  assign y10536 = ~n34350 ;
  assign y10537 = ~1'b0 ;
  assign y10538 = ~n34352 ;
  assign y10539 = n34358 ;
  assign y10540 = ~n34359 ;
  assign y10541 = n34361 ;
  assign y10542 = ~n34362 ;
  assign y10543 = ~n34363 ;
  assign y10544 = n34365 ;
  assign y10545 = ~1'b0 ;
  assign y10546 = ~1'b0 ;
  assign y10547 = ~n34366 ;
  assign y10548 = n34369 ;
  assign y10549 = n34371 ;
  assign y10550 = ~n34373 ;
  assign y10551 = n34375 ;
  assign y10552 = n34379 ;
  assign y10553 = ~n34380 ;
  assign y10554 = n34385 ;
  assign y10555 = n34388 ;
  assign y10556 = n34390 ;
  assign y10557 = ~n34396 ;
  assign y10558 = ~n34397 ;
  assign y10559 = ~n34399 ;
  assign y10560 = ~n34401 ;
  assign y10561 = n34403 ;
  assign y10562 = n34406 ;
  assign y10563 = ~n34407 ;
  assign y10564 = n34413 ;
  assign y10565 = n34415 ;
  assign y10566 = n34426 ;
  assign y10567 = n34428 ;
  assign y10568 = n34430 ;
  assign y10569 = n34434 ;
  assign y10570 = ~n34435 ;
  assign y10571 = ~n34440 ;
  assign y10572 = ~n18776 ;
  assign y10573 = 1'b0 ;
  assign y10574 = ~n34444 ;
  assign y10575 = ~n34446 ;
  assign y10576 = n34449 ;
  assign y10577 = ~1'b0 ;
  assign y10578 = ~n34455 ;
  assign y10579 = ~n34461 ;
  assign y10580 = ~n34463 ;
  assign y10581 = ~n34464 ;
  assign y10582 = ~n34474 ;
  assign y10583 = ~n34476 ;
  assign y10584 = ~1'b0 ;
  assign y10585 = ~n34483 ;
  assign y10586 = n34485 ;
  assign y10587 = n34488 ;
  assign y10588 = n34490 ;
  assign y10589 = n34494 ;
  assign y10590 = ~n34498 ;
  assign y10591 = n34499 ;
  assign y10592 = ~n34502 ;
  assign y10593 = ~n34516 ;
  assign y10594 = ~n34521 ;
  assign y10595 = n34526 ;
  assign y10596 = ~1'b0 ;
  assign y10597 = ~n34531 ;
  assign y10598 = ~n34532 ;
  assign y10599 = ~n13505 ;
  assign y10600 = n7118 ;
  assign y10601 = n34544 ;
  assign y10602 = ~n34547 ;
  assign y10603 = n34549 ;
  assign y10604 = n34551 ;
  assign y10605 = n34552 ;
  assign y10606 = n34554 ;
  assign y10607 = ~n5994 ;
  assign y10608 = n34555 ;
  assign y10609 = ~1'b0 ;
  assign y10610 = ~n34556 ;
  assign y10611 = ~1'b0 ;
  assign y10612 = ~1'b0 ;
  assign y10613 = n34557 ;
  assign y10614 = n34561 ;
  assign y10615 = n34563 ;
  assign y10616 = ~n34566 ;
  assign y10617 = ~n34569 ;
  assign y10618 = n34575 ;
  assign y10619 = ~1'b0 ;
  assign y10620 = ~n34577 ;
  assign y10621 = n34578 ;
  assign y10622 = ~n34582 ;
  assign y10623 = n34584 ;
  assign y10624 = ~1'b0 ;
  assign y10625 = n34585 ;
  assign y10626 = n34587 ;
  assign y10627 = n34588 ;
  assign y10628 = ~n34593 ;
  assign y10629 = ~n34596 ;
  assign y10630 = ~n34597 ;
  assign y10631 = ~n34603 ;
  assign y10632 = ~n34608 ;
  assign y10633 = n34609 ;
  assign y10634 = n34611 ;
  assign y10635 = n34618 ;
  assign y10636 = ~n34621 ;
  assign y10637 = n34623 ;
  assign y10638 = ~1'b0 ;
  assign y10639 = n34628 ;
  assign y10640 = n34629 ;
  assign y10641 = n34631 ;
  assign y10642 = ~n34632 ;
  assign y10643 = ~n34634 ;
  assign y10644 = ~n34635 ;
  assign y10645 = n34641 ;
  assign y10646 = n34643 ;
  assign y10647 = ~n34650 ;
  assign y10648 = ~n34651 ;
  assign y10649 = n34657 ;
  assign y10650 = n34660 ;
  assign y10651 = n34661 ;
  assign y10652 = ~n34664 ;
  assign y10653 = ~n34666 ;
  assign y10654 = n34667 ;
  assign y10655 = ~1'b0 ;
  assign y10656 = ~n34671 ;
  assign y10657 = ~1'b0 ;
  assign y10658 = ~n34678 ;
  assign y10659 = ~n34679 ;
  assign y10660 = n34684 ;
  assign y10661 = n34686 ;
  assign y10662 = n34688 ;
  assign y10663 = n34690 ;
  assign y10664 = n34692 ;
  assign y10665 = n34693 ;
  assign y10666 = n34696 ;
  assign y10667 = ~n34699 ;
  assign y10668 = ~n34701 ;
  assign y10669 = n34704 ;
  assign y10670 = ~n4431 ;
  assign y10671 = ~n34705 ;
  assign y10672 = ~n34710 ;
  assign y10673 = ~n34712 ;
  assign y10674 = ~n34714 ;
  assign y10675 = n34717 ;
  assign y10676 = ~1'b0 ;
  assign y10677 = ~n34718 ;
  assign y10678 = ~n34719 ;
  assign y10679 = n34721 ;
  assign y10680 = n34722 ;
  assign y10681 = n34723 ;
  assign y10682 = ~n34725 ;
  assign y10683 = n34727 ;
  assign y10684 = n34728 ;
  assign y10685 = ~n34730 ;
  assign y10686 = n34732 ;
  assign y10687 = ~n34735 ;
  assign y10688 = ~n34736 ;
  assign y10689 = n34738 ;
  assign y10690 = ~1'b0 ;
  assign y10691 = n34739 ;
  assign y10692 = ~n34741 ;
  assign y10693 = n34742 ;
  assign y10694 = ~n34747 ;
  assign y10695 = ~1'b0 ;
  assign y10696 = n34755 ;
  assign y10697 = n34757 ;
  assign y10698 = ~n34759 ;
  assign y10699 = ~n34761 ;
  assign y10700 = n34762 ;
  assign y10701 = n34763 ;
  assign y10702 = n34767 ;
  assign y10703 = ~n34769 ;
  assign y10704 = n34770 ;
  assign y10705 = ~n34774 ;
  assign y10706 = ~n34775 ;
  assign y10707 = ~n34776 ;
  assign y10708 = 1'b0 ;
  assign y10709 = n34782 ;
  assign y10710 = ~n34789 ;
  assign y10711 = n34792 ;
  assign y10712 = n34794 ;
  assign y10713 = n34795 ;
  assign y10714 = ~n34799 ;
  assign y10715 = n34800 ;
  assign y10716 = ~n34803 ;
  assign y10717 = ~1'b0 ;
  assign y10718 = ~1'b0 ;
  assign y10719 = ~n34809 ;
  assign y10720 = n34815 ;
  assign y10721 = ~n388 ;
  assign y10722 = n34816 ;
  assign y10723 = ~n34819 ;
  assign y10724 = n34821 ;
  assign y10725 = n34823 ;
  assign y10726 = n34824 ;
  assign y10727 = ~n34826 ;
  assign y10728 = n34827 ;
  assign y10729 = n34831 ;
  assign y10730 = n34836 ;
  assign y10731 = n34839 ;
  assign y10732 = n34840 ;
  assign y10733 = ~n34849 ;
  assign y10734 = ~n34854 ;
  assign y10735 = ~1'b0 ;
  assign y10736 = ~n34857 ;
  assign y10737 = ~n34858 ;
  assign y10738 = ~n34863 ;
  assign y10739 = n34864 ;
  assign y10740 = n34866 ;
  assign y10741 = n34868 ;
  assign y10742 = ~n34870 ;
  assign y10743 = ~n34871 ;
  assign y10744 = ~1'b0 ;
  assign y10745 = n34873 ;
  assign y10746 = n34877 ;
  assign y10747 = n34878 ;
  assign y10748 = ~n34888 ;
  assign y10749 = ~n34889 ;
  assign y10750 = n34893 ;
  assign y10751 = ~n34896 ;
  assign y10752 = ~n34898 ;
  assign y10753 = n34902 ;
  assign y10754 = ~n34904 ;
  assign y10755 = n34905 ;
  assign y10756 = ~n34906 ;
  assign y10757 = ~n34907 ;
  assign y10758 = ~1'b0 ;
  assign y10759 = n34910 ;
  assign y10760 = ~n34912 ;
  assign y10761 = ~n34913 ;
  assign y10762 = ~n34915 ;
  assign y10763 = n34918 ;
  assign y10764 = ~n34921 ;
  assign y10765 = ~n34924 ;
  assign y10766 = n34926 ;
  assign y10767 = ~n34929 ;
  assign y10768 = n34939 ;
  assign y10769 = ~n34945 ;
  assign y10770 = ~n34946 ;
  assign y10771 = ~n34948 ;
  assign y10772 = n34950 ;
  assign y10773 = n34951 ;
  assign y10774 = n34953 ;
  assign y10775 = ~n34956 ;
  assign y10776 = ~n34957 ;
  assign y10777 = n34964 ;
  assign y10778 = ~n34967 ;
  assign y10779 = n34968 ;
  assign y10780 = ~n34971 ;
  assign y10781 = ~n34976 ;
  assign y10782 = n34979 ;
  assign y10783 = n4424 ;
  assign y10784 = n34980 ;
  assign y10785 = n34986 ;
  assign y10786 = ~n34990 ;
  assign y10787 = n34995 ;
  assign y10788 = ~n34997 ;
  assign y10789 = n34998 ;
  assign y10790 = n35001 ;
  assign y10791 = n35008 ;
  assign y10792 = ~1'b0 ;
  assign y10793 = ~n35012 ;
  assign y10794 = ~n35014 ;
  assign y10795 = ~n35017 ;
  assign y10796 = ~1'b0 ;
  assign y10797 = n35021 ;
  assign y10798 = n35026 ;
  assign y10799 = ~n35029 ;
  assign y10800 = n35031 ;
  assign y10801 = n35034 ;
  assign y10802 = ~n35038 ;
  assign y10803 = n35044 ;
  assign y10804 = n35051 ;
  assign y10805 = n35054 ;
  assign y10806 = ~n35056 ;
  assign y10807 = n35057 ;
  assign y10808 = ~n35059 ;
  assign y10809 = n35060 ;
  assign y10810 = ~n35064 ;
  assign y10811 = n35065 ;
  assign y10812 = n35068 ;
  assign y10813 = ~n35072 ;
  assign y10814 = ~1'b0 ;
  assign y10815 = ~n35074 ;
  assign y10816 = ~n35077 ;
  assign y10817 = ~n17696 ;
  assign y10818 = ~n35079 ;
  assign y10819 = ~n35080 ;
  assign y10820 = ~n35082 ;
  assign y10821 = n35083 ;
  assign y10822 = ~n35090 ;
  assign y10823 = ~n35103 ;
  assign y10824 = ~n35105 ;
  assign y10825 = n35110 ;
  assign y10826 = ~n35116 ;
  assign y10827 = ~n35118 ;
  assign y10828 = ~1'b0 ;
  assign y10829 = ~n35119 ;
  assign y10830 = 1'b0 ;
  assign y10831 = n35123 ;
  assign y10832 = ~n35125 ;
  assign y10833 = ~n35128 ;
  assign y10834 = n35130 ;
  assign y10835 = ~n35132 ;
  assign y10836 = ~n35136 ;
  assign y10837 = ~n35138 ;
  assign y10838 = ~n35139 ;
  assign y10839 = ~n35145 ;
  assign y10840 = n35147 ;
  assign y10841 = n35151 ;
  assign y10842 = ~n35152 ;
  assign y10843 = ~n35153 ;
  assign y10844 = n35160 ;
  assign y10845 = ~n35164 ;
  assign y10846 = ~n35165 ;
  assign y10847 = n35168 ;
  assign y10848 = ~n35171 ;
  assign y10849 = ~1'b0 ;
  assign y10850 = ~n35173 ;
  assign y10851 = ~1'b0 ;
  assign y10852 = n35174 ;
  assign y10853 = n35177 ;
  assign y10854 = ~n35178 ;
  assign y10855 = ~n35179 ;
  assign y10856 = ~1'b0 ;
  assign y10857 = n35181 ;
  assign y10858 = ~1'b0 ;
  assign y10859 = ~n35182 ;
  assign y10860 = ~n35183 ;
  assign y10861 = n35184 ;
  assign y10862 = n35185 ;
  assign y10863 = n35191 ;
  assign y10864 = n35193 ;
  assign y10865 = n35195 ;
  assign y10866 = ~1'b0 ;
  assign y10867 = ~1'b0 ;
  assign y10868 = n35197 ;
  assign y10869 = ~1'b0 ;
  assign y10870 = n35201 ;
  assign y10871 = ~n35206 ;
  assign y10872 = ~n35207 ;
  assign y10873 = n35208 ;
  assign y10874 = n35209 ;
  assign y10875 = ~1'b0 ;
  assign y10876 = n35211 ;
  assign y10877 = n35218 ;
  assign y10878 = ~n35219 ;
  assign y10879 = n35224 ;
  assign y10880 = n35226 ;
  assign y10881 = ~n35229 ;
  assign y10882 = n35230 ;
  assign y10883 = ~1'b0 ;
  assign y10884 = ~n35233 ;
  assign y10885 = ~n35236 ;
  assign y10886 = n35240 ;
  assign y10887 = n35243 ;
  assign y10888 = n35244 ;
  assign y10889 = ~n35245 ;
  assign y10890 = ~n35247 ;
  assign y10891 = n35249 ;
  assign y10892 = n35254 ;
  assign y10893 = ~n35257 ;
  assign y10894 = n35260 ;
  assign y10895 = ~n35262 ;
  assign y10896 = ~n35263 ;
  assign y10897 = ~n35264 ;
  assign y10898 = ~n35265 ;
  assign y10899 = ~1'b0 ;
  assign y10900 = ~n35267 ;
  assign y10901 = n35271 ;
  assign y10902 = ~1'b0 ;
  assign y10903 = n35273 ;
  assign y10904 = ~n35274 ;
  assign y10905 = ~n35279 ;
  assign y10906 = ~n35282 ;
  assign y10907 = n35289 ;
  assign y10908 = n35290 ;
  assign y10909 = ~n35295 ;
  assign y10910 = ~n35296 ;
  assign y10911 = n35300 ;
  assign y10912 = n35302 ;
  assign y10913 = ~n35303 ;
  assign y10914 = n35304 ;
  assign y10915 = n35307 ;
  assign y10916 = ~n35310 ;
  assign y10917 = n35315 ;
  assign y10918 = ~n35319 ;
  assign y10919 = n35334 ;
  assign y10920 = ~1'b0 ;
  assign y10921 = n35335 ;
  assign y10922 = ~n35339 ;
  assign y10923 = n35342 ;
  assign y10924 = n35345 ;
  assign y10925 = n35349 ;
  assign y10926 = ~1'b0 ;
  assign y10927 = n35353 ;
  assign y10928 = ~n35356 ;
  assign y10929 = ~1'b0 ;
  assign y10930 = ~n35357 ;
  assign y10931 = n35358 ;
  assign y10932 = n35361 ;
  assign y10933 = ~n35364 ;
  assign y10934 = ~n35366 ;
  assign y10935 = ~n35369 ;
  assign y10936 = ~n35371 ;
  assign y10937 = n35376 ;
  assign y10938 = ~n35381 ;
  assign y10939 = ~n35384 ;
  assign y10940 = n35388 ;
  assign y10941 = ~n35394 ;
  assign y10942 = ~1'b0 ;
  assign y10943 = n35395 ;
  assign y10944 = n35397 ;
  assign y10945 = ~1'b0 ;
  assign y10946 = ~1'b0 ;
  assign y10947 = ~n35401 ;
  assign y10948 = n35403 ;
  assign y10949 = n35407 ;
  assign y10950 = n35409 ;
  assign y10951 = ~n35410 ;
  assign y10952 = n35411 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = n35412 ;
  assign y10955 = ~1'b0 ;
  assign y10956 = n35416 ;
  assign y10957 = ~n35419 ;
  assign y10958 = ~n35420 ;
  assign y10959 = ~n35430 ;
  assign y10960 = n35431 ;
  assign y10961 = ~n35433 ;
  assign y10962 = ~n35436 ;
  assign y10963 = n35437 ;
  assign y10964 = n35443 ;
  assign y10965 = ~1'b0 ;
  assign y10966 = n35451 ;
  assign y10967 = ~n35454 ;
  assign y10968 = n35455 ;
  assign y10969 = ~n35456 ;
  assign y10970 = n35458 ;
  assign y10971 = ~n35463 ;
  assign y10972 = ~1'b0 ;
  assign y10973 = 1'b0 ;
  assign y10974 = n35465 ;
  assign y10975 = ~1'b0 ;
  assign y10976 = n35468 ;
  assign y10977 = ~n35469 ;
  assign y10978 = n35472 ;
  assign y10979 = ~n35475 ;
  assign y10980 = n35479 ;
  assign y10981 = ~n35491 ;
  assign y10982 = ~1'b0 ;
  assign y10983 = n35494 ;
  assign y10984 = n35496 ;
  assign y10985 = ~n35498 ;
  assign y10986 = ~n35503 ;
  assign y10987 = ~n35504 ;
  assign y10988 = ~1'b0 ;
  assign y10989 = n35505 ;
  assign y10990 = ~n35506 ;
  assign y10991 = ~n35507 ;
  assign y10992 = ~n35508 ;
  assign y10993 = ~n35509 ;
  assign y10994 = n35515 ;
  assign y10995 = ~1'b0 ;
  assign y10996 = n35524 ;
  assign y10997 = n35529 ;
  assign y10998 = ~n35530 ;
  assign y10999 = ~n35535 ;
  assign y11000 = ~n35536 ;
  assign y11001 = n35538 ;
  assign y11002 = ~n35543 ;
  assign y11003 = n35545 ;
  assign y11004 = ~n35553 ;
  assign y11005 = ~n35556 ;
  assign y11006 = n35558 ;
  assign y11007 = 1'b0 ;
  assign y11008 = n35559 ;
  assign y11009 = n35561 ;
  assign y11010 = ~n29446 ;
  assign y11011 = n35563 ;
  assign y11012 = ~n35564 ;
  assign y11013 = ~n35565 ;
  assign y11014 = ~n35567 ;
  assign y11015 = ~1'b0 ;
  assign y11016 = n35569 ;
  assign y11017 = n35570 ;
  assign y11018 = n35574 ;
  assign y11019 = n35579 ;
  assign y11020 = ~n8819 ;
  assign y11021 = ~n35583 ;
  assign y11022 = n35585 ;
  assign y11023 = n35586 ;
  assign y11024 = n35593 ;
  assign y11025 = n35594 ;
  assign y11026 = n35595 ;
  assign y11027 = ~1'b0 ;
  assign y11028 = ~n35600 ;
  assign y11029 = ~n35603 ;
  assign y11030 = ~n35605 ;
  assign y11031 = ~n35610 ;
  assign y11032 = n35620 ;
  assign y11033 = ~n35622 ;
  assign y11034 = ~1'b0 ;
  assign y11035 = ~n35623 ;
  assign y11036 = n35626 ;
  assign y11037 = ~n35628 ;
  assign y11038 = ~n35630 ;
  assign y11039 = n35632 ;
  assign y11040 = n35637 ;
  assign y11041 = n35640 ;
  assign y11042 = ~n35641 ;
  assign y11043 = n35646 ;
  assign y11044 = ~n35649 ;
  assign y11045 = ~n35650 ;
  assign y11046 = n35653 ;
  assign y11047 = ~n35655 ;
  assign y11048 = ~1'b0 ;
  assign y11049 = n35661 ;
  assign y11050 = n35663 ;
  assign y11051 = n35664 ;
  assign y11052 = n35665 ;
  assign y11053 = ~1'b0 ;
  assign y11054 = ~n35668 ;
  assign y11055 = ~1'b0 ;
  assign y11056 = ~n35671 ;
  assign y11057 = n35672 ;
  assign y11058 = ~n35674 ;
  assign y11059 = n35676 ;
  assign y11060 = ~n35677 ;
  assign y11061 = n35678 ;
  assign y11062 = ~n35682 ;
  assign y11063 = n35683 ;
  assign y11064 = ~n35685 ;
  assign y11065 = ~n35693 ;
  assign y11066 = ~n35695 ;
  assign y11067 = ~n35697 ;
  assign y11068 = ~n35702 ;
  assign y11069 = n35705 ;
  assign y11070 = n35707 ;
  assign y11071 = ~1'b0 ;
  assign y11072 = ~n35717 ;
  assign y11073 = n35725 ;
  assign y11074 = n35727 ;
  assign y11075 = ~n35728 ;
  assign y11076 = ~n35729 ;
  assign y11077 = ~n35730 ;
  assign y11078 = n35735 ;
  assign y11079 = ~n35737 ;
  assign y11080 = ~1'b0 ;
  assign y11081 = 1'b0 ;
  assign y11082 = ~1'b0 ;
  assign y11083 = ~n35740 ;
  assign y11084 = ~n35742 ;
  assign y11085 = n35743 ;
  assign y11086 = ~n35745 ;
  assign y11087 = n35753 ;
  assign y11088 = n35754 ;
  assign y11089 = n35758 ;
  assign y11090 = ~n35761 ;
  assign y11091 = n35762 ;
  assign y11092 = n35764 ;
  assign y11093 = ~n35765 ;
  assign y11094 = ~n35766 ;
  assign y11095 = n35767 ;
  assign y11096 = ~n35772 ;
  assign y11097 = ~n35774 ;
  assign y11098 = ~n35776 ;
  assign y11099 = n35779 ;
  assign y11100 = n35787 ;
  assign y11101 = ~n35788 ;
  assign y11102 = ~n35790 ;
  assign y11103 = ~n35794 ;
  assign y11104 = n35796 ;
  assign y11105 = n35798 ;
  assign y11106 = ~n35800 ;
  assign y11107 = ~n35803 ;
  assign y11108 = n35808 ;
  assign y11109 = n35809 ;
  assign y11110 = n35814 ;
  assign y11111 = n35815 ;
  assign y11112 = ~n35817 ;
  assign y11113 = n35825 ;
  assign y11114 = ~n35831 ;
  assign y11115 = n35834 ;
  assign y11116 = n35837 ;
  assign y11117 = ~n35842 ;
  assign y11118 = ~n35845 ;
  assign y11119 = n35856 ;
  assign y11120 = n35861 ;
  assign y11121 = ~1'b0 ;
  assign y11122 = n35863 ;
  assign y11123 = ~n35866 ;
  assign y11124 = ~n35869 ;
  assign y11125 = ~n35871 ;
  assign y11126 = n35875 ;
  assign y11127 = n35876 ;
  assign y11128 = ~n35878 ;
  assign y11129 = n35880 ;
  assign y11130 = ~n35884 ;
  assign y11131 = n35887 ;
  assign y11132 = n35888 ;
  assign y11133 = ~n35889 ;
  assign y11134 = ~n35890 ;
  assign y11135 = ~n35896 ;
  assign y11136 = ~n35899 ;
  assign y11137 = ~n35901 ;
  assign y11138 = ~1'b0 ;
  assign y11139 = n35903 ;
  assign y11140 = ~n35906 ;
  assign y11141 = ~n35911 ;
  assign y11142 = ~n35918 ;
  assign y11143 = n35928 ;
  assign y11144 = ~n35931 ;
  assign y11145 = n35934 ;
  assign y11146 = n35935 ;
  assign y11147 = n35940 ;
  assign y11148 = n35942 ;
  assign y11149 = n35943 ;
  assign y11150 = n35948 ;
  assign y11151 = n35949 ;
  assign y11152 = n35952 ;
  assign y11153 = ~1'b0 ;
  assign y11154 = n35956 ;
  assign y11155 = ~n35958 ;
  assign y11156 = ~n35962 ;
  assign y11157 = ~n35967 ;
  assign y11158 = ~n35969 ;
  assign y11159 = n35971 ;
  assign y11160 = ~n35973 ;
  assign y11161 = ~1'b0 ;
  assign y11162 = ~n35980 ;
  assign y11163 = n35981 ;
  assign y11164 = n35982 ;
  assign y11165 = ~n35989 ;
  assign y11166 = ~n35993 ;
  assign y11167 = n35997 ;
  assign y11168 = ~1'b0 ;
  assign y11169 = ~1'b0 ;
  assign y11170 = n36001 ;
  assign y11171 = ~n36003 ;
  assign y11172 = ~n36007 ;
  assign y11173 = ~n36010 ;
  assign y11174 = ~n36012 ;
  assign y11175 = n36018 ;
  assign y11176 = n36020 ;
  assign y11177 = ~1'b0 ;
  assign y11178 = ~1'b0 ;
  assign y11179 = ~n36021 ;
  assign y11180 = ~n36026 ;
  assign y11181 = ~n27837 ;
  assign y11182 = ~n36028 ;
  assign y11183 = n36030 ;
  assign y11184 = ~n36032 ;
  assign y11185 = ~1'b0 ;
  assign y11186 = ~1'b0 ;
  assign y11187 = ~n36034 ;
  assign y11188 = n36037 ;
  assign y11189 = n36040 ;
  assign y11190 = n36043 ;
  assign y11191 = n36044 ;
  assign y11192 = ~n36047 ;
  assign y11193 = n36052 ;
  assign y11194 = ~n36054 ;
  assign y11195 = n36057 ;
  assign y11196 = n36059 ;
  assign y11197 = ~n36061 ;
  assign y11198 = ~n36062 ;
  assign y11199 = n36066 ;
  assign y11200 = n36067 ;
  assign y11201 = ~n36069 ;
  assign y11202 = ~n36074 ;
  assign y11203 = n36080 ;
  assign y11204 = n36084 ;
  assign y11205 = ~1'b0 ;
  assign y11206 = ~n36091 ;
  assign y11207 = n36098 ;
  assign y11208 = ~n36104 ;
  assign y11209 = ~n36105 ;
  assign y11210 = ~n36109 ;
  assign y11211 = n36111 ;
  assign y11212 = ~n36115 ;
  assign y11213 = n36119 ;
  assign y11214 = ~1'b0 ;
  assign y11215 = ~n36120 ;
  assign y11216 = n36122 ;
  assign y11217 = n36123 ;
  assign y11218 = n36125 ;
  assign y11219 = ~n36129 ;
  assign y11220 = ~n36132 ;
  assign y11221 = n36134 ;
  assign y11222 = ~n36136 ;
  assign y11223 = ~1'b0 ;
  assign y11224 = ~n36144 ;
  assign y11225 = n36145 ;
  assign y11226 = n36146 ;
  assign y11227 = ~n36150 ;
  assign y11228 = n36155 ;
  assign y11229 = ~1'b0 ;
  assign y11230 = ~n36156 ;
  assign y11231 = ~n36157 ;
  assign y11232 = n36159 ;
  assign y11233 = ~n36163 ;
  assign y11234 = ~n36166 ;
  assign y11235 = n36171 ;
  assign y11236 = n36174 ;
  assign y11237 = ~n36178 ;
  assign y11238 = n36181 ;
  assign y11239 = ~n36185 ;
  assign y11240 = ~n36186 ;
  assign y11241 = n36188 ;
  assign y11242 = n36193 ;
  assign y11243 = n36195 ;
  assign y11244 = n36196 ;
  assign y11245 = n36202 ;
  assign y11246 = ~n36205 ;
  assign y11247 = n36207 ;
  assign y11248 = ~1'b0 ;
  assign y11249 = ~n36210 ;
  assign y11250 = n36214 ;
  assign y11251 = n36221 ;
  assign y11252 = n36222 ;
  assign y11253 = n36223 ;
  assign y11254 = n36225 ;
  assign y11255 = n36226 ;
  assign y11256 = n19435 ;
  assign y11257 = ~n36227 ;
  assign y11258 = ~n36230 ;
  assign y11259 = ~n36231 ;
  assign y11260 = ~n36239 ;
  assign y11261 = ~n36242 ;
  assign y11262 = n36244 ;
  assign y11263 = ~1'b0 ;
  assign y11264 = ~n36245 ;
  assign y11265 = ~n36249 ;
  assign y11266 = ~n36251 ;
  assign y11267 = n36253 ;
  assign y11268 = ~1'b0 ;
  assign y11269 = ~n36257 ;
  assign y11270 = ~n36260 ;
  assign y11271 = n36264 ;
  assign y11272 = n36265 ;
  assign y11273 = n36267 ;
  assign y11274 = n28735 ;
  assign y11275 = ~1'b0 ;
  assign y11276 = n36268 ;
  assign y11277 = ~n36273 ;
  assign y11278 = ~n36278 ;
  assign y11279 = ~n36282 ;
  assign y11280 = ~1'b0 ;
  assign y11281 = ~1'b0 ;
  assign y11282 = ~1'b0 ;
  assign y11283 = ~n36284 ;
  assign y11284 = ~n36288 ;
  assign y11285 = ~n36289 ;
  assign y11286 = ~n36290 ;
  assign y11287 = ~n36296 ;
  assign y11288 = 1'b0 ;
  assign y11289 = ~n36297 ;
  assign y11290 = n36299 ;
  assign y11291 = ~n36302 ;
  assign y11292 = n30635 ;
  assign y11293 = ~n8268 ;
  assign y11294 = ~n36306 ;
  assign y11295 = ~n36307 ;
  assign y11296 = ~1'b0 ;
  assign y11297 = ~1'b0 ;
  assign y11298 = ~n36309 ;
  assign y11299 = n36313 ;
  assign y11300 = ~n36316 ;
  assign y11301 = n36320 ;
  assign y11302 = ~n36322 ;
  assign y11303 = n36323 ;
  assign y11304 = ~n36325 ;
  assign y11305 = n36326 ;
  assign y11306 = n36328 ;
  assign y11307 = n36330 ;
  assign y11308 = ~1'b0 ;
  assign y11309 = n36333 ;
  assign y11310 = ~n36334 ;
  assign y11311 = ~n36336 ;
  assign y11312 = ~1'b0 ;
  assign y11313 = n36337 ;
  assign y11314 = n36345 ;
  assign y11315 = ~n36347 ;
  assign y11316 = n36349 ;
  assign y11317 = ~1'b0 ;
  assign y11318 = n36352 ;
  assign y11319 = n36355 ;
  assign y11320 = ~n36356 ;
  assign y11321 = ~1'b0 ;
  assign y11322 = ~1'b0 ;
  assign y11323 = ~n36364 ;
  assign y11324 = ~n36366 ;
  assign y11325 = ~n36367 ;
  assign y11326 = ~n36380 ;
  assign y11327 = ~1'b0 ;
  assign y11328 = n36388 ;
  assign y11329 = n36390 ;
  assign y11330 = ~n36391 ;
  assign y11331 = ~n36393 ;
  assign y11332 = n36394 ;
  assign y11333 = n36398 ;
  assign y11334 = n36401 ;
  assign y11335 = n36409 ;
  assign y11336 = ~1'b0 ;
  assign y11337 = ~n36417 ;
  assign y11338 = n36418 ;
  assign y11339 = n36419 ;
  assign y11340 = n36425 ;
  assign y11341 = ~n36428 ;
  assign y11342 = n36431 ;
  assign y11343 = ~n36432 ;
  assign y11344 = ~n36435 ;
  assign y11345 = ~n36436 ;
  assign y11346 = ~n36439 ;
  assign y11347 = ~n36442 ;
  assign y11348 = ~n36446 ;
  assign y11349 = ~n36447 ;
  assign y11350 = ~n36452 ;
  assign y11351 = n36460 ;
  assign y11352 = n36462 ;
  assign y11353 = n36464 ;
  assign y11354 = n36467 ;
  assign y11355 = ~n36469 ;
  assign y11356 = n36471 ;
  assign y11357 = ~n36473 ;
  assign y11358 = n36474 ;
  assign y11359 = ~1'b0 ;
  assign y11360 = ~1'b0 ;
  assign y11361 = n36480 ;
  assign y11362 = ~n36484 ;
  assign y11363 = n36488 ;
  assign y11364 = n36493 ;
  assign y11365 = n36494 ;
  assign y11366 = n36500 ;
  assign y11367 = ~n36502 ;
  assign y11368 = ~1'b0 ;
  assign y11369 = n36505 ;
  assign y11370 = ~n36509 ;
  assign y11371 = ~n36513 ;
  assign y11372 = n36515 ;
  assign y11373 = n36516 ;
  assign y11374 = n36517 ;
  assign y11375 = ~n36521 ;
  assign y11376 = n36522 ;
  assign y11377 = ~n36528 ;
  assign y11378 = n36534 ;
  assign y11379 = ~1'b0 ;
  assign y11380 = ~n36535 ;
  assign y11381 = n36536 ;
  assign y11382 = ~n36537 ;
  assign y11383 = ~1'b0 ;
  assign y11384 = n36542 ;
  assign y11385 = n36544 ;
  assign y11386 = ~n36547 ;
  assign y11387 = n36548 ;
  assign y11388 = ~1'b0 ;
  assign y11389 = n36549 ;
  assign y11390 = ~n36556 ;
  assign y11391 = ~n36558 ;
  assign y11392 = ~n36567 ;
  assign y11393 = n36570 ;
  assign y11394 = n36572 ;
  assign y11395 = ~n36579 ;
  assign y11396 = ~n36582 ;
  assign y11397 = ~n36588 ;
  assign y11398 = n36589 ;
  assign y11399 = ~1'b0 ;
  assign y11400 = ~1'b0 ;
  assign y11401 = ~n36591 ;
  assign y11402 = n36593 ;
  assign y11403 = n36594 ;
  assign y11404 = n36596 ;
  assign y11405 = ~n36598 ;
  assign y11406 = ~1'b0 ;
  assign y11407 = n15444 ;
  assign y11408 = ~n36599 ;
  assign y11409 = ~1'b0 ;
  assign y11410 = ~n36607 ;
  assign y11411 = ~n36609 ;
  assign y11412 = n36611 ;
  assign y11413 = n36613 ;
  assign y11414 = ~n36617 ;
  assign y11415 = n36623 ;
  assign y11416 = ~n36624 ;
  assign y11417 = ~n36626 ;
  assign y11418 = ~n36629 ;
  assign y11419 = ~n36630 ;
  assign y11420 = ~n36635 ;
  assign y11421 = n36639 ;
  assign y11422 = ~n36641 ;
  assign y11423 = n20368 ;
  assign y11424 = n36642 ;
  assign y11425 = n36643 ;
  assign y11426 = ~n36648 ;
  assign y11427 = n36652 ;
  assign y11428 = ~n36655 ;
  assign y11429 = ~1'b0 ;
  assign y11430 = ~n36657 ;
  assign y11431 = ~n36662 ;
  assign y11432 = ~n36664 ;
  assign y11433 = n36669 ;
  assign y11434 = ~1'b0 ;
  assign y11435 = n36673 ;
  assign y11436 = 1'b0 ;
  assign y11437 = ~n36675 ;
  assign y11438 = n36677 ;
  assign y11439 = n36678 ;
  assign y11440 = n36681 ;
  assign y11441 = ~n23429 ;
  assign y11442 = n36682 ;
  assign y11443 = ~n36683 ;
  assign y11444 = ~n36688 ;
  assign y11445 = ~1'b0 ;
  assign y11446 = ~n36692 ;
  assign y11447 = ~n36694 ;
  assign y11448 = ~n36695 ;
  assign y11449 = n36696 ;
  assign y11450 = n36698 ;
  assign y11451 = ~n36702 ;
  assign y11452 = ~n36705 ;
  assign y11453 = n36707 ;
  assign y11454 = n36709 ;
  assign y11455 = n36711 ;
  assign y11456 = n36715 ;
  assign y11457 = n36718 ;
  assign y11458 = ~n36721 ;
  assign y11459 = n36725 ;
  assign y11460 = ~1'b0 ;
  assign y11461 = n36726 ;
  assign y11462 = n36728 ;
  assign y11463 = ~n36732 ;
  assign y11464 = n36735 ;
  assign y11465 = ~n36739 ;
  assign y11466 = ~n36741 ;
  assign y11467 = n36742 ;
  assign y11468 = ~n36743 ;
  assign y11469 = n36750 ;
  assign y11470 = ~n36755 ;
  assign y11471 = ~n36764 ;
  assign y11472 = n36765 ;
  assign y11473 = ~n36767 ;
  assign y11474 = ~n36769 ;
  assign y11475 = ~n36770 ;
  assign y11476 = ~n36773 ;
  assign y11477 = n36775 ;
  assign y11478 = ~n36778 ;
  assign y11479 = ~n36782 ;
  assign y11480 = ~n36785 ;
  assign y11481 = n36793 ;
  assign y11482 = n36796 ;
  assign y11483 = n36799 ;
  assign y11484 = ~n36800 ;
  assign y11485 = n36804 ;
  assign y11486 = ~1'b0 ;
  assign y11487 = n36806 ;
  assign y11488 = n36811 ;
  assign y11489 = n36812 ;
  assign y11490 = ~n36813 ;
  assign y11491 = n36816 ;
  assign y11492 = n36820 ;
  assign y11493 = ~n32892 ;
  assign y11494 = ~n36826 ;
  assign y11495 = ~n36830 ;
  assign y11496 = ~1'b0 ;
  assign y11497 = ~1'b0 ;
  assign y11498 = ~1'b0 ;
  assign y11499 = n36833 ;
  assign y11500 = ~n36837 ;
  assign y11501 = n36841 ;
  assign y11502 = ~n36842 ;
  assign y11503 = ~n36850 ;
  assign y11504 = ~n36852 ;
  assign y11505 = ~n36856 ;
  assign y11506 = n36858 ;
  assign y11507 = n36863 ;
  assign y11508 = ~1'b0 ;
  assign y11509 = ~n36865 ;
  assign y11510 = n36871 ;
  assign y11511 = ~n36873 ;
  assign y11512 = ~n36874 ;
  assign y11513 = ~n36875 ;
  assign y11514 = ~n36879 ;
  assign y11515 = n36883 ;
  assign y11516 = ~n36885 ;
  assign y11517 = n36891 ;
  assign y11518 = ~n36892 ;
  assign y11519 = ~n36898 ;
  assign y11520 = ~n36899 ;
  assign y11521 = n36903 ;
  assign y11522 = ~1'b0 ;
  assign y11523 = ~1'b0 ;
  assign y11524 = ~n36908 ;
  assign y11525 = n36909 ;
  assign y11526 = n36580 ;
  assign y11527 = n36911 ;
  assign y11528 = ~n36912 ;
  assign y11529 = ~n36913 ;
  assign y11530 = n36920 ;
  assign y11531 = ~n36921 ;
  assign y11532 = ~n36923 ;
  assign y11533 = ~n36924 ;
  assign y11534 = n36925 ;
  assign y11535 = n36929 ;
  assign y11536 = ~n36930 ;
  assign y11537 = n36932 ;
  assign y11538 = ~1'b0 ;
  assign y11539 = n36936 ;
  assign y11540 = ~n36937 ;
  assign y11541 = ~n36938 ;
  assign y11542 = ~n36939 ;
  assign y11543 = n36941 ;
  assign y11544 = n36945 ;
  assign y11545 = n36950 ;
  assign y11546 = ~n36954 ;
  assign y11547 = ~n36959 ;
  assign y11548 = ~n36963 ;
  assign y11549 = n36965 ;
  assign y11550 = ~n36969 ;
  assign y11551 = n36971 ;
  assign y11552 = ~n36973 ;
  assign y11553 = ~n2147 ;
  assign y11554 = n36977 ;
  assign y11555 = n36980 ;
  assign y11556 = n36984 ;
  assign y11557 = n36985 ;
  assign y11558 = ~n36989 ;
  assign y11559 = ~1'b0 ;
  assign y11560 = ~1'b0 ;
  assign y11561 = n36995 ;
  assign y11562 = n36996 ;
  assign y11563 = n10440 ;
  assign y11564 = ~n36997 ;
  assign y11565 = n36999 ;
  assign y11566 = ~n37000 ;
  assign y11567 = n37001 ;
  assign y11568 = ~n37003 ;
  assign y11569 = n37011 ;
  assign y11570 = ~n37015 ;
  assign y11571 = n37016 ;
  assign y11572 = n37019 ;
  assign y11573 = ~n37020 ;
  assign y11574 = n37023 ;
  assign y11575 = n37026 ;
  assign y11576 = ~n37029 ;
  assign y11577 = ~n37031 ;
  assign y11578 = ~1'b0 ;
  assign y11579 = ~n37033 ;
  assign y11580 = ~n37038 ;
  assign y11581 = n37045 ;
  assign y11582 = ~1'b0 ;
  assign y11583 = ~n37047 ;
  assign y11584 = ~n20491 ;
  assign y11585 = n37053 ;
  assign y11586 = n37055 ;
  assign y11587 = ~n37056 ;
  assign y11588 = ~1'b0 ;
  assign y11589 = n37058 ;
  assign y11590 = ~n37061 ;
  assign y11591 = n37063 ;
  assign y11592 = ~n37064 ;
  assign y11593 = n37069 ;
  assign y11594 = n37070 ;
  assign y11595 = n37072 ;
  assign y11596 = ~n37073 ;
  assign y11597 = ~n37075 ;
  assign y11598 = ~n37076 ;
  assign y11599 = ~n30363 ;
  assign y11600 = ~n37082 ;
  assign y11601 = n37084 ;
  assign y11602 = ~n37086 ;
  assign y11603 = n37088 ;
  assign y11604 = ~n37094 ;
  assign y11605 = ~n37098 ;
  assign y11606 = ~n37099 ;
  assign y11607 = n37100 ;
  assign y11608 = n37102 ;
  assign y11609 = ~1'b0 ;
  assign y11610 = ~n37105 ;
  assign y11611 = ~n37106 ;
  assign y11612 = n37109 ;
  assign y11613 = n37111 ;
  assign y11614 = ~n37112 ;
  assign y11615 = ~n37114 ;
  assign y11616 = n37116 ;
  assign y11617 = ~n37117 ;
  assign y11618 = n37120 ;
  assign y11619 = n37121 ;
  assign y11620 = n37122 ;
  assign y11621 = n21585 ;
  assign y11622 = ~n37129 ;
  assign y11623 = ~n37133 ;
  assign y11624 = ~n37135 ;
  assign y11625 = ~n37138 ;
  assign y11626 = n37143 ;
  assign y11627 = n37146 ;
  assign y11628 = ~n37148 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = 1'b0 ;
  assign y11631 = ~n37151 ;
  assign y11632 = n37153 ;
  assign y11633 = n37156 ;
  assign y11634 = ~n37157 ;
  assign y11635 = n30727 ;
  assign y11636 = ~n37170 ;
  assign y11637 = ~n37178 ;
  assign y11638 = ~n37179 ;
  assign y11639 = n37180 ;
  assign y11640 = ~n37183 ;
  assign y11641 = n37185 ;
  assign y11642 = ~n37188 ;
  assign y11643 = ~1'b0 ;
  assign y11644 = ~n37189 ;
  assign y11645 = ~n37197 ;
  assign y11646 = ~n37199 ;
  assign y11647 = ~n37202 ;
  assign y11648 = ~n37204 ;
  assign y11649 = n37206 ;
  assign y11650 = ~1'b0 ;
  assign y11651 = ~n37214 ;
  assign y11652 = ~n37215 ;
  assign y11653 = n37216 ;
  assign y11654 = ~n22028 ;
  assign y11655 = n37221 ;
  assign y11656 = ~n37225 ;
  assign y11657 = ~1'b0 ;
  assign y11658 = n26257 ;
  assign y11659 = n37226 ;
  assign y11660 = n37228 ;
  assign y11661 = ~n37230 ;
  assign y11662 = n37231 ;
  assign y11663 = n37236 ;
  assign y11664 = ~1'b0 ;
  assign y11665 = ~1'b0 ;
  assign y11666 = n37240 ;
  assign y11667 = ~n37241 ;
  assign y11668 = ~n37242 ;
  assign y11669 = n37245 ;
  assign y11670 = ~n37247 ;
  assign y11671 = ~n37249 ;
  assign y11672 = n37250 ;
  assign y11673 = ~n37263 ;
  assign y11674 = ~n37265 ;
  assign y11675 = ~n36399 ;
  assign y11676 = ~n37270 ;
  assign y11677 = n37277 ;
  assign y11678 = n37278 ;
  assign y11679 = ~n37280 ;
  assign y11680 = n37281 ;
  assign y11681 = n10114 ;
  assign y11682 = ~n37283 ;
  assign y11683 = ~n37285 ;
  assign y11684 = ~1'b0 ;
  assign y11685 = ~n37286 ;
  assign y11686 = ~n37287 ;
  assign y11687 = ~n11830 ;
  assign y11688 = n37288 ;
  assign y11689 = ~n37291 ;
  assign y11690 = ~n37296 ;
  assign y11691 = n37299 ;
  assign y11692 = ~n37303 ;
  assign y11693 = ~1'b0 ;
  assign y11694 = n37307 ;
  assign y11695 = n37309 ;
  assign y11696 = ~n37316 ;
  assign y11697 = ~1'b0 ;
  assign y11698 = ~n37317 ;
  assign y11699 = n37318 ;
  assign y11700 = n37329 ;
  assign y11701 = ~n37332 ;
  assign y11702 = ~n37333 ;
  assign y11703 = n37337 ;
  assign y11704 = ~n37341 ;
  assign y11705 = n37344 ;
  assign y11706 = ~n37346 ;
  assign y11707 = n37347 ;
  assign y11708 = ~1'b0 ;
  assign y11709 = n37350 ;
  assign y11710 = ~n37362 ;
  assign y11711 = n37366 ;
  assign y11712 = ~n37367 ;
  assign y11713 = ~n37368 ;
  assign y11714 = n37371 ;
  assign y11715 = n37379 ;
  assign y11716 = ~n37380 ;
  assign y11717 = ~1'b0 ;
  assign y11718 = ~n37381 ;
  assign y11719 = n37390 ;
  assign y11720 = n37394 ;
  assign y11721 = ~n37395 ;
  assign y11722 = n37397 ;
  assign y11723 = ~n37399 ;
  assign y11724 = ~1'b0 ;
  assign y11725 = ~n37401 ;
  assign y11726 = n37402 ;
  assign y11727 = ~n25094 ;
  assign y11728 = ~n37403 ;
  assign y11729 = n37405 ;
  assign y11730 = ~n37407 ;
  assign y11731 = n37408 ;
  assign y11732 = n37413 ;
  assign y11733 = ~n37414 ;
  assign y11734 = ~n37417 ;
  assign y11735 = ~n37418 ;
  assign y11736 = n37422 ;
  assign y11737 = ~n37427 ;
  assign y11738 = ~1'b0 ;
  assign y11739 = ~1'b0 ;
  assign y11740 = ~n37431 ;
  assign y11741 = ~n37432 ;
  assign y11742 = ~n37437 ;
  assign y11743 = ~n37441 ;
  assign y11744 = n37446 ;
  assign y11745 = ~1'b0 ;
  assign y11746 = ~1'b0 ;
  assign y11747 = ~n37448 ;
  assign y11748 = n37452 ;
  assign y11749 = ~n37453 ;
  assign y11750 = ~n37459 ;
  assign y11751 = n37461 ;
  assign y11752 = ~1'b0 ;
  assign y11753 = ~n37466 ;
  assign y11754 = n37467 ;
  assign y11755 = n37470 ;
  assign y11756 = n37471 ;
  assign y11757 = ~n37475 ;
  assign y11758 = n37480 ;
  assign y11759 = n37482 ;
  assign y11760 = ~1'b0 ;
  assign y11761 = ~n37484 ;
  assign y11762 = ~n37488 ;
  assign y11763 = ~1'b0 ;
  assign y11764 = ~n37492 ;
  assign y11765 = ~n37494 ;
  assign y11766 = n37497 ;
  assign y11767 = ~1'b0 ;
  assign y11768 = n37500 ;
  assign y11769 = ~n37504 ;
  assign y11770 = n37506 ;
  assign y11771 = ~n37508 ;
  assign y11772 = ~n37510 ;
  assign y11773 = ~1'b0 ;
  assign y11774 = n37512 ;
  assign y11775 = n37516 ;
  assign y11776 = ~n37519 ;
  assign y11777 = n37523 ;
  assign y11778 = ~n37526 ;
  assign y11779 = n37527 ;
  assign y11780 = n37531 ;
  assign y11781 = n37534 ;
  assign y11782 = n37536 ;
  assign y11783 = ~1'b0 ;
  assign y11784 = ~n37539 ;
  assign y11785 = ~n37542 ;
  assign y11786 = n37544 ;
  assign y11787 = ~n37546 ;
  assign y11788 = ~n37547 ;
  assign y11789 = n37548 ;
  assign y11790 = n37550 ;
  assign y11791 = n37552 ;
  assign y11792 = ~1'b0 ;
  assign y11793 = ~1'b0 ;
  assign y11794 = ~n37558 ;
  assign y11795 = n37560 ;
  assign y11796 = n37564 ;
  assign y11797 = ~n37567 ;
  assign y11798 = ~1'b0 ;
  assign y11799 = ~1'b0 ;
  assign y11800 = ~1'b0 ;
  assign y11801 = ~n37568 ;
  assign y11802 = ~n37573 ;
  assign y11803 = ~n37580 ;
  assign y11804 = ~n37581 ;
  assign y11805 = n37582 ;
  assign y11806 = ~n37587 ;
  assign y11807 = ~1'b0 ;
  assign y11808 = n37590 ;
  assign y11809 = ~n37592 ;
  assign y11810 = ~n37595 ;
  assign y11811 = ~n37597 ;
  assign y11812 = n37598 ;
  assign y11813 = n37599 ;
  assign y11814 = ~n37604 ;
  assign y11815 = n37605 ;
  assign y11816 = ~n37609 ;
  assign y11817 = ~n37611 ;
  assign y11818 = n37612 ;
  assign y11819 = ~1'b0 ;
  assign y11820 = n37623 ;
  assign y11821 = ~n37624 ;
  assign y11822 = ~n37626 ;
  assign y11823 = ~1'b0 ;
  assign y11824 = n37627 ;
  assign y11825 = n37631 ;
  assign y11826 = ~1'b0 ;
  assign y11827 = n37642 ;
  assign y11828 = n37651 ;
  assign y11829 = n37653 ;
  assign y11830 = n37655 ;
  assign y11831 = ~n37658 ;
  assign y11832 = n37664 ;
  assign y11833 = ~1'b0 ;
  assign y11834 = ~n37666 ;
  assign y11835 = ~n37671 ;
  assign y11836 = ~n37672 ;
  assign y11837 = ~n37689 ;
  assign y11838 = ~n37697 ;
  assign y11839 = n37699 ;
  assign y11840 = 1'b0 ;
  assign y11841 = ~1'b0 ;
  assign y11842 = n37703 ;
  assign y11843 = n37710 ;
  assign y11844 = ~n37714 ;
  assign y11845 = ~n37716 ;
  assign y11846 = ~n37719 ;
  assign y11847 = ~1'b0 ;
  assign y11848 = ~n37724 ;
  assign y11849 = ~n37725 ;
  assign y11850 = ~n37731 ;
  assign y11851 = n37732 ;
  assign y11852 = n37739 ;
  assign y11853 = n37741 ;
  assign y11854 = ~n37747 ;
  assign y11855 = n37750 ;
  assign y11856 = ~n37757 ;
  assign y11857 = ~n37763 ;
  assign y11858 = n37767 ;
  assign y11859 = n37770 ;
  assign y11860 = ~n37772 ;
  assign y11861 = ~n37774 ;
  assign y11862 = n37777 ;
  assign y11863 = n37779 ;
  assign y11864 = n37780 ;
  assign y11865 = ~n37781 ;
  assign y11866 = ~n37786 ;
  assign y11867 = ~n37789 ;
  assign y11868 = n37794 ;
  assign y11869 = ~n37797 ;
  assign y11870 = ~n37799 ;
  assign y11871 = ~n37803 ;
  assign y11872 = ~n37807 ;
  assign y11873 = n37810 ;
  assign y11874 = n37812 ;
  assign y11875 = n37820 ;
  assign y11876 = n37821 ;
  assign y11877 = n37826 ;
  assign y11878 = n37832 ;
  assign y11879 = n37833 ;
  assign y11880 = n37835 ;
  assign y11881 = ~n37837 ;
  assign y11882 = n37842 ;
  assign y11883 = ~n37844 ;
  assign y11884 = ~n37847 ;
  assign y11885 = ~1'b0 ;
  assign y11886 = ~n37849 ;
  assign y11887 = ~n37851 ;
  assign y11888 = n37855 ;
  assign y11889 = ~n37857 ;
  assign y11890 = ~1'b0 ;
  assign y11891 = ~1'b0 ;
  assign y11892 = n37860 ;
  assign y11893 = ~1'b0 ;
  assign y11894 = ~n37863 ;
  assign y11895 = n37864 ;
  assign y11896 = n29581 ;
  assign y11897 = ~n37865 ;
  assign y11898 = n37867 ;
  assign y11899 = ~n37870 ;
  assign y11900 = n37872 ;
  assign y11901 = n37874 ;
  assign y11902 = ~1'b0 ;
  assign y11903 = ~n37877 ;
  assign y11904 = ~n37881 ;
  assign y11905 = ~n37885 ;
  assign y11906 = ~n37886 ;
  assign y11907 = n37889 ;
  assign y11908 = ~n37892 ;
  assign y11909 = n37894 ;
  assign y11910 = ~n32137 ;
  assign y11911 = n37898 ;
  assign y11912 = ~n37901 ;
  assign y11913 = n37904 ;
  assign y11914 = ~n37910 ;
  assign y11915 = ~n37912 ;
  assign y11916 = n37915 ;
  assign y11917 = ~1'b0 ;
  assign y11918 = n37919 ;
  assign y11919 = n37924 ;
  assign y11920 = ~n37927 ;
  assign y11921 = n37928 ;
  assign y11922 = n37931 ;
  assign y11923 = ~1'b0 ;
  assign y11924 = ~n37933 ;
  assign y11925 = ~1'b0 ;
  assign y11926 = n37935 ;
  assign y11927 = ~n37936 ;
  assign y11928 = ~n37941 ;
  assign y11929 = n37942 ;
  assign y11930 = ~n37948 ;
  assign y11931 = ~n37952 ;
  assign y11932 = n37956 ;
  assign y11933 = ~1'b0 ;
  assign y11934 = ~1'b0 ;
  assign y11935 = ~1'b0 ;
  assign y11936 = ~n15892 ;
  assign y11937 = n37957 ;
  assign y11938 = n37959 ;
  assign y11939 = ~1'b0 ;
  assign y11940 = ~n37960 ;
  assign y11941 = ~n37962 ;
  assign y11942 = ~n28357 ;
  assign y11943 = n37965 ;
  assign y11944 = ~1'b0 ;
  assign y11945 = n37968 ;
  assign y11946 = ~n37974 ;
  assign y11947 = n37975 ;
  assign y11948 = ~1'b0 ;
  assign y11949 = n37977 ;
  assign y11950 = ~n37982 ;
  assign y11951 = ~n37983 ;
  assign y11952 = ~n37988 ;
  assign y11953 = n37990 ;
  assign y11954 = ~n11510 ;
  assign y11955 = n37994 ;
  assign y11956 = ~1'b0 ;
  assign y11957 = ~n32914 ;
  assign y11958 = n37998 ;
  assign y11959 = ~n38003 ;
  assign y11960 = n38004 ;
  assign y11961 = n38007 ;
  assign y11962 = n38011 ;
  assign y11963 = ~1'b0 ;
  assign y11964 = ~n38012 ;
  assign y11965 = n17787 ;
  assign y11966 = ~n38015 ;
  assign y11967 = ~n38017 ;
  assign y11968 = n38023 ;
  assign y11969 = ~n38026 ;
  assign y11970 = ~n38028 ;
  assign y11971 = n38029 ;
  assign y11972 = ~n38030 ;
  assign y11973 = ~n38042 ;
  assign y11974 = ~n38044 ;
  assign y11975 = ~n38045 ;
  assign y11976 = ~1'b0 ;
  assign y11977 = ~1'b0 ;
  assign y11978 = ~n18765 ;
  assign y11979 = n38046 ;
  assign y11980 = ~n38047 ;
  assign y11981 = n38052 ;
  assign y11982 = n38055 ;
  assign y11983 = n38057 ;
  assign y11984 = ~n38059 ;
  assign y11985 = ~1'b0 ;
  assign y11986 = ~1'b0 ;
  assign y11987 = ~1'b0 ;
  assign y11988 = ~n38060 ;
  assign y11989 = ~n38065 ;
  assign y11990 = ~n38066 ;
  assign y11991 = n38068 ;
  assign y11992 = ~n38069 ;
  assign y11993 = ~n38071 ;
  assign y11994 = ~n38072 ;
  assign y11995 = ~1'b0 ;
  assign y11996 = ~n38074 ;
  assign y11997 = ~n38077 ;
  assign y11998 = n38080 ;
  assign y11999 = n38082 ;
  assign y12000 = ~n38087 ;
  assign y12001 = ~1'b0 ;
  assign y12002 = n38091 ;
  assign y12003 = ~n38092 ;
  assign y12004 = n38093 ;
  assign y12005 = n38095 ;
  assign y12006 = ~1'b0 ;
  assign y12007 = ~n38097 ;
  assign y12008 = n38100 ;
  assign y12009 = n38101 ;
  assign y12010 = ~n38104 ;
  assign y12011 = n38107 ;
  assign y12012 = ~1'b0 ;
  assign y12013 = n38109 ;
  assign y12014 = ~n38111 ;
  assign y12015 = ~n38114 ;
  assign y12016 = ~n38120 ;
  assign y12017 = n38122 ;
  assign y12018 = n38123 ;
  assign y12019 = n38125 ;
  assign y12020 = ~n38126 ;
  assign y12021 = n38128 ;
  assign y12022 = ~n38130 ;
  assign y12023 = ~n38134 ;
  assign y12024 = n38142 ;
  assign y12025 = n38144 ;
  assign y12026 = ~n38149 ;
  assign y12027 = n38155 ;
  assign y12028 = n38165 ;
  assign y12029 = n38166 ;
  assign y12030 = ~1'b0 ;
  assign y12031 = ~n38168 ;
  assign y12032 = n38171 ;
  assign y12033 = n38173 ;
  assign y12034 = ~n38174 ;
  assign y12035 = ~n38175 ;
  assign y12036 = ~n38182 ;
  assign y12037 = ~n38184 ;
  assign y12038 = n38187 ;
  assign y12039 = n38191 ;
  assign y12040 = ~1'b0 ;
  assign y12041 = ~n38192 ;
  assign y12042 = n38193 ;
  assign y12043 = ~n38194 ;
  assign y12044 = ~n38195 ;
  assign y12045 = ~n38196 ;
  assign y12046 = ~n38198 ;
  assign y12047 = ~n38200 ;
  assign y12048 = ~n38204 ;
  assign y12049 = ~n38209 ;
  assign y12050 = ~n38214 ;
  assign y12051 = ~n38217 ;
  assign y12052 = ~n38220 ;
  assign y12053 = ~n38222 ;
  assign y12054 = n38226 ;
  assign y12055 = n38227 ;
  assign y12056 = n38228 ;
  assign y12057 = ~n38231 ;
  assign y12058 = ~n38233 ;
  assign y12059 = n38234 ;
  assign y12060 = n38236 ;
  assign y12061 = ~1'b0 ;
  assign y12062 = n38245 ;
  assign y12063 = ~n38247 ;
  assign y12064 = n11519 ;
  assign y12065 = ~n38251 ;
  assign y12066 = n38252 ;
  assign y12067 = ~n38254 ;
  assign y12068 = ~n38260 ;
  assign y12069 = ~n38261 ;
  assign y12070 = n38262 ;
  assign y12071 = n38263 ;
  assign y12072 = n38264 ;
  assign y12073 = n38267 ;
  assign y12074 = ~n38269 ;
  assign y12075 = ~n38270 ;
  assign y12076 = ~1'b0 ;
  assign y12077 = n38273 ;
  assign y12078 = ~n38274 ;
  assign y12079 = n38277 ;
  assign y12080 = n38279 ;
  assign y12081 = ~n38280 ;
  assign y12082 = n38286 ;
  assign y12083 = ~n38287 ;
  assign y12084 = ~n38294 ;
  assign y12085 = n38295 ;
  assign y12086 = ~n38296 ;
  assign y12087 = ~n38299 ;
  assign y12088 = n38300 ;
  assign y12089 = n38301 ;
  assign y12090 = ~1'b0 ;
  assign y12091 = ~n38303 ;
  assign y12092 = ~n38304 ;
  assign y12093 = n24120 ;
  assign y12094 = ~n38307 ;
  assign y12095 = ~1'b0 ;
  assign y12096 = ~n38309 ;
  assign y12097 = ~n38312 ;
  assign y12098 = ~n38313 ;
  assign y12099 = ~n38314 ;
  assign y12100 = n38315 ;
  assign y12101 = ~n38322 ;
  assign y12102 = n38323 ;
  assign y12103 = ~1'b0 ;
  assign y12104 = 1'b0 ;
  assign y12105 = n38324 ;
  assign y12106 = ~n38330 ;
  assign y12107 = ~n38332 ;
  assign y12108 = n38333 ;
  assign y12109 = n38337 ;
  assign y12110 = ~n38340 ;
  assign y12111 = ~1'b0 ;
  assign y12112 = ~n38341 ;
  assign y12113 = n38344 ;
  assign y12114 = n38346 ;
  assign y12115 = n38348 ;
  assign y12116 = n38353 ;
  assign y12117 = n38358 ;
  assign y12118 = n38359 ;
  assign y12119 = n38361 ;
  assign y12120 = ~n38362 ;
  assign y12121 = n38371 ;
  assign y12122 = n38377 ;
  assign y12123 = ~n38385 ;
  assign y12124 = ~n38387 ;
  assign y12125 = ~n38390 ;
  assign y12126 = n38391 ;
  assign y12127 = n38393 ;
  assign y12128 = ~n38394 ;
  assign y12129 = ~1'b0 ;
  assign y12130 = ~n38398 ;
  assign y12131 = n11353 ;
  assign y12132 = n38402 ;
  assign y12133 = ~n38403 ;
  assign y12134 = n38408 ;
  assign y12135 = ~1'b0 ;
  assign y12136 = ~n38409 ;
  assign y12137 = n38411 ;
  assign y12138 = n38414 ;
  assign y12139 = n38420 ;
  assign y12140 = n38421 ;
  assign y12141 = ~1'b0 ;
  assign y12142 = ~1'b0 ;
  assign y12143 = ~n38422 ;
  assign y12144 = ~n38432 ;
  assign y12145 = ~n38435 ;
  assign y12146 = ~1'b0 ;
  assign y12147 = n38436 ;
  assign y12148 = n38437 ;
  assign y12149 = n38446 ;
  assign y12150 = ~n38448 ;
  assign y12151 = ~n38451 ;
  assign y12152 = n38454 ;
  assign y12153 = ~1'b0 ;
  assign y12154 = ~n38456 ;
  assign y12155 = n38457 ;
  assign y12156 = ~n38459 ;
  assign y12157 = ~n38461 ;
  assign y12158 = ~n38463 ;
  assign y12159 = ~n38465 ;
  assign y12160 = n38468 ;
  assign y12161 = ~n38470 ;
  assign y12162 = n38472 ;
  assign y12163 = n38473 ;
  assign y12164 = n38483 ;
  assign y12165 = ~n38489 ;
  assign y12166 = n38490 ;
  assign y12167 = n38491 ;
  assign y12168 = ~n38497 ;
  assign y12169 = n38503 ;
  assign y12170 = n38507 ;
  assign y12171 = ~n38512 ;
  assign y12172 = ~n38517 ;
  assign y12173 = ~n38520 ;
  assign y12174 = n38521 ;
  assign y12175 = ~n38524 ;
  assign y12176 = ~n38525 ;
  assign y12177 = ~n38531 ;
  assign y12178 = n38538 ;
  assign y12179 = ~n38540 ;
  assign y12180 = ~1'b0 ;
  assign y12181 = n38541 ;
  assign y12182 = n38542 ;
  assign y12183 = n38543 ;
  assign y12184 = n38544 ;
  assign y12185 = n38547 ;
  assign y12186 = ~n38549 ;
  assign y12187 = n17785 ;
  assign y12188 = n38550 ;
  assign y12189 = n38551 ;
  assign y12190 = n38553 ;
  assign y12191 = n38559 ;
  assign y12192 = ~n38560 ;
  assign y12193 = n38564 ;
  assign y12194 = n38566 ;
  assign y12195 = n38568 ;
  assign y12196 = ~n38573 ;
  assign y12197 = n38576 ;
  assign y12198 = ~n38577 ;
  assign y12199 = n38582 ;
  assign y12200 = n38583 ;
  assign y12201 = ~n38585 ;
  assign y12202 = ~n38588 ;
  assign y12203 = ~1'b0 ;
  assign y12204 = n38590 ;
  assign y12205 = ~n38593 ;
  assign y12206 = ~n38595 ;
  assign y12207 = n38596 ;
  assign y12208 = n38597 ;
  assign y12209 = ~n38602 ;
  assign y12210 = n38605 ;
  assign y12211 = ~n38607 ;
  assign y12212 = n38609 ;
  assign y12213 = ~n38613 ;
  assign y12214 = n38616 ;
  assign y12215 = n38620 ;
  assign y12216 = n38626 ;
  assign y12217 = ~n38627 ;
  assign y12218 = n38636 ;
  assign y12219 = n38640 ;
  assign y12220 = n38641 ;
  assign y12221 = n38642 ;
  assign y12222 = ~n38645 ;
  assign y12223 = n38647 ;
  assign y12224 = n38650 ;
  assign y12225 = ~n38653 ;
  assign y12226 = n38654 ;
  assign y12227 = ~1'b0 ;
  assign y12228 = ~n38656 ;
  assign y12229 = ~n38657 ;
  assign y12230 = ~1'b0 ;
  assign y12231 = ~n38660 ;
  assign y12232 = ~n38665 ;
  assign y12233 = n38667 ;
  assign y12234 = ~n38668 ;
  assign y12235 = ~n38669 ;
  assign y12236 = ~n38671 ;
  assign y12237 = ~1'b0 ;
  assign y12238 = ~n38675 ;
  assign y12239 = n38676 ;
  assign y12240 = ~n38678 ;
  assign y12241 = ~n38685 ;
  assign y12242 = n38686 ;
  assign y12243 = ~n38690 ;
  assign y12244 = ~1'b0 ;
  assign y12245 = ~n38696 ;
  assign y12246 = ~n38699 ;
  assign y12247 = ~1'b0 ;
  assign y12248 = ~n38700 ;
  assign y12249 = n38701 ;
  assign y12250 = n38706 ;
  assign y12251 = ~n38708 ;
  assign y12252 = ~n38715 ;
  assign y12253 = n38716 ;
  assign y12254 = ~1'b0 ;
  assign y12255 = ~1'b0 ;
  assign y12256 = ~n38719 ;
  assign y12257 = ~n38721 ;
  assign y12258 = ~n38726 ;
  assign y12259 = n38728 ;
  assign y12260 = ~n38733 ;
  assign y12261 = n38738 ;
  assign y12262 = ~n38740 ;
  assign y12263 = ~n38741 ;
  assign y12264 = n38742 ;
  assign y12265 = ~n38743 ;
  assign y12266 = ~1'b0 ;
  assign y12267 = ~1'b0 ;
  assign y12268 = ~n38748 ;
  assign y12269 = ~n38749 ;
  assign y12270 = ~n38750 ;
  assign y12271 = ~n38754 ;
  assign y12272 = n38756 ;
  assign y12273 = n38760 ;
  assign y12274 = n38762 ;
  assign y12275 = n38765 ;
  assign y12276 = n38767 ;
  assign y12277 = ~n38768 ;
  assign y12278 = ~n38771 ;
  assign y12279 = n38774 ;
  assign y12280 = ~n38777 ;
  assign y12281 = n38783 ;
  assign y12282 = ~n38789 ;
  assign y12283 = n38791 ;
  assign y12284 = ~1'b0 ;
  assign y12285 = ~n38796 ;
  assign y12286 = ~1'b0 ;
  assign y12287 = ~1'b0 ;
  assign y12288 = ~n38797 ;
  assign y12289 = n38800 ;
  assign y12290 = ~n38805 ;
  assign y12291 = ~n38806 ;
  assign y12292 = ~n38813 ;
  assign y12293 = ~n38815 ;
  assign y12294 = ~n38816 ;
  assign y12295 = n38817 ;
  assign y12296 = ~n38820 ;
  assign y12297 = n38822 ;
  assign y12298 = n38823 ;
  assign y12299 = ~n38825 ;
  assign y12300 = n38827 ;
  assign y12301 = ~n38829 ;
  assign y12302 = ~n38833 ;
  assign y12303 = n38837 ;
  assign y12304 = ~n38839 ;
  assign y12305 = ~1'b0 ;
  assign y12306 = n38840 ;
  assign y12307 = ~n38842 ;
  assign y12308 = n38843 ;
  assign y12309 = ~n38845 ;
  assign y12310 = n38851 ;
  assign y12311 = n38855 ;
  assign y12312 = ~1'b0 ;
  assign y12313 = ~n38857 ;
  assign y12314 = ~1'b0 ;
  assign y12315 = ~n38870 ;
  assign y12316 = n38874 ;
  assign y12317 = n38877 ;
  assign y12318 = ~n38878 ;
  assign y12319 = ~n38881 ;
  assign y12320 = ~n38882 ;
  assign y12321 = ~1'b0 ;
  assign y12322 = ~n38884 ;
  assign y12323 = n38890 ;
  assign y12324 = n38891 ;
  assign y12325 = ~n38899 ;
  assign y12326 = n38900 ;
  assign y12327 = ~n38901 ;
  assign y12328 = ~n38905 ;
  assign y12329 = n38908 ;
  assign y12330 = ~1'b0 ;
  assign y12331 = ~n38912 ;
  assign y12332 = ~1'b0 ;
  assign y12333 = ~n38916 ;
  assign y12334 = ~n38917 ;
  assign y12335 = ~n38920 ;
  assign y12336 = ~1'b0 ;
  assign y12337 = ~1'b0 ;
  assign y12338 = ~n38922 ;
  assign y12339 = ~n38923 ;
  assign y12340 = ~n38924 ;
  assign y12341 = ~n38926 ;
  assign y12342 = ~1'b0 ;
  assign y12343 = ~1'b0 ;
  assign y12344 = ~n38937 ;
  assign y12345 = ~n38938 ;
  assign y12346 = ~n38940 ;
  assign y12347 = ~n38942 ;
  assign y12348 = ~1'b0 ;
  assign y12349 = ~n38944 ;
  assign y12350 = ~n38952 ;
  assign y12351 = ~n38953 ;
  assign y12352 = ~n38954 ;
  assign y12353 = ~n38956 ;
  assign y12354 = ~n38959 ;
  assign y12355 = ~n38961 ;
  assign y12356 = n38965 ;
  assign y12357 = n38967 ;
  assign y12358 = ~n38968 ;
  assign y12359 = ~n38970 ;
  assign y12360 = n38972 ;
  assign y12361 = ~n38974 ;
  assign y12362 = n38977 ;
  assign y12363 = n38982 ;
  assign y12364 = ~n38987 ;
  assign y12365 = ~n38991 ;
  assign y12366 = n38992 ;
  assign y12367 = n38994 ;
  assign y12368 = ~n38998 ;
  assign y12369 = ~n38999 ;
  assign y12370 = n39003 ;
  assign y12371 = n39005 ;
  assign y12372 = n39009 ;
  assign y12373 = n39010 ;
  assign y12374 = n39013 ;
  assign y12375 = n39016 ;
  assign y12376 = ~n39017 ;
  assign y12377 = n39019 ;
  assign y12378 = ~1'b0 ;
  assign y12379 = ~n39021 ;
  assign y12380 = n39024 ;
  assign y12381 = ~n39026 ;
  assign y12382 = n39027 ;
  assign y12383 = n39039 ;
  assign y12384 = ~1'b0 ;
  assign y12385 = ~n39043 ;
  assign y12386 = n39048 ;
  assign y12387 = ~n39049 ;
  assign y12388 = ~n39052 ;
  assign y12389 = n39053 ;
  assign y12390 = ~n39055 ;
  assign y12391 = ~n39056 ;
  assign y12392 = ~n39058 ;
  assign y12393 = ~n39060 ;
  assign y12394 = ~n39062 ;
  assign y12395 = n39063 ;
  assign y12396 = n39066 ;
  assign y12397 = ~n39069 ;
  assign y12398 = ~1'b0 ;
  assign y12399 = n39071 ;
  assign y12400 = n39073 ;
  assign y12401 = ~1'b0 ;
  assign y12402 = n39074 ;
  assign y12403 = n39076 ;
  assign y12404 = ~n39080 ;
  assign y12405 = n39081 ;
  assign y12406 = ~n39084 ;
  assign y12407 = ~n39085 ;
  assign y12408 = ~n39087 ;
  assign y12409 = ~n39089 ;
  assign y12410 = n39090 ;
  assign y12411 = n39092 ;
  assign y12412 = ~n39094 ;
  assign y12413 = ~n39095 ;
  assign y12414 = ~n39098 ;
  assign y12415 = ~n39103 ;
  assign y12416 = ~1'b0 ;
  assign y12417 = ~n39107 ;
  assign y12418 = ~n39108 ;
  assign y12419 = n39110 ;
  assign y12420 = ~n39113 ;
  assign y12421 = n39116 ;
  assign y12422 = n39118 ;
  assign y12423 = n39119 ;
  assign y12424 = n39128 ;
  assign y12425 = ~n39134 ;
  assign y12426 = n39136 ;
  assign y12427 = n39141 ;
  assign y12428 = ~n39142 ;
  assign y12429 = ~1'b0 ;
  assign y12430 = n39143 ;
  assign y12431 = n39148 ;
  assign y12432 = ~1'b0 ;
  assign y12433 = ~1'b0 ;
  assign y12434 = n39152 ;
  assign y12435 = n39153 ;
  assign y12436 = ~n39157 ;
  assign y12437 = n39166 ;
  assign y12438 = ~n39174 ;
  assign y12439 = n39177 ;
  assign y12440 = ~1'b0 ;
  assign y12441 = n39178 ;
  assign y12442 = ~n39180 ;
  assign y12443 = n39184 ;
  assign y12444 = n39185 ;
  assign y12445 = n39186 ;
  assign y12446 = n39191 ;
  assign y12447 = ~1'b0 ;
  assign y12448 = n39192 ;
  assign y12449 = ~n39193 ;
  assign y12450 = ~n39194 ;
  assign y12451 = ~n39196 ;
  assign y12452 = n39202 ;
  assign y12453 = ~1'b0 ;
  assign y12454 = n39207 ;
  assign y12455 = ~n39210 ;
  assign y12456 = n39218 ;
  assign y12457 = ~n39219 ;
  assign y12458 = ~n39221 ;
  assign y12459 = ~n39222 ;
  assign y12460 = n39226 ;
  assign y12461 = n39229 ;
  assign y12462 = n39235 ;
  assign y12463 = n39239 ;
  assign y12464 = n39240 ;
  assign y12465 = ~n39243 ;
  assign y12466 = ~n39245 ;
  assign y12467 = ~n39247 ;
  assign y12468 = ~1'b0 ;
  assign y12469 = ~n39250 ;
  assign y12470 = n39251 ;
  assign y12471 = n39252 ;
  assign y12472 = ~n39256 ;
  assign y12473 = ~n39259 ;
  assign y12474 = n39262 ;
  assign y12475 = n39265 ;
  assign y12476 = ~n39271 ;
  assign y12477 = ~n39276 ;
  assign y12478 = n39280 ;
  assign y12479 = n39282 ;
  assign y12480 = ~n39286 ;
  assign y12481 = ~1'b0 ;
  assign y12482 = n39287 ;
  assign y12483 = ~n39291 ;
  assign y12484 = n39293 ;
  assign y12485 = n39300 ;
  assign y12486 = ~n39302 ;
  assign y12487 = ~n39307 ;
  assign y12488 = ~1'b0 ;
  assign y12489 = ~n39309 ;
  assign y12490 = n39311 ;
  assign y12491 = ~n39312 ;
  assign y12492 = n39316 ;
  assign y12493 = n39317 ;
  assign y12494 = ~n39325 ;
  assign y12495 = n39326 ;
  assign y12496 = n39327 ;
  assign y12497 = ~1'b0 ;
  assign y12498 = ~n39329 ;
  assign y12499 = n39330 ;
  assign y12500 = ~n39337 ;
  assign y12501 = ~n39343 ;
  assign y12502 = ~n39344 ;
  assign y12503 = n39345 ;
  assign y12504 = ~n39347 ;
  assign y12505 = ~n39348 ;
  assign y12506 = n39350 ;
  assign y12507 = ~n39351 ;
  assign y12508 = ~n39353 ;
  assign y12509 = n39354 ;
  assign y12510 = n39356 ;
  assign y12511 = ~n39359 ;
  assign y12512 = ~n39361 ;
  assign y12513 = n39364 ;
  assign y12514 = n39368 ;
  assign y12515 = n39370 ;
  assign y12516 = n39371 ;
  assign y12517 = ~n39373 ;
  assign y12518 = n39374 ;
  assign y12519 = ~1'b0 ;
  assign y12520 = n39375 ;
  assign y12521 = ~n39377 ;
  assign y12522 = ~n39380 ;
  assign y12523 = ~1'b0 ;
  assign y12524 = ~n39381 ;
  assign y12525 = ~n39383 ;
  assign y12526 = n39384 ;
  assign y12527 = n39386 ;
  assign y12528 = ~1'b0 ;
  assign y12529 = ~n39387 ;
  assign y12530 = ~n39389 ;
  assign y12531 = ~n39390 ;
  assign y12532 = ~1'b0 ;
  assign y12533 = ~n39392 ;
  assign y12534 = n39396 ;
  assign y12535 = ~n39398 ;
  assign y12536 = n39400 ;
  assign y12537 = ~n39407 ;
  assign y12538 = n39411 ;
  assign y12539 = n39413 ;
  assign y12540 = ~1'b0 ;
  assign y12541 = n39419 ;
  assign y12542 = ~n39421 ;
  assign y12543 = ~n39427 ;
  assign y12544 = ~n39428 ;
  assign y12545 = n39433 ;
  assign y12546 = ~n39439 ;
  assign y12547 = ~n39442 ;
  assign y12548 = n39444 ;
  assign y12549 = ~n39446 ;
  assign y12550 = ~1'b0 ;
  assign y12551 = ~n39449 ;
  assign y12552 = n39452 ;
  assign y12553 = n31802 ;
  assign y12554 = n39453 ;
  assign y12555 = n39455 ;
  assign y12556 = ~n39461 ;
  assign y12557 = n39462 ;
  assign y12558 = ~n39466 ;
  assign y12559 = ~n39467 ;
  assign y12560 = ~n39479 ;
  assign y12561 = ~n39483 ;
  assign y12562 = n39489 ;
  assign y12563 = n39490 ;
  assign y12564 = ~1'b0 ;
  assign y12565 = ~1'b0 ;
  assign y12566 = ~1'b0 ;
  assign y12567 = ~n39494 ;
  assign y12568 = ~n39497 ;
  assign y12569 = ~n39498 ;
  assign y12570 = ~n39501 ;
  assign y12571 = ~n39502 ;
  assign y12572 = ~n39506 ;
  assign y12573 = ~n39507 ;
  assign y12574 = ~n39508 ;
  assign y12575 = n39511 ;
  assign y12576 = ~n39512 ;
  assign y12577 = n39516 ;
  assign y12578 = ~n39517 ;
  assign y12579 = ~n39526 ;
  assign y12580 = ~1'b0 ;
  assign y12581 = n39527 ;
  assign y12582 = ~n39528 ;
  assign y12583 = n39531 ;
  assign y12584 = ~1'b0 ;
  assign y12585 = n39533 ;
  assign y12586 = ~1'b0 ;
  assign y12587 = ~1'b0 ;
  assign y12588 = n39534 ;
  assign y12589 = ~n39536 ;
  assign y12590 = ~n39537 ;
  assign y12591 = ~n39542 ;
  assign y12592 = ~n39547 ;
  assign y12593 = n39549 ;
  assign y12594 = ~1'b0 ;
  assign y12595 = ~n39553 ;
  assign y12596 = n39556 ;
  assign y12597 = n39559 ;
  assign y12598 = n39562 ;
  assign y12599 = ~n39573 ;
  assign y12600 = ~n39576 ;
  assign y12601 = n39582 ;
  assign y12602 = ~1'b0 ;
  assign y12603 = n39586 ;
  assign y12604 = n39588 ;
  assign y12605 = ~n39593 ;
  assign y12606 = n39595 ;
  assign y12607 = ~n39596 ;
  assign y12608 = n39600 ;
  assign y12609 = ~n39603 ;
  assign y12610 = ~n39607 ;
  assign y12611 = ~n39608 ;
  assign y12612 = ~n39622 ;
  assign y12613 = n39623 ;
  assign y12614 = n39625 ;
  assign y12615 = ~n39629 ;
  assign y12616 = ~1'b0 ;
  assign y12617 = n9672 ;
  assign y12618 = n39631 ;
  assign y12619 = ~n39632 ;
  assign y12620 = ~n39638 ;
  assign y12621 = ~n39639 ;
  assign y12622 = ~n39640 ;
  assign y12623 = ~n39643 ;
  assign y12624 = ~n39646 ;
  assign y12625 = ~n39651 ;
  assign y12626 = ~n39658 ;
  assign y12627 = ~n39660 ;
  assign y12628 = n39663 ;
  assign y12629 = n39668 ;
  assign y12630 = n39669 ;
  assign y12631 = ~n39671 ;
  assign y12632 = n39673 ;
  assign y12633 = ~n39675 ;
  assign y12634 = ~n39679 ;
  assign y12635 = n39680 ;
  assign y12636 = ~n39681 ;
  assign y12637 = n39682 ;
  assign y12638 = n39683 ;
  assign y12639 = ~n39687 ;
  assign y12640 = n39689 ;
  assign y12641 = ~n39690 ;
  assign y12642 = n39696 ;
  assign y12643 = ~n39698 ;
  assign y12644 = n39702 ;
  assign y12645 = n39705 ;
  assign y12646 = n39709 ;
  assign y12647 = ~n39711 ;
  assign y12648 = n39714 ;
  assign y12649 = ~n5844 ;
  assign y12650 = n39717 ;
  assign y12651 = n39719 ;
  assign y12652 = n39724 ;
  assign y12653 = n39725 ;
  assign y12654 = ~1'b0 ;
  assign y12655 = ~n39726 ;
  assign y12656 = ~n39729 ;
  assign y12657 = ~n39732 ;
  assign y12658 = ~n39734 ;
  assign y12659 = n39735 ;
  assign y12660 = ~1'b0 ;
  assign y12661 = n39737 ;
  assign y12662 = ~1'b0 ;
  assign y12663 = ~n39741 ;
  assign y12664 = n39743 ;
  assign y12665 = ~n39745 ;
  assign y12666 = n39747 ;
  assign y12667 = ~n39749 ;
  assign y12668 = ~1'b0 ;
  assign y12669 = n1941 ;
  assign y12670 = ~n39753 ;
  assign y12671 = ~n39757 ;
  assign y12672 = n39760 ;
  assign y12673 = n39764 ;
  assign y12674 = ~n39765 ;
  assign y12675 = n39768 ;
  assign y12676 = ~n39769 ;
  assign y12677 = ~1'b0 ;
  assign y12678 = ~1'b0 ;
  assign y12679 = ~n39771 ;
  assign y12680 = ~n39772 ;
  assign y12681 = ~n39773 ;
  assign y12682 = n39781 ;
  assign y12683 = n39783 ;
  assign y12684 = ~n39784 ;
  assign y12685 = n39786 ;
  assign y12686 = ~n39791 ;
  assign y12687 = n39793 ;
  assign y12688 = n39801 ;
  assign y12689 = ~n39804 ;
  assign y12690 = n39807 ;
  assign y12691 = n39810 ;
  assign y12692 = ~n39811 ;
  assign y12693 = n39813 ;
  assign y12694 = ~n39817 ;
  assign y12695 = n39821 ;
  assign y12696 = n39822 ;
  assign y12697 = ~n39823 ;
  assign y12698 = n39826 ;
  assign y12699 = n39829 ;
  assign y12700 = ~n39832 ;
  assign y12701 = n39833 ;
  assign y12702 = ~n39834 ;
  assign y12703 = n39836 ;
  assign y12704 = n39840 ;
  assign y12705 = ~n39841 ;
  assign y12706 = n39844 ;
  assign y12707 = n39846 ;
  assign y12708 = ~n39847 ;
  assign y12709 = ~1'b0 ;
  assign y12710 = ~n39849 ;
  assign y12711 = n39852 ;
  assign y12712 = n39857 ;
  assign y12713 = ~n39859 ;
  assign y12714 = ~n39860 ;
  assign y12715 = n39868 ;
  assign y12716 = ~n39869 ;
  assign y12717 = ~n39873 ;
  assign y12718 = ~n39874 ;
  assign y12719 = ~1'b0 ;
  assign y12720 = ~n39875 ;
  assign y12721 = n39878 ;
  assign y12722 = ~1'b0 ;
  assign y12723 = ~1'b0 ;
  assign y12724 = ~1'b0 ;
  assign y12725 = ~n39879 ;
  assign y12726 = n39880 ;
  assign y12727 = n39888 ;
  assign y12728 = ~1'b0 ;
  assign y12729 = ~1'b0 ;
  assign y12730 = ~n39890 ;
  assign y12731 = ~n39895 ;
  assign y12732 = ~1'b0 ;
  assign y12733 = ~n39898 ;
  assign y12734 = ~n39900 ;
  assign y12735 = ~n39903 ;
  assign y12736 = ~n39905 ;
  assign y12737 = ~n39907 ;
  assign y12738 = ~n39910 ;
  assign y12739 = ~n39911 ;
  assign y12740 = ~n39914 ;
  assign y12741 = ~1'b0 ;
  assign y12742 = ~1'b0 ;
  assign y12743 = n39917 ;
  assign y12744 = ~n39920 ;
  assign y12745 = ~n39921 ;
  assign y12746 = n39922 ;
  assign y12747 = ~n39923 ;
  assign y12748 = ~n703 ;
  assign y12749 = ~n39927 ;
  assign y12750 = ~n39929 ;
  assign y12751 = ~1'b0 ;
  assign y12752 = ~1'b0 ;
  assign y12753 = ~n39932 ;
  assign y12754 = ~n39943 ;
  assign y12755 = ~n39946 ;
  assign y12756 = n39948 ;
  assign y12757 = n39949 ;
  assign y12758 = n39951 ;
  assign y12759 = ~n39954 ;
  assign y12760 = ~n39955 ;
  assign y12761 = n36198 ;
  assign y12762 = n39956 ;
  assign y12763 = ~1'b0 ;
  assign y12764 = n39958 ;
  assign y12765 = ~1'b0 ;
  assign y12766 = ~n39962 ;
  assign y12767 = ~n39963 ;
  assign y12768 = ~n39964 ;
  assign y12769 = n39968 ;
  assign y12770 = n39970 ;
  assign y12771 = n39973 ;
  assign y12772 = n39975 ;
  assign y12773 = n39978 ;
  assign y12774 = n39981 ;
  assign y12775 = n39982 ;
  assign y12776 = n39985 ;
  assign y12777 = ~n39987 ;
  assign y12778 = n39988 ;
  assign y12779 = ~n39991 ;
  assign y12780 = n39995 ;
  assign y12781 = n39997 ;
  assign y12782 = ~1'b0 ;
  assign y12783 = ~n39998 ;
  assign y12784 = ~1'b0 ;
  assign y12785 = n39999 ;
  assign y12786 = n40002 ;
  assign y12787 = n40004 ;
  assign y12788 = ~n40007 ;
  assign y12789 = ~n40008 ;
  assign y12790 = n40015 ;
  assign y12791 = n40016 ;
  assign y12792 = ~n40018 ;
  assign y12793 = ~1'b0 ;
  assign y12794 = ~1'b0 ;
  assign y12795 = ~n40022 ;
  assign y12796 = ~n40034 ;
  assign y12797 = n40035 ;
  assign y12798 = ~n40045 ;
  assign y12799 = ~n40050 ;
  assign y12800 = ~n40052 ;
  assign y12801 = n40054 ;
  assign y12802 = ~n40060 ;
  assign y12803 = ~n40062 ;
  assign y12804 = ~n40066 ;
  assign y12805 = n40067 ;
  assign y12806 = ~n40068 ;
  assign y12807 = n40071 ;
  assign y12808 = ~n40072 ;
  assign y12809 = ~1'b0 ;
  assign y12810 = ~n40074 ;
  assign y12811 = ~n40075 ;
  assign y12812 = ~1'b0 ;
  assign y12813 = ~n40076 ;
  assign y12814 = n40077 ;
  assign y12815 = n40078 ;
  assign y12816 = n40081 ;
  assign y12817 = ~n40083 ;
  assign y12818 = ~1'b0 ;
  assign y12819 = ~1'b0 ;
  assign y12820 = ~1'b0 ;
  assign y12821 = ~n40084 ;
  assign y12822 = n40085 ;
  assign y12823 = ~n40091 ;
  assign y12824 = n40098 ;
  assign y12825 = ~n40102 ;
  assign y12826 = n40106 ;
  assign y12827 = ~1'b0 ;
  assign y12828 = ~n40108 ;
  assign y12829 = n40110 ;
  assign y12830 = ~n40114 ;
  assign y12831 = n40115 ;
  assign y12832 = ~n40117 ;
  assign y12833 = ~n40118 ;
  assign y12834 = ~1'b0 ;
  assign y12835 = n40122 ;
  assign y12836 = ~n40126 ;
  assign y12837 = n40129 ;
  assign y12838 = ~n40132 ;
  assign y12839 = n40133 ;
  assign y12840 = ~n40139 ;
  assign y12841 = n40145 ;
  assign y12842 = ~1'b0 ;
  assign y12843 = ~1'b0 ;
  assign y12844 = ~1'b0 ;
  assign y12845 = n40150 ;
  assign y12846 = n16905 ;
  assign y12847 = ~n40151 ;
  assign y12848 = n40152 ;
  assign y12849 = ~n40157 ;
  assign y12850 = ~1'b0 ;
  assign y12851 = ~1'b0 ;
  assign y12852 = ~1'b0 ;
  assign y12853 = n40160 ;
  assign y12854 = n40162 ;
  assign y12855 = n40167 ;
  assign y12856 = ~n40171 ;
  assign y12857 = n40173 ;
  assign y12858 = n40175 ;
  assign y12859 = n40177 ;
  assign y12860 = n40182 ;
  assign y12861 = n40184 ;
  assign y12862 = n40185 ;
  assign y12863 = n40188 ;
  assign y12864 = ~n40194 ;
  assign y12865 = n40197 ;
  assign y12866 = ~n40200 ;
  assign y12867 = ~1'b0 ;
  assign y12868 = ~n40211 ;
  assign y12869 = ~n40214 ;
  assign y12870 = n40215 ;
  assign y12871 = ~n40220 ;
  assign y12872 = ~n40224 ;
  assign y12873 = n40226 ;
  assign y12874 = n40232 ;
  assign y12875 = ~n40235 ;
  assign y12876 = ~n40236 ;
  assign y12877 = ~n40237 ;
  assign y12878 = n40238 ;
  assign y12879 = n40243 ;
  assign y12880 = ~n40244 ;
  assign y12881 = n40245 ;
  assign y12882 = n40248 ;
  assign y12883 = ~n40250 ;
  assign y12884 = ~n40252 ;
  assign y12885 = n40254 ;
  assign y12886 = n40260 ;
  assign y12887 = n40261 ;
  assign y12888 = ~n40263 ;
  assign y12889 = n40266 ;
  assign y12890 = n40268 ;
  assign y12891 = ~1'b0 ;
  assign y12892 = ~n40269 ;
  assign y12893 = n40270 ;
  assign y12894 = n40273 ;
  assign y12895 = n40276 ;
  assign y12896 = ~n40280 ;
  assign y12897 = n40282 ;
  assign y12898 = n40283 ;
  assign y12899 = n40294 ;
  assign y12900 = n40295 ;
  assign y12901 = n40299 ;
  assign y12902 = ~1'b0 ;
  assign y12903 = n40300 ;
  assign y12904 = n40302 ;
  assign y12905 = ~1'b0 ;
  assign y12906 = ~n40308 ;
  assign y12907 = n40314 ;
  assign y12908 = ~n40315 ;
  assign y12909 = ~n40322 ;
  assign y12910 = ~n40325 ;
  assign y12911 = ~1'b0 ;
  assign y12912 = ~n40326 ;
  assign y12913 = ~n40328 ;
  assign y12914 = n40329 ;
  assign y12915 = ~n40330 ;
  assign y12916 = n40334 ;
  assign y12917 = ~1'b0 ;
  assign y12918 = ~n40335 ;
  assign y12919 = ~1'b0 ;
  assign y12920 = ~n40340 ;
  assign y12921 = n40344 ;
  assign y12922 = ~n40346 ;
  assign y12923 = ~n40349 ;
  assign y12924 = ~n40350 ;
  assign y12925 = ~n40352 ;
  assign y12926 = ~1'b0 ;
  assign y12927 = ~n40354 ;
  assign y12928 = n40355 ;
  assign y12929 = n40359 ;
  assign y12930 = ~n40361 ;
  assign y12931 = ~1'b0 ;
  assign y12932 = n40366 ;
  assign y12933 = ~n40374 ;
  assign y12934 = n40376 ;
  assign y12935 = ~n40378 ;
  assign y12936 = ~n40379 ;
  assign y12937 = ~1'b0 ;
  assign y12938 = n40384 ;
  assign y12939 = ~n40386 ;
  assign y12940 = n40387 ;
  assign y12941 = ~n40389 ;
  assign y12942 = ~n40390 ;
  assign y12943 = ~n40394 ;
  assign y12944 = n40397 ;
  assign y12945 = n40399 ;
  assign y12946 = ~1'b0 ;
  assign y12947 = n40401 ;
  assign y12948 = ~1'b0 ;
  assign y12949 = ~n40403 ;
  assign y12950 = ~n40404 ;
  assign y12951 = ~n40406 ;
  assign y12952 = n40414 ;
  assign y12953 = ~n40425 ;
  assign y12954 = ~n40428 ;
  assign y12955 = n40430 ;
  assign y12956 = ~1'b0 ;
  assign y12957 = ~n40434 ;
  assign y12958 = n40436 ;
  assign y12959 = n40437 ;
  assign y12960 = n40445 ;
  assign y12961 = ~n40447 ;
  assign y12962 = ~n40451 ;
  assign y12963 = n40452 ;
  assign y12964 = ~n40455 ;
  assign y12965 = ~n40456 ;
  assign y12966 = ~1'b0 ;
  assign y12967 = n40457 ;
  assign y12968 = n40461 ;
  assign y12969 = ~n40467 ;
  assign y12970 = n40468 ;
  assign y12971 = ~n40469 ;
  assign y12972 = ~n40470 ;
  assign y12973 = ~1'b0 ;
  assign y12974 = n40471 ;
  assign y12975 = n40475 ;
  assign y12976 = n40476 ;
  assign y12977 = n40480 ;
  assign y12978 = ~n40484 ;
  assign y12979 = ~n40486 ;
  assign y12980 = ~n40488 ;
  assign y12981 = ~1'b0 ;
  assign y12982 = n40491 ;
  assign y12983 = ~1'b0 ;
  assign y12984 = n40496 ;
  assign y12985 = ~n40503 ;
  assign y12986 = n40506 ;
  assign y12987 = n40509 ;
  assign y12988 = ~n40515 ;
  assign y12989 = ~n40516 ;
  assign y12990 = ~n40519 ;
  assign y12991 = n40523 ;
  assign y12992 = n40528 ;
  assign y12993 = ~n40529 ;
  assign y12994 = ~n40530 ;
  assign y12995 = n40532 ;
  assign y12996 = ~n40535 ;
  assign y12997 = ~n40537 ;
  assign y12998 = n40542 ;
  assign y12999 = ~n40544 ;
  assign y13000 = ~n40546 ;
  assign y13001 = n40550 ;
  assign y13002 = ~n40555 ;
  assign y13003 = n40557 ;
  assign y13004 = ~n40558 ;
  assign y13005 = ~n40565 ;
  assign y13006 = ~1'b0 ;
  assign y13007 = ~n40568 ;
  assign y13008 = n40572 ;
  assign y13009 = n40577 ;
  assign y13010 = n40578 ;
  assign y13011 = ~n40588 ;
  assign y13012 = n40589 ;
  assign y13013 = n20279 ;
  assign y13014 = ~n40592 ;
  assign y13015 = n40594 ;
  assign y13016 = ~1'b0 ;
  assign y13017 = ~n40597 ;
  assign y13018 = n40598 ;
  assign y13019 = n40600 ;
  assign y13020 = ~n40601 ;
  assign y13021 = n40606 ;
  assign y13022 = n40609 ;
  assign y13023 = n40611 ;
  assign y13024 = ~n40613 ;
  assign y13025 = ~n40616 ;
  assign y13026 = ~n40622 ;
  assign y13027 = n40627 ;
  assign y13028 = n40631 ;
  assign y13029 = n40639 ;
  assign y13030 = n40643 ;
  assign y13031 = n1751 ;
  assign y13032 = n40645 ;
  assign y13033 = ~n40648 ;
  assign y13034 = ~n40651 ;
  assign y13035 = ~n40656 ;
  assign y13036 = ~n40657 ;
  assign y13037 = ~n40660 ;
  assign y13038 = n40662 ;
  assign y13039 = n40668 ;
  assign y13040 = n40673 ;
  assign y13041 = ~n40677 ;
  assign y13042 = ~n40679 ;
  assign y13043 = ~1'b0 ;
  assign y13044 = n40684 ;
  assign y13045 = ~n40693 ;
  assign y13046 = n40696 ;
  assign y13047 = n40698 ;
  assign y13048 = ~n40702 ;
  assign y13049 = n40707 ;
  assign y13050 = ~n40712 ;
  assign y13051 = ~n40716 ;
  assign y13052 = n40717 ;
  assign y13053 = ~n40718 ;
  assign y13054 = ~n40720 ;
  assign y13055 = ~n40723 ;
  assign y13056 = n40725 ;
  assign y13057 = ~1'b0 ;
  assign y13058 = n40730 ;
  assign y13059 = ~n40735 ;
  assign y13060 = n40740 ;
  assign y13061 = n40749 ;
  assign y13062 = n40751 ;
  assign y13063 = ~1'b0 ;
  assign y13064 = ~n40753 ;
  assign y13065 = ~n40755 ;
  assign y13066 = ~n40757 ;
  assign y13067 = ~n40761 ;
  assign y13068 = ~n40762 ;
  assign y13069 = ~n40763 ;
  assign y13070 = ~n40767 ;
  assign y13071 = ~n40770 ;
  assign y13072 = ~1'b0 ;
  assign y13073 = n40780 ;
  assign y13074 = ~n40782 ;
  assign y13075 = ~n40783 ;
  assign y13076 = n40786 ;
  assign y13077 = ~n40789 ;
  assign y13078 = ~n40795 ;
  assign y13079 = ~1'b0 ;
  assign y13080 = ~n40797 ;
  assign y13081 = n40802 ;
  assign y13082 = ~n40803 ;
  assign y13083 = ~n1732 ;
  assign y13084 = ~n40806 ;
  assign y13085 = ~n40809 ;
  assign y13086 = ~n40810 ;
  assign y13087 = n40814 ;
  assign y13088 = ~n40820 ;
  assign y13089 = n40826 ;
  assign y13090 = ~n7474 ;
  assign y13091 = ~n40829 ;
  assign y13092 = n40830 ;
  assign y13093 = n40831 ;
  assign y13094 = n40835 ;
  assign y13095 = ~1'b0 ;
  assign y13096 = ~n40836 ;
  assign y13097 = n40839 ;
  assign y13098 = n40840 ;
  assign y13099 = ~n40848 ;
  assign y13100 = n40852 ;
  assign y13101 = n40855 ;
  assign y13102 = n40858 ;
  assign y13103 = n40859 ;
  assign y13104 = n40863 ;
  assign y13105 = ~n40864 ;
  assign y13106 = ~1'b0 ;
  assign y13107 = ~n40865 ;
  assign y13108 = n40867 ;
  assign y13109 = n40869 ;
  assign y13110 = ~n40872 ;
  assign y13111 = n40875 ;
  assign y13112 = ~n40878 ;
  assign y13113 = ~1'b0 ;
  assign y13114 = n40883 ;
  assign y13115 = ~1'b0 ;
  assign y13116 = ~n40886 ;
  assign y13117 = n40895 ;
  assign y13118 = n40896 ;
  assign y13119 = ~n40898 ;
  assign y13120 = n40900 ;
  assign y13121 = n40905 ;
  assign y13122 = n40907 ;
  assign y13123 = ~n40913 ;
  assign y13124 = ~n40916 ;
  assign y13125 = ~n40920 ;
  assign y13126 = ~n40922 ;
  assign y13127 = ~n40925 ;
  assign y13128 = n40926 ;
  assign y13129 = n40928 ;
  assign y13130 = ~n40929 ;
  assign y13131 = ~n40931 ;
  assign y13132 = ~n40933 ;
  assign y13133 = ~1'b0 ;
  assign y13134 = ~1'b0 ;
  assign y13135 = ~n40935 ;
  assign y13136 = n40936 ;
  assign y13137 = n40937 ;
  assign y13138 = ~n40938 ;
  assign y13139 = n40940 ;
  assign y13140 = ~n40947 ;
  assign y13141 = ~n30195 ;
  assign y13142 = n40951 ;
  assign y13143 = ~1'b0 ;
  assign y13144 = ~1'b0 ;
  assign y13145 = ~n40954 ;
  assign y13146 = n40955 ;
  assign y13147 = ~n40957 ;
  assign y13148 = ~n40960 ;
  assign y13149 = ~n40966 ;
  assign y13150 = ~1'b0 ;
  assign y13151 = ~1'b0 ;
  assign y13152 = n40971 ;
  assign y13153 = ~n40974 ;
  assign y13154 = ~n40975 ;
  assign y13155 = ~n4702 ;
  assign y13156 = n40976 ;
  assign y13157 = n40982 ;
  assign y13158 = n40984 ;
  assign y13159 = ~n40988 ;
  assign y13160 = ~1'b0 ;
  assign y13161 = n40990 ;
  assign y13162 = ~n40991 ;
  assign y13163 = n40996 ;
  assign y13164 = ~1'b0 ;
  assign y13165 = ~1'b0 ;
  assign y13166 = n40998 ;
  assign y13167 = n41000 ;
  assign y13168 = ~n41002 ;
  assign y13169 = n41003 ;
  assign y13170 = n41005 ;
  assign y13171 = n6761 ;
  assign y13172 = n41007 ;
  assign y13173 = ~n41009 ;
  assign y13174 = ~n41012 ;
  assign y13175 = ~1'b0 ;
  assign y13176 = ~1'b0 ;
  assign y13177 = n41013 ;
  assign y13178 = n41014 ;
  assign y13179 = n41015 ;
  assign y13180 = n41016 ;
  assign y13181 = ~n15454 ;
  assign y13182 = ~1'b0 ;
  assign y13183 = n41018 ;
  assign y13184 = ~n41021 ;
  assign y13185 = ~n41026 ;
  assign y13186 = ~n41027 ;
  assign y13187 = ~n41028 ;
  assign y13188 = n41030 ;
  assign y13189 = n41031 ;
  assign y13190 = ~n41034 ;
  assign y13191 = ~n41040 ;
  assign y13192 = ~n41042 ;
  assign y13193 = ~n41044 ;
  assign y13194 = ~n41046 ;
  assign y13195 = ~n41051 ;
  assign y13196 = n41052 ;
  assign y13197 = n41054 ;
  assign y13198 = n41058 ;
  assign y13199 = n41059 ;
  assign y13200 = ~n41066 ;
  assign y13201 = n41068 ;
  assign y13202 = n41069 ;
  assign y13203 = n41070 ;
  assign y13204 = ~n41072 ;
  assign y13205 = n41075 ;
  assign y13206 = ~1'b0 ;
  assign y13207 = ~n41078 ;
  assign y13208 = ~n41080 ;
  assign y13209 = n41083 ;
  assign y13210 = n41084 ;
  assign y13211 = n41086 ;
  assign y13212 = ~n41094 ;
  assign y13213 = n41097 ;
  assign y13214 = n41100 ;
  assign y13215 = ~n41104 ;
  assign y13216 = n41105 ;
  assign y13217 = ~n41108 ;
  assign y13218 = ~n41110 ;
  assign y13219 = ~1'b0 ;
  assign y13220 = ~1'b0 ;
  assign y13221 = ~1'b0 ;
  assign y13222 = ~1'b0 ;
  assign y13223 = ~n41112 ;
  assign y13224 = ~n41117 ;
  assign y13225 = ~n41123 ;
  assign y13226 = ~n41125 ;
  assign y13227 = ~n41126 ;
  assign y13228 = ~n41128 ;
  assign y13229 = ~n41134 ;
  assign y13230 = n41135 ;
  assign y13231 = ~n41137 ;
  assign y13232 = ~1'b0 ;
  assign y13233 = n41139 ;
  assign y13234 = ~n41145 ;
  assign y13235 = ~n41149 ;
  assign y13236 = ~n41154 ;
  assign y13237 = n41163 ;
  assign y13238 = ~n41164 ;
  assign y13239 = ~1'b0 ;
  assign y13240 = ~n41166 ;
  assign y13241 = n41167 ;
  assign y13242 = n41175 ;
  assign y13243 = ~n41176 ;
  assign y13244 = ~n41177 ;
  assign y13245 = ~1'b0 ;
  assign y13246 = n41184 ;
  assign y13247 = ~n41186 ;
  assign y13248 = ~n41190 ;
  assign y13249 = ~n41195 ;
  assign y13250 = ~n41196 ;
  assign y13251 = n41200 ;
  assign y13252 = n5254 ;
  assign y13253 = ~n41202 ;
  assign y13254 = n41209 ;
  assign y13255 = ~n41213 ;
  assign y13256 = n41217 ;
  assign y13257 = ~1'b0 ;
  assign y13258 = ~n41223 ;
  assign y13259 = ~1'b0 ;
  assign y13260 = ~n41224 ;
  assign y13261 = ~n41227 ;
  assign y13262 = n41229 ;
  assign y13263 = n41239 ;
  assign y13264 = n41242 ;
  assign y13265 = ~1'b0 ;
  assign y13266 = ~n41249 ;
  assign y13267 = n41254 ;
  assign y13268 = ~n41257 ;
  assign y13269 = n41259 ;
  assign y13270 = n41260 ;
  assign y13271 = n41262 ;
  assign y13272 = ~n41263 ;
  assign y13273 = ~n41266 ;
  assign y13274 = n41273 ;
  assign y13275 = ~n41274 ;
  assign y13276 = ~n41275 ;
  assign y13277 = n41281 ;
  assign y13278 = n41283 ;
  assign y13279 = n41286 ;
  assign y13280 = n41287 ;
  assign y13281 = n41288 ;
  assign y13282 = ~1'b0 ;
  assign y13283 = n41290 ;
  assign y13284 = ~1'b0 ;
  assign y13285 = n41292 ;
  assign y13286 = n41299 ;
  assign y13287 = ~n41303 ;
  assign y13288 = ~n41306 ;
  assign y13289 = n41308 ;
  assign y13290 = ~n41309 ;
  assign y13291 = ~n41311 ;
  assign y13292 = ~n36137 ;
  assign y13293 = n41312 ;
  assign y13294 = ~n41313 ;
  assign y13295 = ~n41317 ;
  assign y13296 = ~n41318 ;
  assign y13297 = ~n41333 ;
  assign y13298 = ~n41337 ;
  assign y13299 = ~n41338 ;
  assign y13300 = ~n41340 ;
  assign y13301 = n41344 ;
  assign y13302 = n41345 ;
  assign y13303 = ~n41346 ;
  assign y13304 = n41353 ;
  assign y13305 = n41354 ;
  assign y13306 = n41355 ;
  assign y13307 = n41358 ;
  assign y13308 = n41361 ;
  assign y13309 = ~1'b0 ;
  assign y13310 = ~n41369 ;
  assign y13311 = ~n41371 ;
  assign y13312 = ~1'b0 ;
  assign y13313 = ~n41372 ;
  assign y13314 = ~n41373 ;
  assign y13315 = ~n41381 ;
  assign y13316 = n41383 ;
  assign y13317 = ~1'b0 ;
  assign y13318 = ~1'b0 ;
  assign y13319 = ~1'b0 ;
  assign y13320 = ~1'b0 ;
  assign y13321 = ~n41387 ;
  assign y13322 = n41391 ;
  assign y13323 = ~1'b0 ;
  assign y13324 = ~n41393 ;
  assign y13325 = ~n41395 ;
  assign y13326 = ~n41398 ;
  assign y13327 = ~n41400 ;
  assign y13328 = n41402 ;
  assign y13329 = ~n41409 ;
  assign y13330 = ~n41410 ;
  assign y13331 = ~1'b0 ;
  assign y13332 = n41415 ;
  assign y13333 = n41419 ;
  assign y13334 = n41425 ;
  assign y13335 = n41427 ;
  assign y13336 = n41429 ;
  assign y13337 = ~n41436 ;
  assign y13338 = ~1'b0 ;
  assign y13339 = n41437 ;
  assign y13340 = n41438 ;
  assign y13341 = n41439 ;
  assign y13342 = n41441 ;
  assign y13343 = n41446 ;
  assign y13344 = n41448 ;
  assign y13345 = ~n41454 ;
  assign y13346 = n41456 ;
  assign y13347 = ~1'b0 ;
  assign y13348 = ~1'b0 ;
  assign y13349 = ~n41459 ;
  assign y13350 = n41462 ;
  assign y13351 = ~n41463 ;
  assign y13352 = ~n41464 ;
  assign y13353 = n41465 ;
  assign y13354 = n41466 ;
  assign y13355 = ~n41467 ;
  assign y13356 = ~n41472 ;
  assign y13357 = ~n41476 ;
  assign y13358 = n41479 ;
  assign y13359 = ~n41481 ;
  assign y13360 = n41486 ;
  assign y13361 = ~n41487 ;
  assign y13362 = ~n41490 ;
  assign y13363 = ~n41493 ;
  assign y13364 = ~n41494 ;
  assign y13365 = n41497 ;
  assign y13366 = n41498 ;
  assign y13367 = n33033 ;
  assign y13368 = ~n41499 ;
  assign y13369 = ~n41503 ;
  assign y13370 = ~n41507 ;
  assign y13371 = ~n41511 ;
  assign y13372 = ~n41512 ;
  assign y13373 = n41515 ;
  assign y13374 = ~n41517 ;
  assign y13375 = n41518 ;
  assign y13376 = ~1'b0 ;
  assign y13377 = n41519 ;
  assign y13378 = n41521 ;
  assign y13379 = ~n41524 ;
  assign y13380 = n41528 ;
  assign y13381 = ~n41529 ;
  assign y13382 = n41532 ;
  assign y13383 = ~n41537 ;
  assign y13384 = ~n33025 ;
  assign y13385 = ~1'b0 ;
  assign y13386 = ~n41540 ;
  assign y13387 = ~n41541 ;
  assign y13388 = n41542 ;
  assign y13389 = n41544 ;
  assign y13390 = ~n41545 ;
  assign y13391 = n41546 ;
  assign y13392 = ~1'b0 ;
  assign y13393 = n41554 ;
  assign y13394 = n41555 ;
  assign y13395 = ~n41556 ;
  assign y13396 = ~n41563 ;
  assign y13397 = n41566 ;
  assign y13398 = n41570 ;
  assign y13399 = ~n41576 ;
  assign y13400 = ~1'b0 ;
  assign y13401 = n41584 ;
  assign y13402 = n41585 ;
  assign y13403 = n41587 ;
  assign y13404 = n41595 ;
  assign y13405 = n41597 ;
  assign y13406 = ~n41598 ;
  assign y13407 = ~1'b0 ;
  assign y13408 = ~n41600 ;
  assign y13409 = n41602 ;
  assign y13410 = ~n41603 ;
  assign y13411 = ~n41609 ;
  assign y13412 = ~n41610 ;
  assign y13413 = ~n41611 ;
  assign y13414 = n41615 ;
  assign y13415 = n41617 ;
  assign y13416 = ~n41625 ;
  assign y13417 = ~n41627 ;
  assign y13418 = ~1'b0 ;
  assign y13419 = ~n41628 ;
  assign y13420 = n41629 ;
  assign y13421 = n41633 ;
  assign y13422 = ~n41637 ;
  assign y13423 = n41639 ;
  assign y13424 = ~n41643 ;
  assign y13425 = n41645 ;
  assign y13426 = ~1'b0 ;
  assign y13427 = ~n41648 ;
  assign y13428 = n41649 ;
  assign y13429 = ~n41650 ;
  assign y13430 = ~n41653 ;
  assign y13431 = ~n41654 ;
  assign y13432 = ~n41657 ;
  assign y13433 = n41662 ;
  assign y13434 = ~1'b0 ;
  assign y13435 = ~n41667 ;
  assign y13436 = ~n41670 ;
  assign y13437 = n41674 ;
  assign y13438 = ~n41675 ;
  assign y13439 = n41676 ;
  assign y13440 = ~1'b0 ;
  assign y13441 = n41679 ;
  assign y13442 = n41680 ;
  assign y13443 = ~n1196 ;
  assign y13444 = n41684 ;
  assign y13445 = ~n41687 ;
  assign y13446 = n41690 ;
  assign y13447 = ~n41691 ;
  assign y13448 = n41693 ;
  assign y13449 = n34707 ;
  assign y13450 = n41696 ;
  assign y13451 = n41698 ;
  assign y13452 = ~n41700 ;
  assign y13453 = n41704 ;
  assign y13454 = ~n41705 ;
  assign y13455 = ~n41707 ;
  assign y13456 = n41708 ;
  assign y13457 = n41710 ;
  assign y13458 = ~1'b0 ;
  assign y13459 = ~1'b0 ;
  assign y13460 = ~n41711 ;
  assign y13461 = ~1'b0 ;
  assign y13462 = ~n41714 ;
  assign y13463 = ~n41715 ;
  assign y13464 = ~n41717 ;
  assign y13465 = ~1'b0 ;
  assign y13466 = ~1'b0 ;
  assign y13467 = ~1'b0 ;
  assign y13468 = n41720 ;
  assign y13469 = ~n41725 ;
  assign y13470 = ~n41728 ;
  assign y13471 = n41730 ;
  assign y13472 = ~n41731 ;
  assign y13473 = ~1'b0 ;
  assign y13474 = ~n41736 ;
  assign y13475 = n41738 ;
  assign y13476 = ~1'b0 ;
  assign y13477 = ~n41740 ;
  assign y13478 = ~n41744 ;
  assign y13479 = n41748 ;
  assign y13480 = ~n41751 ;
  assign y13481 = ~n41755 ;
  assign y13482 = n41758 ;
  assign y13483 = ~1'b0 ;
  assign y13484 = ~1'b0 ;
  assign y13485 = ~n41764 ;
  assign y13486 = n41766 ;
  assign y13487 = ~n41769 ;
  assign y13488 = n41771 ;
  assign y13489 = ~n41776 ;
  assign y13490 = n41781 ;
  assign y13491 = ~n41783 ;
  assign y13492 = ~n41787 ;
  assign y13493 = ~n41790 ;
  assign y13494 = n41792 ;
  assign y13495 = ~n41793 ;
  assign y13496 = n41794 ;
  assign y13497 = n41795 ;
  assign y13498 = n41796 ;
  assign y13499 = n41799 ;
  assign y13500 = ~n41804 ;
  assign y13501 = ~n41807 ;
  assign y13502 = ~1'b0 ;
  assign y13503 = ~n41809 ;
  assign y13504 = ~n41812 ;
  assign y13505 = ~n41817 ;
  assign y13506 = n41818 ;
  assign y13507 = n41821 ;
  assign y13508 = ~n41824 ;
  assign y13509 = ~1'b0 ;
  assign y13510 = ~n41825 ;
  assign y13511 = ~n41826 ;
  assign y13512 = ~1'b0 ;
  assign y13513 = ~n41830 ;
  assign y13514 = ~n41832 ;
  assign y13515 = n41839 ;
  assign y13516 = ~n41840 ;
  assign y13517 = ~1'b0 ;
  assign y13518 = n41844 ;
  assign y13519 = ~n41848 ;
  assign y13520 = ~n41851 ;
  assign y13521 = n41855 ;
  assign y13522 = ~n41860 ;
  assign y13523 = ~n41862 ;
  assign y13524 = ~n41863 ;
  assign y13525 = n41864 ;
  assign y13526 = ~n41867 ;
  assign y13527 = ~1'b0 ;
  assign y13528 = ~1'b0 ;
  assign y13529 = n41869 ;
  assign y13530 = ~n41871 ;
  assign y13531 = n41872 ;
  assign y13532 = ~n41876 ;
  assign y13533 = n41884 ;
  assign y13534 = ~n41888 ;
  assign y13535 = ~n41895 ;
  assign y13536 = ~n41897 ;
  assign y13537 = ~1'b0 ;
  assign y13538 = ~n41899 ;
  assign y13539 = ~n41901 ;
  assign y13540 = ~n41902 ;
  assign y13541 = n41903 ;
  assign y13542 = n41904 ;
  assign y13543 = ~1'b0 ;
  assign y13544 = ~n41906 ;
  assign y13545 = n41907 ;
  assign y13546 = n41913 ;
  assign y13547 = n41914 ;
  assign y13548 = ~n41916 ;
  assign y13549 = n41917 ;
  assign y13550 = n41920 ;
  assign y13551 = ~n41922 ;
  assign y13552 = ~n41927 ;
  assign y13553 = ~n41928 ;
  assign y13554 = ~n41931 ;
  assign y13555 = n41932 ;
  assign y13556 = n41938 ;
  assign y13557 = ~n41944 ;
  assign y13558 = n41950 ;
  assign y13559 = ~n41954 ;
  assign y13560 = n41955 ;
  assign y13561 = n41957 ;
  assign y13562 = ~n41958 ;
  assign y13563 = n41960 ;
  assign y13564 = ~n41964 ;
  assign y13565 = ~n41970 ;
  assign y13566 = n41971 ;
  assign y13567 = ~n41977 ;
  assign y13568 = ~1'b0 ;
  assign y13569 = ~n41979 ;
  assign y13570 = n41981 ;
  assign y13571 = ~n41982 ;
  assign y13572 = n41984 ;
  assign y13573 = ~n41985 ;
  assign y13574 = n41994 ;
  assign y13575 = n41995 ;
  assign y13576 = ~n42000 ;
  assign y13577 = n42005 ;
  assign y13578 = ~n42008 ;
  assign y13579 = ~n42009 ;
  assign y13580 = n42010 ;
  assign y13581 = ~n42013 ;
  assign y13582 = n42016 ;
  assign y13583 = ~n42019 ;
  assign y13584 = n42022 ;
  assign y13585 = ~1'b0 ;
  assign y13586 = n42025 ;
  assign y13587 = n35895 ;
  assign y13588 = ~n42026 ;
  assign y13589 = ~n42031 ;
  assign y13590 = ~n42034 ;
  assign y13591 = ~n42035 ;
  assign y13592 = ~1'b0 ;
  assign y13593 = ~1'b0 ;
  assign y13594 = ~1'b0 ;
  assign y13595 = ~1'b0 ;
  assign y13596 = ~n42037 ;
  assign y13597 = ~n42038 ;
  assign y13598 = ~n42041 ;
  assign y13599 = ~n24620 ;
  assign y13600 = n42045 ;
  assign y13601 = ~n42048 ;
  assign y13602 = ~1'b0 ;
  assign y13603 = ~n42050 ;
  assign y13604 = n42052 ;
  assign y13605 = ~n42053 ;
  assign y13606 = n42058 ;
  assign y13607 = ~n42062 ;
  assign y13608 = n42063 ;
  assign y13609 = ~n42067 ;
  assign y13610 = ~1'b0 ;
  assign y13611 = ~n42068 ;
  assign y13612 = n42069 ;
  assign y13613 = ~n42075 ;
  assign y13614 = n42080 ;
  assign y13615 = n42083 ;
  assign y13616 = n42085 ;
  assign y13617 = ~n42087 ;
  assign y13618 = 1'b0 ;
  assign y13619 = ~n42089 ;
  assign y13620 = ~1'b0 ;
  assign y13621 = n42090 ;
  assign y13622 = ~n42092 ;
  assign y13623 = ~n42094 ;
  assign y13624 = ~n42097 ;
  assign y13625 = ~n42098 ;
  assign y13626 = ~n42106 ;
  assign y13627 = n36071 ;
  assign y13628 = ~n42110 ;
  assign y13629 = n42111 ;
  assign y13630 = ~n42112 ;
  assign y13631 = n42113 ;
  assign y13632 = ~n42114 ;
  assign y13633 = ~n42119 ;
  assign y13634 = n42122 ;
  assign y13635 = n42126 ;
  assign y13636 = ~1'b0 ;
  assign y13637 = n42130 ;
  assign y13638 = n42132 ;
  assign y13639 = n42133 ;
  assign y13640 = ~n42135 ;
  assign y13641 = n42136 ;
  assign y13642 = ~n42137 ;
  assign y13643 = ~n42138 ;
  assign y13644 = ~1'b0 ;
  assign y13645 = n42140 ;
  assign y13646 = n42143 ;
  assign y13647 = ~1'b0 ;
  assign y13648 = ~n42149 ;
  assign y13649 = ~n42152 ;
  assign y13650 = n42153 ;
  assign y13651 = n42155 ;
  assign y13652 = ~n42156 ;
  assign y13653 = ~n42157 ;
  assign y13654 = ~1'b0 ;
  assign y13655 = n42158 ;
  assign y13656 = n42165 ;
  assign y13657 = ~1'b0 ;
  assign y13658 = ~n42169 ;
  assign y13659 = n42171 ;
  assign y13660 = ~n42174 ;
  assign y13661 = ~n42177 ;
  assign y13662 = n42180 ;
  assign y13663 = ~n42182 ;
  assign y13664 = n42184 ;
  assign y13665 = n3978 ;
  assign y13666 = ~n42185 ;
  assign y13667 = ~n42189 ;
  assign y13668 = n42191 ;
  assign y13669 = ~1'b0 ;
  assign y13670 = n42192 ;
  assign y13671 = ~n42194 ;
  assign y13672 = ~1'b0 ;
  assign y13673 = ~n42197 ;
  assign y13674 = n42198 ;
  assign y13675 = n42203 ;
  assign y13676 = n42204 ;
  assign y13677 = ~n42205 ;
  assign y13678 = ~1'b0 ;
  assign y13679 = n42209 ;
  assign y13680 = ~n42211 ;
  assign y13681 = ~1'b0 ;
  assign y13682 = ~n42217 ;
  assign y13683 = n42219 ;
  assign y13684 = n42220 ;
  assign y13685 = ~n42231 ;
  assign y13686 = n42236 ;
  assign y13687 = n42237 ;
  assign y13688 = ~1'b0 ;
  assign y13689 = ~n42247 ;
  assign y13690 = ~n42248 ;
  assign y13691 = ~n42250 ;
  assign y13692 = ~n42252 ;
  assign y13693 = ~n42253 ;
  assign y13694 = n42254 ;
  assign y13695 = n42255 ;
  assign y13696 = n42257 ;
  assign y13697 = n42258 ;
  assign y13698 = ~1'b0 ;
  assign y13699 = n42261 ;
  assign y13700 = ~n42262 ;
  assign y13701 = n42263 ;
  assign y13702 = n42264 ;
  assign y13703 = ~n42268 ;
  assign y13704 = n42269 ;
  assign y13705 = ~n42271 ;
  assign y13706 = ~n42274 ;
  assign y13707 = n42277 ;
  assign y13708 = ~1'b0 ;
  assign y13709 = ~n42284 ;
  assign y13710 = ~n42289 ;
  assign y13711 = n42291 ;
  assign y13712 = n42292 ;
  assign y13713 = n42293 ;
  assign y13714 = n42297 ;
  assign y13715 = ~n42300 ;
  assign y13716 = n644 ;
  assign y13717 = ~n42303 ;
  assign y13718 = ~n42307 ;
  assign y13719 = n42309 ;
  assign y13720 = n42310 ;
  assign y13721 = ~n42314 ;
  assign y13722 = ~n42315 ;
  assign y13723 = ~n2801 ;
  assign y13724 = n42318 ;
  assign y13725 = ~n42321 ;
  assign y13726 = n42330 ;
  assign y13727 = ~n42335 ;
  assign y13728 = n42339 ;
  assign y13729 = ~n42340 ;
  assign y13730 = n42344 ;
  assign y13731 = ~1'b0 ;
  assign y13732 = ~n42347 ;
  assign y13733 = ~n12574 ;
  assign y13734 = ~1'b0 ;
  assign y13735 = n42350 ;
  assign y13736 = ~n42355 ;
  assign y13737 = ~n24926 ;
  assign y13738 = n42356 ;
  assign y13739 = n42358 ;
  assign y13740 = ~1'b0 ;
  assign y13741 = n42361 ;
  assign y13742 = n42365 ;
  assign y13743 = n42366 ;
  assign y13744 = n42370 ;
  assign y13745 = ~n42375 ;
  assign y13746 = ~1'b0 ;
  assign y13747 = ~1'b0 ;
  assign y13748 = n42378 ;
  assign y13749 = n42382 ;
  assign y13750 = ~n42383 ;
  assign y13751 = n42385 ;
  assign y13752 = n42390 ;
  assign y13753 = n42393 ;
  assign y13754 = n42396 ;
  assign y13755 = ~1'b0 ;
  assign y13756 = ~1'b0 ;
  assign y13757 = ~n42397 ;
  assign y13758 = ~n42402 ;
  assign y13759 = n42405 ;
  assign y13760 = ~n42407 ;
  assign y13761 = ~1'b0 ;
  assign y13762 = n42408 ;
  assign y13763 = n42411 ;
  assign y13764 = 1'b0 ;
  assign y13765 = ~n42413 ;
  assign y13766 = n42414 ;
  assign y13767 = n42417 ;
  assign y13768 = ~n42418 ;
  assign y13769 = ~n42420 ;
  assign y13770 = ~n42423 ;
  assign y13771 = ~n42430 ;
  assign y13772 = n42432 ;
  assign y13773 = n42433 ;
  assign y13774 = ~n42435 ;
  assign y13775 = ~n42436 ;
  assign y13776 = ~n42437 ;
  assign y13777 = ~1'b0 ;
  assign y13778 = ~n42439 ;
  assign y13779 = ~n42441 ;
  assign y13780 = ~n42445 ;
  assign y13781 = ~1'b0 ;
  assign y13782 = n42448 ;
  assign y13783 = n42452 ;
  assign y13784 = ~n42456 ;
  assign y13785 = n42457 ;
  assign y13786 = ~n42458 ;
  assign y13787 = ~n42459 ;
  assign y13788 = n42461 ;
  assign y13789 = ~n42464 ;
  assign y13790 = ~1'b0 ;
  assign y13791 = ~1'b0 ;
  assign y13792 = ~n42465 ;
  assign y13793 = n42466 ;
  assign y13794 = ~n42467 ;
  assign y13795 = ~n42469 ;
  assign y13796 = ~n42471 ;
  assign y13797 = ~n42475 ;
  assign y13798 = ~n42476 ;
  assign y13799 = n42478 ;
  assign y13800 = n42480 ;
  assign y13801 = 1'b0 ;
  assign y13802 = ~n42486 ;
  assign y13803 = ~n42496 ;
  assign y13804 = n42498 ;
  assign y13805 = ~n42502 ;
  assign y13806 = n42504 ;
  assign y13807 = ~n42505 ;
  assign y13808 = n42506 ;
  assign y13809 = ~n42514 ;
  assign y13810 = ~n42517 ;
  assign y13811 = ~n42519 ;
  assign y13812 = ~1'b0 ;
  assign y13813 = ~n42520 ;
  assign y13814 = ~1'b0 ;
  assign y13815 = 1'b0 ;
  assign y13816 = ~n42521 ;
  assign y13817 = ~n42524 ;
  assign y13818 = n42526 ;
  assign y13819 = ~1'b0 ;
  assign y13820 = ~1'b0 ;
  assign y13821 = ~n42530 ;
  assign y13822 = ~n42535 ;
  assign y13823 = ~n42536 ;
  assign y13824 = n42540 ;
  assign y13825 = ~n42543 ;
  assign y13826 = ~1'b0 ;
  assign y13827 = ~n42545 ;
  assign y13828 = ~n42550 ;
  assign y13829 = ~n42557 ;
  assign y13830 = n42561 ;
  assign y13831 = n42563 ;
  assign y13832 = n42564 ;
  assign y13833 = ~1'b0 ;
  assign y13834 = ~n42566 ;
  assign y13835 = ~n42567 ;
  assign y13836 = n42570 ;
  assign y13837 = n42576 ;
  assign y13838 = ~n42577 ;
  assign y13839 = n42579 ;
  assign y13840 = ~n42582 ;
  assign y13841 = ~n42584 ;
  assign y13842 = ~1'b0 ;
  assign y13843 = ~n42587 ;
  assign y13844 = ~n42590 ;
  assign y13845 = ~n42591 ;
  assign y13846 = n42592 ;
  assign y13847 = ~n42594 ;
  assign y13848 = n42595 ;
  assign y13849 = n42596 ;
  assign y13850 = ~1'b0 ;
  assign y13851 = ~n42599 ;
  assign y13852 = ~1'b0 ;
  assign y13853 = ~1'b0 ;
  assign y13854 = n42601 ;
  assign y13855 = n42610 ;
  assign y13856 = ~n42613 ;
  assign y13857 = n42614 ;
  assign y13858 = n42618 ;
  assign y13859 = ~n42622 ;
  assign y13860 = ~n42624 ;
  assign y13861 = ~n42628 ;
  assign y13862 = ~1'b0 ;
  assign y13863 = n42629 ;
  assign y13864 = ~n42630 ;
  assign y13865 = ~n42631 ;
  assign y13866 = n42634 ;
  assign y13867 = n42639 ;
  assign y13868 = ~1'b0 ;
  assign y13869 = ~1'b0 ;
  assign y13870 = ~n42643 ;
  assign y13871 = n42644 ;
  assign y13872 = ~n42645 ;
  assign y13873 = ~n42646 ;
  assign y13874 = n42647 ;
  assign y13875 = n42649 ;
  assign y13876 = n42651 ;
  assign y13877 = ~1'b0 ;
  assign y13878 = n42653 ;
  assign y13879 = ~n42654 ;
  assign y13880 = n42656 ;
  assign y13881 = ~n42659 ;
  assign y13882 = ~n42663 ;
  assign y13883 = ~1'b0 ;
  assign y13884 = n42665 ;
  assign y13885 = ~1'b0 ;
  assign y13886 = ~n42669 ;
  assign y13887 = ~n42675 ;
  assign y13888 = n42677 ;
  assign y13889 = n42683 ;
  assign y13890 = ~n42685 ;
  assign y13891 = ~1'b0 ;
  assign y13892 = ~n42686 ;
  assign y13893 = n42688 ;
  assign y13894 = n42690 ;
  assign y13895 = ~n42693 ;
  assign y13896 = n42699 ;
  assign y13897 = ~n42701 ;
  assign y13898 = ~1'b0 ;
  assign y13899 = ~1'b0 ;
  assign y13900 = ~n42702 ;
  assign y13901 = ~n28543 ;
  assign y13902 = n42703 ;
  assign y13903 = ~n42707 ;
  assign y13904 = ~1'b0 ;
  assign y13905 = ~n42713 ;
  assign y13906 = n42714 ;
  assign y13907 = ~n42715 ;
  assign y13908 = ~n42720 ;
  assign y13909 = n42723 ;
  assign y13910 = ~n42726 ;
  assign y13911 = ~1'b0 ;
  assign y13912 = n42729 ;
  assign y13913 = n42731 ;
  assign y13914 = ~n42732 ;
  assign y13915 = ~n42735 ;
  assign y13916 = n42737 ;
  assign y13917 = n42738 ;
  assign y13918 = ~n42740 ;
  assign y13919 = ~1'b0 ;
  assign y13920 = n42743 ;
  assign y13921 = ~n42746 ;
  assign y13922 = n42747 ;
  assign y13923 = n42748 ;
  assign y13924 = ~n27084 ;
  assign y13925 = n42750 ;
  assign y13926 = ~n42754 ;
  assign y13927 = n42756 ;
  assign y13928 = ~n42760 ;
  assign y13929 = n42764 ;
  assign y13930 = ~1'b0 ;
  assign y13931 = n42766 ;
  assign y13932 = n42771 ;
  assign y13933 = ~n42772 ;
  assign y13934 = n42774 ;
  assign y13935 = n42777 ;
  assign y13936 = ~n42778 ;
  assign y13937 = n42786 ;
  assign y13938 = ~1'b0 ;
  assign y13939 = ~n42795 ;
  assign y13940 = n42796 ;
  assign y13941 = ~n42805 ;
  assign y13942 = n42806 ;
  assign y13943 = n42811 ;
  assign y13944 = ~n42815 ;
  assign y13945 = ~n42817 ;
  assign y13946 = n42819 ;
  assign y13947 = n42825 ;
  assign y13948 = ~1'b0 ;
  assign y13949 = ~n42833 ;
  assign y13950 = ~n42834 ;
  assign y13951 = ~n42835 ;
  assign y13952 = ~1'b0 ;
  assign y13953 = n42837 ;
  assign y13954 = ~n42840 ;
  assign y13955 = ~n42846 ;
  assign y13956 = ~1'b0 ;
  assign y13957 = n42860 ;
  assign y13958 = ~n42861 ;
  assign y13959 = ~n42862 ;
  assign y13960 = ~n42863 ;
  assign y13961 = ~n42865 ;
  assign y13962 = n42870 ;
  assign y13963 = ~1'b0 ;
  assign y13964 = n34475 ;
  assign y13965 = ~n42871 ;
  assign y13966 = n42889 ;
  assign y13967 = n42890 ;
  assign y13968 = ~1'b0 ;
  assign y13969 = n42893 ;
  assign y13970 = ~n42895 ;
  assign y13971 = n25003 ;
  assign y13972 = ~n42896 ;
  assign y13973 = ~n42900 ;
  assign y13974 = n42901 ;
  assign y13975 = ~n42905 ;
  assign y13976 = n42906 ;
  assign y13977 = n42912 ;
  assign y13978 = ~n42917 ;
  assign y13979 = ~1'b0 ;
  assign y13980 = ~n42918 ;
  assign y13981 = n27741 ;
  assign y13982 = ~n42921 ;
  assign y13983 = n42922 ;
  assign y13984 = n42924 ;
  assign y13985 = ~1'b0 ;
  assign y13986 = ~1'b0 ;
  assign y13987 = ~n42928 ;
  assign y13988 = n42933 ;
  assign y13989 = ~n42934 ;
  assign y13990 = ~n42935 ;
  assign y13991 = ~n42938 ;
  assign y13992 = n42941 ;
  assign y13993 = ~1'b0 ;
  assign y13994 = ~n42943 ;
  assign y13995 = n42944 ;
  assign y13996 = n42945 ;
  assign y13997 = ~n42946 ;
  assign y13998 = n42949 ;
  assign y13999 = ~n42950 ;
  assign y14000 = ~1'b0 ;
  assign y14001 = ~n18963 ;
  assign y14002 = ~n42951 ;
  assign y14003 = n42952 ;
  assign y14004 = n42953 ;
  assign y14005 = n42957 ;
  assign y14006 = n42962 ;
  assign y14007 = ~n42965 ;
  assign y14008 = n42967 ;
  assign y14009 = ~n42968 ;
  assign y14010 = n42969 ;
  assign y14011 = ~n42970 ;
  assign y14012 = ~n42971 ;
  assign y14013 = n42974 ;
  assign y14014 = n42975 ;
  assign y14015 = n42976 ;
  assign y14016 = n42978 ;
  assign y14017 = n42980 ;
  assign y14018 = ~n42982 ;
  assign y14019 = ~1'b0 ;
  assign y14020 = ~n42992 ;
  assign y14021 = ~n43004 ;
  assign y14022 = ~n41997 ;
  assign y14023 = n43010 ;
  assign y14024 = n43014 ;
  assign y14025 = ~n43015 ;
  assign y14026 = ~n43016 ;
  assign y14027 = n43018 ;
  assign y14028 = ~n43020 ;
  assign y14029 = n43025 ;
  assign y14030 = ~1'b0 ;
  assign y14031 = ~n43028 ;
  assign y14032 = ~n43032 ;
  assign y14033 = n43033 ;
  assign y14034 = n43034 ;
  assign y14035 = ~n43035 ;
  assign y14036 = n43044 ;
  assign y14037 = ~n2720 ;
  assign y14038 = ~n43050 ;
  assign y14039 = n43053 ;
  assign y14040 = n43055 ;
  assign y14041 = ~n43059 ;
  assign y14042 = n23199 ;
  assign y14043 = n43062 ;
  assign y14044 = ~n43064 ;
  assign y14045 = n43067 ;
  assign y14046 = ~n43068 ;
  assign y14047 = ~n43069 ;
  assign y14048 = ~n43080 ;
  assign y14049 = ~1'b0 ;
  assign y14050 = n43086 ;
  assign y14051 = ~n43090 ;
  assign y14052 = ~n43094 ;
  assign y14053 = n43095 ;
  assign y14054 = ~n43099 ;
  assign y14055 = n43101 ;
  assign y14056 = n43104 ;
  assign y14057 = n43105 ;
  assign y14058 = n43106 ;
  assign y14059 = n43107 ;
  assign y14060 = ~n43109 ;
  assign y14061 = n43111 ;
  assign y14062 = ~1'b0 ;
  assign y14063 = ~1'b0 ;
  assign y14064 = ~n43114 ;
  assign y14065 = n43115 ;
  assign y14066 = ~n31019 ;
  assign y14067 = ~n43117 ;
  assign y14068 = ~n43119 ;
  assign y14069 = n43122 ;
  assign y14070 = n43129 ;
  assign y14071 = ~n43130 ;
  assign y14072 = ~n43135 ;
  assign y14073 = ~n30008 ;
  assign y14074 = ~n43136 ;
  assign y14075 = n43138 ;
  assign y14076 = ~1'b0 ;
  assign y14077 = ~1'b0 ;
  assign y14078 = ~n43140 ;
  assign y14079 = ~n43141 ;
  assign y14080 = ~n43142 ;
  assign y14081 = n43149 ;
  assign y14082 = n43156 ;
  assign y14083 = ~1'b0 ;
  assign y14084 = ~n43160 ;
  assign y14085 = ~n43161 ;
  assign y14086 = n28283 ;
  assign y14087 = ~n43166 ;
  assign y14088 = ~n43167 ;
  assign y14089 = n43169 ;
  assign y14090 = ~1'b0 ;
  assign y14091 = ~n43177 ;
  assign y14092 = n43180 ;
  assign y14093 = n43181 ;
  assign y14094 = n43182 ;
  assign y14095 = n43185 ;
  assign y14096 = n43189 ;
  assign y14097 = ~n1791 ;
  assign y14098 = ~1'b0 ;
  assign y14099 = n43191 ;
  assign y14100 = ~1'b0 ;
  assign y14101 = ~n43197 ;
  assign y14102 = n43199 ;
  assign y14103 = n43207 ;
  assign y14104 = ~n43216 ;
  assign y14105 = n43217 ;
  assign y14106 = n43220 ;
  assign y14107 = n43221 ;
  assign y14108 = n43224 ;
  assign y14109 = ~n43225 ;
  assign y14110 = ~n10724 ;
  assign y14111 = n43226 ;
  assign y14112 = n43227 ;
  assign y14113 = ~n43231 ;
  assign y14114 = ~n43232 ;
  assign y14115 = ~1'b0 ;
  assign y14116 = n11329 ;
  assign y14117 = ~n43236 ;
  assign y14118 = ~n43247 ;
  assign y14119 = n43250 ;
  assign y14120 = n43252 ;
  assign y14121 = n43255 ;
  assign y14122 = n43259 ;
  assign y14123 = ~1'b0 ;
  assign y14124 = n43261 ;
  assign y14125 = n43262 ;
  assign y14126 = ~n43263 ;
  assign y14127 = ~n43269 ;
  assign y14128 = n43270 ;
  assign y14129 = ~n43272 ;
  assign y14130 = ~1'b0 ;
  assign y14131 = ~n43276 ;
  assign y14132 = n43278 ;
  assign y14133 = n43283 ;
  assign y14134 = ~n43284 ;
  assign y14135 = ~n43287 ;
  assign y14136 = n43289 ;
  assign y14137 = ~n43292 ;
  assign y14138 = ~1'b0 ;
  assign y14139 = n43293 ;
  assign y14140 = n43298 ;
  assign y14141 = ~n43301 ;
  assign y14142 = ~n43307 ;
  assign y14143 = ~n43308 ;
  assign y14144 = n43310 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = n43312 ;
  assign y14147 = ~n43314 ;
  assign y14148 = ~n43316 ;
  assign y14149 = n43320 ;
  assign y14150 = ~n43321 ;
  assign y14151 = n43328 ;
  assign y14152 = ~n43329 ;
  assign y14153 = ~1'b0 ;
  assign y14154 = ~n43330 ;
  assign y14155 = n43338 ;
  assign y14156 = ~n43342 ;
  assign y14157 = n43348 ;
  assign y14158 = n43349 ;
  assign y14159 = n43350 ;
  assign y14160 = ~n43351 ;
  assign y14161 = ~1'b0 ;
  assign y14162 = n43354 ;
  assign y14163 = ~1'b0 ;
  assign y14164 = ~n43357 ;
  assign y14165 = ~n43360 ;
  assign y14166 = ~n43365 ;
  assign y14167 = n43366 ;
  assign y14168 = n43368 ;
  assign y14169 = n43373 ;
  assign y14170 = ~n43374 ;
  assign y14171 = n43375 ;
  assign y14172 = n43377 ;
  assign y14173 = n43378 ;
  assign y14174 = ~n43380 ;
  assign y14175 = ~n43381 ;
  assign y14176 = ~n43382 ;
  assign y14177 = ~n43387 ;
  assign y14178 = 1'b0 ;
  assign y14179 = n43389 ;
  assign y14180 = ~1'b0 ;
  assign y14181 = n43392 ;
  assign y14182 = n43399 ;
  assign y14183 = ~n43400 ;
  assign y14184 = n43404 ;
  assign y14185 = ~n43409 ;
  assign y14186 = n43415 ;
  assign y14187 = ~1'b0 ;
  assign y14188 = n43419 ;
  assign y14189 = ~1'b0 ;
  assign y14190 = ~n43422 ;
  assign y14191 = ~n43423 ;
  assign y14192 = n43426 ;
  assign y14193 = n43428 ;
  assign y14194 = ~n43429 ;
  assign y14195 = ~1'b0 ;
  assign y14196 = ~n43432 ;
  assign y14197 = n43437 ;
  assign y14198 = ~n43439 ;
  assign y14199 = ~n43440 ;
  assign y14200 = ~1'b0 ;
  assign y14201 = n43443 ;
  assign y14202 = ~n43445 ;
  assign y14203 = ~n43447 ;
  assign y14204 = n43451 ;
  assign y14205 = n39912 ;
  assign y14206 = n43452 ;
  assign y14207 = ~1'b0 ;
  assign y14208 = ~1'b0 ;
  assign y14209 = ~1'b0 ;
  assign y14210 = ~1'b0 ;
  assign y14211 = n43454 ;
  assign y14212 = ~n43455 ;
  assign y14213 = ~n43458 ;
  assign y14214 = ~n43463 ;
  assign y14215 = ~n43467 ;
  assign y14216 = ~1'b0 ;
  assign y14217 = ~1'b0 ;
  assign y14218 = n43468 ;
  assign y14219 = n43470 ;
  assign y14220 = n43471 ;
  assign y14221 = ~n43473 ;
  assign y14222 = ~n43475 ;
  assign y14223 = ~n43477 ;
  assign y14224 = n43478 ;
  assign y14225 = n43480 ;
  assign y14226 = n43488 ;
  assign y14227 = ~n43489 ;
  assign y14228 = ~n43490 ;
  assign y14229 = n43492 ;
  assign y14230 = ~n43493 ;
  assign y14231 = ~n43496 ;
  assign y14232 = ~n43498 ;
  assign y14233 = n43500 ;
  assign y14234 = n43503 ;
  assign y14235 = ~n43504 ;
  assign y14236 = ~n43505 ;
  assign y14237 = n43507 ;
  assign y14238 = n43509 ;
  assign y14239 = n43510 ;
  assign y14240 = ~1'b0 ;
  assign y14241 = ~n43513 ;
  assign y14242 = n43517 ;
  assign y14243 = ~n43518 ;
  assign y14244 = ~n43521 ;
  assign y14245 = n43523 ;
  assign y14246 = n43526 ;
  assign y14247 = ~n43529 ;
  assign y14248 = n43530 ;
  assign y14249 = ~n43531 ;
  assign y14250 = n43536 ;
  assign y14251 = n43538 ;
  assign y14252 = ~1'b0 ;
  assign y14253 = ~n43539 ;
  assign y14254 = n43541 ;
  assign y14255 = n43542 ;
  assign y14256 = n43543 ;
  assign y14257 = n43545 ;
  assign y14258 = ~1'b0 ;
  assign y14259 = ~n43547 ;
  assign y14260 = n43549 ;
  assign y14261 = ~n43550 ;
  assign y14262 = ~1'b0 ;
  assign y14263 = n43551 ;
  assign y14264 = ~n43553 ;
  assign y14265 = ~n43554 ;
  assign y14266 = ~n43555 ;
  assign y14267 = ~n43556 ;
  assign y14268 = n43557 ;
  assign y14269 = ~n43560 ;
  assign y14270 = n18672 ;
  assign y14271 = ~1'b0 ;
  assign y14272 = n43562 ;
  assign y14273 = n43564 ;
  assign y14274 = n43565 ;
  assign y14275 = ~n43567 ;
  assign y14276 = ~n43570 ;
  assign y14277 = n43572 ;
  assign y14278 = ~n43575 ;
  assign y14279 = ~n43577 ;
  assign y14280 = ~n43580 ;
  assign y14281 = ~n43582 ;
  assign y14282 = n43583 ;
  assign y14283 = ~n43584 ;
  assign y14284 = n43585 ;
  assign y14285 = n43590 ;
  assign y14286 = n43591 ;
  assign y14287 = n43593 ;
  assign y14288 = n43597 ;
  assign y14289 = ~n43599 ;
  assign y14290 = n43603 ;
  assign y14291 = n43606 ;
  assign y14292 = ~n43610 ;
  assign y14293 = n43613 ;
  assign y14294 = n43617 ;
  assign y14295 = n43620 ;
  assign y14296 = n43622 ;
  assign y14297 = n43625 ;
  assign y14298 = n43629 ;
  assign y14299 = n43635 ;
  assign y14300 = ~n43639 ;
  assign y14301 = ~n43643 ;
  assign y14302 = ~1'b0 ;
  assign y14303 = ~n43644 ;
  assign y14304 = ~n43645 ;
  assign y14305 = ~n43647 ;
  assign y14306 = n43651 ;
  assign y14307 = n43652 ;
  assign y14308 = n43653 ;
  assign y14309 = n43655 ;
  assign y14310 = n43656 ;
  assign y14311 = n43658 ;
  assign y14312 = ~1'b0 ;
  assign y14313 = ~1'b0 ;
  assign y14314 = ~n43661 ;
  assign y14315 = ~n43662 ;
  assign y14316 = n43663 ;
  assign y14317 = n43664 ;
  assign y14318 = ~n43665 ;
  assign y14319 = n43667 ;
  assign y14320 = ~n43668 ;
  assign y14321 = ~1'b0 ;
  assign y14322 = n43669 ;
  assign y14323 = ~n43671 ;
  assign y14324 = n25531 ;
  assign y14325 = ~1'b0 ;
  assign y14326 = ~n43674 ;
  assign y14327 = n43676 ;
  assign y14328 = ~n43679 ;
  assign y14329 = ~n43680 ;
  assign y14330 = ~1'b0 ;
  assign y14331 = ~n43682 ;
  assign y14332 = ~n43684 ;
  assign y14333 = n43691 ;
  assign y14334 = n43694 ;
  assign y14335 = ~n43695 ;
  assign y14336 = n43699 ;
  assign y14337 = ~n43703 ;
  assign y14338 = ~n43705 ;
  assign y14339 = ~1'b0 ;
  assign y14340 = ~n40821 ;
  assign y14341 = n43706 ;
  assign y14342 = n43707 ;
  assign y14343 = n43710 ;
  assign y14344 = n43716 ;
  assign y14345 = n43717 ;
  assign y14346 = n43721 ;
  assign y14347 = ~n43726 ;
  assign y14348 = ~n43730 ;
  assign y14349 = ~n43732 ;
  assign y14350 = ~n43736 ;
  assign y14351 = ~n43738 ;
  assign y14352 = ~n43739 ;
  assign y14353 = n43742 ;
  assign y14354 = ~n43743 ;
  assign y14355 = ~n43745 ;
  assign y14356 = n43750 ;
  assign y14357 = n43751 ;
  assign y14358 = ~n43754 ;
  assign y14359 = n43758 ;
  assign y14360 = ~n35421 ;
  assign y14361 = n43759 ;
  assign y14362 = ~n43761 ;
  assign y14363 = n43763 ;
  assign y14364 = ~n43767 ;
  assign y14365 = n43769 ;
  assign y14366 = ~n43771 ;
  assign y14367 = n43773 ;
  assign y14368 = n43776 ;
  assign y14369 = ~n43777 ;
  assign y14370 = n43778 ;
  assign y14371 = n43779 ;
  assign y14372 = n43781 ;
  assign y14373 = n16195 ;
  assign y14374 = ~n43783 ;
  assign y14375 = ~n43786 ;
  assign y14376 = n43795 ;
  assign y14377 = ~1'b0 ;
  assign y14378 = n43806 ;
  assign y14379 = ~n43808 ;
  assign y14380 = n43811 ;
  assign y14381 = n43812 ;
  assign y14382 = n43814 ;
  assign y14383 = ~n43816 ;
  assign y14384 = ~n43818 ;
  assign y14385 = n43827 ;
  assign y14386 = ~n43829 ;
  assign y14387 = n43830 ;
  assign y14388 = n43833 ;
  assign y14389 = ~n43836 ;
  assign y14390 = ~n43838 ;
  assign y14391 = n43839 ;
  assign y14392 = n43841 ;
  assign y14393 = n43844 ;
  assign y14394 = ~n43848 ;
  assign y14395 = ~n43850 ;
  assign y14396 = ~1'b0 ;
  assign y14397 = n43852 ;
  assign y14398 = n43855 ;
  assign y14399 = ~n43856 ;
  assign y14400 = ~n43857 ;
  assign y14401 = n43858 ;
  assign y14402 = ~n43860 ;
  assign y14403 = ~n43862 ;
  assign y14404 = ~1'b0 ;
  assign y14405 = 1'b0 ;
  assign y14406 = ~n17439 ;
  assign y14407 = n43863 ;
  assign y14408 = ~n43866 ;
  assign y14409 = n43868 ;
  assign y14410 = n43873 ;
  assign y14411 = ~1'b0 ;
  assign y14412 = ~n43877 ;
  assign y14413 = n43879 ;
  assign y14414 = n43883 ;
  assign y14415 = ~n43885 ;
  assign y14416 = ~n43890 ;
  assign y14417 = n43891 ;
  assign y14418 = n43895 ;
  assign y14419 = ~1'b0 ;
  assign y14420 = ~n43898 ;
  assign y14421 = ~n43899 ;
  assign y14422 = ~n43900 ;
  assign y14423 = ~n43901 ;
  assign y14424 = n43902 ;
  assign y14425 = n43903 ;
  assign y14426 = n43904 ;
  assign y14427 = ~n43906 ;
  assign y14428 = ~1'b0 ;
  assign y14429 = ~1'b0 ;
  assign y14430 = n43908 ;
  assign y14431 = ~n43913 ;
  assign y14432 = ~n43914 ;
  assign y14433 = ~1'b0 ;
  assign y14434 = ~1'b0 ;
  assign y14435 = n43916 ;
  assign y14436 = ~n43920 ;
  assign y14437 = ~n43923 ;
  assign y14438 = ~n43925 ;
  assign y14439 = n43927 ;
  assign y14440 = ~n39892 ;
  assign y14441 = n43928 ;
  assign y14442 = ~1'b0 ;
  assign y14443 = ~1'b0 ;
  assign y14444 = n43930 ;
  assign y14445 = n43933 ;
  assign y14446 = n43934 ;
  assign y14447 = n43935 ;
  assign y14448 = n43936 ;
  assign y14449 = ~n43938 ;
  assign y14450 = ~1'b0 ;
  assign y14451 = n43939 ;
  assign y14452 = ~1'b0 ;
  assign y14453 = ~n12870 ;
  assign y14454 = n43946 ;
  assign y14455 = ~n43948 ;
  assign y14456 = ~n43949 ;
  assign y14457 = n43950 ;
  assign y14458 = ~n43954 ;
  assign y14459 = n43955 ;
  assign y14460 = ~1'b0 ;
  assign y14461 = ~1'b0 ;
  assign y14462 = n43961 ;
  assign y14463 = n43964 ;
  assign y14464 = ~n43965 ;
  assign y14465 = ~n43966 ;
  assign y14466 = n43971 ;
  assign y14467 = ~n43975 ;
  assign y14468 = n43983 ;
  assign y14469 = ~1'b0 ;
  assign y14470 = ~1'b0 ;
  assign y14471 = n43985 ;
  assign y14472 = ~n43991 ;
  assign y14473 = ~n43995 ;
  assign y14474 = n43997 ;
  assign y14475 = ~n43999 ;
  assign y14476 = ~n44000 ;
  assign y14477 = ~n44002 ;
  assign y14478 = ~n44004 ;
  assign y14479 = ~n44012 ;
  assign y14480 = n44015 ;
  assign y14481 = ~n44016 ;
  assign y14482 = ~n11170 ;
  assign y14483 = n44019 ;
  assign y14484 = n44020 ;
  assign y14485 = ~n44022 ;
  assign y14486 = ~n44028 ;
  assign y14487 = ~n44033 ;
  assign y14488 = ~n44035 ;
  assign y14489 = ~1'b0 ;
  assign y14490 = ~1'b0 ;
  assign y14491 = ~n44036 ;
  assign y14492 = n44040 ;
  assign y14493 = ~n24671 ;
  assign y14494 = n44041 ;
  assign y14495 = ~n44043 ;
  assign y14496 = n44052 ;
  assign y14497 = n44055 ;
  assign y14498 = n44056 ;
  assign y14499 = n44057 ;
  assign y14500 = ~n44060 ;
  assign y14501 = ~n44062 ;
  assign y14502 = ~n44066 ;
  assign y14503 = ~n44071 ;
  assign y14504 = ~1'b0 ;
  assign y14505 = n44076 ;
  assign y14506 = ~n44080 ;
  assign y14507 = ~n44082 ;
  assign y14508 = n44084 ;
  assign y14509 = ~1'b0 ;
  assign y14510 = ~n44086 ;
  assign y14511 = n44087 ;
  assign y14512 = ~n44088 ;
  assign y14513 = ~n38482 ;
  assign y14514 = n44089 ;
  assign y14515 = ~n44092 ;
  assign y14516 = n44097 ;
  assign y14517 = n44101 ;
  assign y14518 = ~n44102 ;
  assign y14519 = ~n42606 ;
  assign y14520 = ~n44103 ;
  assign y14521 = ~n44105 ;
  assign y14522 = ~1'b0 ;
  assign y14523 = ~1'b0 ;
  assign y14524 = n44106 ;
  assign y14525 = n44109 ;
  assign y14526 = ~n44110 ;
  assign y14527 = ~n44113 ;
  assign y14528 = n44114 ;
  assign y14529 = ~1'b0 ;
  assign y14530 = ~n44117 ;
  assign y14531 = ~n44118 ;
  assign y14532 = ~1'b0 ;
  assign y14533 = n44122 ;
  assign y14534 = n44124 ;
  assign y14535 = n44130 ;
  assign y14536 = n44132 ;
  assign y14537 = n44135 ;
  assign y14538 = n44136 ;
  assign y14539 = n44137 ;
  assign y14540 = ~1'b0 ;
  assign y14541 = n44141 ;
  assign y14542 = n44142 ;
  assign y14543 = ~n44150 ;
  assign y14544 = n44153 ;
  assign y14545 = ~n44154 ;
  assign y14546 = n44158 ;
  assign y14547 = n44161 ;
  assign y14548 = ~1'b0 ;
  assign y14549 = ~n44163 ;
  assign y14550 = ~n44164 ;
  assign y14551 = n44165 ;
  assign y14552 = n44166 ;
  assign y14553 = n44169 ;
  assign y14554 = ~n44174 ;
  assign y14555 = n44175 ;
  assign y14556 = ~n44178 ;
  assign y14557 = n44179 ;
  assign y14558 = ~n44181 ;
  assign y14559 = ~1'b0 ;
  assign y14560 = ~n44184 ;
  assign y14561 = ~n44189 ;
  assign y14562 = ~n44190 ;
  assign y14563 = ~n44191 ;
  assign y14564 = n44198 ;
  assign y14565 = ~1'b0 ;
  assign y14566 = n44203 ;
  assign y14567 = n44204 ;
  assign y14568 = n44208 ;
  assign y14569 = n44209 ;
  assign y14570 = ~n44212 ;
  assign y14571 = n44216 ;
  assign y14572 = n44217 ;
  assign y14573 = ~1'b0 ;
  assign y14574 = n44219 ;
  assign y14575 = n44221 ;
  assign y14576 = ~n44222 ;
  assign y14577 = ~n44228 ;
  assign y14578 = ~n44232 ;
  assign y14579 = ~n44234 ;
  assign y14580 = ~n44235 ;
  assign y14581 = ~n44241 ;
  assign y14582 = ~n44244 ;
  assign y14583 = ~n44246 ;
  assign y14584 = ~1'b0 ;
  assign y14585 = ~n44249 ;
  assign y14586 = n44250 ;
  assign y14587 = n44252 ;
  assign y14588 = n44254 ;
  assign y14589 = ~n44257 ;
  assign y14590 = n44258 ;
  assign y14591 = ~n44262 ;
  assign y14592 = ~n44266 ;
  assign y14593 = ~n44267 ;
  assign y14594 = ~n44270 ;
  assign y14595 = n44274 ;
  assign y14596 = ~n44275 ;
  assign y14597 = ~n44279 ;
  assign y14598 = ~n44282 ;
  assign y14599 = ~n44286 ;
  assign y14600 = ~1'b0 ;
  assign y14601 = ~1'b0 ;
  assign y14602 = ~n44290 ;
  assign y14603 = ~n44291 ;
  assign y14604 = ~n44292 ;
  assign y14605 = ~n44294 ;
  assign y14606 = ~n44295 ;
  assign y14607 = ~n44296 ;
  assign y14608 = ~1'b0 ;
  assign y14609 = n44297 ;
  assign y14610 = ~n44299 ;
  assign y14611 = ~1'b0 ;
  assign y14612 = n44305 ;
  assign y14613 = n44308 ;
  assign y14614 = ~n44310 ;
  assign y14615 = ~n44312 ;
  assign y14616 = ~n44314 ;
  assign y14617 = ~n44318 ;
  assign y14618 = n44320 ;
  assign y14619 = n44324 ;
  assign y14620 = ~n44325 ;
  assign y14621 = ~n44326 ;
  assign y14622 = ~n44330 ;
  assign y14623 = ~1'b0 ;
  assign y14624 = ~1'b0 ;
  assign y14625 = ~n7223 ;
  assign y14626 = n44331 ;
  assign y14627 = ~n44334 ;
  assign y14628 = n44337 ;
  assign y14629 = ~n44338 ;
  assign y14630 = ~n44341 ;
  assign y14631 = n44342 ;
  assign y14632 = ~1'b0 ;
  assign y14633 = ~n44349 ;
  assign y14634 = ~1'b0 ;
  assign y14635 = ~1'b0 ;
  assign y14636 = n44350 ;
  assign y14637 = ~n44355 ;
  assign y14638 = n44363 ;
  assign y14639 = ~n44365 ;
  assign y14640 = ~n44366 ;
  assign y14641 = ~1'b0 ;
  assign y14642 = n44371 ;
  assign y14643 = n10838 ;
  assign y14644 = ~n44372 ;
  assign y14645 = ~n44374 ;
  assign y14646 = ~n44376 ;
  assign y14647 = ~n44380 ;
  assign y14648 = n44382 ;
  assign y14649 = ~1'b0 ;
  assign y14650 = n44385 ;
  assign y14651 = ~n44387 ;
  assign y14652 = n44389 ;
  assign y14653 = ~n44390 ;
  assign y14654 = n22451 ;
  assign y14655 = n44394 ;
  assign y14656 = n44397 ;
  assign y14657 = ~1'b0 ;
  assign y14658 = ~1'b0 ;
  assign y14659 = n44400 ;
  assign y14660 = ~n44403 ;
  assign y14661 = ~n44406 ;
  assign y14662 = n44408 ;
  assign y14663 = ~n44413 ;
  assign y14664 = ~1'b0 ;
  assign y14665 = ~1'b0 ;
  assign y14666 = ~n44416 ;
  assign y14667 = n44420 ;
  assign y14668 = n44422 ;
  assign y14669 = ~n44423 ;
  assign y14670 = n44424 ;
  assign y14671 = ~n44432 ;
  assign y14672 = ~1'b0 ;
  assign y14673 = ~n4681 ;
  assign y14674 = ~n44434 ;
  assign y14675 = n44436 ;
  assign y14676 = n44439 ;
  assign y14677 = ~n44440 ;
  assign y14678 = n44443 ;
  assign y14679 = ~n44444 ;
  assign y14680 = n44448 ;
  assign y14681 = ~1'b0 ;
  assign y14682 = n44449 ;
  assign y14683 = ~1'b0 ;
  assign y14684 = ~1'b0 ;
  assign y14685 = ~1'b0 ;
  assign y14686 = ~n44452 ;
  assign y14687 = n44458 ;
  assign y14688 = n44463 ;
  assign y14689 = n44465 ;
  assign y14690 = ~n44467 ;
  assign y14691 = ~n44468 ;
  assign y14692 = n44469 ;
  assign y14693 = ~n8119 ;
  assign y14694 = ~n44470 ;
  assign y14695 = n44474 ;
  assign y14696 = ~1'b0 ;
  assign y14697 = ~n44477 ;
  assign y14698 = ~n44480 ;
  assign y14699 = ~n44482 ;
  assign y14700 = n44483 ;
  assign y14701 = ~n44485 ;
  assign y14702 = ~n44486 ;
  assign y14703 = ~n44488 ;
  assign y14704 = n44489 ;
  assign y14705 = n44493 ;
  assign y14706 = n9474 ;
  assign y14707 = ~1'b0 ;
  assign y14708 = n44501 ;
  assign y14709 = n44502 ;
  assign y14710 = n44504 ;
  assign y14711 = n44506 ;
  assign y14712 = ~n44508 ;
  assign y14713 = ~1'b0 ;
  assign y14714 = ~n44512 ;
  assign y14715 = ~1'b0 ;
  assign y14716 = n44514 ;
  assign y14717 = ~n44516 ;
  assign y14718 = n44517 ;
  assign y14719 = n44518 ;
  assign y14720 = n44519 ;
  assign y14721 = n44522 ;
  assign y14722 = n44523 ;
  assign y14723 = ~n44526 ;
  assign y14724 = n44531 ;
  assign y14725 = ~n44532 ;
  assign y14726 = ~n44537 ;
  assign y14727 = n44539 ;
  assign y14728 = n44540 ;
  assign y14729 = n44541 ;
  assign y14730 = n44544 ;
  assign y14731 = ~n44545 ;
  assign y14732 = ~1'b0 ;
  assign y14733 = ~n44546 ;
  assign y14734 = ~1'b0 ;
  assign y14735 = ~1'b0 ;
  assign y14736 = n44549 ;
  assign y14737 = ~n44551 ;
  assign y14738 = ~n44553 ;
  assign y14739 = ~n44554 ;
  assign y14740 = ~n44555 ;
  assign y14741 = ~n44558 ;
  assign y14742 = n44561 ;
  assign y14743 = ~n44562 ;
  assign y14744 = ~n44563 ;
  assign y14745 = n44565 ;
  assign y14746 = ~n44566 ;
  assign y14747 = ~n44567 ;
  assign y14748 = ~1'b0 ;
  assign y14749 = ~1'b0 ;
  assign y14750 = n44570 ;
  assign y14751 = n44573 ;
  assign y14752 = n4173 ;
  assign y14753 = ~n44575 ;
  assign y14754 = ~n44583 ;
  assign y14755 = n44584 ;
  assign y14756 = n44587 ;
  assign y14757 = n44589 ;
  assign y14758 = ~n44591 ;
  assign y14759 = ~n13273 ;
  assign y14760 = ~n44594 ;
  assign y14761 = ~n44597 ;
  assign y14762 = n44598 ;
  assign y14763 = ~n44601 ;
  assign y14764 = ~n44603 ;
  assign y14765 = ~n44605 ;
  assign y14766 = ~n44606 ;
  assign y14767 = ~n44607 ;
  assign y14768 = ~n44610 ;
  assign y14769 = ~n44611 ;
  assign y14770 = n44613 ;
  assign y14771 = n44617 ;
  assign y14772 = n44618 ;
  assign y14773 = ~n44620 ;
  assign y14774 = n44622 ;
  assign y14775 = ~1'b0 ;
  assign y14776 = ~1'b0 ;
  assign y14777 = n44624 ;
  assign y14778 = ~n44625 ;
  assign y14779 = n44627 ;
  assign y14780 = ~n44628 ;
  assign y14781 = n44631 ;
  assign y14782 = ~n44633 ;
  assign y14783 = n44639 ;
  assign y14784 = n44642 ;
  assign y14785 = ~1'b0 ;
  assign y14786 = n44643 ;
  assign y14787 = ~n44649 ;
  assign y14788 = ~n44650 ;
  assign y14789 = n44651 ;
  assign y14790 = n44654 ;
  assign y14791 = n44657 ;
  assign y14792 = ~n44659 ;
  assign y14793 = n44662 ;
  assign y14794 = n44663 ;
  assign y14795 = n35234 ;
  assign y14796 = ~n44666 ;
  assign y14797 = n44667 ;
  assign y14798 = n44670 ;
  assign y14799 = ~n44671 ;
  assign y14800 = n44674 ;
  assign y14801 = n44676 ;
  assign y14802 = ~1'b0 ;
  assign y14803 = ~1'b0 ;
  assign y14804 = n44679 ;
  assign y14805 = n44682 ;
  assign y14806 = n44686 ;
  assign y14807 = ~n44688 ;
  assign y14808 = n44689 ;
  assign y14809 = ~n44692 ;
  assign y14810 = ~n44694 ;
  assign y14811 = n44696 ;
  assign y14812 = ~n44698 ;
  assign y14813 = ~1'b0 ;
  assign y14814 = ~n44701 ;
  assign y14815 = n44703 ;
  assign y14816 = ~n44706 ;
  assign y14817 = ~n44708 ;
  assign y14818 = ~n44709 ;
  assign y14819 = ~1'b0 ;
  assign y14820 = ~1'b0 ;
  assign y14821 = ~1'b0 ;
  assign y14822 = ~n44711 ;
  assign y14823 = n44712 ;
  assign y14824 = ~n44719 ;
  assign y14825 = n44726 ;
  assign y14826 = ~n44727 ;
  assign y14827 = ~n44728 ;
  assign y14828 = n44730 ;
  assign y14829 = n44731 ;
  assign y14830 = ~n44733 ;
  assign y14831 = n7171 ;
  assign y14832 = n44735 ;
  assign y14833 = ~n44740 ;
  assign y14834 = n44741 ;
  assign y14835 = n44748 ;
  assign y14836 = ~n44750 ;
  assign y14837 = n44754 ;
  assign y14838 = n44761 ;
  assign y14839 = ~1'b0 ;
  assign y14840 = ~n44762 ;
  assign y14841 = ~n44764 ;
  assign y14842 = ~1'b0 ;
  assign y14843 = ~n44411 ;
  assign y14844 = n44766 ;
  assign y14845 = ~n44772 ;
  assign y14846 = ~n44781 ;
  assign y14847 = ~n44782 ;
  assign y14848 = n44783 ;
  assign y14849 = ~n44784 ;
  assign y14850 = ~n44788 ;
  assign y14851 = ~1'b0 ;
  assign y14852 = n44791 ;
  assign y14853 = ~n44793 ;
  assign y14854 = ~1'b0 ;
  assign y14855 = ~n44795 ;
  assign y14856 = n44798 ;
  assign y14857 = n44799 ;
  assign y14858 = n44803 ;
  assign y14859 = n44809 ;
  assign y14860 = ~n44812 ;
  assign y14861 = ~1'b0 ;
  assign y14862 = ~n44814 ;
  assign y14863 = n44816 ;
  assign y14864 = n44819 ;
  assign y14865 = ~n44821 ;
  assign y14866 = ~n44826 ;
  assign y14867 = n44828 ;
  assign y14868 = ~n44829 ;
  assign y14869 = ~n44830 ;
  assign y14870 = ~n44833 ;
  assign y14871 = n44835 ;
  assign y14872 = n44838 ;
  assign y14873 = ~1'b0 ;
  assign y14874 = ~1'b0 ;
  assign y14875 = n44841 ;
  assign y14876 = n44846 ;
  assign y14877 = ~n44849 ;
  assign y14878 = ~n44852 ;
  assign y14879 = ~1'b0 ;
  assign y14880 = n44854 ;
  assign y14881 = ~n44856 ;
  assign y14882 = ~1'b0 ;
  assign y14883 = n44857 ;
  assign y14884 = ~n44861 ;
  assign y14885 = n44865 ;
  assign y14886 = ~n44866 ;
  assign y14887 = ~n44870 ;
  assign y14888 = n44873 ;
  assign y14889 = ~1'b0 ;
  assign y14890 = ~n44875 ;
  assign y14891 = ~n44879 ;
  assign y14892 = ~1'b0 ;
  assign y14893 = ~n44883 ;
  assign y14894 = n44885 ;
  assign y14895 = ~n44893 ;
  assign y14896 = ~n44896 ;
  assign y14897 = ~n44901 ;
  assign y14898 = n44902 ;
  assign y14899 = ~1'b0 ;
  assign y14900 = ~n44903 ;
  assign y14901 = ~1'b0 ;
  assign y14902 = n44905 ;
  assign y14903 = n44910 ;
  assign y14904 = n44911 ;
  assign y14905 = n44914 ;
  assign y14906 = ~n44915 ;
  assign y14907 = n44917 ;
  assign y14908 = n44918 ;
  assign y14909 = ~n44919 ;
  assign y14910 = ~n44921 ;
  assign y14911 = ~n44922 ;
  assign y14912 = ~n44923 ;
  assign y14913 = ~n44927 ;
  assign y14914 = ~1'b0 ;
  assign y14915 = ~n44932 ;
  assign y14916 = ~1'b0 ;
  assign y14917 = ~n44934 ;
  assign y14918 = ~n44935 ;
  assign y14919 = ~n44939 ;
  assign y14920 = ~n44940 ;
  assign y14921 = ~n44941 ;
  assign y14922 = ~1'b0 ;
  assign y14923 = ~n44942 ;
  assign y14924 = ~1'b0 ;
  assign y14925 = ~n44944 ;
  assign y14926 = ~1'b0 ;
  assign y14927 = n44948 ;
  assign y14928 = n44949 ;
  assign y14929 = n44952 ;
  assign y14930 = n44953 ;
  assign y14931 = ~n44954 ;
  assign y14932 = ~n44955 ;
  assign y14933 = ~n44956 ;
  assign y14934 = n44957 ;
  assign y14935 = ~1'b0 ;
  assign y14936 = ~n44958 ;
  assign y14937 = n44960 ;
  assign y14938 = ~n44966 ;
  assign y14939 = ~n44969 ;
  assign y14940 = n44972 ;
  assign y14941 = ~1'b0 ;
  assign y14942 = ~n44975 ;
  assign y14943 = ~1'b0 ;
  assign y14944 = n44977 ;
  assign y14945 = n44978 ;
  assign y14946 = ~n44981 ;
  assign y14947 = n44982 ;
  assign y14948 = ~n44983 ;
  assign y14949 = n44985 ;
  assign y14950 = n44987 ;
  assign y14951 = n44990 ;
  assign y14952 = ~n44992 ;
  assign y14953 = ~n44993 ;
  assign y14954 = ~n44994 ;
  assign y14955 = ~n44998 ;
  assign y14956 = ~n45001 ;
  assign y14957 = n45002 ;
  assign y14958 = n26295 ;
  assign y14959 = ~1'b0 ;
  assign y14960 = n45004 ;
  assign y14961 = n45006 ;
  assign y14962 = n45007 ;
  assign y14963 = ~n45010 ;
  assign y14964 = ~n45012 ;
  assign y14965 = ~n45016 ;
  assign y14966 = ~n45017 ;
  assign y14967 = ~1'b0 ;
  assign y14968 = ~1'b0 ;
  assign y14969 = ~n45019 ;
  assign y14970 = n45022 ;
  assign y14971 = ~n45026 ;
  assign y14972 = n45028 ;
  assign y14973 = n45032 ;
  assign y14974 = n45033 ;
  assign y14975 = ~1'b0 ;
  assign y14976 = ~1'b0 ;
  assign y14977 = n45034 ;
  assign y14978 = n45035 ;
  assign y14979 = n45037 ;
  assign y14980 = ~n45041 ;
  assign y14981 = ~n45042 ;
  assign y14982 = ~n45043 ;
  assign y14983 = ~n45045 ;
  assign y14984 = n45046 ;
  assign y14985 = ~n45048 ;
  assign y14986 = ~n45053 ;
  assign y14987 = n45054 ;
  assign y14988 = n45055 ;
  assign y14989 = n45057 ;
  assign y14990 = ~n45064 ;
  assign y14991 = n45066 ;
  assign y14992 = n45069 ;
  assign y14993 = ~n45071 ;
  assign y14994 = ~n45072 ;
  assign y14995 = ~n45077 ;
  assign y14996 = ~n45078 ;
  assign y14997 = ~n45079 ;
  assign y14998 = n45081 ;
  assign y14999 = ~n45086 ;
  assign y15000 = ~1'b0 ;
  assign y15001 = n45091 ;
  assign y15002 = n45092 ;
  assign y15003 = n45094 ;
  assign y15004 = ~n45098 ;
  assign y15005 = ~n45099 ;
  assign y15006 = n45100 ;
  assign y15007 = ~n45102 ;
  assign y15008 = ~n45103 ;
  assign y15009 = ~n45104 ;
  assign y15010 = ~1'b0 ;
  assign y15011 = ~1'b0 ;
  assign y15012 = ~n45107 ;
  assign y15013 = ~n45113 ;
  assign y15014 = n45115 ;
  assign y15015 = ~n45118 ;
  assign y15016 = ~n45125 ;
  assign y15017 = ~n45126 ;
  assign y15018 = n45131 ;
  assign y15019 = 1'b0 ;
  assign y15020 = ~n45133 ;
  assign y15021 = ~1'b0 ;
  assign y15022 = n45135 ;
  assign y15023 = ~n45143 ;
  assign y15024 = n45144 ;
  assign y15025 = ~n45145 ;
  assign y15026 = ~n45146 ;
  assign y15027 = n45151 ;
  assign y15028 = n45155 ;
  assign y15029 = n45156 ;
  assign y15030 = ~1'b0 ;
  assign y15031 = ~n45159 ;
  assign y15032 = n45161 ;
  assign y15033 = ~n45166 ;
  assign y15034 = ~1'b0 ;
  assign y15035 = n45168 ;
  assign y15036 = n45169 ;
  assign y15037 = ~n45176 ;
  assign y15038 = ~n45177 ;
  assign y15039 = ~n45178 ;
  assign y15040 = ~n45179 ;
  assign y15041 = n45182 ;
  assign y15042 = n45184 ;
  assign y15043 = ~n45186 ;
  assign y15044 = ~n45191 ;
  assign y15045 = ~n45193 ;
  assign y15046 = n45197 ;
  assign y15047 = n45200 ;
  assign y15048 = ~n45201 ;
  assign y15049 = ~n45206 ;
  assign y15050 = ~1'b0 ;
  assign y15051 = ~n45207 ;
  assign y15052 = n45209 ;
  assign y15053 = n45217 ;
  assign y15054 = n45218 ;
  assign y15055 = n45219 ;
  assign y15056 = n45220 ;
  assign y15057 = ~n45225 ;
  assign y15058 = ~n45227 ;
  assign y15059 = ~1'b0 ;
  assign y15060 = ~1'b0 ;
  assign y15061 = ~n45228 ;
  assign y15062 = n45231 ;
  assign y15063 = n45232 ;
  assign y15064 = n45236 ;
  assign y15065 = ~n45239 ;
  assign y15066 = ~n45242 ;
  assign y15067 = n45251 ;
  assign y15068 = ~1'b0 ;
  assign y15069 = ~n19097 ;
  assign y15070 = ~n45254 ;
  assign y15071 = n45255 ;
  assign y15072 = n45257 ;
  assign y15073 = n45259 ;
  assign y15074 = ~1'b0 ;
  assign y15075 = ~n45261 ;
  assign y15076 = ~n45266 ;
  assign y15077 = ~n45268 ;
  assign y15078 = n45271 ;
  assign y15079 = ~n45274 ;
  assign y15080 = ~n45275 ;
  assign y15081 = ~1'b0 ;
  assign y15082 = ~1'b0 ;
  assign y15083 = ~n45277 ;
  assign y15084 = n45285 ;
  assign y15085 = ~n45287 ;
  assign y15086 = ~n45288 ;
  assign y15087 = n45289 ;
  assign y15088 = n45290 ;
  assign y15089 = n45295 ;
  assign y15090 = ~1'b0 ;
  assign y15091 = ~n45296 ;
  assign y15092 = n33818 ;
  assign y15093 = n45298 ;
  assign y15094 = ~n45300 ;
  assign y15095 = n45302 ;
  assign y15096 = ~n45303 ;
  assign y15097 = n45307 ;
  assign y15098 = ~n45310 ;
  assign y15099 = ~n37205 ;
  assign y15100 = n45312 ;
  assign y15101 = n45317 ;
  assign y15102 = ~n45318 ;
  assign y15103 = n45319 ;
  assign y15104 = n45321 ;
  assign y15105 = n45326 ;
  assign y15106 = ~n45328 ;
  assign y15107 = n45330 ;
  assign y15108 = n45331 ;
  assign y15109 = ~1'b0 ;
  assign y15110 = n45332 ;
  assign y15111 = ~n4376 ;
  assign y15112 = ~n45337 ;
  assign y15113 = ~n45340 ;
  assign y15114 = n45343 ;
  assign y15115 = n45344 ;
  assign y15116 = ~n45346 ;
  assign y15117 = ~1'b0 ;
  assign y15118 = n45348 ;
  assign y15119 = n45349 ;
  assign y15120 = ~1'b0 ;
  assign y15121 = n45353 ;
  assign y15122 = ~n45356 ;
  assign y15123 = ~n45359 ;
  assign y15124 = ~n45361 ;
  assign y15125 = n45365 ;
  assign y15126 = n45367 ;
  assign y15127 = ~1'b0 ;
  assign y15128 = ~n45370 ;
  assign y15129 = n45372 ;
  assign y15130 = ~n45375 ;
  assign y15131 = n45376 ;
  assign y15132 = n45378 ;
  assign y15133 = ~n45380 ;
  assign y15134 = ~n45381 ;
  assign y15135 = ~n45383 ;
  assign y15136 = ~n45385 ;
  assign y15137 = ~1'b0 ;
  assign y15138 = ~1'b0 ;
  assign y15139 = ~n45386 ;
  assign y15140 = n45390 ;
  assign y15141 = ~1'b0 ;
  assign y15142 = ~n45391 ;
  assign y15143 = ~1'b0 ;
  assign y15144 = n45393 ;
  assign y15145 = ~1'b0 ;
  assign y15146 = n45397 ;
  assign y15147 = ~n45400 ;
  assign y15148 = ~n45404 ;
  assign y15149 = ~n45405 ;
  assign y15150 = n45409 ;
  assign y15151 = ~1'b0 ;
  assign y15152 = ~n45412 ;
  assign y15153 = n45414 ;
  assign y15154 = ~1'b0 ;
  assign y15155 = ~n45418 ;
  assign y15156 = n45422 ;
  assign y15157 = n45432 ;
  assign y15158 = n45438 ;
  assign y15159 = n45440 ;
  assign y15160 = ~n45441 ;
  assign y15161 = ~n45442 ;
  assign y15162 = n45444 ;
  assign y15163 = n45445 ;
  assign y15164 = n45450 ;
  assign y15165 = n45451 ;
  assign y15166 = ~n45453 ;
  assign y15167 = n45454 ;
  assign y15168 = n45456 ;
  assign y15169 = ~1'b0 ;
  assign y15170 = ~n45457 ;
  assign y15171 = ~1'b0 ;
  assign y15172 = n45458 ;
  assign y15173 = ~n45463 ;
  assign y15174 = ~n45467 ;
  assign y15175 = ~n45472 ;
  assign y15176 = ~n45473 ;
  assign y15177 = n45474 ;
  assign y15178 = n45482 ;
  assign y15179 = ~n45483 ;
  assign y15180 = ~1'b0 ;
  assign y15181 = n45486 ;
  assign y15182 = ~1'b0 ;
  assign y15183 = 1'b0 ;
  assign y15184 = ~n45487 ;
  assign y15185 = ~n45489 ;
  assign y15186 = n45491 ;
  assign y15187 = ~n45492 ;
  assign y15188 = ~n45496 ;
  assign y15189 = ~n45497 ;
  assign y15190 = n45499 ;
  assign y15191 = n45501 ;
  assign y15192 = ~n45504 ;
  assign y15193 = n45505 ;
  assign y15194 = ~n45511 ;
  assign y15195 = n45515 ;
  assign y15196 = ~1'b0 ;
  assign y15197 = n45517 ;
  assign y15198 = n45519 ;
  assign y15199 = ~n45521 ;
  assign y15200 = ~n45524 ;
  assign y15201 = ~n43872 ;
  assign y15202 = n45525 ;
  assign y15203 = n45526 ;
  assign y15204 = n45530 ;
  assign y15205 = ~n45531 ;
  assign y15206 = ~n45534 ;
  assign y15207 = ~n45536 ;
  assign y15208 = ~1'b0 ;
  assign y15209 = ~1'b0 ;
  assign y15210 = ~n45538 ;
  assign y15211 = ~n45541 ;
  assign y15212 = n45545 ;
  assign y15213 = n45547 ;
  assign y15214 = ~n45557 ;
  assign y15215 = n45562 ;
  assign y15216 = ~1'b0 ;
  assign y15217 = ~n45564 ;
  assign y15218 = n45567 ;
  assign y15219 = ~1'b0 ;
  assign y15220 = ~1'b0 ;
  assign y15221 = ~n45568 ;
  assign y15222 = ~n45569 ;
  assign y15223 = n45571 ;
  assign y15224 = n45572 ;
  assign y15225 = n45575 ;
  assign y15226 = ~n45577 ;
  assign y15227 = ~n45579 ;
  assign y15228 = ~n45581 ;
  assign y15229 = ~n45585 ;
  assign y15230 = ~n45586 ;
  assign y15231 = ~n45587 ;
  assign y15232 = ~n45590 ;
  assign y15233 = ~n45591 ;
  assign y15234 = ~n11452 ;
  assign y15235 = n45592 ;
  assign y15236 = n45593 ;
  assign y15237 = ~1'b0 ;
  assign y15238 = n45598 ;
  assign y15239 = ~n45603 ;
  assign y15240 = n45604 ;
  assign y15241 = ~n45607 ;
  assign y15242 = ~n45608 ;
  assign y15243 = ~n45610 ;
  assign y15244 = ~n45613 ;
  assign y15245 = n22004 ;
  assign y15246 = ~n45618 ;
  assign y15247 = ~n45620 ;
  assign y15248 = ~n45621 ;
  assign y15249 = n45623 ;
  assign y15250 = ~n45624 ;
  assign y15251 = n45625 ;
  assign y15252 = n45626 ;
  assign y15253 = ~n45628 ;
  assign y15254 = ~1'b0 ;
  assign y15255 = ~n45630 ;
  assign y15256 = n45634 ;
  assign y15257 = n45637 ;
  assign y15258 = n45639 ;
  assign y15259 = n45643 ;
  assign y15260 = ~n45645 ;
  assign y15261 = ~n45647 ;
  assign y15262 = ~n45648 ;
  assign y15263 = ~n45652 ;
  assign y15264 = n45655 ;
  assign y15265 = ~1'b0 ;
  assign y15266 = ~n45659 ;
  assign y15267 = n45661 ;
  assign y15268 = ~n45664 ;
  assign y15269 = ~n45673 ;
  assign y15270 = n45674 ;
  assign y15271 = n45678 ;
  assign y15272 = n45679 ;
  assign y15273 = n45680 ;
  assign y15274 = ~1'b0 ;
  assign y15275 = ~1'b0 ;
  assign y15276 = ~1'b0 ;
  assign y15277 = ~n45681 ;
  assign y15278 = n45682 ;
  assign y15279 = n45683 ;
  assign y15280 = n45685 ;
  assign y15281 = ~n45689 ;
  assign y15282 = ~n45695 ;
  assign y15283 = ~1'b0 ;
  assign y15284 = ~n45701 ;
  assign y15285 = ~1'b0 ;
  assign y15286 = n45705 ;
  assign y15287 = ~n45711 ;
  assign y15288 = n45713 ;
  assign y15289 = ~n45717 ;
  assign y15290 = n45719 ;
  assign y15291 = ~1'b0 ;
  assign y15292 = ~1'b0 ;
  assign y15293 = n45721 ;
  assign y15294 = ~1'b0 ;
  assign y15295 = n45722 ;
  assign y15296 = n45724 ;
  assign y15297 = ~n45726 ;
  assign y15298 = ~n45730 ;
  assign y15299 = ~n45731 ;
  assign y15300 = ~n45732 ;
  assign y15301 = ~1'b0 ;
  assign y15302 = ~n45735 ;
  assign y15303 = n45737 ;
  assign y15304 = n5459 ;
  assign y15305 = n45739 ;
  assign y15306 = n45741 ;
  assign y15307 = ~n45742 ;
  assign y15308 = n45743 ;
  assign y15309 = ~n45745 ;
  assign y15310 = n45746 ;
  assign y15311 = ~n45747 ;
  assign y15312 = ~n45749 ;
  assign y15313 = ~1'b0 ;
  assign y15314 = ~n45751 ;
  assign y15315 = ~n45756 ;
  assign y15316 = ~n45757 ;
  assign y15317 = ~n45758 ;
  assign y15318 = n45760 ;
  assign y15319 = ~n45762 ;
  assign y15320 = ~n45764 ;
  assign y15321 = n45766 ;
  assign y15322 = ~n45768 ;
  assign y15323 = n45774 ;
  assign y15324 = ~1'b0 ;
  assign y15325 = n45780 ;
  assign y15326 = ~n45784 ;
  assign y15327 = ~n45787 ;
  assign y15328 = n45789 ;
  assign y15329 = ~n45791 ;
  assign y15330 = ~n45795 ;
  assign y15331 = ~n45798 ;
  assign y15332 = ~n45800 ;
  assign y15333 = ~n45801 ;
  assign y15334 = n45804 ;
  assign y15335 = ~n45806 ;
  assign y15336 = n45808 ;
  assign y15337 = n45809 ;
  assign y15338 = ~n45810 ;
  assign y15339 = ~n45812 ;
  assign y15340 = ~n45815 ;
  assign y15341 = ~n45820 ;
  assign y15342 = n45822 ;
  assign y15343 = ~1'b0 ;
  assign y15344 = ~n45824 ;
  assign y15345 = n45825 ;
  assign y15346 = n45832 ;
  assign y15347 = ~n45835 ;
  assign y15348 = n45836 ;
  assign y15349 = ~n45841 ;
  assign y15350 = ~n45843 ;
  assign y15351 = ~1'b0 ;
  assign y15352 = n45845 ;
  assign y15353 = n45847 ;
  assign y15354 = ~1'b0 ;
  assign y15355 = n45848 ;
  assign y15356 = n45849 ;
  assign y15357 = ~n45850 ;
  assign y15358 = ~n45852 ;
  assign y15359 = n45854 ;
  assign y15360 = ~1'b0 ;
  assign y15361 = n45856 ;
  assign y15362 = ~n45859 ;
  assign y15363 = ~1'b0 ;
  assign y15364 = ~n45862 ;
  assign y15365 = ~n45864 ;
  assign y15366 = n45867 ;
  assign y15367 = n45869 ;
  assign y15368 = n45875 ;
  assign y15369 = ~n45876 ;
  assign y15370 = ~n45879 ;
  assign y15371 = ~n45881 ;
  assign y15372 = n45890 ;
  assign y15373 = n45892 ;
  assign y15374 = n45893 ;
  assign y15375 = n45894 ;
  assign y15376 = ~1'b0 ;
  assign y15377 = ~1'b0 ;
  assign y15378 = n45896 ;
  assign y15379 = n45900 ;
  assign y15380 = n45902 ;
  assign y15381 = ~n45906 ;
  assign y15382 = n45907 ;
  assign y15383 = ~n45909 ;
  assign y15384 = n45911 ;
  assign y15385 = ~n45916 ;
  assign y15386 = ~n45918 ;
  assign y15387 = ~n45920 ;
  assign y15388 = ~n45923 ;
  assign y15389 = n45925 ;
  assign y15390 = n45926 ;
  assign y15391 = n45928 ;
  assign y15392 = n45929 ;
  assign y15393 = ~n45933 ;
  assign y15394 = ~n45935 ;
  assign y15395 = ~n45937 ;
  assign y15396 = ~1'b0 ;
  assign y15397 = n45939 ;
  assign y15398 = ~1'b0 ;
  assign y15399 = ~1'b0 ;
  assign y15400 = n45941 ;
  assign y15401 = ~n45944 ;
  assign y15402 = n45945 ;
  assign y15403 = n45948 ;
  assign y15404 = n45951 ;
  assign y15405 = ~1'b0 ;
  assign y15406 = n45953 ;
  assign y15407 = n45956 ;
  assign y15408 = n45957 ;
  assign y15409 = ~n45958 ;
  assign y15410 = n45959 ;
  assign y15411 = ~n45960 ;
  assign y15412 = ~n45832 ;
  assign y15413 = n45963 ;
  assign y15414 = n45964 ;
  assign y15415 = ~n45967 ;
  assign y15416 = n45969 ;
  assign y15417 = n45975 ;
  assign y15418 = n45977 ;
  assign y15419 = ~n45979 ;
  assign y15420 = n45984 ;
  assign y15421 = n45985 ;
  assign y15422 = ~n45986 ;
  assign y15423 = n45987 ;
  assign y15424 = ~1'b0 ;
  assign y15425 = ~n45989 ;
  assign y15426 = ~n45990 ;
  assign y15427 = n45991 ;
  assign y15428 = n45995 ;
  assign y15429 = ~n45996 ;
  assign y15430 = n45997 ;
  assign y15431 = n32298 ;
  assign y15432 = n46000 ;
  assign y15433 = n46004 ;
  assign y15434 = n46007 ;
  assign y15435 = n46008 ;
  assign y15436 = n46009 ;
  assign y15437 = ~n46010 ;
  assign y15438 = ~n46016 ;
  assign y15439 = ~n46017 ;
  assign y15440 = n46018 ;
  assign y15441 = ~n46019 ;
  assign y15442 = ~1'b0 ;
  assign y15443 = ~n46022 ;
  assign y15444 = ~1'b0 ;
  assign y15445 = ~n46023 ;
  assign y15446 = n46025 ;
  assign y15447 = ~n46028 ;
  assign y15448 = n46029 ;
  assign y15449 = ~n46031 ;
  assign y15450 = n46032 ;
  assign y15451 = ~1'b0 ;
  assign y15452 = n46034 ;
  assign y15453 = ~n46042 ;
  assign y15454 = n46044 ;
  assign y15455 = n46045 ;
  assign y15456 = n41023 ;
  assign y15457 = n46046 ;
  assign y15458 = ~n46054 ;
  assign y15459 = ~n21666 ;
  assign y15460 = ~1'b0 ;
  assign y15461 = ~n46055 ;
  assign y15462 = ~n46062 ;
  assign y15463 = n46063 ;
  assign y15464 = ~n46064 ;
  assign y15465 = ~1'b0 ;
  assign y15466 = ~n46066 ;
  assign y15467 = n46068 ;
  assign y15468 = n46069 ;
  assign y15469 = ~n46071 ;
  assign y15470 = n46073 ;
  assign y15471 = ~n46081 ;
  assign y15472 = ~n46085 ;
  assign y15473 = ~n46087 ;
  assign y15474 = n46091 ;
  assign y15475 = n46093 ;
  assign y15476 = n46094 ;
  assign y15477 = n46098 ;
  assign y15478 = ~n46102 ;
  assign y15479 = ~n46103 ;
  assign y15480 = ~n46105 ;
  assign y15481 = ~1'b0 ;
  assign y15482 = ~1'b0 ;
  assign y15483 = ~n46107 ;
  assign y15484 = n46109 ;
  assign y15485 = n46113 ;
  assign y15486 = n46117 ;
  assign y15487 = n46120 ;
  assign y15488 = ~n46121 ;
  assign y15489 = ~n46122 ;
  assign y15490 = ~n24543 ;
  assign y15491 = ~1'b0 ;
  assign y15492 = n46124 ;
  assign y15493 = ~n46126 ;
  assign y15494 = n46128 ;
  assign y15495 = n46133 ;
  assign y15496 = n46134 ;
  assign y15497 = ~n46136 ;
  assign y15498 = ~1'b0 ;
  assign y15499 = ~1'b0 ;
  assign y15500 = ~1'b0 ;
  assign y15501 = n46138 ;
  assign y15502 = ~n46147 ;
  assign y15503 = n46150 ;
  assign y15504 = ~n46154 ;
  assign y15505 = ~n46161 ;
  assign y15506 = n46163 ;
  assign y15507 = n46164 ;
  assign y15508 = n46169 ;
  assign y15509 = n46170 ;
  assign y15510 = ~1'b0 ;
  assign y15511 = ~n46172 ;
  assign y15512 = ~n46177 ;
  assign y15513 = ~n46179 ;
  assign y15514 = ~n46182 ;
  assign y15515 = ~n46186 ;
  assign y15516 = ~n46187 ;
  assign y15517 = ~1'b0 ;
  assign y15518 = ~n46189 ;
  assign y15519 = n46192 ;
  assign y15520 = ~n46196 ;
  assign y15521 = n46197 ;
  assign y15522 = n46198 ;
  assign y15523 = ~n46202 ;
  assign y15524 = ~n46205 ;
  assign y15525 = ~n46206 ;
  assign y15526 = ~n46208 ;
  assign y15527 = ~n46210 ;
  assign y15528 = n46215 ;
  assign y15529 = ~n46216 ;
  assign y15530 = n46219 ;
  assign y15531 = ~n46220 ;
  assign y15532 = n46221 ;
  assign y15533 = n8757 ;
  assign y15534 = ~n46223 ;
  assign y15535 = ~n46225 ;
  assign y15536 = ~n46227 ;
  assign y15537 = ~1'b0 ;
  assign y15538 = n46228 ;
  assign y15539 = n46229 ;
  assign y15540 = ~n46230 ;
  assign y15541 = ~1'b0 ;
  assign y15542 = ~n46231 ;
  assign y15543 = ~n46233 ;
  assign y15544 = ~1'b0 ;
  assign y15545 = ~1'b0 ;
  assign y15546 = ~n46236 ;
  assign y15547 = ~n46239 ;
  assign y15548 = n46240 ;
  assign y15549 = ~n46246 ;
  assign y15550 = ~n46247 ;
  assign y15551 = ~n46250 ;
  assign y15552 = n46251 ;
  assign y15553 = ~n46254 ;
  assign y15554 = n46256 ;
  assign y15555 = ~1'b0 ;
  assign y15556 = n46260 ;
  assign y15557 = ~1'b0 ;
  assign y15558 = ~n46261 ;
  assign y15559 = ~n46262 ;
  assign y15560 = n46263 ;
  assign y15561 = ~n46265 ;
  assign y15562 = n46266 ;
  assign y15563 = n46268 ;
  assign y15564 = n46270 ;
  assign y15565 = ~1'b0 ;
  assign y15566 = ~n46275 ;
  assign y15567 = n46276 ;
  assign y15568 = ~n46277 ;
  assign y15569 = n46278 ;
  assign y15570 = n19316 ;
  assign y15571 = n46279 ;
  assign y15572 = ~n46281 ;
  assign y15573 = n46286 ;
  assign y15574 = ~1'b0 ;
  assign y15575 = n46289 ;
  assign y15576 = ~n46291 ;
  assign y15577 = n46295 ;
  assign y15578 = ~n46296 ;
  assign y15579 = ~1'b0 ;
  assign y15580 = ~1'b0 ;
  assign y15581 = ~n46299 ;
  assign y15582 = ~n46302 ;
  assign y15583 = ~n46303 ;
  assign y15584 = n46304 ;
  assign y15585 = n46307 ;
  assign y15586 = n46308 ;
  assign y15587 = ~n46309 ;
  assign y15588 = ~1'b0 ;
  assign y15589 = ~1'b0 ;
  assign y15590 = n46311 ;
  assign y15591 = n46313 ;
  assign y15592 = ~n46314 ;
  assign y15593 = ~n46316 ;
  assign y15594 = ~n46319 ;
  assign y15595 = ~n46320 ;
  assign y15596 = n46324 ;
  assign y15597 = ~n46325 ;
  assign y15598 = ~1'b0 ;
  assign y15599 = n46326 ;
  assign y15600 = ~1'b0 ;
  assign y15601 = ~n46327 ;
  assign y15602 = ~n46328 ;
  assign y15603 = n46330 ;
  assign y15604 = n46333 ;
  assign y15605 = ~1'b0 ;
  assign y15606 = ~n46335 ;
  assign y15607 = n46340 ;
  assign y15608 = ~n46343 ;
  assign y15609 = ~n46346 ;
  assign y15610 = n46348 ;
  assign y15611 = n46350 ;
  assign y15612 = ~n46351 ;
  assign y15613 = n46352 ;
  assign y15614 = ~1'b0 ;
  assign y15615 = n46354 ;
  assign y15616 = ~1'b0 ;
  assign y15617 = ~n46356 ;
  assign y15618 = ~n46360 ;
  assign y15619 = ~n46361 ;
  assign y15620 = ~n46362 ;
  assign y15621 = ~1'b0 ;
  assign y15622 = ~1'b0 ;
  assign y15623 = ~n46363 ;
  assign y15624 = ~1'b0 ;
  assign y15625 = n46364 ;
  assign y15626 = n46371 ;
  assign y15627 = n11578 ;
  assign y15628 = n46372 ;
  assign y15629 = n46375 ;
  assign y15630 = ~n46377 ;
  assign y15631 = ~1'b0 ;
  assign y15632 = ~n46384 ;
  assign y15633 = ~1'b0 ;
  assign y15634 = n46386 ;
  assign y15635 = n46390 ;
  assign y15636 = n46392 ;
  assign y15637 = ~n46394 ;
  assign y15638 = n46399 ;
  assign y15639 = ~n46400 ;
  assign y15640 = n46402 ;
  assign y15641 = ~n46405 ;
  assign y15642 = ~n46410 ;
  assign y15643 = ~n46412 ;
  assign y15644 = ~n46414 ;
  assign y15645 = n46418 ;
  assign y15646 = ~n46419 ;
  assign y15647 = ~n46424 ;
  assign y15648 = ~n46427 ;
  assign y15649 = n46430 ;
  assign y15650 = n46432 ;
  assign y15651 = ~n46435 ;
  assign y15652 = ~1'b0 ;
  assign y15653 = n46436 ;
  assign y15654 = ~n46440 ;
  assign y15655 = ~n46444 ;
  assign y15656 = ~1'b0 ;
  assign y15657 = ~n46447 ;
  assign y15658 = ~n46452 ;
  assign y15659 = ~n24089 ;
  assign y15660 = n46454 ;
  assign y15661 = n46455 ;
  assign y15662 = ~n46457 ;
  assign y15663 = ~1'b0 ;
  assign y15664 = ~n46460 ;
  assign y15665 = ~n46461 ;
  assign y15666 = ~n46462 ;
  assign y15667 = ~n46465 ;
  assign y15668 = ~n46467 ;
  assign y15669 = ~1'b0 ;
  assign y15670 = ~n46472 ;
  assign y15671 = ~1'b0 ;
  assign y15672 = ~n46475 ;
  assign y15673 = n46476 ;
  assign y15674 = n46477 ;
  assign y15675 = n46479 ;
  assign y15676 = ~n46481 ;
  assign y15677 = n46485 ;
  assign y15678 = n46486 ;
  assign y15679 = ~1'b0 ;
  assign y15680 = ~n46489 ;
  assign y15681 = ~n46490 ;
  assign y15682 = n46491 ;
  assign y15683 = n46497 ;
  assign y15684 = n46498 ;
  assign y15685 = ~n46499 ;
  assign y15686 = n46502 ;
  assign y15687 = ~n46505 ;
  assign y15688 = ~1'b0 ;
  assign y15689 = ~n46509 ;
  assign y15690 = ~1'b0 ;
  assign y15691 = ~n46513 ;
  assign y15692 = ~n46519 ;
  assign y15693 = ~n46520 ;
  assign y15694 = ~n46524 ;
  assign y15695 = n46525 ;
  assign y15696 = ~n17370 ;
  assign y15697 = ~1'b0 ;
  assign y15698 = n25594 ;
  assign y15699 = n46529 ;
  assign y15700 = ~1'b0 ;
  assign y15701 = ~n46530 ;
  assign y15702 = n46531 ;
  assign y15703 = ~n46533 ;
  assign y15704 = n46534 ;
  assign y15705 = ~n46538 ;
  assign y15706 = ~n46540 ;
  assign y15707 = n46542 ;
  assign y15708 = ~n46545 ;
  assign y15709 = ~n46547 ;
  assign y15710 = ~n46552 ;
  assign y15711 = ~n46556 ;
  assign y15712 = ~n46557 ;
  assign y15713 = ~n46560 ;
  assign y15714 = ~n46561 ;
  assign y15715 = n46564 ;
  assign y15716 = n46566 ;
  assign y15717 = ~n46568 ;
  assign y15718 = n46576 ;
  assign y15719 = ~n46580 ;
  assign y15720 = ~n46583 ;
  assign y15721 = n46585 ;
  assign y15722 = ~n46589 ;
  assign y15723 = ~n46590 ;
  assign y15724 = n46597 ;
  assign y15725 = n46600 ;
  assign y15726 = ~n15504 ;
  assign y15727 = n46603 ;
  assign y15728 = n46604 ;
  assign y15729 = n46607 ;
  assign y15730 = n46614 ;
  assign y15731 = ~1'b0 ;
  assign y15732 = n46618 ;
  assign y15733 = ~n46620 ;
  assign y15734 = ~n46621 ;
  assign y15735 = ~n46622 ;
  assign y15736 = n46623 ;
  assign y15737 = ~n46625 ;
  assign y15738 = ~n46632 ;
  assign y15739 = n46635 ;
  assign y15740 = n46638 ;
  assign y15741 = ~n46639 ;
  assign y15742 = n46645 ;
  assign y15743 = n46646 ;
  assign y15744 = n46647 ;
  assign y15745 = n46653 ;
  assign y15746 = n46655 ;
  assign y15747 = ~1'b0 ;
  assign y15748 = n46659 ;
  assign y15749 = ~n46662 ;
  assign y15750 = n46663 ;
  assign y15751 = n46665 ;
  assign y15752 = ~n46668 ;
  assign y15753 = ~n46669 ;
  assign y15754 = n46672 ;
  assign y15755 = ~1'b0 ;
  assign y15756 = ~1'b0 ;
  assign y15757 = ~n46679 ;
  assign y15758 = n46680 ;
  assign y15759 = n46682 ;
  assign y15760 = n46683 ;
  assign y15761 = ~n46684 ;
  assign y15762 = ~n46685 ;
  assign y15763 = n46688 ;
  assign y15764 = ~n46691 ;
  assign y15765 = ~n46696 ;
  assign y15766 = n46697 ;
  assign y15767 = n46699 ;
  assign y15768 = ~n46702 ;
  assign y15769 = n46703 ;
  assign y15770 = ~n46704 ;
  assign y15771 = n46705 ;
  assign y15772 = n46708 ;
  assign y15773 = ~1'b0 ;
  assign y15774 = ~1'b0 ;
  assign y15775 = ~n46710 ;
  assign y15776 = ~1'b0 ;
  assign y15777 = ~n46712 ;
  assign y15778 = n46718 ;
  assign y15779 = ~n46721 ;
  assign y15780 = n46726 ;
  assign y15781 = n46727 ;
  assign y15782 = n46730 ;
  assign y15783 = n46731 ;
  assign y15784 = ~n46733 ;
  assign y15785 = ~n46735 ;
  assign y15786 = ~n46737 ;
  assign y15787 = ~n46739 ;
  assign y15788 = n46740 ;
  assign y15789 = n46742 ;
  assign y15790 = ~n46743 ;
  assign y15791 = ~n46745 ;
  assign y15792 = ~n46747 ;
  assign y15793 = ~1'b0 ;
  assign y15794 = ~n46749 ;
  assign y15795 = ~1'b0 ;
  assign y15796 = n46751 ;
  assign y15797 = n46753 ;
  assign y15798 = n46754 ;
  assign y15799 = n46755 ;
  assign y15800 = n46757 ;
  assign y15801 = ~n46758 ;
  assign y15802 = n46760 ;
  assign y15803 = n46763 ;
  assign y15804 = ~1'b0 ;
  assign y15805 = n46765 ;
  assign y15806 = ~1'b0 ;
  assign y15807 = n46766 ;
  assign y15808 = n46771 ;
  assign y15809 = ~n46775 ;
  assign y15810 = ~n46780 ;
  assign y15811 = ~n46788 ;
  assign y15812 = ~n46794 ;
  assign y15813 = ~1'b0 ;
  assign y15814 = ~1'b0 ;
  assign y15815 = ~n46795 ;
  assign y15816 = ~1'b0 ;
  assign y15817 = n46798 ;
  assign y15818 = ~n46801 ;
  assign y15819 = n46802 ;
  assign y15820 = n46803 ;
  assign y15821 = n46806 ;
  assign y15822 = ~n46807 ;
  assign y15823 = ~n46812 ;
  assign y15824 = ~n46813 ;
  assign y15825 = ~1'b0 ;
  assign y15826 = ~1'b0 ;
  assign y15827 = ~n46814 ;
  assign y15828 = n46816 ;
  assign y15829 = ~n46819 ;
  assign y15830 = n46822 ;
  assign y15831 = ~n46825 ;
  assign y15832 = ~n46826 ;
  assign y15833 = ~n46831 ;
  assign y15834 = n46835 ;
  assign y15835 = ~1'b0 ;
  assign y15836 = ~n46836 ;
  assign y15837 = ~n46839 ;
  assign y15838 = n46840 ;
  assign y15839 = n46841 ;
  assign y15840 = n46844 ;
  assign y15841 = n46848 ;
  assign y15842 = ~n46849 ;
  assign y15843 = n46851 ;
  assign y15844 = n46854 ;
  assign y15845 = ~1'b0 ;
  assign y15846 = n46855 ;
  assign y15847 = ~n46857 ;
  assign y15848 = ~n46859 ;
  assign y15849 = n46860 ;
  assign y15850 = n46864 ;
  assign y15851 = n46866 ;
  assign y15852 = n46870 ;
  assign y15853 = ~n46873 ;
  assign y15854 = ~n46876 ;
  assign y15855 = ~n46880 ;
  assign y15856 = ~n46881 ;
  assign y15857 = n46882 ;
  assign y15858 = ~n46886 ;
  assign y15859 = ~n46887 ;
  assign y15860 = ~n46892 ;
  assign y15861 = ~1'b0 ;
  assign y15862 = ~1'b0 ;
  assign y15863 = ~n46894 ;
  assign y15864 = ~n46896 ;
  assign y15865 = ~n46897 ;
  assign y15866 = ~n46899 ;
  assign y15867 = n46901 ;
  assign y15868 = ~1'b0 ;
  assign y15869 = ~n46902 ;
  assign y15870 = ~n46907 ;
  assign y15871 = n46910 ;
  assign y15872 = n46912 ;
  assign y15873 = n46913 ;
  assign y15874 = n46916 ;
  assign y15875 = n46925 ;
  assign y15876 = ~n46931 ;
  assign y15877 = ~n46934 ;
  assign y15878 = n46938 ;
  assign y15879 = ~n46939 ;
  assign y15880 = n46942 ;
  assign y15881 = n46943 ;
  assign y15882 = n46944 ;
  assign y15883 = n46946 ;
  assign y15884 = n46948 ;
  assign y15885 = ~n46950 ;
  assign y15886 = ~n46951 ;
  assign y15887 = n46952 ;
  assign y15888 = n46961 ;
  assign y15889 = n46965 ;
  assign y15890 = n46966 ;
  assign y15891 = n46968 ;
  assign y15892 = ~n46969 ;
  assign y15893 = n46972 ;
  assign y15894 = n46974 ;
  assign y15895 = ~n46976 ;
  assign y15896 = n46982 ;
  assign y15897 = ~n46987 ;
  assign y15898 = ~n46989 ;
  assign y15899 = n46992 ;
  assign y15900 = ~n46994 ;
  assign y15901 = ~n46995 ;
  assign y15902 = ~n47011 ;
  assign y15903 = ~n47020 ;
  assign y15904 = ~1'b0 ;
  assign y15905 = ~n47022 ;
  assign y15906 = ~n47032 ;
  assign y15907 = n47033 ;
  assign y15908 = n47034 ;
  assign y15909 = n47036 ;
  assign y15910 = ~n47038 ;
  assign y15911 = n47043 ;
  assign y15912 = ~n47044 ;
  assign y15913 = ~n47047 ;
  assign y15914 = ~1'b0 ;
  assign y15915 = n47049 ;
  assign y15916 = n47050 ;
  assign y15917 = ~n47052 ;
  assign y15918 = ~n47054 ;
  assign y15919 = n47055 ;
  assign y15920 = ~n47056 ;
  assign y15921 = ~n47059 ;
  assign y15922 = ~n47064 ;
  assign y15923 = ~1'b0 ;
  assign y15924 = ~n35322 ;
  assign y15925 = n47066 ;
  assign y15926 = ~n47068 ;
  assign y15927 = n47072 ;
  assign y15928 = n47076 ;
  assign y15929 = ~n47077 ;
  assign y15930 = n47083 ;
  assign y15931 = n47084 ;
  assign y15932 = n47090 ;
  assign y15933 = n47092 ;
  assign y15934 = ~1'b0 ;
  assign y15935 = ~1'b0 ;
  assign y15936 = n47094 ;
  assign y15937 = ~n47096 ;
  assign y15938 = ~n47097 ;
  assign y15939 = ~n47098 ;
  assign y15940 = n47100 ;
  assign y15941 = ~n9569 ;
  assign y15942 = n47105 ;
  assign y15943 = ~n47107 ;
  assign y15944 = ~n47110 ;
  assign y15945 = ~n47112 ;
  assign y15946 = ~n47116 ;
  assign y15947 = ~n47119 ;
  assign y15948 = n47120 ;
  assign y15949 = ~n47121 ;
  assign y15950 = n47122 ;
  assign y15951 = ~n47132 ;
  assign y15952 = ~n47133 ;
  assign y15953 = ~1'b0 ;
  assign y15954 = ~1'b0 ;
  assign y15955 = ~n47135 ;
  assign y15956 = ~1'b0 ;
  assign y15957 = n47137 ;
  assign y15958 = n47138 ;
  assign y15959 = n47139 ;
  assign y15960 = ~n47140 ;
  assign y15961 = ~n47143 ;
  assign y15962 = n47147 ;
  assign y15963 = ~1'b0 ;
  assign y15964 = ~1'b0 ;
  assign y15965 = ~1'b0 ;
  assign y15966 = n47150 ;
  assign y15967 = ~n47153 ;
  assign y15968 = ~n47154 ;
  assign y15969 = n47159 ;
  assign y15970 = ~n47160 ;
  assign y15971 = ~n47163 ;
  assign y15972 = ~n47164 ;
  assign y15973 = ~1'b0 ;
  assign y15974 = ~n47166 ;
  assign y15975 = n47173 ;
  assign y15976 = ~n47178 ;
  assign y15977 = n47183 ;
  assign y15978 = ~n47184 ;
  assign y15979 = ~n47187 ;
  assign y15980 = ~n47188 ;
  assign y15981 = ~1'b0 ;
  assign y15982 = ~n47191 ;
  assign y15983 = ~n47193 ;
  assign y15984 = ~n47195 ;
  assign y15985 = ~n47197 ;
  assign y15986 = n47199 ;
  assign y15987 = ~n47200 ;
  assign y15988 = ~n47201 ;
  assign y15989 = n47204 ;
  assign y15990 = n47208 ;
  assign y15991 = ~n47209 ;
  assign y15992 = n47215 ;
  assign y15993 = n47216 ;
  assign y15994 = ~n47218 ;
  assign y15995 = n47221 ;
  assign y15996 = ~n47222 ;
  assign y15997 = ~n47223 ;
  assign y15998 = ~n47225 ;
  assign y15999 = n47226 ;
  assign y16000 = n47230 ;
  assign y16001 = ~1'b0 ;
  assign y16002 = n47233 ;
  assign y16003 = ~n47234 ;
  assign y16004 = n47235 ;
  assign y16005 = ~n47236 ;
  assign y16006 = ~n40680 ;
  assign y16007 = ~n47241 ;
  assign y16008 = ~n47243 ;
  assign y16009 = n47246 ;
  assign y16010 = ~1'b0 ;
  assign y16011 = n47248 ;
  assign y16012 = n47249 ;
  assign y16013 = n47251 ;
  assign y16014 = ~n47253 ;
  assign y16015 = ~n47255 ;
  assign y16016 = n47257 ;
  assign y16017 = ~n47258 ;
  assign y16018 = n47260 ;
  assign y16019 = ~1'b0 ;
  assign y16020 = ~n47263 ;
  assign y16021 = n47266 ;
  assign y16022 = n47267 ;
  assign y16023 = ~n47268 ;
  assign y16024 = ~n47271 ;
  assign y16025 = ~n47272 ;
  assign y16026 = n47276 ;
  assign y16027 = ~n47277 ;
  assign y16028 = ~n47280 ;
  assign y16029 = ~n47283 ;
  assign y16030 = ~n47287 ;
  assign y16031 = n47288 ;
  assign y16032 = ~n47290 ;
  assign y16033 = n47292 ;
  assign y16034 = ~n47293 ;
  assign y16035 = n47294 ;
  assign y16036 = n47295 ;
  assign y16037 = ~n47296 ;
  assign y16038 = n47297 ;
  assign y16039 = ~1'b0 ;
  assign y16040 = 1'b0 ;
  assign y16041 = n47301 ;
  assign y16042 = n47303 ;
  assign y16043 = ~n47304 ;
  assign y16044 = n47307 ;
  assign y16045 = ~n47308 ;
  assign y16046 = n47310 ;
  assign y16047 = ~n47313 ;
  assign y16048 = ~n6027 ;
  assign y16049 = ~1'b0 ;
  assign y16050 = n47316 ;
  assign y16051 = ~n47318 ;
  assign y16052 = n47319 ;
  assign y16053 = ~n47320 ;
  assign y16054 = n47322 ;
  assign y16055 = ~n47323 ;
  assign y16056 = n47327 ;
  assign y16057 = n47328 ;
  assign y16058 = ~n47332 ;
  assign y16059 = ~1'b0 ;
  assign y16060 = n47337 ;
  assign y16061 = ~n44203 ;
  assign y16062 = ~n47338 ;
  assign y16063 = n47341 ;
  assign y16064 = ~n47342 ;
  assign y16065 = ~n47343 ;
  assign y16066 = ~n47345 ;
  assign y16067 = n47346 ;
  assign y16068 = ~n47348 ;
  assign y16069 = n47351 ;
  assign y16070 = ~n47356 ;
  assign y16071 = ~1'b0 ;
  assign y16072 = ~1'b0 ;
  assign y16073 = n47359 ;
  assign y16074 = ~n47361 ;
  assign y16075 = n47362 ;
  assign y16076 = ~n47367 ;
  assign y16077 = ~n47368 ;
  assign y16078 = ~n47371 ;
  assign y16079 = ~n47372 ;
  assign y16080 = ~1'b0 ;
  assign y16081 = ~n47374 ;
  assign y16082 = ~1'b0 ;
  assign y16083 = n47378 ;
  assign y16084 = ~n47379 ;
  assign y16085 = n47380 ;
  assign y16086 = ~n33862 ;
  assign y16087 = n47382 ;
  assign y16088 = ~n47383 ;
  assign y16089 = ~n47386 ;
  assign y16090 = ~1'b0 ;
  assign y16091 = ~n47391 ;
  assign y16092 = ~1'b0 ;
  assign y16093 = n47393 ;
  assign y16094 = ~n47396 ;
  assign y16095 = n47398 ;
  assign y16096 = n47401 ;
  assign y16097 = ~n47402 ;
  assign y16098 = n47406 ;
  assign y16099 = n47408 ;
  assign y16100 = n47410 ;
  assign y16101 = n47413 ;
  assign y16102 = ~n47415 ;
  assign y16103 = ~1'b0 ;
  assign y16104 = ~1'b0 ;
  assign y16105 = ~n47421 ;
  assign y16106 = ~n47422 ;
  assign y16107 = ~n47425 ;
  assign y16108 = n47428 ;
  assign y16109 = n47430 ;
  assign y16110 = ~n47431 ;
  assign y16111 = ~n47438 ;
  assign y16112 = ~1'b0 ;
  assign y16113 = n47440 ;
  assign y16114 = ~1'b0 ;
  assign y16115 = n47444 ;
  assign y16116 = n47445 ;
  assign y16117 = ~n47446 ;
  assign y16118 = ~n47447 ;
  assign y16119 = ~n47448 ;
  assign y16120 = ~n47449 ;
  assign y16121 = ~1'b0 ;
  assign y16122 = ~n47451 ;
  assign y16123 = n47455 ;
  assign y16124 = n47459 ;
  assign y16125 = ~1'b0 ;
  assign y16126 = n47465 ;
  assign y16127 = ~n47466 ;
  assign y16128 = n47472 ;
  assign y16129 = n47473 ;
  assign y16130 = n47477 ;
  assign y16131 = n47479 ;
  assign y16132 = ~1'b0 ;
  assign y16133 = n47480 ;
  assign y16134 = ~1'b0 ;
  assign y16135 = ~n47481 ;
  assign y16136 = ~n47482 ;
  assign y16137 = ~n47483 ;
  assign y16138 = n47484 ;
  assign y16139 = ~n47485 ;
  assign y16140 = ~1'b0 ;
  assign y16141 = ~n47490 ;
  assign y16142 = ~1'b0 ;
  assign y16143 = ~n47493 ;
  assign y16144 = n47495 ;
  assign y16145 = n47496 ;
  assign y16146 = ~n47498 ;
  assign y16147 = n47499 ;
  assign y16148 = ~n47505 ;
  assign y16149 = ~n47511 ;
  assign y16150 = ~1'b0 ;
  assign y16151 = ~n47512 ;
  assign y16152 = n47513 ;
  assign y16153 = ~n47514 ;
  assign y16154 = n47517 ;
  assign y16155 = n47522 ;
  assign y16156 = ~n47525 ;
  assign y16157 = ~n47526 ;
  assign y16158 = ~n47527 ;
  assign y16159 = ~n47529 ;
  assign y16160 = n47532 ;
  assign y16161 = n47535 ;
  assign y16162 = ~1'b0 ;
  assign y16163 = ~n47538 ;
  assign y16164 = ~n47541 ;
  assign y16165 = n47543 ;
  assign y16166 = n47545 ;
  assign y16167 = ~n47555 ;
  assign y16168 = ~1'b0 ;
  assign y16169 = ~n47557 ;
  assign y16170 = n47558 ;
  assign y16171 = n47565 ;
  assign y16172 = ~n47567 ;
  assign y16173 = ~n47571 ;
  assign y16174 = ~n22830 ;
  assign y16175 = n47572 ;
  assign y16176 = ~n47573 ;
  assign y16177 = n47576 ;
  assign y16178 = n47580 ;
  assign y16179 = ~n47583 ;
  assign y16180 = ~1'b0 ;
  assign y16181 = ~n47586 ;
  assign y16182 = ~1'b0 ;
  assign y16183 = ~n47587 ;
  assign y16184 = ~n47590 ;
  assign y16185 = n47592 ;
  assign y16186 = n47596 ;
  assign y16187 = ~n47597 ;
  assign y16188 = n47598 ;
  assign y16189 = 1'b0 ;
  assign y16190 = ~n47600 ;
  assign y16191 = n47604 ;
  assign y16192 = ~1'b0 ;
  assign y16193 = n47606 ;
  assign y16194 = n47608 ;
  assign y16195 = ~n47610 ;
  assign y16196 = n47614 ;
  assign y16197 = n47618 ;
  assign y16198 = 1'b0 ;
  assign y16199 = ~n47619 ;
  assign y16200 = ~1'b0 ;
  assign y16201 = ~1'b0 ;
  assign y16202 = ~1'b0 ;
  assign y16203 = n47624 ;
  assign y16204 = ~n47630 ;
  assign y16205 = ~n47631 ;
  assign y16206 = n47632 ;
  assign y16207 = ~n47633 ;
  assign y16208 = ~n47637 ;
  assign y16209 = ~1'b0 ;
  assign y16210 = ~n47644 ;
  assign y16211 = ~1'b0 ;
  assign y16212 = ~1'b0 ;
  assign y16213 = ~n47653 ;
  assign y16214 = n47654 ;
  assign y16215 = ~n47655 ;
  assign y16216 = ~n47660 ;
  assign y16217 = ~n47662 ;
  assign y16218 = ~n47664 ;
  assign y16219 = n47667 ;
  assign y16220 = ~n47670 ;
  assign y16221 = ~n47672 ;
  assign y16222 = ~n47675 ;
  assign y16223 = n47677 ;
  assign y16224 = n47678 ;
  assign y16225 = n47681 ;
  assign y16226 = ~n47684 ;
  assign y16227 = ~n47687 ;
  assign y16228 = n47689 ;
  assign y16229 = n47690 ;
  assign y16230 = ~n47692 ;
  assign y16231 = n47695 ;
  assign y16232 = ~1'b0 ;
  assign y16233 = ~1'b0 ;
  assign y16234 = ~n47699 ;
  assign y16235 = n47700 ;
  assign y16236 = ~n47704 ;
  assign y16237 = n47709 ;
  assign y16238 = ~n47711 ;
  assign y16239 = ~n47713 ;
  assign y16240 = n47715 ;
  assign y16241 = ~1'b0 ;
  assign y16242 = n47717 ;
  assign y16243 = ~n47719 ;
  assign y16244 = n47722 ;
  assign y16245 = ~n47723 ;
  assign y16246 = n47725 ;
  assign y16247 = ~n47726 ;
  assign y16248 = ~n47729 ;
  assign y16249 = ~n47736 ;
  assign y16250 = n47739 ;
  assign y16251 = n47740 ;
  assign y16252 = n47742 ;
  assign y16253 = n47749 ;
  assign y16254 = n47753 ;
  assign y16255 = ~n47755 ;
  assign y16256 = ~n47757 ;
  assign y16257 = n47758 ;
  assign y16258 = n47763 ;
  assign y16259 = ~n47764 ;
  assign y16260 = n47773 ;
  assign y16261 = n47778 ;
  assign y16262 = n47780 ;
  assign y16263 = n47782 ;
  assign y16264 = ~n47783 ;
  assign y16265 = ~n47785 ;
  assign y16266 = ~n47788 ;
  assign y16267 = ~n47791 ;
  assign y16268 = n47800 ;
  assign y16269 = ~n47802 ;
  assign y16270 = n47803 ;
  assign y16271 = n47810 ;
  assign y16272 = ~n47812 ;
  assign y16273 = n47813 ;
  assign y16274 = ~1'b0 ;
  assign y16275 = ~n47817 ;
  assign y16276 = n47819 ;
  assign y16277 = ~n47821 ;
  assign y16278 = ~n47823 ;
  assign y16279 = n47825 ;
  assign y16280 = n47828 ;
  assign y16281 = ~n47829 ;
  assign y16282 = n47832 ;
  assign y16283 = n47837 ;
  assign y16284 = ~1'b0 ;
  assign y16285 = n47842 ;
  assign y16286 = ~n47845 ;
  assign y16287 = n47847 ;
  assign y16288 = n47848 ;
  assign y16289 = ~n47852 ;
  assign y16290 = ~n47854 ;
  assign y16291 = n47855 ;
  assign y16292 = ~n47856 ;
  assign y16293 = n47860 ;
  assign y16294 = ~x85 ;
  assign y16295 = n47862 ;
  assign y16296 = ~1'b0 ;
  assign y16297 = ~n47864 ;
  assign y16298 = n47867 ;
  assign y16299 = ~n47870 ;
  assign y16300 = ~n47871 ;
  assign y16301 = ~n47877 ;
  assign y16302 = n47881 ;
  assign y16303 = ~n47884 ;
  assign y16304 = ~1'b0 ;
  assign y16305 = ~1'b0 ;
  assign y16306 = n47887 ;
  assign y16307 = ~n47888 ;
  assign y16308 = ~n47889 ;
  assign y16309 = ~n47891 ;
  assign y16310 = ~n47892 ;
  assign y16311 = ~n47895 ;
  assign y16312 = n47896 ;
  assign y16313 = ~1'b0 ;
  assign y16314 = n47898 ;
  assign y16315 = ~n47901 ;
  assign y16316 = n47902 ;
  assign y16317 = ~n47904 ;
  assign y16318 = ~n47907 ;
  assign y16319 = ~n47908 ;
  assign y16320 = n47909 ;
  assign y16321 = n47910 ;
  assign y16322 = ~n47916 ;
  assign y16323 = ~n47918 ;
  assign y16324 = n47925 ;
  assign y16325 = n47926 ;
  assign y16326 = ~n47929 ;
  assign y16327 = n47936 ;
  assign y16328 = n47939 ;
  assign y16329 = ~n47942 ;
  assign y16330 = ~n47945 ;
  assign y16331 = ~n47947 ;
  assign y16332 = n47948 ;
  assign y16333 = ~n47950 ;
  assign y16334 = ~1'b0 ;
  assign y16335 = ~n47951 ;
  assign y16336 = n47953 ;
  assign y16337 = ~n47965 ;
  assign y16338 = ~n47968 ;
  assign y16339 = n47969 ;
  assign y16340 = n47970 ;
  assign y16341 = ~n47974 ;
  assign y16342 = n47981 ;
  assign y16343 = ~1'b0 ;
  assign y16344 = n47983 ;
  assign y16345 = n47984 ;
  assign y16346 = ~n47985 ;
  assign y16347 = ~n47986 ;
  assign y16348 = n47988 ;
  assign y16349 = ~n47989 ;
  assign y16350 = ~1'b0 ;
  assign y16351 = ~n47990 ;
  assign y16352 = ~1'b0 ;
  assign y16353 = ~1'b0 ;
  assign y16354 = ~n47991 ;
  assign y16355 = n47992 ;
  assign y16356 = n47993 ;
  assign y16357 = ~1'b0 ;
  assign y16358 = ~n47994 ;
  assign y16359 = ~n47995 ;
  assign y16360 = ~n47997 ;
  assign y16361 = ~1'b0 ;
  assign y16362 = n47998 ;
  assign y16363 = ~n47999 ;
  assign y16364 = ~n48000 ;
  assign y16365 = ~n48003 ;
  assign y16366 = ~n48005 ;
  assign y16367 = ~n48006 ;
  assign y16368 = ~n48010 ;
  assign y16369 = n48012 ;
  assign y16370 = ~1'b0 ;
  assign y16371 = n48014 ;
  assign y16372 = ~1'b0 ;
  assign y16373 = ~n48015 ;
  assign y16374 = n48018 ;
  assign y16375 = n48019 ;
  assign y16376 = n48020 ;
  assign y16377 = n48021 ;
  assign y16378 = ~1'b0 ;
  assign y16379 = ~1'b0 ;
  assign y16380 = ~n48025 ;
  assign y16381 = ~n48026 ;
  assign y16382 = ~n48030 ;
  assign y16383 = ~1'b0 ;
  assign y16384 = ~n48031 ;
  assign y16385 = n48034 ;
  assign y16386 = n48037 ;
  assign y16387 = ~n48039 ;
  assign y16388 = ~1'b0 ;
  assign y16389 = ~n48042 ;
  assign y16390 = ~n48043 ;
  assign y16391 = ~n48045 ;
  assign y16392 = n45693 ;
  assign y16393 = n48051 ;
  assign y16394 = n48054 ;
  assign y16395 = n48055 ;
  assign y16396 = ~1'b0 ;
  assign y16397 = ~1'b0 ;
  assign y16398 = ~1'b0 ;
  assign y16399 = ~n48056 ;
  assign y16400 = n48061 ;
  assign y16401 = ~n48063 ;
  assign y16402 = n48066 ;
  assign y16403 = n48067 ;
  assign y16404 = n48074 ;
  assign y16405 = n48076 ;
  assign y16406 = ~n48077 ;
  assign y16407 = ~n48079 ;
  assign y16408 = ~1'b0 ;
  assign y16409 = ~1'b0 ;
  assign y16410 = ~n48080 ;
  assign y16411 = n510 ;
  assign y16412 = n48081 ;
  assign y16413 = ~n48090 ;
  assign y16414 = n48092 ;
  assign y16415 = ~1'b0 ;
  assign y16416 = ~1'b0 ;
  assign y16417 = ~1'b0 ;
  assign y16418 = ~n48099 ;
  assign y16419 = n48102 ;
  assign y16420 = ~n48104 ;
  assign y16421 = n48106 ;
  assign y16422 = ~1'b0 ;
  assign y16423 = n48113 ;
  assign y16424 = ~n48116 ;
  assign y16425 = n48119 ;
  assign y16426 = ~n48121 ;
  assign y16427 = ~n48122 ;
  assign y16428 = ~n48123 ;
  assign y16429 = ~n48124 ;
  assign y16430 = ~n48127 ;
  assign y16431 = ~1'b0 ;
  assign y16432 = ~1'b0 ;
  assign y16433 = ~n48129 ;
  assign y16434 = ~n48135 ;
  assign y16435 = n48137 ;
  assign y16436 = n48140 ;
  assign y16437 = ~n48141 ;
  assign y16438 = n48146 ;
  assign y16439 = ~n48150 ;
  assign y16440 = ~n48153 ;
  assign y16441 = ~n48154 ;
  assign y16442 = ~n48155 ;
  assign y16443 = ~n48156 ;
  assign y16444 = ~n48158 ;
  assign y16445 = ~n48159 ;
  assign y16446 = ~1'b0 ;
  assign y16447 = ~n48162 ;
  assign y16448 = n48163 ;
  assign y16449 = ~n48164 ;
  assign y16450 = ~n48165 ;
  assign y16451 = n48168 ;
  assign y16452 = ~n48170 ;
  assign y16453 = ~n48171 ;
  assign y16454 = ~n48177 ;
  assign y16455 = ~n48178 ;
  assign y16456 = n48179 ;
  assign y16457 = n48181 ;
  assign y16458 = ~n48182 ;
  assign y16459 = ~n48187 ;
  assign y16460 = n48189 ;
  assign y16461 = ~n48190 ;
  assign y16462 = n48191 ;
  assign y16463 = n48192 ;
  assign y16464 = n48194 ;
  assign y16465 = ~1'b0 ;
  assign y16466 = ~n48195 ;
  assign y16467 = ~1'b0 ;
  assign y16468 = ~n48197 ;
  assign y16469 = n48198 ;
  assign y16470 = n48199 ;
  assign y16471 = ~n48201 ;
  assign y16472 = n48149 ;
  assign y16473 = n48203 ;
  assign y16474 = ~n48205 ;
  assign y16475 = n48209 ;
  assign y16476 = n48210 ;
  assign y16477 = ~n48217 ;
  assign y16478 = ~1'b0 ;
  assign y16479 = n48224 ;
  assign y16480 = n48225 ;
  assign y16481 = n48227 ;
  assign y16482 = n48229 ;
  assign y16483 = ~n48232 ;
  assign y16484 = n48234 ;
  assign y16485 = ~1'b0 ;
  assign y16486 = ~n48241 ;
  assign y16487 = n48246 ;
  assign y16488 = ~n48252 ;
  assign y16489 = ~n48254 ;
  assign y16490 = ~n48256 ;
  assign y16491 = n48257 ;
  assign y16492 = ~n47701 ;
  assign y16493 = n48258 ;
  assign y16494 = ~n48259 ;
  assign y16495 = ~n48263 ;
  assign y16496 = ~1'b0 ;
  assign y16497 = ~1'b0 ;
  assign y16498 = ~n48276 ;
  assign y16499 = ~n48283 ;
  assign y16500 = ~n48293 ;
  assign y16501 = n48295 ;
  assign y16502 = ~n48297 ;
  assign y16503 = n48300 ;
  assign y16504 = n48310 ;
  assign y16505 = n48312 ;
  assign y16506 = ~n48314 ;
  assign y16507 = ~n48317 ;
  assign y16508 = ~1'b0 ;
  assign y16509 = ~n48318 ;
  assign y16510 = ~n48319 ;
  assign y16511 = n48320 ;
  assign y16512 = ~n48321 ;
  assign y16513 = n48324 ;
  assign y16514 = n48325 ;
  assign y16515 = ~n48330 ;
  assign y16516 = ~n48331 ;
  assign y16517 = ~1'b0 ;
  assign y16518 = n48333 ;
  assign y16519 = ~n48339 ;
  assign y16520 = ~n48340 ;
  assign y16521 = ~1'b0 ;
  assign y16522 = n48341 ;
  assign y16523 = ~n48342 ;
  assign y16524 = n48343 ;
  assign y16525 = ~n48345 ;
  assign y16526 = ~n48348 ;
  assign y16527 = ~1'b0 ;
  assign y16528 = n48350 ;
  assign y16529 = n48351 ;
  assign y16530 = ~n48352 ;
  assign y16531 = n48353 ;
  assign y16532 = n48354 ;
  assign y16533 = n48355 ;
  assign y16534 = ~1'b0 ;
  assign y16535 = ~1'b0 ;
  assign y16536 = ~n48356 ;
  assign y16537 = ~n48360 ;
  assign y16538 = ~n48363 ;
  assign y16539 = ~n48366 ;
  assign y16540 = n48367 ;
  assign y16541 = ~n48368 ;
  assign y16542 = n48373 ;
  assign y16543 = n48376 ;
  assign y16544 = n48378 ;
  assign y16545 = ~1'b0 ;
  assign y16546 = n48379 ;
  assign y16547 = n48381 ;
  assign y16548 = n48382 ;
  assign y16549 = n48383 ;
  assign y16550 = n48386 ;
  assign y16551 = ~1'b0 ;
  assign y16552 = ~n48392 ;
  assign y16553 = ~1'b0 ;
  assign y16554 = ~n48393 ;
  assign y16555 = n48395 ;
  assign y16556 = ~n48396 ;
  assign y16557 = n48397 ;
  assign y16558 = n48398 ;
  assign y16559 = n48399 ;
  assign y16560 = ~n48400 ;
  assign y16561 = ~n48404 ;
  assign y16562 = ~n48406 ;
  assign y16563 = ~n48408 ;
  assign y16564 = ~n48411 ;
  assign y16565 = n48412 ;
  assign y16566 = ~n48414 ;
  assign y16567 = ~n48415 ;
  assign y16568 = n48417 ;
  assign y16569 = ~n48423 ;
  assign y16570 = ~1'b0 ;
  assign y16571 = n48428 ;
  assign y16572 = n48430 ;
  assign y16573 = n48434 ;
  assign y16574 = n48436 ;
  assign y16575 = ~n48437 ;
  assign y16576 = n48443 ;
  assign y16577 = n48444 ;
  assign y16578 = ~1'b0 ;
  assign y16579 = n48449 ;
  assign y16580 = ~1'b0 ;
  assign y16581 = ~n48454 ;
  assign y16582 = n48456 ;
  assign y16583 = ~n48458 ;
  assign y16584 = ~n48459 ;
  assign y16585 = ~n48462 ;
  assign y16586 = n48465 ;
  assign y16587 = n48466 ;
  assign y16588 = ~n48468 ;
  assign y16589 = n48470 ;
  assign y16590 = ~n48473 ;
  assign y16591 = ~1'b0 ;
  assign y16592 = ~1'b0 ;
  assign y16593 = 1'b0 ;
  assign y16594 = n48474 ;
  assign y16595 = n48477 ;
  assign y16596 = n48478 ;
  assign y16597 = ~n16220 ;
  assign y16598 = ~n48479 ;
  assign y16599 = n48480 ;
  assign y16600 = ~n48481 ;
  assign y16601 = ~1'b0 ;
  assign y16602 = ~1'b0 ;
  assign y16603 = n48482 ;
  assign y16604 = ~n21399 ;
  assign y16605 = n48483 ;
  assign y16606 = ~n48484 ;
  assign y16607 = ~n48485 ;
  assign y16608 = ~n48486 ;
  assign y16609 = ~1'b0 ;
  assign y16610 = ~n48488 ;
  assign y16611 = n48491 ;
  assign y16612 = ~n48495 ;
  assign y16613 = ~1'b0 ;
  assign y16614 = n48497 ;
  assign y16615 = n48500 ;
  assign y16616 = ~n48501 ;
  assign y16617 = n48503 ;
  assign y16618 = n48507 ;
  assign y16619 = n48508 ;
  assign y16620 = ~1'b0 ;
  assign y16621 = ~1'b0 ;
  assign y16622 = ~1'b0 ;
  assign y16623 = ~n48513 ;
  assign y16624 = ~n48518 ;
  assign y16625 = ~n48519 ;
  assign y16626 = ~n31866 ;
  assign y16627 = ~n48524 ;
  assign y16628 = n48526 ;
  assign y16629 = n48527 ;
  assign y16630 = ~1'b0 ;
  assign y16631 = ~n48532 ;
  assign y16632 = n48533 ;
  assign y16633 = n48534 ;
  assign y16634 = ~n48538 ;
  assign y16635 = n48539 ;
  assign y16636 = ~n48540 ;
  assign y16637 = ~n48541 ;
  assign y16638 = ~1'b0 ;
  assign y16639 = ~n48543 ;
  assign y16640 = ~n48545 ;
  assign y16641 = n48547 ;
  assign y16642 = n48549 ;
  assign y16643 = n48551 ;
  assign y16644 = ~n48553 ;
  assign y16645 = ~n48557 ;
  assign y16646 = n48558 ;
  assign y16647 = ~n48559 ;
  assign y16648 = n48561 ;
  assign y16649 = 1'b0 ;
  assign y16650 = ~n48565 ;
  assign y16651 = n48569 ;
  assign y16652 = n48574 ;
  assign y16653 = ~n48576 ;
  assign y16654 = ~n48577 ;
  assign y16655 = ~n48579 ;
  assign y16656 = ~n48582 ;
  assign y16657 = ~n48584 ;
  assign y16658 = ~n48587 ;
  assign y16659 = n48588 ;
  assign y16660 = ~1'b0 ;
  assign y16661 = n48589 ;
  assign y16662 = ~1'b0 ;
  assign y16663 = ~1'b0 ;
  assign y16664 = ~1'b0 ;
  assign y16665 = ~n48590 ;
  assign y16666 = ~n48594 ;
  assign y16667 = n48595 ;
  assign y16668 = n48596 ;
  assign y16669 = n48601 ;
  assign y16670 = ~n48603 ;
  assign y16671 = n48608 ;
  assign y16672 = n48610 ;
  assign y16673 = ~n48612 ;
  assign y16674 = ~n48613 ;
  assign y16675 = ~n48614 ;
  assign y16676 = ~n48615 ;
  assign y16677 = n46165 ;
  assign y16678 = n48619 ;
  assign y16679 = ~n48624 ;
  assign y16680 = n48630 ;
  assign y16681 = n48632 ;
  assign y16682 = n48636 ;
  assign y16683 = n48639 ;
  assign y16684 = n48640 ;
  assign y16685 = ~n48641 ;
  assign y16686 = ~n48642 ;
  assign y16687 = n48644 ;
  assign y16688 = ~n48645 ;
  assign y16689 = n48648 ;
  assign y16690 = ~1'b0 ;
  assign y16691 = ~1'b0 ;
  assign y16692 = ~1'b0 ;
  assign y16693 = ~n48649 ;
  assign y16694 = n48657 ;
  assign y16695 = ~n48658 ;
  assign y16696 = ~n48660 ;
  assign y16697 = ~n48661 ;
  assign y16698 = ~n48662 ;
  assign y16699 = n48665 ;
  assign y16700 = ~1'b0 ;
  assign y16701 = n48666 ;
  assign y16702 = ~1'b0 ;
  assign y16703 = ~n48673 ;
  assign y16704 = n48674 ;
  assign y16705 = ~n48677 ;
  assign y16706 = n48679 ;
  assign y16707 = ~n48683 ;
  assign y16708 = n48686 ;
  assign y16709 = n48687 ;
  assign y16710 = n48689 ;
  assign y16711 = ~1'b0 ;
  assign y16712 = n48692 ;
  assign y16713 = ~n48694 ;
  assign y16714 = ~1'b0 ;
  assign y16715 = n48695 ;
  assign y16716 = n48697 ;
  assign y16717 = ~n48698 ;
  assign y16718 = ~n48701 ;
  assign y16719 = n48704 ;
  assign y16720 = ~n48706 ;
  assign y16721 = ~1'b0 ;
  assign y16722 = n48708 ;
  assign y16723 = ~1'b0 ;
  assign y16724 = ~1'b0 ;
  assign y16725 = n48713 ;
  assign y16726 = n48714 ;
  assign y16727 = ~n48715 ;
  assign y16728 = n48719 ;
  assign y16729 = ~n48721 ;
  assign y16730 = ~n48726 ;
  assign y16731 = n48729 ;
  assign y16732 = n48731 ;
  assign y16733 = n48735 ;
  assign y16734 = n48739 ;
  assign y16735 = n48748 ;
  assign y16736 = n48749 ;
  assign y16737 = ~n48755 ;
  assign y16738 = n48759 ;
  assign y16739 = n48761 ;
  assign y16740 = ~n48763 ;
  assign y16741 = ~1'b0 ;
  assign y16742 = ~1'b0 ;
  assign y16743 = n48764 ;
  assign y16744 = ~n48765 ;
  assign y16745 = n48767 ;
  assign y16746 = ~n48772 ;
  assign y16747 = ~n48778 ;
  assign y16748 = ~n48781 ;
  assign y16749 = n48783 ;
  assign y16750 = ~n48785 ;
  assign y16751 = ~n48788 ;
  assign y16752 = ~1'b0 ;
  assign y16753 = ~n48789 ;
  assign y16754 = ~n48790 ;
  assign y16755 = ~n48792 ;
  assign y16756 = ~n48797 ;
  assign y16757 = ~n48798 ;
  assign y16758 = n48799 ;
  assign y16759 = ~1'b0 ;
  assign y16760 = n48800 ;
  assign y16761 = ~n48804 ;
  assign y16762 = ~n48806 ;
  assign y16763 = n48807 ;
  assign y16764 = ~n48808 ;
  assign y16765 = ~n48811 ;
  assign y16766 = n48812 ;
  assign y16767 = n11717 ;
  assign y16768 = ~n48813 ;
  assign y16769 = ~n48814 ;
  assign y16770 = ~1'b0 ;
  assign y16771 = n48817 ;
  assign y16772 = ~1'b0 ;
  assign y16773 = ~n48819 ;
  assign y16774 = ~n48821 ;
  assign y16775 = n48823 ;
  assign y16776 = n48828 ;
  assign y16777 = n48831 ;
  assign y16778 = ~n48832 ;
  assign y16779 = ~n48838 ;
  assign y16780 = ~n7335 ;
  assign y16781 = ~1'b0 ;
  assign y16782 = n48840 ;
  assign y16783 = ~n48842 ;
  assign y16784 = ~n48844 ;
  assign y16785 = n48846 ;
  assign y16786 = ~n48848 ;
  assign y16787 = ~n48851 ;
  assign y16788 = ~n48852 ;
  assign y16789 = ~1'b0 ;
  assign y16790 = ~1'b0 ;
  assign y16791 = n48854 ;
  assign y16792 = ~1'b0 ;
  assign y16793 = ~1'b0 ;
  assign y16794 = n48859 ;
  assign y16795 = ~n48861 ;
  assign y16796 = ~n48862 ;
  assign y16797 = ~n48870 ;
  assign y16798 = ~n48871 ;
  assign y16799 = n48876 ;
  assign y16800 = ~1'b0 ;
  assign y16801 = ~n48878 ;
  assign y16802 = ~1'b0 ;
  assign y16803 = n48883 ;
  assign y16804 = ~n48884 ;
  assign y16805 = n48885 ;
  assign y16806 = n48888 ;
  assign y16807 = ~n48889 ;
  assign y16808 = ~n48892 ;
  assign y16809 = n48900 ;
  assign y16810 = n48905 ;
  assign y16811 = ~n48909 ;
  assign y16812 = ~1'b0 ;
  assign y16813 = ~n48911 ;
  assign y16814 = ~n48913 ;
  assign y16815 = n48918 ;
  assign y16816 = ~n48919 ;
  assign y16817 = ~n48920 ;
  assign y16818 = n48922 ;
  assign y16819 = ~n48923 ;
  assign y16820 = ~1'b0 ;
  assign y16821 = n48926 ;
  assign y16822 = n48929 ;
  assign y16823 = ~n48931 ;
  assign y16824 = n48932 ;
  assign y16825 = ~n48933 ;
  assign y16826 = ~n48935 ;
  assign y16827 = n48936 ;
  assign y16828 = n48938 ;
  assign y16829 = n48939 ;
  assign y16830 = ~n48942 ;
  assign y16831 = ~n48944 ;
  assign y16832 = ~n48948 ;
  assign y16833 = ~n48952 ;
  assign y16834 = n48955 ;
  assign y16835 = n48960 ;
  assign y16836 = ~n48961 ;
  assign y16837 = ~n48962 ;
  assign y16838 = ~n48965 ;
  assign y16839 = ~n48966 ;
  assign y16840 = ~n48967 ;
  assign y16841 = ~n48971 ;
  assign y16842 = ~n48973 ;
  assign y16843 = ~n48976 ;
  assign y16844 = ~1'b0 ;
  assign y16845 = n48978 ;
  assign y16846 = n48980 ;
  assign y16847 = ~n48987 ;
  assign y16848 = n48988 ;
  assign y16849 = n48989 ;
  assign y16850 = ~n48995 ;
  assign y16851 = n48999 ;
  assign y16852 = ~n49001 ;
  assign y16853 = n49004 ;
  assign y16854 = ~n49008 ;
  assign y16855 = ~n49009 ;
  assign y16856 = ~n49012 ;
  assign y16857 = n49013 ;
  assign y16858 = ~n49014 ;
  assign y16859 = n49016 ;
  assign y16860 = ~n43344 ;
  assign y16861 = n49017 ;
  assign y16862 = ~1'b0 ;
  assign y16863 = n49018 ;
  assign y16864 = n49028 ;
  assign y16865 = ~1'b0 ;
  assign y16866 = ~n49030 ;
  assign y16867 = ~n49031 ;
  assign y16868 = ~n49035 ;
  assign y16869 = n49040 ;
  assign y16870 = ~n49041 ;
  assign y16871 = n49042 ;
  assign y16872 = ~1'b0 ;
  assign y16873 = ~n49046 ;
  assign y16874 = ~1'b0 ;
  assign y16875 = ~n49049 ;
  assign y16876 = n49051 ;
  assign y16877 = n49053 ;
  assign y16878 = n49058 ;
  assign y16879 = n49059 ;
  assign y16880 = n49060 ;
  assign y16881 = n49061 ;
  assign y16882 = ~n49062 ;
  assign y16883 = ~1'b0 ;
  assign y16884 = n49067 ;
  assign y16885 = ~1'b0 ;
  assign y16886 = ~n49068 ;
  assign y16887 = ~1'b0 ;
  assign y16888 = n49069 ;
  assign y16889 = n49070 ;
  assign y16890 = ~n49072 ;
  assign y16891 = n49076 ;
  assign y16892 = n49077 ;
  assign y16893 = n49078 ;
  assign y16894 = n49081 ;
  assign y16895 = ~n49088 ;
  assign y16896 = ~1'b0 ;
  assign y16897 = ~1'b0 ;
  assign y16898 = ~n49089 ;
  assign y16899 = n49090 ;
  assign y16900 = n49092 ;
  assign y16901 = ~n49096 ;
  assign y16902 = n49098 ;
  assign y16903 = ~n49100 ;
  assign y16904 = ~1'b0 ;
  assign y16905 = ~1'b0 ;
  assign y16906 = n49101 ;
  assign y16907 = n49103 ;
  assign y16908 = ~n49104 ;
  assign y16909 = ~n49107 ;
  assign y16910 = ~n49108 ;
  assign y16911 = n49109 ;
  assign y16912 = n49122 ;
  assign y16913 = ~n49123 ;
  assign y16914 = ~n49124 ;
  assign y16915 = ~n49125 ;
  assign y16916 = ~1'b0 ;
  assign y16917 = ~n49130 ;
  assign y16918 = ~1'b0 ;
  assign y16919 = ~n49131 ;
  assign y16920 = ~n49132 ;
  assign y16921 = n49135 ;
  assign y16922 = ~n49136 ;
  assign y16923 = ~n49137 ;
  assign y16924 = ~1'b0 ;
  assign y16925 = ~n49140 ;
  assign y16926 = n49143 ;
  assign y16927 = n49146 ;
  assign y16928 = ~n49147 ;
  assign y16929 = n49149 ;
  assign y16930 = ~n49150 ;
  assign y16931 = n49152 ;
  assign y16932 = n49155 ;
  assign y16933 = n49158 ;
  assign y16934 = ~n49164 ;
  assign y16935 = ~n49166 ;
  assign y16936 = ~1'b0 ;
  assign y16937 = n49167 ;
  assign y16938 = ~n49171 ;
  assign y16939 = n49172 ;
  assign y16940 = n49173 ;
  assign y16941 = n49174 ;
  assign y16942 = n49175 ;
  assign y16943 = ~n49176 ;
  assign y16944 = n49178 ;
  assign y16945 = ~1'b0 ;
  assign y16946 = n49182 ;
  assign y16947 = ~n49184 ;
  assign y16948 = ~n49186 ;
  assign y16949 = ~n49187 ;
  assign y16950 = ~n49190 ;
  assign y16951 = n49192 ;
  assign y16952 = ~n49193 ;
  assign y16953 = n49197 ;
  assign y16954 = n49198 ;
  assign y16955 = ~1'b0 ;
  assign y16956 = ~n49200 ;
  assign y16957 = n49202 ;
  assign y16958 = ~1'b0 ;
  assign y16959 = ~n49205 ;
  assign y16960 = ~n49208 ;
  assign y16961 = n49210 ;
  assign y16962 = n49213 ;
  assign y16963 = ~n49215 ;
  assign y16964 = n49216 ;
  assign y16965 = ~n49217 ;
  assign y16966 = ~n49219 ;
  assign y16967 = ~1'b0 ;
  assign y16968 = ~n49227 ;
  assign y16969 = ~n49228 ;
  assign y16970 = n49230 ;
  assign y16971 = n49231 ;
  assign y16972 = ~n49238 ;
  assign y16973 = n49239 ;
  assign y16974 = ~n49244 ;
  assign y16975 = ~1'b0 ;
  assign y16976 = ~n49246 ;
  assign y16977 = ~n49247 ;
  assign y16978 = n49250 ;
  assign y16979 = n49253 ;
  assign y16980 = ~n49254 ;
  assign y16981 = ~n49263 ;
  assign y16982 = ~1'b0 ;
  assign y16983 = ~1'b0 ;
  assign y16984 = ~n49265 ;
  assign y16985 = ~1'b0 ;
  assign y16986 = ~n49266 ;
  assign y16987 = ~n49267 ;
  assign y16988 = ~n49271 ;
  assign y16989 = n49274 ;
  assign y16990 = ~n49275 ;
  assign y16991 = ~n1786 ;
  assign y16992 = n49277 ;
  assign y16993 = ~n49279 ;
  assign y16994 = n49280 ;
  assign y16995 = n49282 ;
  assign y16996 = ~n49283 ;
  assign y16997 = ~n49284 ;
  assign y16998 = n49286 ;
  assign y16999 = n49295 ;
  assign y17000 = n49298 ;
  assign y17001 = ~1'b0 ;
  assign y17002 = ~n49300 ;
  assign y17003 = ~n49304 ;
  assign y17004 = ~1'b0 ;
  assign y17005 = ~n49306 ;
  assign y17006 = ~n36088 ;
  assign y17007 = n49307 ;
  assign y17008 = ~n49308 ;
  assign y17009 = n49309 ;
  assign y17010 = n49311 ;
  assign y17011 = n49315 ;
  assign y17012 = ~n49317 ;
  assign y17013 = ~n49319 ;
  assign y17014 = ~1'b0 ;
  assign y17015 = ~n49324 ;
  assign y17016 = ~n49326 ;
  assign y17017 = n49334 ;
  assign y17018 = ~n49335 ;
  assign y17019 = ~n49339 ;
  assign y17020 = ~n49341 ;
  assign y17021 = n49344 ;
  assign y17022 = ~1'b0 ;
  assign y17023 = ~1'b0 ;
  assign y17024 = ~n16405 ;
  assign y17025 = ~n49345 ;
  assign y17026 = ~n49346 ;
  assign y17027 = n49347 ;
  assign y17028 = ~n49349 ;
  assign y17029 = ~n49350 ;
  assign y17030 = ~n49354 ;
  assign y17031 = ~1'b0 ;
  assign y17032 = ~1'b0 ;
  assign y17033 = ~n49355 ;
  assign y17034 = n49356 ;
  assign y17035 = ~n49362 ;
  assign y17036 = n49363 ;
  assign y17037 = ~n49364 ;
  assign y17038 = ~n49366 ;
  assign y17039 = n49370 ;
  assign y17040 = ~1'b0 ;
  assign y17041 = ~n49372 ;
  assign y17042 = ~n49375 ;
  assign y17043 = n49384 ;
  assign y17044 = ~n49385 ;
  assign y17045 = ~n49387 ;
  assign y17046 = n49394 ;
  assign y17047 = ~n49395 ;
  assign y17048 = n49396 ;
  assign y17049 = ~1'b0 ;
  assign y17050 = n49398 ;
  assign y17051 = ~1'b0 ;
  assign y17052 = ~1'b0 ;
  assign y17053 = ~n49400 ;
  assign y17054 = n49402 ;
  assign y17055 = ~n49408 ;
  assign y17056 = n49410 ;
  assign y17057 = ~n49413 ;
  assign y17058 = n49414 ;
  assign y17059 = ~n49415 ;
  assign y17060 = n49419 ;
  assign y17061 = n49422 ;
  assign y17062 = n49425 ;
  assign y17063 = ~n49427 ;
  assign y17064 = ~n49428 ;
  assign y17065 = n49430 ;
  assign y17066 = ~n49431 ;
  assign y17067 = ~n49434 ;
  assign y17068 = ~n49436 ;
  assign y17069 = ~n49437 ;
  assign y17070 = ~n49438 ;
  assign y17071 = n49439 ;
  assign y17072 = ~n49443 ;
  assign y17073 = ~n49444 ;
  assign y17074 = ~n49445 ;
  assign y17075 = ~n49448 ;
  assign y17076 = n49449 ;
  assign y17077 = ~n49450 ;
  assign y17078 = ~n49452 ;
  assign y17079 = ~n49457 ;
  assign y17080 = n2144 ;
  assign y17081 = n49463 ;
  assign y17082 = n49465 ;
  assign y17083 = n49467 ;
  assign y17084 = n49469 ;
  assign y17085 = ~n49470 ;
  assign y17086 = ~n49471 ;
  assign y17087 = n49472 ;
  assign y17088 = n49474 ;
  assign y17089 = n30197 ;
  assign y17090 = ~1'b0 ;
  assign y17091 = n49479 ;
  assign y17092 = ~n49482 ;
  assign y17093 = n49483 ;
  assign y17094 = n49485 ;
  assign y17095 = n49487 ;
  assign y17096 = ~n49489 ;
  assign y17097 = ~n49491 ;
  assign y17098 = ~n49494 ;
  assign y17099 = ~n49505 ;
  assign y17100 = n49506 ;
  assign y17101 = n49507 ;
  assign y17102 = ~n49513 ;
  assign y17103 = ~1'b0 ;
  assign y17104 = n49515 ;
  assign y17105 = ~1'b0 ;
  assign y17106 = n49517 ;
  assign y17107 = ~n49519 ;
  assign y17108 = ~n49520 ;
  assign y17109 = ~n49521 ;
  assign y17110 = n49525 ;
  assign y17111 = n49528 ;
  assign y17112 = ~1'b0 ;
  assign y17113 = ~1'b0 ;
  assign y17114 = ~1'b0 ;
  assign y17115 = ~n49529 ;
  assign y17116 = n49531 ;
  assign y17117 = n49534 ;
  assign y17118 = ~n49535 ;
  assign y17119 = n49537 ;
  assign y17120 = n49540 ;
  assign y17121 = ~n49542 ;
  assign y17122 = ~n49545 ;
  assign y17123 = n49546 ;
  assign y17124 = n49548 ;
  assign y17125 = n49549 ;
  assign y17126 = n49553 ;
  assign y17127 = ~n49554 ;
  assign y17128 = n49555 ;
  assign y17129 = ~n49556 ;
  assign y17130 = ~n49557 ;
  assign y17131 = ~n49560 ;
  assign y17132 = n49562 ;
  assign y17133 = ~1'b0 ;
  assign y17134 = ~n49565 ;
  assign y17135 = ~1'b0 ;
  assign y17136 = ~n49568 ;
  assign y17137 = n49571 ;
  assign y17138 = ~n49572 ;
  assign y17139 = ~n49575 ;
  assign y17140 = n49578 ;
  assign y17141 = ~1'b0 ;
  assign y17142 = n49582 ;
  assign y17143 = n49584 ;
  assign y17144 = n49587 ;
  assign y17145 = ~n49590 ;
  assign y17146 = n49594 ;
  assign y17147 = ~n49597 ;
  assign y17148 = ~n49599 ;
  assign y17149 = ~1'b0 ;
  assign y17150 = ~n49601 ;
  assign y17151 = ~1'b0 ;
  assign y17152 = ~1'b0 ;
  assign y17153 = ~n49612 ;
  assign y17154 = n49613 ;
  assign y17155 = ~n49616 ;
  assign y17156 = ~n49617 ;
  assign y17157 = n49623 ;
  assign y17158 = n49626 ;
  assign y17159 = n49628 ;
  assign y17160 = n49630 ;
  assign y17161 = ~n49632 ;
  assign y17162 = ~n49633 ;
  assign y17163 = ~n49636 ;
  assign y17164 = n49638 ;
  assign y17165 = n49639 ;
  assign y17166 = n49640 ;
  assign y17167 = n49644 ;
  assign y17168 = ~1'b0 ;
  assign y17169 = ~1'b0 ;
  assign y17170 = ~1'b0 ;
  assign y17171 = n49648 ;
  assign y17172 = n49649 ;
  assign y17173 = n49650 ;
  assign y17174 = ~n49653 ;
  assign y17175 = n49654 ;
  assign y17176 = n49659 ;
  assign y17177 = n49660 ;
  assign y17178 = n49663 ;
  assign y17179 = ~n49665 ;
  assign y17180 = ~n49668 ;
  assign y17181 = ~n49673 ;
  assign y17182 = n49676 ;
  assign y17183 = ~n2095 ;
  assign y17184 = ~n49680 ;
  assign y17185 = ~n49681 ;
  assign y17186 = n49682 ;
  assign y17187 = ~n49683 ;
  assign y17188 = ~1'b0 ;
  assign y17189 = n49684 ;
  assign y17190 = ~n49685 ;
  assign y17191 = n49687 ;
  assign y17192 = ~n49688 ;
  assign y17193 = ~n49692 ;
  assign y17194 = ~n1309 ;
  assign y17195 = ~n49693 ;
  assign y17196 = n49697 ;
  assign y17197 = n49700 ;
  assign y17198 = ~n49703 ;
  assign y17199 = ~n49707 ;
  assign y17200 = ~1'b0 ;
  assign y17201 = ~n49708 ;
  assign y17202 = n49709 ;
  assign y17203 = n49711 ;
  assign y17204 = ~n49712 ;
  assign y17205 = ~n49718 ;
  assign y17206 = n49722 ;
  assign y17207 = n49723 ;
  assign y17208 = ~n49726 ;
  assign y17209 = ~n49728 ;
  assign y17210 = ~n49729 ;
  assign y17211 = ~n49732 ;
  assign y17212 = n49733 ;
  assign y17213 = ~n49740 ;
  assign y17214 = ~n49742 ;
  assign y17215 = ~1'b0 ;
  assign y17216 = n49746 ;
  assign y17217 = ~1'b0 ;
  assign y17218 = ~n49747 ;
  assign y17219 = ~n49748 ;
  assign y17220 = ~n19268 ;
  assign y17221 = n49749 ;
  assign y17222 = n49750 ;
  assign y17223 = ~n49751 ;
  assign y17224 = ~1'b0 ;
  assign y17225 = n49753 ;
  assign y17226 = ~n49754 ;
  assign y17227 = ~n49756 ;
  assign y17228 = n49761 ;
  assign y17229 = ~n49763 ;
  assign y17230 = n49766 ;
  assign y17231 = n49769 ;
  assign y17232 = n49770 ;
  assign y17233 = n49771 ;
  assign y17234 = ~n49773 ;
  assign y17235 = ~1'b0 ;
  assign y17236 = ~n49777 ;
  assign y17237 = ~n49783 ;
  assign y17238 = ~n49787 ;
  assign y17239 = ~n49788 ;
  assign y17240 = ~n49793 ;
  assign y17241 = n49794 ;
  assign y17242 = ~n49795 ;
  assign y17243 = ~n49801 ;
  assign y17244 = n49803 ;
  assign y17245 = ~1'b0 ;
  assign y17246 = n49804 ;
  assign y17247 = n49807 ;
  assign y17248 = ~n49809 ;
  assign y17249 = n49816 ;
  assign y17250 = n49817 ;
  assign y17251 = ~n49821 ;
  assign y17252 = ~n49823 ;
  assign y17253 = n49826 ;
  assign y17254 = ~n49828 ;
  assign y17255 = ~n49830 ;
  assign y17256 = n49831 ;
  assign y17257 = ~n49835 ;
  assign y17258 = ~1'b0 ;
  assign y17259 = ~n49836 ;
  assign y17260 = ~n49839 ;
  assign y17261 = n49842 ;
  assign y17262 = ~n49846 ;
  assign y17263 = ~n49848 ;
  assign y17264 = n49850 ;
  assign y17265 = ~n49853 ;
  assign y17266 = ~n49854 ;
  assign y17267 = ~1'b0 ;
  assign y17268 = ~1'b0 ;
  assign y17269 = n49856 ;
  assign y17270 = n49857 ;
  assign y17271 = ~n49858 ;
  assign y17272 = n49859 ;
  assign y17273 = n49860 ;
  assign y17274 = ~n49862 ;
  assign y17275 = ~1'b0 ;
  assign y17276 = ~1'b0 ;
  assign y17277 = n49864 ;
  assign y17278 = n49868 ;
  assign y17279 = n26226 ;
  assign y17280 = n49871 ;
  assign y17281 = n49872 ;
  assign y17282 = n49875 ;
  assign y17283 = ~n49882 ;
  assign y17284 = ~n49885 ;
  assign y17285 = n49887 ;
  assign y17286 = ~n49892 ;
  assign y17287 = n49893 ;
  assign y17288 = n49898 ;
  assign y17289 = ~n49899 ;
  assign y17290 = ~n49906 ;
  assign y17291 = ~n49907 ;
  assign y17292 = ~n49909 ;
  assign y17293 = ~1'b0 ;
  assign y17294 = n26469 ;
  assign y17295 = ~n49911 ;
  assign y17296 = n49915 ;
  assign y17297 = n49919 ;
  assign y17298 = ~n49921 ;
  assign y17299 = ~n49924 ;
  assign y17300 = n49936 ;
  assign y17301 = n49938 ;
  assign y17302 = ~n49939 ;
  assign y17303 = ~1'b0 ;
  assign y17304 = ~1'b0 ;
  assign y17305 = n49940 ;
  assign y17306 = n49943 ;
  assign y17307 = n49944 ;
  assign y17308 = ~n49947 ;
  assign y17309 = n49950 ;
  assign y17310 = n49951 ;
  assign y17311 = ~n49952 ;
  assign y17312 = n49955 ;
  assign y17313 = n49957 ;
  assign y17314 = n49960 ;
  assign y17315 = n49962 ;
  assign y17316 = ~1'b0 ;
  assign y17317 = n49971 ;
  assign y17318 = n49973 ;
  assign y17319 = ~n49977 ;
  assign y17320 = ~n49979 ;
  assign y17321 = n49985 ;
  assign y17322 = ~n49987 ;
  assign y17323 = ~n49988 ;
  assign y17324 = ~1'b0 ;
  assign y17325 = ~n49990 ;
  assign y17326 = ~1'b0 ;
  assign y17327 = ~n49994 ;
  assign y17328 = ~1'b0 ;
  assign y17329 = n49996 ;
  assign y17330 = n49999 ;
  assign y17331 = n50001 ;
  assign y17332 = ~n50004 ;
  assign y17333 = ~n50005 ;
  assign y17334 = n50008 ;
  assign y17335 = n50013 ;
  assign y17336 = n50014 ;
  assign y17337 = ~n50019 ;
  assign y17338 = n50023 ;
  assign y17339 = n50024 ;
  assign y17340 = n50025 ;
  assign y17341 = ~n50028 ;
  assign y17342 = n50029 ;
  assign y17343 = ~n50031 ;
  assign y17344 = ~n50033 ;
  assign y17345 = ~n50035 ;
  assign y17346 = ~n50037 ;
  assign y17347 = ~n50040 ;
  assign y17348 = ~n50041 ;
  assign y17349 = n50044 ;
  assign y17350 = ~n50045 ;
  assign y17351 = ~n50046 ;
  assign y17352 = n50047 ;
  assign y17353 = n50048 ;
  assign y17354 = n50050 ;
  assign y17355 = ~1'b0 ;
  assign y17356 = n50051 ;
  assign y17357 = ~1'b0 ;
  assign y17358 = ~1'b0 ;
  assign y17359 = n50052 ;
  assign y17360 = ~n50054 ;
  assign y17361 = ~n50055 ;
  assign y17362 = ~n50056 ;
  assign y17363 = ~n50059 ;
  assign y17364 = ~n50062 ;
  assign y17365 = ~n50065 ;
  assign y17366 = ~n50067 ;
  assign y17367 = ~1'b0 ;
  assign y17368 = ~n50069 ;
  assign y17369 = ~1'b0 ;
  assign y17370 = ~n50073 ;
  assign y17371 = n10713 ;
  assign y17372 = ~n50083 ;
  assign y17373 = n50089 ;
  assign y17374 = n50090 ;
  assign y17375 = n50092 ;
  assign y17376 = n50098 ;
  assign y17377 = ~1'b0 ;
  assign y17378 = n50101 ;
  assign y17379 = n50102 ;
  assign y17380 = ~1'b0 ;
  assign y17381 = n50106 ;
  assign y17382 = n50107 ;
  assign y17383 = ~n50112 ;
  assign y17384 = ~n50117 ;
  assign y17385 = n50119 ;
  assign y17386 = ~n50124 ;
  assign y17387 = ~1'b0 ;
  assign y17388 = ~1'b0 ;
  assign y17389 = ~n50126 ;
  assign y17390 = n50129 ;
  assign y17391 = ~n7337 ;
  assign y17392 = ~n50134 ;
  assign y17393 = ~n50140 ;
  assign y17394 = ~n50141 ;
  assign y17395 = ~n50142 ;
  assign y17396 = n50143 ;
  assign y17397 = n50147 ;
  assign y17398 = ~1'b0 ;
  assign y17399 = ~n50148 ;
  assign y17400 = ~n50149 ;
  assign y17401 = ~n50151 ;
  assign y17402 = n50155 ;
  assign y17403 = ~n50157 ;
  assign y17404 = n50158 ;
  assign y17405 = ~n50160 ;
  assign y17406 = ~n50162 ;
  assign y17407 = n50169 ;
  assign y17408 = n50170 ;
  assign y17409 = ~1'b0 ;
  assign y17410 = ~n50171 ;
  assign y17411 = n50173 ;
  assign y17412 = ~n50175 ;
  assign y17413 = n50178 ;
  assign y17414 = n50180 ;
  assign y17415 = n50182 ;
  assign y17416 = n50185 ;
  assign y17417 = n50186 ;
  assign y17418 = n50187 ;
  assign y17419 = n50190 ;
  assign y17420 = ~n50191 ;
  assign y17421 = ~1'b0 ;
  assign y17422 = ~n50193 ;
  assign y17423 = ~n50195 ;
  assign y17424 = n50197 ;
  assign y17425 = n50201 ;
  assign y17426 = ~n50205 ;
  assign y17427 = n50209 ;
  assign y17428 = n50215 ;
  assign y17429 = ~n50219 ;
  assign y17430 = ~n50221 ;
  assign y17431 = ~n50225 ;
  assign y17432 = ~n50226 ;
  assign y17433 = ~n50229 ;
  assign y17434 = ~n50233 ;
  assign y17435 = ~n50234 ;
  assign y17436 = ~n50235 ;
  assign y17437 = ~n50237 ;
  assign y17438 = n50239 ;
  assign y17439 = n50241 ;
  assign y17440 = ~1'b0 ;
  assign y17441 = ~1'b0 ;
  assign y17442 = ~n50245 ;
  assign y17443 = ~n50247 ;
  assign y17444 = ~n50249 ;
  assign y17445 = n50250 ;
  assign y17446 = n50256 ;
  assign y17447 = ~n50258 ;
  assign y17448 = ~n50259 ;
  assign y17449 = ~n50263 ;
  assign y17450 = ~n50271 ;
  assign y17451 = ~n50272 ;
  assign y17452 = ~n50275 ;
  assign y17453 = ~n50281 ;
  assign y17454 = ~n50289 ;
  assign y17455 = n50292 ;
  assign y17456 = ~n50294 ;
  assign y17457 = ~n50295 ;
  assign y17458 = ~n50296 ;
  assign y17459 = ~1'b0 ;
  assign y17460 = n50297 ;
  assign y17461 = ~n50298 ;
  assign y17462 = n50300 ;
  assign y17463 = n50303 ;
  assign y17464 = ~n50304 ;
  assign y17465 = n50307 ;
  assign y17466 = n50309 ;
  assign y17467 = n50310 ;
  assign y17468 = n50312 ;
  assign y17469 = ~n50313 ;
  assign y17470 = n50315 ;
  assign y17471 = n50319 ;
  assign y17472 = ~1'b0 ;
  assign y17473 = ~n50322 ;
  assign y17474 = ~1'b0 ;
  assign y17475 = ~n50323 ;
  assign y17476 = n50324 ;
  assign y17477 = ~n50326 ;
  assign y17478 = ~n50328 ;
  assign y17479 = n50334 ;
  assign y17480 = n50338 ;
  assign y17481 = ~1'b0 ;
  assign y17482 = ~1'b0 ;
  assign y17483 = n50340 ;
  assign y17484 = n50342 ;
  assign y17485 = ~n50344 ;
  assign y17486 = n15798 ;
  assign y17487 = ~n50348 ;
  assign y17488 = ~n50349 ;
  assign y17489 = n49473 ;
  assign y17490 = ~n50350 ;
  assign y17491 = n50354 ;
  assign y17492 = ~n50357 ;
  assign y17493 = ~n50360 ;
  assign y17494 = ~n50361 ;
  assign y17495 = ~n50363 ;
  assign y17496 = n50364 ;
  assign y17497 = n50370 ;
  assign y17498 = n50371 ;
  assign y17499 = ~n50372 ;
  assign y17500 = n50376 ;
  assign y17501 = ~n50382 ;
  assign y17502 = n50386 ;
  assign y17503 = ~n19209 ;
  assign y17504 = ~n50388 ;
  assign y17505 = ~1'b0 ;
  assign y17506 = n50395 ;
  assign y17507 = n50401 ;
  assign y17508 = ~n50402 ;
  assign y17509 = ~n50403 ;
  assign y17510 = n50405 ;
  assign y17511 = ~n50406 ;
  assign y17512 = ~n50407 ;
  assign y17513 = n50408 ;
  assign y17514 = ~1'b0 ;
  assign y17515 = n50411 ;
  assign y17516 = ~n50414 ;
  assign y17517 = ~1'b0 ;
  assign y17518 = ~n50415 ;
  assign y17519 = n50417 ;
  assign y17520 = n50421 ;
  assign y17521 = n50424 ;
  assign y17522 = n50431 ;
  assign y17523 = ~n50432 ;
  assign y17524 = ~n50434 ;
  assign y17525 = n50435 ;
  assign y17526 = ~1'b0 ;
  assign y17527 = ~n50437 ;
  assign y17528 = n50439 ;
  assign y17529 = ~n50442 ;
  assign y17530 = ~n50443 ;
  assign y17531 = n50447 ;
  assign y17532 = n50449 ;
  assign y17533 = ~n50455 ;
  assign y17534 = n50456 ;
  assign y17535 = n50458 ;
  assign y17536 = ~n50460 ;
  assign y17537 = ~1'b0 ;
  assign y17538 = ~n50464 ;
  assign y17539 = ~n50465 ;
  assign y17540 = n50467 ;
  assign y17541 = n50470 ;
  assign y17542 = ~n50471 ;
  assign y17543 = n50473 ;
  assign y17544 = ~n50477 ;
  assign y17545 = n50478 ;
  assign y17546 = n50479 ;
  assign y17547 = ~n50481 ;
  assign y17548 = ~n50487 ;
  assign y17549 = n50493 ;
  assign y17550 = n50495 ;
  assign y17551 = n50498 ;
  assign y17552 = n50500 ;
  assign y17553 = n21318 ;
  assign y17554 = ~n50502 ;
  assign y17555 = n50506 ;
  assign y17556 = ~n50514 ;
  assign y17557 = ~1'b0 ;
  assign y17558 = n50516 ;
  assign y17559 = ~n4760 ;
  assign y17560 = ~n50519 ;
  assign y17561 = ~n50520 ;
  assign y17562 = n50523 ;
  assign y17563 = ~n50527 ;
  assign y17564 = n50531 ;
  assign y17565 = n50534 ;
  assign y17566 = ~n50537 ;
  assign y17567 = n18400 ;
  assign y17568 = ~n50539 ;
  assign y17569 = n50543 ;
  assign y17570 = ~n50544 ;
  assign y17571 = n50545 ;
  assign y17572 = n50547 ;
  assign y17573 = ~n50549 ;
  assign y17574 = n50552 ;
  assign y17575 = ~n50553 ;
  assign y17576 = n50554 ;
  assign y17577 = ~n50556 ;
  assign y17578 = ~n50557 ;
  assign y17579 = ~n50559 ;
  assign y17580 = ~1'b0 ;
  assign y17581 = n50561 ;
  assign y17582 = ~n50562 ;
  assign y17583 = ~n50567 ;
  assign y17584 = n50568 ;
  assign y17585 = n50570 ;
  assign y17586 = n50571 ;
  assign y17587 = n50573 ;
  assign y17588 = n50575 ;
  assign y17589 = ~n50577 ;
  assign y17590 = ~n19868 ;
  assign y17591 = n50580 ;
  assign y17592 = ~n50584 ;
  assign y17593 = n50585 ;
  assign y17594 = n50592 ;
  assign y17595 = ~n50594 ;
  assign y17596 = n50595 ;
  assign y17597 = ~n50601 ;
  assign y17598 = ~n50607 ;
  assign y17599 = ~1'b0 ;
  assign y17600 = ~1'b0 ;
  assign y17601 = ~1'b0 ;
  assign y17602 = n50609 ;
  assign y17603 = ~n50611 ;
  assign y17604 = ~n50613 ;
  assign y17605 = ~n50615 ;
  assign y17606 = ~n50616 ;
  assign y17607 = ~1'b0 ;
  assign y17608 = ~1'b0 ;
  assign y17609 = n50618 ;
  assign y17610 = ~n50620 ;
  assign y17611 = ~n50622 ;
  assign y17612 = n50623 ;
  assign y17613 = n50625 ;
  assign y17614 = ~n50627 ;
  assign y17615 = n50628 ;
  assign y17616 = ~n50630 ;
  assign y17617 = n50633 ;
  assign y17618 = ~n50637 ;
  assign y17619 = ~n50643 ;
  assign y17620 = ~n50645 ;
  assign y17621 = n50646 ;
  assign y17622 = ~n50647 ;
  assign y17623 = ~n50649 ;
  assign y17624 = n50652 ;
  assign y17625 = ~n50653 ;
  assign y17626 = ~n50654 ;
  assign y17627 = ~n50658 ;
  assign y17628 = n50663 ;
  assign y17629 = n50666 ;
  assign y17630 = ~n50667 ;
  assign y17631 = n50676 ;
  assign y17632 = ~n48435 ;
  assign y17633 = ~n50678 ;
  assign y17634 = ~n50679 ;
  assign y17635 = ~1'b0 ;
  assign y17636 = ~1'b0 ;
  assign y17637 = ~n50681 ;
  assign y17638 = n50685 ;
  assign y17639 = ~1'b0 ;
  assign y17640 = ~n50687 ;
  assign y17641 = n50692 ;
  assign y17642 = ~n50696 ;
  assign y17643 = ~n50698 ;
  assign y17644 = ~n50700 ;
  assign y17645 = ~n50701 ;
  assign y17646 = n50703 ;
  assign y17647 = ~1'b0 ;
  assign y17648 = ~n50705 ;
  assign y17649 = n50707 ;
  assign y17650 = ~n50712 ;
  assign y17651 = ~n50721 ;
  assign y17652 = n50728 ;
  assign y17653 = n50730 ;
  assign y17654 = ~n50731 ;
  assign y17655 = n50734 ;
  assign y17656 = ~n50735 ;
  assign y17657 = ~n50741 ;
  assign y17658 = n50742 ;
  assign y17659 = ~n50745 ;
  assign y17660 = n50747 ;
  assign y17661 = n50748 ;
  assign y17662 = n50749 ;
  assign y17663 = n50751 ;
  assign y17664 = n50752 ;
  assign y17665 = ~1'b0 ;
  assign y17666 = n50753 ;
  assign y17667 = ~n50754 ;
  assign y17668 = n50757 ;
  assign y17669 = n50759 ;
  assign y17670 = n50760 ;
  assign y17671 = ~n50762 ;
  assign y17672 = ~n11432 ;
  assign y17673 = ~n50763 ;
  assign y17674 = ~n50764 ;
  assign y17675 = ~1'b0 ;
  assign y17676 = ~n50765 ;
  assign y17677 = ~n50767 ;
  assign y17678 = n50769 ;
  assign y17679 = ~n50774 ;
  assign y17680 = n50784 ;
  assign y17681 = n50786 ;
  assign y17682 = n50787 ;
  assign y17683 = n50789 ;
  assign y17684 = ~n50791 ;
  assign y17685 = ~n50793 ;
  assign y17686 = ~n50797 ;
  assign y17687 = ~n50800 ;
  assign y17688 = ~n50802 ;
  assign y17689 = n50803 ;
  assign y17690 = n50806 ;
  assign y17691 = n50808 ;
  assign y17692 = ~n50810 ;
  assign y17693 = ~n50815 ;
  assign y17694 = ~n50818 ;
  assign y17695 = ~n17755 ;
  assign y17696 = n50820 ;
  assign y17697 = ~1'b0 ;
  assign y17698 = ~1'b0 ;
  assign y17699 = n50826 ;
  assign y17700 = n50831 ;
  assign y17701 = ~n50832 ;
  assign y17702 = n50834 ;
  assign y17703 = n50837 ;
  assign y17704 = ~n50839 ;
  assign y17705 = n50844 ;
  assign y17706 = n50846 ;
  assign y17707 = ~1'b0 ;
  assign y17708 = ~n50848 ;
  assign y17709 = ~n50850 ;
  assign y17710 = n50851 ;
  assign y17711 = n50852 ;
  assign y17712 = ~n50856 ;
  assign y17713 = ~n50860 ;
  assign y17714 = n50866 ;
  assign y17715 = ~n50867 ;
  assign y17716 = ~n50872 ;
  assign y17717 = ~1'b0 ;
  assign y17718 = ~1'b0 ;
  assign y17719 = n50876 ;
  assign y17720 = ~n50879 ;
  assign y17721 = ~n50882 ;
  assign y17722 = n50883 ;
  assign y17723 = n50885 ;
  assign y17724 = n50886 ;
  assign y17725 = ~n50891 ;
  assign y17726 = n50894 ;
  assign y17727 = n50902 ;
  assign y17728 = ~n50904 ;
  assign y17729 = ~1'b0 ;
  assign y17730 = n50905 ;
  assign y17731 = ~n50906 ;
  assign y17732 = ~n50908 ;
  assign y17733 = ~n50909 ;
  assign y17734 = ~1'b0 ;
  assign y17735 = ~n50912 ;
  assign y17736 = n50915 ;
  assign y17737 = ~n50916 ;
  assign y17738 = ~n50920 ;
  assign y17739 = n50921 ;
  assign y17740 = n50922 ;
  assign y17741 = n50924 ;
  assign y17742 = ~n50926 ;
  assign y17743 = ~n50927 ;
  assign y17744 = n50930 ;
  assign y17745 = n50931 ;
  assign y17746 = ~n50933 ;
  assign y17747 = ~n50935 ;
  assign y17748 = n50939 ;
  assign y17749 = ~1'b0 ;
  assign y17750 = ~n50945 ;
  assign y17751 = ~1'b0 ;
  assign y17752 = n50952 ;
  assign y17753 = n50955 ;
  assign y17754 = ~n50959 ;
  assign y17755 = ~1'b0 ;
  assign y17756 = n50960 ;
  assign y17757 = n50966 ;
  assign y17758 = ~n50967 ;
  assign y17759 = ~1'b0 ;
  assign y17760 = ~1'b0 ;
  assign y17761 = ~1'b0 ;
  assign y17762 = ~1'b0 ;
  assign y17763 = ~n50970 ;
  assign y17764 = n50971 ;
  assign y17765 = n50973 ;
  assign y17766 = n50975 ;
  assign y17767 = ~n50976 ;
  assign y17768 = n50978 ;
  assign y17769 = n50979 ;
  assign y17770 = n50981 ;
  assign y17771 = n50983 ;
  assign y17772 = n50985 ;
  assign y17773 = ~1'b0 ;
  assign y17774 = ~n50988 ;
  assign y17775 = n50991 ;
  assign y17776 = n50992 ;
  assign y17777 = ~n50995 ;
  assign y17778 = ~n50998 ;
  assign y17779 = ~n50999 ;
  assign y17780 = n51002 ;
  assign y17781 = ~n51004 ;
  assign y17782 = ~1'b0 ;
  assign y17783 = ~n51010 ;
  assign y17784 = n51012 ;
  assign y17785 = ~1'b0 ;
  assign y17786 = n51013 ;
  assign y17787 = n51014 ;
  assign y17788 = ~n51015 ;
  assign y17789 = n51016 ;
  assign y17790 = n51018 ;
  assign y17791 = n51025 ;
  assign y17792 = ~1'b0 ;
  assign y17793 = ~n51027 ;
  assign y17794 = n51033 ;
  assign y17795 = n51035 ;
  assign y17796 = n51038 ;
  assign y17797 = n51040 ;
  assign y17798 = ~n51045 ;
  assign y17799 = n51049 ;
  assign y17800 = n51050 ;
  assign y17801 = ~n51053 ;
  assign y17802 = ~n51055 ;
  assign y17803 = ~1'b0 ;
  assign y17804 = n51057 ;
  assign y17805 = ~n51059 ;
  assign y17806 = ~1'b0 ;
  assign y17807 = ~n51060 ;
  assign y17808 = ~n51061 ;
  assign y17809 = n51065 ;
  assign y17810 = n51067 ;
  assign y17811 = ~n51070 ;
  assign y17812 = ~n51072 ;
  assign y17813 = ~1'b0 ;
  assign y17814 = n51074 ;
  assign y17815 = ~n51075 ;
  assign y17816 = ~n51078 ;
  assign y17817 = 1'b0 ;
  assign y17818 = ~n51083 ;
  assign y17819 = ~n29761 ;
  assign y17820 = n51085 ;
  assign y17821 = ~n51088 ;
  assign y17822 = ~n51091 ;
  assign y17823 = ~n51094 ;
  assign y17824 = n51096 ;
  assign y17825 = ~n51100 ;
  assign y17826 = ~n51102 ;
  assign y17827 = n51104 ;
  assign y17828 = ~n51106 ;
  assign y17829 = ~n51112 ;
  assign y17830 = ~n51114 ;
  assign y17831 = ~n51116 ;
  assign y17832 = ~n51117 ;
  assign y17833 = ~n51118 ;
  assign y17834 = ~n51119 ;
  assign y17835 = n51125 ;
  assign y17836 = ~1'b0 ;
  assign y17837 = ~1'b0 ;
  assign y17838 = ~n51126 ;
  assign y17839 = n16339 ;
  assign y17840 = ~1'b0 ;
  assign y17841 = ~n51130 ;
  assign y17842 = n51131 ;
  assign y17843 = n51134 ;
  assign y17844 = ~n51137 ;
  assign y17845 = ~1'b0 ;
  assign y17846 = ~n51138 ;
  assign y17847 = ~n51142 ;
  assign y17848 = n51143 ;
  assign y17849 = ~n51145 ;
  assign y17850 = n51146 ;
  assign y17851 = ~n51147 ;
  assign y17852 = ~n51148 ;
  assign y17853 = n51149 ;
  assign y17854 = n51150 ;
  assign y17855 = ~n51152 ;
  assign y17856 = ~1'b0 ;
  assign y17857 = n51155 ;
  assign y17858 = ~1'b0 ;
  assign y17859 = ~1'b0 ;
  assign y17860 = n51156 ;
  assign y17861 = ~n51157 ;
  assign y17862 = n51158 ;
  assign y17863 = n51163 ;
  assign y17864 = ~n51165 ;
  assign y17865 = n51167 ;
  assign y17866 = ~n51171 ;
  assign y17867 = n51173 ;
  assign y17868 = ~n51176 ;
  assign y17869 = ~n51178 ;
  assign y17870 = n26945 ;
  assign y17871 = ~n51184 ;
  assign y17872 = n51191 ;
  assign y17873 = n51192 ;
  assign y17874 = n51193 ;
  assign y17875 = ~n51195 ;
  assign y17876 = n51197 ;
  assign y17877 = ~1'b0 ;
  assign y17878 = ~n51200 ;
  assign y17879 = ~n51202 ;
  assign y17880 = ~n51204 ;
  assign y17881 = n51206 ;
  assign y17882 = n51209 ;
  assign y17883 = n51210 ;
  assign y17884 = ~n51211 ;
  assign y17885 = n51214 ;
  assign y17886 = ~n51217 ;
  assign y17887 = ~n51219 ;
  assign y17888 = ~n51223 ;
  assign y17889 = ~1'b0 ;
  assign y17890 = ~n51225 ;
  assign y17891 = n51227 ;
  assign y17892 = ~n51228 ;
  assign y17893 = ~n51229 ;
  assign y17894 = ~n51234 ;
  assign y17895 = n51235 ;
  assign y17896 = ~n51236 ;
  assign y17897 = ~n51241 ;
  assign y17898 = ~n51243 ;
  assign y17899 = ~n51251 ;
  assign y17900 = n30995 ;
  assign y17901 = ~n15289 ;
  assign y17902 = n51254 ;
  assign y17903 = n51257 ;
  assign y17904 = ~n51258 ;
  assign y17905 = n51259 ;
  assign y17906 = ~n51260 ;
  assign y17907 = n51261 ;
  assign y17908 = n6322 ;
  assign y17909 = n51264 ;
  assign y17910 = n51267 ;
  assign y17911 = n51268 ;
  assign y17912 = n51269 ;
  assign y17913 = ~n51274 ;
  assign y17914 = n51275 ;
  assign y17915 = ~n51277 ;
  assign y17916 = n51281 ;
  assign y17917 = n51282 ;
  assign y17918 = n51286 ;
  assign y17919 = ~n51288 ;
  assign y17920 = n51293 ;
  assign y17921 = n51295 ;
  assign y17922 = n51301 ;
  assign y17923 = ~n51304 ;
  assign y17924 = ~n51310 ;
  assign y17925 = ~n51311 ;
  assign y17926 = n51313 ;
  assign y17927 = n51314 ;
  assign y17928 = ~n51315 ;
  assign y17929 = ~1'b0 ;
  assign y17930 = ~n51317 ;
  assign y17931 = ~1'b0 ;
  assign y17932 = ~n51321 ;
  assign y17933 = n51326 ;
  assign y17934 = ~n51327 ;
  assign y17935 = ~n51328 ;
  assign y17936 = ~n51333 ;
  assign y17937 = ~1'b0 ;
  assign y17938 = ~n51335 ;
  assign y17939 = ~n34949 ;
  assign y17940 = n51337 ;
  assign y17941 = ~n51338 ;
  assign y17942 = n51341 ;
  assign y17943 = ~n51342 ;
  assign y17944 = n51343 ;
  assign y17945 = n51344 ;
  assign y17946 = ~n51345 ;
  assign y17947 = n51349 ;
  assign y17948 = ~n51351 ;
  assign y17949 = ~1'b0 ;
  assign y17950 = ~1'b0 ;
  assign y17951 = ~n51352 ;
  assign y17952 = ~n51362 ;
  assign y17953 = n51365 ;
  assign y17954 = n51366 ;
  assign y17955 = n51367 ;
  assign y17956 = ~n51372 ;
  assign y17957 = ~n51373 ;
  assign y17958 = ~n51375 ;
  assign y17959 = ~1'b0 ;
  assign y17960 = n51378 ;
  assign y17961 = ~1'b0 ;
  assign y17962 = ~1'b0 ;
  assign y17963 = ~n51380 ;
  assign y17964 = n51381 ;
  assign y17965 = ~n51384 ;
  assign y17966 = ~n51385 ;
  assign y17967 = n51386 ;
  assign y17968 = n51391 ;
  assign y17969 = ~n51392 ;
  assign y17970 = ~1'b0 ;
  assign y17971 = ~n51394 ;
  assign y17972 = n51395 ;
  assign y17973 = ~n51396 ;
  assign y17974 = ~n51400 ;
  assign y17975 = ~n51401 ;
  assign y17976 = n51403 ;
  assign y17977 = n51404 ;
  assign y17978 = n51409 ;
  assign y17979 = ~n51414 ;
  assign y17980 = n51415 ;
  assign y17981 = n51417 ;
  assign y17982 = ~n51420 ;
  assign y17983 = n51421 ;
  assign y17984 = ~n51425 ;
  assign y17985 = n51428 ;
  assign y17986 = n51429 ;
  assign y17987 = n51430 ;
  assign y17988 = n51436 ;
  assign y17989 = ~n51440 ;
  assign y17990 = ~n51442 ;
  assign y17991 = ~n51448 ;
  assign y17992 = ~1'b0 ;
  assign y17993 = ~n51450 ;
  assign y17994 = ~n51451 ;
  assign y17995 = ~n51456 ;
  assign y17996 = ~n51459 ;
  assign y17997 = ~n51464 ;
  assign y17998 = n51466 ;
  assign y17999 = ~n51471 ;
  assign y18000 = ~n51472 ;
  assign y18001 = n51477 ;
  assign y18002 = ~1'b0 ;
  assign y18003 = ~n51481 ;
  assign y18004 = ~1'b0 ;
  assign y18005 = ~1'b0 ;
  assign y18006 = n51485 ;
  assign y18007 = ~n51486 ;
  assign y18008 = n51487 ;
  assign y18009 = n51491 ;
  assign y18010 = n51493 ;
  assign y18011 = n51494 ;
  assign y18012 = ~1'b0 ;
  assign y18013 = ~1'b0 ;
  assign y18014 = ~1'b0 ;
  assign y18015 = n51495 ;
  assign y18016 = n51498 ;
  assign y18017 = ~n51501 ;
  assign y18018 = n51506 ;
  assign y18019 = n51508 ;
  assign y18020 = ~n51512 ;
  assign y18021 = ~n51513 ;
  assign y18022 = ~n50179 ;
  assign y18023 = ~1'b0 ;
  assign y18024 = ~n51514 ;
  assign y18025 = ~n51516 ;
  assign y18026 = ~n51522 ;
  assign y18027 = n51523 ;
  assign y18028 = ~n51524 ;
  assign y18029 = ~n51529 ;
  assign y18030 = ~n51533 ;
  assign y18031 = n51535 ;
  assign y18032 = ~n51538 ;
  assign y18033 = ~1'b0 ;
  assign y18034 = ~n51540 ;
  assign y18035 = ~n51547 ;
  assign y18036 = n51549 ;
  assign y18037 = n51550 ;
  assign y18038 = ~n51551 ;
  assign y18039 = ~n51552 ;
  assign y18040 = ~n51553 ;
  assign y18041 = ~n51555 ;
  assign y18042 = n51557 ;
  assign y18043 = ~n51560 ;
  assign y18044 = n51562 ;
  assign y18045 = n51564 ;
  assign y18046 = ~n51566 ;
  assign y18047 = n51567 ;
  assign y18048 = n51571 ;
  assign y18049 = n51575 ;
  assign y18050 = ~n51577 ;
  assign y18051 = ~n51578 ;
  assign y18052 = ~n51581 ;
  assign y18053 = ~n51582 ;
  assign y18054 = ~n51583 ;
  assign y18055 = ~1'b0 ;
  assign y18056 = ~n51584 ;
  assign y18057 = n51585 ;
  assign y18058 = ~n51586 ;
  assign y18059 = ~n51590 ;
  assign y18060 = n51591 ;
  assign y18061 = ~n51594 ;
  assign y18062 = ~n51597 ;
  assign y18063 = n51599 ;
  assign y18064 = ~n51609 ;
  assign y18065 = ~n51614 ;
  assign y18066 = n51618 ;
  assign y18067 = n51620 ;
  assign y18068 = ~n51621 ;
  assign y18069 = ~n51626 ;
  assign y18070 = ~n51635 ;
  assign y18071 = ~n51636 ;
  assign y18072 = ~n51638 ;
  assign y18073 = n51640 ;
  assign y18074 = ~n51641 ;
  assign y18075 = n51642 ;
  assign y18076 = n51643 ;
  assign y18077 = n51644 ;
  assign y18078 = ~n51645 ;
  assign y18079 = n51646 ;
  assign y18080 = n51647 ;
  assign y18081 = ~n51648 ;
  assign y18082 = ~1'b0 ;
  assign y18083 = ~1'b0 ;
  assign y18084 = ~n51650 ;
  assign y18085 = ~1'b0 ;
  assign y18086 = n51651 ;
  assign y18087 = ~n51653 ;
  assign y18088 = ~n51655 ;
  assign y18089 = ~n51656 ;
  assign y18090 = n51658 ;
  assign y18091 = n51659 ;
  assign y18092 = ~1'b0 ;
  assign y18093 = ~n51662 ;
  assign y18094 = ~n51665 ;
  assign y18095 = ~n51666 ;
  assign y18096 = n51667 ;
  assign y18097 = n51670 ;
  assign y18098 = n51672 ;
  assign y18099 = ~n51675 ;
  assign y18100 = ~1'b0 ;
  assign y18101 = ~1'b0 ;
  assign y18102 = ~n51679 ;
  assign y18103 = ~n51681 ;
  assign y18104 = ~n51683 ;
  assign y18105 = ~n51687 ;
  assign y18106 = n51690 ;
  assign y18107 = ~n51691 ;
  assign y18108 = ~n51693 ;
  assign y18109 = n51695 ;
  assign y18110 = n51696 ;
  assign y18111 = n51697 ;
  assign y18112 = n51701 ;
  assign y18113 = n51711 ;
  assign y18114 = n51712 ;
  assign y18115 = ~n51713 ;
  assign y18116 = n51714 ;
  assign y18117 = n51715 ;
  assign y18118 = n3329 ;
  assign y18119 = ~n51716 ;
  assign y18120 = ~n51720 ;
  assign y18121 = ~1'b0 ;
  assign y18122 = ~n51721 ;
  assign y18123 = n51723 ;
  assign y18124 = n51724 ;
  assign y18125 = ~n51725 ;
  assign y18126 = n51726 ;
  assign y18127 = ~n51727 ;
  assign y18128 = ~n51732 ;
  assign y18129 = ~n51736 ;
  assign y18130 = ~1'b0 ;
  assign y18131 = n51739 ;
  assign y18132 = ~1'b0 ;
  assign y18133 = n51740 ;
  assign y18134 = ~1'b0 ;
  assign y18135 = ~n51741 ;
  assign y18136 = n51744 ;
  assign y18137 = n51748 ;
  assign y18138 = ~n51754 ;
  assign y18139 = ~n51755 ;
  assign y18140 = ~n51757 ;
  assign y18141 = ~n51760 ;
  assign y18142 = n32674 ;
  assign y18143 = ~n51764 ;
  assign y18144 = ~1'b0 ;
  assign y18145 = n51765 ;
  assign y18146 = ~n51766 ;
  assign y18147 = ~n51767 ;
  assign y18148 = n51768 ;
  assign y18149 = n51773 ;
  assign y18150 = n51774 ;
  assign y18151 = ~n51776 ;
  assign y18152 = n51780 ;
  assign y18153 = ~n51782 ;
  assign y18154 = ~1'b0 ;
  assign y18155 = n51783 ;
  assign y18156 = ~n51790 ;
  assign y18157 = ~n51791 ;
  assign y18158 = ~n51795 ;
  assign y18159 = n51796 ;
  assign y18160 = ~n51798 ;
  assign y18161 = ~n51801 ;
  assign y18162 = ~n51804 ;
  assign y18163 = ~1'b0 ;
  assign y18164 = ~n51806 ;
  assign y18165 = ~n51807 ;
  assign y18166 = n51808 ;
  assign y18167 = ~n51812 ;
  assign y18168 = n51814 ;
  assign y18169 = n51821 ;
  assign y18170 = n51822 ;
  assign y18171 = ~n51826 ;
  assign y18172 = ~n51829 ;
  assign y18173 = ~1'b0 ;
  assign y18174 = n51833 ;
  assign y18175 = n51835 ;
  assign y18176 = ~n51839 ;
  assign y18177 = n51844 ;
  assign y18178 = ~n51847 ;
  assign y18179 = ~n51848 ;
  assign y18180 = n51849 ;
  assign y18181 = n51850 ;
  assign y18182 = ~n51854 ;
  assign y18183 = n51859 ;
  assign y18184 = ~n4413 ;
  assign y18185 = n51861 ;
  assign y18186 = ~1'b0 ;
  assign y18187 = n51862 ;
  assign y18188 = ~n51863 ;
  assign y18189 = ~n51866 ;
  assign y18190 = ~n51867 ;
  assign y18191 = n51869 ;
  assign y18192 = ~n51871 ;
  assign y18193 = ~1'b0 ;
  assign y18194 = ~n51874 ;
  assign y18195 = ~n51877 ;
  assign y18196 = n51879 ;
  assign y18197 = n51880 ;
  assign y18198 = n51883 ;
  assign y18199 = ~n51884 ;
  assign y18200 = n51885 ;
  assign y18201 = n51887 ;
  assign y18202 = n51889 ;
  assign y18203 = ~n51891 ;
  assign y18204 = ~n51892 ;
  assign y18205 = n51896 ;
  assign y18206 = ~1'b0 ;
  assign y18207 = ~n51900 ;
  assign y18208 = n51901 ;
  assign y18209 = ~n51904 ;
  assign y18210 = n51907 ;
  assign y18211 = ~n51908 ;
  assign y18212 = ~n51909 ;
  assign y18213 = ~1'b0 ;
  assign y18214 = ~1'b0 ;
  assign y18215 = ~n51913 ;
  assign y18216 = n51916 ;
  assign y18217 = ~1'b0 ;
  assign y18218 = n51918 ;
  assign y18219 = n51920 ;
  assign y18220 = ~n51922 ;
  assign y18221 = n51923 ;
  assign y18222 = n51924 ;
  assign y18223 = ~n51926 ;
  assign y18224 = n51929 ;
  assign y18225 = ~1'b0 ;
  assign y18226 = ~1'b0 ;
  assign y18227 = n51931 ;
  assign y18228 = n51933 ;
  assign y18229 = n51935 ;
  assign y18230 = ~n51937 ;
  assign y18231 = n51940 ;
  assign y18232 = n51941 ;
  assign y18233 = n51943 ;
  assign y18234 = ~n51949 ;
  assign y18235 = ~1'b0 ;
  assign y18236 = ~n51951 ;
  assign y18237 = ~n51957 ;
  assign y18238 = ~1'b0 ;
  assign y18239 = ~1'b0 ;
  assign y18240 = ~n3735 ;
  assign y18241 = ~n51958 ;
  assign y18242 = ~n51960 ;
  assign y18243 = n51961 ;
  assign y18244 = n51962 ;
  assign y18245 = ~n51963 ;
  assign y18246 = ~n51965 ;
  assign y18247 = ~n51966 ;
  assign y18248 = ~1'b0 ;
  assign y18249 = n51969 ;
  assign y18250 = ~1'b0 ;
  assign y18251 = n51970 ;
  assign y18252 = ~n51972 ;
  assign y18253 = n51975 ;
  assign y18254 = ~n51977 ;
  assign y18255 = ~n51978 ;
  assign y18256 = n51981 ;
  assign y18257 = ~1'b0 ;
  assign y18258 = n51984 ;
  assign y18259 = ~1'b0 ;
  assign y18260 = ~n51985 ;
  assign y18261 = ~n51987 ;
  assign y18262 = n51988 ;
  assign y18263 = ~n51989 ;
  assign y18264 = ~n51995 ;
  assign y18265 = n51997 ;
  assign y18266 = n51998 ;
  assign y18267 = ~n51999 ;
  assign y18268 = ~n52001 ;
  assign y18269 = ~n11141 ;
  assign y18270 = ~n52004 ;
  assign y18271 = ~n52005 ;
  assign y18272 = ~n52007 ;
  assign y18273 = ~n52008 ;
  assign y18274 = n52011 ;
  assign y18275 = ~n52012 ;
  assign y18276 = n52015 ;
  assign y18277 = ~n52016 ;
  assign y18278 = ~n52017 ;
  assign y18279 = ~n52019 ;
  assign y18280 = ~1'b0 ;
  assign y18281 = ~1'b0 ;
  assign y18282 = ~n52021 ;
  assign y18283 = n52025 ;
  assign y18284 = ~n52026 ;
  assign y18285 = ~n52028 ;
  assign y18286 = ~n52035 ;
  assign y18287 = n52038 ;
  assign y18288 = n52040 ;
  assign y18289 = ~1'b0 ;
  assign y18290 = ~n52042 ;
  assign y18291 = ~1'b0 ;
  assign y18292 = ~n52045 ;
  assign y18293 = ~n52053 ;
  assign y18294 = n52059 ;
  assign y18295 = n52062 ;
  assign y18296 = ~n52063 ;
  assign y18297 = n52065 ;
  assign y18298 = ~n52072 ;
  assign y18299 = n52073 ;
  assign y18300 = ~n52075 ;
  assign y18301 = n52081 ;
  assign y18302 = ~1'b0 ;
  assign y18303 = ~n52083 ;
  assign y18304 = n52085 ;
  assign y18305 = n52088 ;
  assign y18306 = n52090 ;
  assign y18307 = ~n52091 ;
  assign y18308 = n26411 ;
  assign y18309 = ~n52093 ;
  assign y18310 = n52096 ;
  assign y18311 = ~n52098 ;
  assign y18312 = ~1'b0 ;
  assign y18313 = n52100 ;
  assign y18314 = n52104 ;
  assign y18315 = n52107 ;
  assign y18316 = n52110 ;
  assign y18317 = ~n52115 ;
  assign y18318 = ~n52116 ;
  assign y18319 = n52118 ;
  assign y18320 = ~n52121 ;
  assign y18321 = ~n52123 ;
  assign y18322 = ~n52129 ;
  assign y18323 = ~n52131 ;
  assign y18324 = ~n52135 ;
  assign y18325 = ~n52137 ;
  assign y18326 = ~1'b0 ;
  assign y18327 = ~n52138 ;
  assign y18328 = ~n52142 ;
  assign y18329 = n52153 ;
  assign y18330 = ~n52156 ;
  assign y18331 = ~n52160 ;
  assign y18332 = n52161 ;
  assign y18333 = n52165 ;
  assign y18334 = ~1'b0 ;
  assign y18335 = ~n52167 ;
  assign y18336 = ~1'b0 ;
  assign y18337 = ~n52172 ;
  assign y18338 = n52176 ;
  assign y18339 = n52181 ;
  assign y18340 = n52182 ;
  assign y18341 = ~n52184 ;
  assign y18342 = ~n52185 ;
  assign y18343 = n52188 ;
  assign y18344 = n52189 ;
  assign y18345 = ~n52195 ;
  assign y18346 = ~n52196 ;
  assign y18347 = ~n52198 ;
  assign y18348 = ~1'b0 ;
  assign y18349 = ~n52199 ;
  assign y18350 = ~n52200 ;
  assign y18351 = ~n52203 ;
  assign y18352 = n52205 ;
  assign y18353 = n52206 ;
  assign y18354 = ~n52207 ;
  assign y18355 = ~1'b0 ;
  assign y18356 = n52210 ;
  assign y18357 = ~1'b0 ;
  assign y18358 = n52217 ;
  assign y18359 = ~1'b0 ;
  assign y18360 = ~n52221 ;
  assign y18361 = ~n52223 ;
  assign y18362 = ~n52225 ;
  assign y18363 = ~n52226 ;
  assign y18364 = ~n52227 ;
  assign y18365 = ~n52230 ;
  assign y18366 = n52237 ;
  assign y18367 = n52244 ;
  assign y18368 = ~n20602 ;
  assign y18369 = ~1'b0 ;
  assign y18370 = ~n52252 ;
  assign y18371 = n52253 ;
  assign y18372 = ~n52259 ;
  assign y18373 = n52260 ;
  assign y18374 = ~n52261 ;
  assign y18375 = n52263 ;
  assign y18376 = ~n52264 ;
  assign y18377 = ~n52266 ;
  assign y18378 = n52268 ;
  assign y18379 = ~n52271 ;
  assign y18380 = ~1'b0 ;
  assign y18381 = n52275 ;
  assign y18382 = ~n52278 ;
  assign y18383 = ~n52282 ;
  assign y18384 = ~n52284 ;
  assign y18385 = n52285 ;
  assign y18386 = ~n52286 ;
  assign y18387 = n52289 ;
  assign y18388 = ~1'b0 ;
  assign y18389 = ~n52291 ;
  assign y18390 = ~1'b0 ;
  assign y18391 = ~n52293 ;
  assign y18392 = ~n52295 ;
  assign y18393 = n52297 ;
  assign y18394 = n52298 ;
  assign y18395 = ~n52301 ;
  assign y18396 = ~n52303 ;
  assign y18397 = n52304 ;
  assign y18398 = n52306 ;
  assign y18399 = ~1'b0 ;
  assign y18400 = ~1'b0 ;
  assign y18401 = ~n52308 ;
  assign y18402 = ~n52309 ;
  assign y18403 = ~n52311 ;
  assign y18404 = n52313 ;
  assign y18405 = n52315 ;
  assign y18406 = n52318 ;
  assign y18407 = ~n52319 ;
  assign y18408 = n52324 ;
  assign y18409 = ~1'b0 ;
  assign y18410 = ~n52326 ;
  assign y18411 = n52327 ;
  assign y18412 = n52329 ;
  assign y18413 = n52330 ;
  assign y18414 = ~n52331 ;
  assign y18415 = n52334 ;
  assign y18416 = n52343 ;
  assign y18417 = ~n52348 ;
  assign y18418 = n52350 ;
  assign y18419 = ~n52351 ;
  assign y18420 = n52352 ;
  assign y18421 = n52354 ;
  assign y18422 = ~n52355 ;
  assign y18423 = n52357 ;
  assign y18424 = ~n52361 ;
  assign y18425 = n52362 ;
  assign y18426 = n52364 ;
  assign y18427 = n52372 ;
  assign y18428 = n52374 ;
  assign y18429 = ~n52375 ;
  assign y18430 = ~n52376 ;
  assign y18431 = ~n52380 ;
  assign y18432 = ~1'b0 ;
  assign y18433 = ~n52382 ;
  assign y18434 = ~1'b0 ;
  assign y18435 = ~n52383 ;
  assign y18436 = n52388 ;
  assign y18437 = ~n52391 ;
  assign y18438 = ~n52392 ;
  assign y18439 = n52395 ;
  assign y18440 = ~n52396 ;
  assign y18441 = ~n52397 ;
  assign y18442 = ~n52399 ;
  assign y18443 = ~1'b0 ;
  assign y18444 = ~n52403 ;
  assign y18445 = ~n52405 ;
  assign y18446 = ~n52406 ;
  assign y18447 = ~n52407 ;
  assign y18448 = n52408 ;
  assign y18449 = ~n52411 ;
  assign y18450 = ~n52412 ;
  assign y18451 = n52415 ;
  assign y18452 = ~n52419 ;
  assign y18453 = ~n52421 ;
  assign y18454 = n52423 ;
  assign y18455 = ~n16123 ;
  assign y18456 = ~n52425 ;
  assign y18457 = ~n27145 ;
  assign y18458 = n52426 ;
  assign y18459 = n52427 ;
  assign y18460 = n52431 ;
  assign y18461 = ~n52434 ;
  assign y18462 = ~1'b0 ;
  assign y18463 = ~n52440 ;
  assign y18464 = n52442 ;
  assign y18465 = ~n52443 ;
  assign y18466 = ~n52448 ;
  assign y18467 = ~n52449 ;
  assign y18468 = n52452 ;
  assign y18469 = n52453 ;
  assign y18470 = ~n52454 ;
  assign y18471 = n52462 ;
  assign y18472 = ~1'b0 ;
  assign y18473 = ~n52466 ;
  assign y18474 = ~1'b0 ;
  assign y18475 = ~1'b0 ;
  assign y18476 = ~n52467 ;
  assign y18477 = n52468 ;
  assign y18478 = ~n52469 ;
  assign y18479 = n52475 ;
  assign y18480 = n52478 ;
  assign y18481 = ~n52479 ;
  assign y18482 = ~n52486 ;
  assign y18483 = ~n52487 ;
  assign y18484 = n52488 ;
  assign y18485 = ~n52490 ;
  assign y18486 = ~n52493 ;
  assign y18487 = n52494 ;
  assign y18488 = ~n52495 ;
  assign y18489 = ~n52497 ;
  assign y18490 = ~n52499 ;
  assign y18491 = n52503 ;
  assign y18492 = n52505 ;
  assign y18493 = n52507 ;
  assign y18494 = ~1'b0 ;
  assign y18495 = ~1'b0 ;
  assign y18496 = ~n52508 ;
  assign y18497 = ~n52509 ;
  assign y18498 = ~n52513 ;
  assign y18499 = ~n52517 ;
  assign y18500 = n52520 ;
  assign y18501 = n52522 ;
  assign y18502 = ~1'b0 ;
  assign y18503 = ~1'b0 ;
  assign y18504 = ~n52525 ;
  assign y18505 = n52532 ;
  assign y18506 = ~n52533 ;
  assign y18507 = ~n52537 ;
  assign y18508 = ~n52538 ;
  assign y18509 = n46744 ;
  assign y18510 = n52539 ;
  assign y18511 = ~n52540 ;
  assign y18512 = n52544 ;
  assign y18513 = n52546 ;
  assign y18514 = ~1'b0 ;
  assign y18515 = ~n52548 ;
  assign y18516 = ~1'b0 ;
  assign y18517 = ~1'b0 ;
  assign y18518 = ~n52549 ;
  assign y18519 = ~n52551 ;
  assign y18520 = ~n52552 ;
  assign y18521 = n52553 ;
  assign y18522 = n52563 ;
  assign y18523 = n52567 ;
  assign y18524 = n52569 ;
  assign y18525 = n52572 ;
  assign y18526 = ~n52575 ;
  assign y18527 = n52576 ;
  assign y18528 = ~n52580 ;
  assign y18529 = n52585 ;
  assign y18530 = n52587 ;
  assign y18531 = ~n52591 ;
  assign y18532 = n52594 ;
  assign y18533 = ~n52596 ;
  assign y18534 = ~n12102 ;
  assign y18535 = n52597 ;
  assign y18536 = ~n52599 ;
  assign y18537 = ~n52604 ;
  assign y18538 = ~n52605 ;
  assign y18539 = ~n52607 ;
  assign y18540 = ~n23007 ;
  assign y18541 = ~n52608 ;
  assign y18542 = n52610 ;
  assign y18543 = ~n52611 ;
  assign y18544 = ~n52612 ;
  assign y18545 = ~n52614 ;
  assign y18546 = n52616 ;
  assign y18547 = ~1'b0 ;
  assign y18548 = ~1'b0 ;
  assign y18549 = ~n52625 ;
  assign y18550 = n52632 ;
  assign y18551 = ~n52634 ;
  assign y18552 = n52641 ;
  assign y18553 = n52644 ;
  assign y18554 = n52645 ;
  assign y18555 = n52647 ;
  assign y18556 = n52656 ;
  assign y18557 = ~n52658 ;
  assign y18558 = ~n52660 ;
  assign y18559 = ~n52661 ;
  assign y18560 = n52663 ;
  assign y18561 = ~n52665 ;
  assign y18562 = n52667 ;
  assign y18563 = ~n52669 ;
  assign y18564 = ~n52670 ;
  assign y18565 = ~n52674 ;
  assign y18566 = ~1'b0 ;
  assign y18567 = n52680 ;
  assign y18568 = ~n52686 ;
  assign y18569 = ~n52691 ;
  assign y18570 = ~n52692 ;
  assign y18571 = ~n52697 ;
  assign y18572 = n52700 ;
  assign y18573 = n52710 ;
  assign y18574 = n52711 ;
  assign y18575 = ~n52713 ;
  assign y18576 = ~1'b0 ;
  assign y18577 = ~n52717 ;
  assign y18578 = n52718 ;
  assign y18579 = ~n52719 ;
  assign y18580 = ~n52723 ;
  assign y18581 = ~n52724 ;
  assign y18582 = n52729 ;
  assign y18583 = ~n52732 ;
  assign y18584 = ~n52733 ;
  assign y18585 = ~n52734 ;
  assign y18586 = ~n52738 ;
  assign y18587 = ~1'b0 ;
  assign y18588 = ~n52740 ;
  assign y18589 = ~n52742 ;
  assign y18590 = n52744 ;
  assign y18591 = ~n52747 ;
  assign y18592 = n52748 ;
  assign y18593 = ~n52751 ;
  assign y18594 = n52754 ;
  assign y18595 = ~n52755 ;
  assign y18596 = ~1'b0 ;
  assign y18597 = ~1'b0 ;
  assign y18598 = ~1'b0 ;
  assign y18599 = ~n52758 ;
  assign y18600 = n52762 ;
  assign y18601 = ~n52763 ;
  assign y18602 = n52765 ;
  assign y18603 = n52766 ;
  assign y18604 = n52769 ;
  assign y18605 = n52771 ;
  assign y18606 = n52772 ;
  assign y18607 = ~1'b0 ;
  assign y18608 = ~1'b0 ;
  assign y18609 = ~n52776 ;
  assign y18610 = ~n52779 ;
  assign y18611 = ~n52780 ;
  assign y18612 = ~n52783 ;
  assign y18613 = ~n52784 ;
  assign y18614 = ~n52786 ;
  assign y18615 = ~n52787 ;
  assign y18616 = n52788 ;
  assign y18617 = ~n52792 ;
  assign y18618 = ~n52794 ;
  assign y18619 = ~n52796 ;
  assign y18620 = ~n52801 ;
  assign y18621 = n52807 ;
  assign y18622 = n52809 ;
  assign y18623 = ~n52813 ;
  assign y18624 = n52814 ;
  assign y18625 = ~n52816 ;
  assign y18626 = ~n52818 ;
  assign y18627 = ~n52821 ;
  assign y18628 = ~n52824 ;
  assign y18629 = ~n52826 ;
  assign y18630 = ~n52828 ;
  assign y18631 = ~1'b0 ;
  assign y18632 = n52830 ;
  assign y18633 = ~n52838 ;
  assign y18634 = ~n52841 ;
  assign y18635 = n52842 ;
  assign y18636 = n52845 ;
  assign y18637 = n52847 ;
  assign y18638 = ~n52850 ;
  assign y18639 = n52853 ;
  assign y18640 = n52854 ;
  assign y18641 = ~n52856 ;
  assign y18642 = n52860 ;
  assign y18643 = n52865 ;
  assign y18644 = n52869 ;
  assign y18645 = ~n52872 ;
  assign y18646 = n52873 ;
  assign y18647 = ~n52875 ;
  assign y18648 = ~n52876 ;
  assign y18649 = ~1'b0 ;
  assign y18650 = ~n52878 ;
  assign y18651 = n52880 ;
  assign y18652 = ~1'b0 ;
  assign y18653 = ~n52883 ;
  assign y18654 = n52884 ;
  assign y18655 = n52885 ;
  assign y18656 = ~n52887 ;
  assign y18657 = n52892 ;
  assign y18658 = n52897 ;
  assign y18659 = ~n52901 ;
  assign y18660 = n52902 ;
  assign y18661 = ~1'b0 ;
  assign y18662 = n52904 ;
  assign y18663 = n52907 ;
  assign y18664 = ~1'b0 ;
  assign y18665 = n52908 ;
  assign y18666 = n52911 ;
  assign y18667 = n52912 ;
  assign y18668 = ~n52915 ;
  assign y18669 = n52920 ;
  assign y18670 = ~n52922 ;
  assign y18671 = n52924 ;
  assign y18672 = n52929 ;
  assign y18673 = ~n52931 ;
  assign y18674 = ~1'b0 ;
  assign y18675 = ~n52932 ;
  assign y18676 = ~n52937 ;
  assign y18677 = ~n52938 ;
  assign y18678 = ~n52943 ;
  assign y18679 = ~n52947 ;
  assign y18680 = ~n52950 ;
  assign y18681 = ~n52952 ;
  assign y18682 = ~1'b0 ;
  assign y18683 = n52954 ;
  assign y18684 = n52955 ;
  assign y18685 = n52957 ;
  assign y18686 = n52958 ;
  assign y18687 = n52959 ;
  assign y18688 = n52960 ;
  assign y18689 = n52962 ;
  assign y18690 = n52964 ;
  assign y18691 = n52965 ;
  assign y18692 = ~n52967 ;
  assign y18693 = n37457 ;
  assign y18694 = ~1'b0 ;
  assign y18695 = n52971 ;
  assign y18696 = ~1'b0 ;
  assign y18697 = n52974 ;
  assign y18698 = ~n52977 ;
  assign y18699 = ~n52980 ;
  assign y18700 = ~n52981 ;
  assign y18701 = ~n52983 ;
  assign y18702 = ~n52986 ;
  assign y18703 = ~1'b0 ;
  assign y18704 = n52987 ;
  assign y18705 = ~1'b0 ;
  assign y18706 = ~1'b0 ;
  assign y18707 = ~n52990 ;
  assign y18708 = n52991 ;
  assign y18709 = n52992 ;
  assign y18710 = n52994 ;
  assign y18711 = ~n52996 ;
  assign y18712 = n52997 ;
  assign y18713 = ~1'b0 ;
  assign y18714 = n52998 ;
  assign y18715 = ~n53003 ;
  assign y18716 = ~n53005 ;
  assign y18717 = n53007 ;
  assign y18718 = n53010 ;
  assign y18719 = n53011 ;
  assign y18720 = ~n53012 ;
  assign y18721 = ~n53013 ;
  assign y18722 = n53016 ;
  assign y18723 = ~n53017 ;
  assign y18724 = n53018 ;
  assign y18725 = n53022 ;
  assign y18726 = ~n53023 ;
  assign y18727 = n53027 ;
  assign y18728 = n53028 ;
  assign y18729 = n53029 ;
  assign y18730 = ~n53030 ;
  assign y18731 = n53031 ;
  assign y18732 = ~n53035 ;
  assign y18733 = ~n53036 ;
  assign y18734 = n53038 ;
  assign y18735 = n53039 ;
  assign y18736 = ~n53041 ;
  assign y18737 = n53045 ;
  assign y18738 = ~n53047 ;
  assign y18739 = ~n53048 ;
  assign y18740 = ~n53049 ;
  assign y18741 = ~n53050 ;
  assign y18742 = ~n53053 ;
  assign y18743 = n53054 ;
  assign y18744 = ~n53055 ;
  assign y18745 = n53056 ;
  assign y18746 = ~n53058 ;
  assign y18747 = n53062 ;
  assign y18748 = ~1'b0 ;
  assign y18749 = n53066 ;
  assign y18750 = n53067 ;
  assign y18751 = ~n53070 ;
  assign y18752 = n53071 ;
  assign y18753 = ~n53075 ;
  assign y18754 = ~n53076 ;
  assign y18755 = ~n53077 ;
  assign y18756 = ~n53084 ;
  assign y18757 = ~n53088 ;
  assign y18758 = ~1'b0 ;
  assign y18759 = ~1'b0 ;
  assign y18760 = ~n53089 ;
  assign y18761 = ~n53092 ;
  assign y18762 = n53094 ;
  assign y18763 = ~n53095 ;
  assign y18764 = n53096 ;
  assign y18765 = n53097 ;
  assign y18766 = n53098 ;
  assign y18767 = ~1'b0 ;
  assign y18768 = ~n53100 ;
  assign y18769 = ~1'b0 ;
  assign y18770 = ~n53102 ;
  assign y18771 = ~1'b0 ;
  assign y18772 = n53104 ;
  assign y18773 = n53105 ;
  assign y18774 = ~n53108 ;
  assign y18775 = ~n53111 ;
  assign y18776 = n53112 ;
  assign y18777 = n53115 ;
  assign y18778 = ~1'b0 ;
  assign y18779 = n53118 ;
  assign y18780 = ~n53120 ;
  assign y18781 = ~n53122 ;
  assign y18782 = ~n53123 ;
  assign y18783 = ~n53127 ;
  assign y18784 = ~n53128 ;
  assign y18785 = ~n53129 ;
  assign y18786 = n53130 ;
  assign y18787 = n53131 ;
  assign y18788 = ~n53132 ;
  assign y18789 = ~1'b0 ;
  assign y18790 = ~1'b0 ;
  assign y18791 = ~n53136 ;
  assign y18792 = ~n53140 ;
  assign y18793 = ~n53141 ;
  assign y18794 = ~n53145 ;
  assign y18795 = n53147 ;
  assign y18796 = ~n800 ;
  assign y18797 = n53154 ;
  assign y18798 = ~1'b0 ;
  assign y18799 = ~1'b0 ;
  assign y18800 = ~n53160 ;
  assign y18801 = ~n53164 ;
  assign y18802 = ~n53167 ;
  assign y18803 = n32345 ;
  assign y18804 = n53168 ;
  assign y18805 = ~n53171 ;
  assign y18806 = n53172 ;
  assign y18807 = ~n53174 ;
  assign y18808 = ~n53175 ;
  assign y18809 = ~1'b0 ;
  assign y18810 = ~1'b0 ;
  assign y18811 = ~1'b0 ;
  assign y18812 = ~1'b0 ;
  assign y18813 = ~1'b0 ;
  assign y18814 = n53176 ;
  assign y18815 = ~n53178 ;
  assign y18816 = n53179 ;
  assign y18817 = ~n53183 ;
  assign y18818 = ~n53195 ;
  assign y18819 = ~n53197 ;
  assign y18820 = n53199 ;
  assign y18821 = ~n53201 ;
  assign y18822 = n53203 ;
  assign y18823 = n53206 ;
  assign y18824 = ~n53208 ;
  assign y18825 = n53211 ;
  assign y18826 = n53212 ;
  assign y18827 = n53213 ;
  assign y18828 = ~n53214 ;
  assign y18829 = n53215 ;
  assign y18830 = n7790 ;
  assign y18831 = ~1'b0 ;
  assign y18832 = ~n53217 ;
  assign y18833 = ~n53218 ;
  assign y18834 = ~n53220 ;
  assign y18835 = ~n53222 ;
  assign y18836 = ~n53223 ;
  assign y18837 = ~n53224 ;
  assign y18838 = n53229 ;
  assign y18839 = ~n53230 ;
  assign y18840 = n53232 ;
  assign y18841 = n53237 ;
  assign y18842 = n53239 ;
  assign y18843 = ~n53241 ;
  assign y18844 = ~n53246 ;
  assign y18845 = ~n53248 ;
  assign y18846 = ~1'b0 ;
  assign y18847 = n19766 ;
  assign y18848 = ~n53249 ;
  assign y18849 = n53253 ;
  assign y18850 = n53254 ;
  assign y18851 = ~n53255 ;
  assign y18852 = ~n53256 ;
  assign y18853 = n53259 ;
  assign y18854 = ~1'b0 ;
  assign y18855 = ~n53263 ;
  assign y18856 = n53267 ;
  assign y18857 = ~n53269 ;
  assign y18858 = n53270 ;
  assign y18859 = n53271 ;
  assign y18860 = ~n53272 ;
  assign y18861 = n53273 ;
  assign y18862 = n53274 ;
  assign y18863 = ~n53277 ;
  assign y18864 = n53278 ;
  assign y18865 = ~n53280 ;
  assign y18866 = ~n53282 ;
  assign y18867 = n53285 ;
  assign y18868 = ~n53288 ;
  assign y18869 = ~n53289 ;
  assign y18870 = n53292 ;
  assign y18871 = ~n53294 ;
  assign y18872 = n53296 ;
  assign y18873 = n53299 ;
  assign y18874 = ~n53304 ;
  assign y18875 = n53308 ;
  assign y18876 = n53311 ;
  assign y18877 = n53316 ;
  assign y18878 = ~1'b0 ;
  assign y18879 = ~n53320 ;
  assign y18880 = ~n53322 ;
  assign y18881 = ~n53323 ;
  assign y18882 = n53324 ;
  assign y18883 = ~n53325 ;
  assign y18884 = n53326 ;
  assign y18885 = n53327 ;
  assign y18886 = n53333 ;
  assign y18887 = n53335 ;
  assign y18888 = n53337 ;
  assign y18889 = ~n53340 ;
  assign y18890 = ~n53344 ;
  assign y18891 = n53351 ;
  assign y18892 = ~n53353 ;
  assign y18893 = ~n53354 ;
  assign y18894 = n53356 ;
  assign y18895 = n53360 ;
  assign y18896 = ~n53364 ;
  assign y18897 = ~1'b0 ;
  assign y18898 = ~n53370 ;
  assign y18899 = ~n53372 ;
  assign y18900 = n1237 ;
  assign y18901 = n53373 ;
  assign y18902 = ~n53374 ;
  assign y18903 = n53378 ;
  assign y18904 = n53380 ;
  assign y18905 = n53381 ;
  assign y18906 = n53382 ;
  assign y18907 = ~n53384 ;
  assign y18908 = n53386 ;
  assign y18909 = n53388 ;
  assign y18910 = ~n53389 ;
  assign y18911 = ~n53393 ;
  assign y18912 = n53394 ;
  assign y18913 = ~n53397 ;
  assign y18914 = n53400 ;
  assign y18915 = ~n53402 ;
  assign y18916 = n53403 ;
  assign y18917 = ~n53404 ;
  assign y18918 = ~n53406 ;
  assign y18919 = ~1'b0 ;
  assign y18920 = n53407 ;
  assign y18921 = ~1'b0 ;
  assign y18922 = n53408 ;
  assign y18923 = ~n53410 ;
  assign y18924 = ~n53414 ;
  assign y18925 = n53415 ;
  assign y18926 = n53420 ;
  assign y18927 = n53421 ;
  assign y18928 = n53422 ;
  assign y18929 = n53423 ;
  assign y18930 = n19295 ;
  assign y18931 = ~n53425 ;
  assign y18932 = ~1'b0 ;
  assign y18933 = n53427 ;
  assign y18934 = ~n53428 ;
  assign y18935 = n53431 ;
  assign y18936 = n53432 ;
  assign y18937 = ~n53436 ;
  assign y18938 = ~n53438 ;
  assign y18939 = ~n53439 ;
  assign y18940 = ~1'b0 ;
  assign y18941 = ~1'b0 ;
  assign y18942 = ~1'b0 ;
  assign y18943 = n53441 ;
  assign y18944 = ~1'b0 ;
  assign y18945 = n53444 ;
  assign y18946 = ~n53451 ;
  assign y18947 = ~n53452 ;
  assign y18948 = ~n53453 ;
  assign y18949 = n53456 ;
  assign y18950 = n53457 ;
  assign y18951 = ~1'b0 ;
  assign y18952 = ~n53462 ;
  assign y18953 = ~1'b0 ;
  assign y18954 = ~n53464 ;
  assign y18955 = n53469 ;
  assign y18956 = n53470 ;
  assign y18957 = ~n53471 ;
  assign y18958 = ~n53472 ;
  assign y18959 = n53475 ;
  assign y18960 = n53483 ;
  assign y18961 = ~n53485 ;
  assign y18962 = n53489 ;
  assign y18963 = ~n53491 ;
  assign y18964 = ~n53492 ;
  assign y18965 = ~1'b0 ;
  assign y18966 = ~n53493 ;
  assign y18967 = ~n53494 ;
  assign y18968 = ~n53496 ;
  assign y18969 = ~n53500 ;
  assign y18970 = n53502 ;
  assign y18971 = ~n53505 ;
  assign y18972 = ~n53510 ;
  assign y18973 = ~n53512 ;
  assign y18974 = ~n53517 ;
  assign y18975 = ~1'b0 ;
  assign y18976 = ~1'b0 ;
  assign y18977 = ~n53520 ;
  assign y18978 = ~n53525 ;
  assign y18979 = ~n53526 ;
  assign y18980 = n53527 ;
  assign y18981 = n53529 ;
  assign y18982 = ~n53530 ;
  assign y18983 = ~1'b0 ;
  assign y18984 = ~1'b0 ;
  assign y18985 = ~n53532 ;
  assign y18986 = ~1'b0 ;
  assign y18987 = ~1'b0 ;
  assign y18988 = n53533 ;
  assign y18989 = ~n53537 ;
  assign y18990 = ~n53541 ;
  assign y18991 = n53544 ;
  assign y18992 = ~n53545 ;
  assign y18993 = ~n53547 ;
  assign y18994 = ~1'b0 ;
  assign y18995 = ~n53549 ;
  assign y18996 = n53550 ;
  assign y18997 = n53551 ;
  assign y18998 = n53554 ;
  assign y18999 = ~n53557 ;
  assign y19000 = ~n53559 ;
  assign y19001 = n53562 ;
  assign y19002 = n53563 ;
  assign y19003 = ~n53568 ;
  assign y19004 = ~n53573 ;
  assign y19005 = ~n53575 ;
  assign y19006 = ~1'b0 ;
  assign y19007 = ~n53580 ;
  assign y19008 = n53582 ;
  assign y19009 = ~n53584 ;
  assign y19010 = n53585 ;
  assign y19011 = n53586 ;
  assign y19012 = n53587 ;
  assign y19013 = ~n53588 ;
  assign y19014 = n53593 ;
  assign y19015 = ~n53595 ;
  assign y19016 = ~n53597 ;
  assign y19017 = ~1'b0 ;
  assign y19018 = ~n53599 ;
  assign y19019 = ~1'b0 ;
  assign y19020 = 1'b0 ;
  assign y19021 = ~n53602 ;
  assign y19022 = ~n53606 ;
  assign y19023 = n53610 ;
  assign y19024 = ~n53611 ;
  assign y19025 = n53614 ;
  assign y19026 = ~n53619 ;
  assign y19027 = n53622 ;
  assign y19028 = ~1'b0 ;
  assign y19029 = ~n53624 ;
  assign y19030 = n53631 ;
  assign y19031 = n53638 ;
  assign y19032 = ~n53640 ;
  assign y19033 = n53641 ;
  assign y19034 = ~n53642 ;
  assign y19035 = n53644 ;
  assign y19036 = ~n53647 ;
  assign y19037 = ~n53648 ;
  assign y19038 = ~n53649 ;
  assign y19039 = n53650 ;
  assign y19040 = n53656 ;
  assign y19041 = ~1'b0 ;
  assign y19042 = ~1'b0 ;
  assign y19043 = ~n53659 ;
  assign y19044 = n53662 ;
  assign y19045 = n53663 ;
  assign y19046 = n53664 ;
  assign y19047 = n53665 ;
  assign y19048 = ~n53669 ;
  assign y19049 = ~1'b0 ;
  assign y19050 = n53671 ;
  assign y19051 = ~1'b0 ;
  assign y19052 = n53674 ;
  assign y19053 = n53676 ;
  assign y19054 = ~n53681 ;
  assign y19055 = ~n53682 ;
  assign y19056 = n53683 ;
  assign y19057 = n53684 ;
  assign y19058 = n53688 ;
  assign y19059 = n53689 ;
  assign y19060 = ~1'b0 ;
  assign y19061 = ~1'b0 ;
  assign y19062 = ~n53691 ;
  assign y19063 = ~1'b0 ;
  assign y19064 = n53693 ;
  assign y19065 = ~n53695 ;
  assign y19066 = ~n53696 ;
  assign y19067 = n53697 ;
  assign y19068 = ~n53698 ;
  assign y19069 = n53701 ;
  assign y19070 = n53704 ;
  assign y19071 = ~n18088 ;
  assign y19072 = n53706 ;
  assign y19073 = ~n53707 ;
  assign y19074 = ~1'b0 ;
  assign y19075 = n53708 ;
  assign y19076 = n53709 ;
  assign y19077 = ~1'b0 ;
  assign y19078 = n53712 ;
  assign y19079 = ~n53714 ;
  assign y19080 = n53715 ;
  assign y19081 = n53716 ;
  assign y19082 = ~1'b0 ;
  assign y19083 = ~1'b0 ;
  assign y19084 = n53720 ;
  assign y19085 = n53722 ;
  assign y19086 = ~1'b0 ;
  assign y19087 = n53728 ;
  assign y19088 = n53731 ;
  assign y19089 = n53732 ;
  assign y19090 = ~n53734 ;
  assign y19091 = ~n53735 ;
  assign y19092 = ~n53738 ;
  assign y19093 = ~n53742 ;
  assign y19094 = n53747 ;
  assign y19095 = ~1'b0 ;
  assign y19096 = ~n53749 ;
  assign y19097 = ~n53751 ;
  assign y19098 = ~n53752 ;
  assign y19099 = n53753 ;
  assign y19100 = n53757 ;
  assign y19101 = ~n53758 ;
  assign y19102 = ~n53759 ;
  assign y19103 = ~n53763 ;
  assign y19104 = ~n53765 ;
  assign y19105 = n53767 ;
  assign y19106 = n53772 ;
  assign y19107 = n53778 ;
  assign y19108 = ~1'b0 ;
  assign y19109 = n53780 ;
  assign y19110 = n53785 ;
  assign y19111 = n53788 ;
  assign y19112 = ~n53791 ;
  assign y19113 = n53794 ;
  assign y19114 = ~n53796 ;
  assign y19115 = ~1'b0 ;
  assign y19116 = ~1'b0 ;
  assign y19117 = ~1'b0 ;
  assign y19118 = ~n53799 ;
  assign y19119 = n53801 ;
  assign y19120 = ~n53802 ;
  assign y19121 = ~n53803 ;
  assign y19122 = n34300 ;
  assign y19123 = n53807 ;
  assign y19124 = n53808 ;
  assign y19125 = ~n53809 ;
  assign y19126 = ~n53811 ;
  assign y19127 = n53813 ;
  assign y19128 = n53815 ;
  assign y19129 = n53818 ;
  assign y19130 = ~n53821 ;
  assign y19131 = n53827 ;
  assign y19132 = ~n53830 ;
  assign y19133 = ~n53834 ;
  assign y19134 = ~n53835 ;
  assign y19135 = n53839 ;
  assign y19136 = ~n53840 ;
  assign y19137 = ~1'b0 ;
  assign y19138 = ~1'b0 ;
endmodule
