module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n408 , n409 , n410 , n412 , n413 , n414 , n415 , n416 , n417 , n419 , n420 , n421 , n423 , n424 , n425 ;
  assign n8 = x0 & ~x1 ;
  assign n9 = x3 & x4 ;
  assign n10 = n8 & n9 ;
  assign n11 = x1 & x3 ;
  assign n12 = x4 & n11 ;
  assign n13 = ~n10 & ~n12 ;
  assign n14 = ~x2 & ~n13 ;
  assign n15 = ~x1 & x3 ;
  assign n16 = x4 & n15 ;
  assign n17 = ~x3 & ~x4 ;
  assign n18 = ~n9 & ~n17 ;
  assign n19 = x1 & ~n18 ;
  assign n20 = ~n16 & ~n19 ;
  assign n21 = x2 & ~n20 ;
  assign n22 = ~n14 & ~n21 ;
  assign n36 = ~n22 & x7 ;
  assign n23 = ~x0 & x1 ;
  assign n24 = n17 & n23 ;
  assign n25 = ~x1 & ~x3 ;
  assign n26 = ~x4 & n25 ;
  assign n27 = ~n24 & ~n26 ;
  assign n28 = x2 & ~n27 ;
  assign n29 = x1 & ~x3 ;
  assign n30 = ~x4 & n29 ;
  assign n31 = ~x1 & ~n18 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = ~x2 & ~n32 ;
  assign n34 = ~n28 & ~n33 ;
  assign n37 = n34 & ~x7 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = ~x0 & ~n9 ;
  assign n40 = ~x0 & ~n39 ;
  assign n41 = ~x1 & ~n40 ;
  assign n42 = ~x3 & ~n17 ;
  assign n43 = x1 & ~n42 ;
  assign n44 = ~n41 & ~n43 ;
  assign n45 = ~x2 & ~n44 ;
  assign n46 = ~x3 & x4 ;
  assign n47 = ~x3 & ~n46 ;
  assign n48 = x1 & ~n47 ;
  assign n49 = x1 & ~n48 ;
  assign n50 = x2 & ~n49 ;
  assign n51 = ~n45 & ~n50 ;
  assign n66 = n51 & x8 ;
  assign n52 = x0 & ~n17 ;
  assign n53 = x0 & ~n52 ;
  assign n54 = x1 & ~n53 ;
  assign n55 = x3 & ~n9 ;
  assign n56 = ~x1 & ~n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = x2 & ~n57 ;
  assign n59 = x3 & ~x4 ;
  assign n60 = x3 & ~n59 ;
  assign n61 = ~x1 & ~n60 ;
  assign n62 = ~x1 & ~n61 ;
  assign n63 = ~x2 & ~n62 ;
  assign n64 = ~n58 & ~n63 ;
  assign n67 = ~n64 & ~x8 ;
  assign n68 = ~n66 & ~n67 ;
  assign n69 = ~x0 & ~n18 ;
  assign n70 = x0 & ~n55 ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = x1 & ~n71 ;
  assign n73 = ~n41 & ~n72 ;
  assign n74 = ~x2 & ~n73 ;
  assign n75 = ~x2 & ~n74 ;
  assign n84 = n75 & x9 ;
  assign n76 = x0 & ~n18 ;
  assign n77 = ~x0 & ~n42 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = ~x1 & ~n78 ;
  assign n80 = ~n54 & ~n79 ;
  assign n81 = x2 & ~n80 ;
  assign n82 = x2 & ~n81 ;
  assign n85 = ~n82 & ~x9 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = ~x0 & ~x3 ;
  assign n88 = ~n46 & n87 ;
  assign n89 = ~n76 & ~n88 ;
  assign n90 = ~x1 & ~n89 ;
  assign n91 = ~n43 & ~n90 ;
  assign n92 = ~x2 & ~n91 ;
  assign n93 = x2 & ~n42 ;
  assign n94 = ~n92 & ~n93 ;
  assign n104 = n94 & x10 ;
  assign n95 = x0 & x3 ;
  assign n96 = ~n59 & n95 ;
  assign n97 = ~n69 & ~n96 ;
  assign n98 = x1 & ~n97 ;
  assign n99 = ~n56 & ~n98 ;
  assign n100 = x2 & ~n99 ;
  assign n101 = ~x2 & ~n55 ;
  assign n102 = ~n100 & ~n101 ;
  assign n105 = ~n102 & ~x10 ;
  assign n106 = ~n104 & ~n105 ;
  assign n107 = ~x0 & x3 ;
  assign n108 = x4 & x5 ;
  assign n109 = n107 & n108 ;
  assign n110 = x3 & ~x6 ;
  assign n111 = ~n9 & n110 ;
  assign n112 = x3 & ~x5 ;
  assign n113 = ~n9 & n112 ;
  assign n114 = x3 & x5 ;
  assign n115 = ~n113 & ~n114 ;
  assign n116 = x6 & ~n115 ;
  assign n117 = ~n111 & ~n116 ;
  assign n118 = x0 & ~n117 ;
  assign n119 = ~n109 & ~n118 ;
  assign n120 = x1 & ~n119 ;
  assign n121 = ~x2 & ~n120 ;
  assign n122 = x0 & ~n42 ;
  assign n123 = x0 & ~n122 ;
  assign n124 = x2 & ~n123 ;
  assign n125 = ~n121 & ~n124 ;
  assign n146 = n125 & x11 ;
  assign n126 = x0 & ~x3 ;
  assign n127 = ~x4 & ~x5 ;
  assign n128 = n126 & n127 ;
  assign n129 = ~x3 & x6 ;
  assign n130 = ~n17 & n129 ;
  assign n131 = ~x3 & x5 ;
  assign n132 = ~n17 & n131 ;
  assign n133 = ~x3 & ~x5 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = ~x6 & ~n134 ;
  assign n136 = ~n130 & ~n135 ;
  assign n137 = ~x0 & ~n136 ;
  assign n138 = ~n128 & ~n137 ;
  assign n139 = ~x1 & ~n138 ;
  assign n140 = x2 & ~n139 ;
  assign n141 = ~x0 & ~n55 ;
  assign n142 = ~x0 & ~n141 ;
  assign n143 = ~x2 & ~n142 ;
  assign n144 = ~n140 & ~n143 ;
  assign n147 = ~n144 & ~x11 ;
  assign n148 = ~n146 & ~n147 ;
  assign n149 = x3 & x6 ;
  assign n150 = ~n111 & ~n149 ;
  assign n151 = x1 & ~n150 ;
  assign n152 = ~x2 & ~n151 ;
  assign n153 = x1 & ~n43 ;
  assign n154 = x2 & ~n153 ;
  assign n155 = ~n152 & ~n154 ;
  assign n164 = n155 & x12 ;
  assign n156 = ~x3 & ~x6 ;
  assign n157 = ~n130 & ~n156 ;
  assign n158 = ~x1 & ~n157 ;
  assign n159 = x2 & ~n158 ;
  assign n160 = ~x1 & ~n56 ;
  assign n161 = ~x2 & ~n160 ;
  assign n162 = ~n159 & ~n161 ;
  assign n165 = ~n162 & ~x12 ;
  assign n166 = ~n164 & ~n165 ;
  assign n167 = ~x1 & ~n9 ;
  assign n168 = ~n17 & n167 ;
  assign n169 = ~n17 & n39 ;
  assign n170 = x0 & ~n47 ;
  assign n171 = ~n169 & ~n170 ;
  assign n172 = x1 & ~n171 ;
  assign n173 = ~n168 & ~n172 ;
  assign n174 = ~x2 & ~n173 ;
  assign n175 = x2 & x3 ;
  assign n176 = x4 & n175 ;
  assign n177 = ~n174 & ~n176 ;
  assign n190 = ~n177 & x13 ;
  assign n178 = x1 & ~n17 ;
  assign n179 = ~n9 & n178 ;
  assign n180 = ~n9 & n52 ;
  assign n181 = ~x0 & ~n60 ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = ~x1 & ~n182 ;
  assign n184 = ~n179 & ~n183 ;
  assign n185 = x2 & ~n184 ;
  assign n186 = ~x2 & ~x3 ;
  assign n187 = ~x4 & n186 ;
  assign n188 = ~n185 & ~n187 ;
  assign n191 = n188 & ~x13 ;
  assign n192 = ~n190 & ~n191 ;
  assign n193 = ~x1 & ~x2 ;
  assign n194 = ~n41 & n193 ;
  assign n195 = x1 & ~n89 ;
  assign n196 = ~n10 & ~n195 ;
  assign n197 = x2 & ~n196 ;
  assign n198 = ~n194 & ~n197 ;
  assign n206 = ~n198 & x14 ;
  assign n199 = x1 & x2 ;
  assign n200 = ~n54 & n199 ;
  assign n201 = ~x1 & ~n97 ;
  assign n202 = ~n24 & ~n201 ;
  assign n203 = ~x2 & ~n202 ;
  assign n204 = ~n200 & ~n203 ;
  assign n207 = n204 & ~x14 ;
  assign n208 = ~n206 & ~n207 ;
  assign n209 = ~x0 & ~n77 ;
  assign n210 = x1 & ~n209 ;
  assign n211 = x1 & ~x2 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = ~n18 & n199 ;
  assign n214 = ~n212 & ~n213 ;
  assign n222 = ~n214 & x15 ;
  assign n215 = x0 & ~n70 ;
  assign n216 = ~x1 & ~n215 ;
  assign n217 = ~x1 & x2 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = ~n18 & n193 ;
  assign n220 = ~n218 & ~n219 ;
  assign n223 = n220 & ~x15 ;
  assign n224 = ~n222 & ~n223 ;
  assign n225 = ~n167 & ~n210 ;
  assign n226 = ~x2 & ~n225 ;
  assign n227 = ~n50 & ~n226 ;
  assign n232 = n227 & x16 ;
  assign n228 = ~n178 & ~n216 ;
  assign n229 = x2 & ~n228 ;
  assign n230 = ~n63 & ~n229 ;
  assign n233 = ~n230 & ~x16 ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = ~n107 & ~n170 ;
  assign n236 = x1 & ~n235 ;
  assign n237 = ~x2 & ~n168 ;
  assign n238 = ~n236 & n237 ;
  assign n239 = ~n93 & ~n238 ;
  assign n246 = n239 & x17 ;
  assign n240 = ~n126 & ~n181 ;
  assign n241 = ~x1 & ~n240 ;
  assign n242 = x2 & ~n179 ;
  assign n243 = ~n241 & n242 ;
  assign n244 = ~n101 & ~n243 ;
  assign n247 = ~n244 & ~x17 ;
  assign n248 = ~n246 & ~n247 ;
  assign n249 = ~x0 & ~n47 ;
  assign n250 = ~x0 & ~n249 ;
  assign n251 = ~x1 & ~n250 ;
  assign n252 = ~x1 & ~n251 ;
  assign n253 = ~x2 & ~n252 ;
  assign n254 = ~x2 & ~n253 ;
  assign n262 = n254 & x18 ;
  assign n255 = x0 & ~n60 ;
  assign n256 = x0 & ~n255 ;
  assign n257 = x1 & ~n256 ;
  assign n258 = x1 & ~n257 ;
  assign n259 = x2 & ~n258 ;
  assign n260 = x2 & ~n259 ;
  assign n263 = ~n260 & ~x18 ;
  assign n264 = ~n262 & ~n263 ;
  assign n265 = ~x1 & ~n235 ;
  assign n266 = ~n48 & ~n265 ;
  assign n267 = ~x2 & ~n266 ;
  assign n268 = ~x1 & x4 ;
  assign n269 = x1 & ~n55 ;
  assign n270 = ~n268 & ~n269 ;
  assign n271 = x2 & ~n270 ;
  assign n272 = ~n267 & ~n271 ;
  assign n282 = ~n272 & x19 ;
  assign n273 = x1 & ~n240 ;
  assign n274 = ~n61 & ~n273 ;
  assign n275 = x2 & ~n274 ;
  assign n276 = x1 & ~x4 ;
  assign n277 = ~x1 & ~n42 ;
  assign n278 = ~n276 & ~n277 ;
  assign n279 = ~x2 & ~n278 ;
  assign n280 = ~n275 & ~n279 ;
  assign n283 = n280 & ~x19 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = x0 & ~n170 ;
  assign n286 = x2 & ~n285 ;
  assign n287 = x2 & ~n286 ;
  assign n292 = n287 & x20 ;
  assign n288 = ~x0 & ~n181 ;
  assign n289 = ~x2 & ~n288 ;
  assign n290 = ~x2 & ~n289 ;
  assign n293 = ~n290 & ~x20 ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = x2 & ~n250 ;
  assign n296 = x2 & ~n295 ;
  assign n300 = n296 & x21 ;
  assign n297 = ~x2 & ~n256 ;
  assign n298 = ~x2 & ~n297 ;
  assign n301 = ~n298 & ~x21 ;
  assign n302 = ~n300 & ~n301 ;
  assign n303 = ~x1 & ~n142 ;
  assign n304 = ~x1 & ~n303 ;
  assign n305 = x2 & ~n304 ;
  assign n306 = x2 & ~n305 ;
  assign n312 = n306 & x22 ;
  assign n307 = x1 & ~n123 ;
  assign n308 = x1 & ~n307 ;
  assign n309 = ~x2 & ~n308 ;
  assign n310 = ~x2 & ~n309 ;
  assign n313 = ~n310 & ~x22 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = ~x1 & ~n216 ;
  assign n316 = x2 & ~n315 ;
  assign n317 = x2 & ~n316 ;
  assign n322 = n317 & x23 ;
  assign n318 = x1 & ~n210 ;
  assign n319 = ~x2 & ~n318 ;
  assign n320 = ~x2 & ~n319 ;
  assign n323 = ~n320 & ~x23 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = x1 & ~n215 ;
  assign n326 = x1 & ~n325 ;
  assign n327 = x2 & ~n326 ;
  assign n328 = x2 & ~n327 ;
  assign n334 = n328 & x24 ;
  assign n329 = ~x1 & ~n209 ;
  assign n330 = ~x1 & ~n329 ;
  assign n331 = ~x2 & ~n330 ;
  assign n332 = ~x2 & ~n331 ;
  assign n335 = ~n332 & ~x24 ;
  assign n336 = ~n334 & ~n335 ;
  assign n337 = x1 & ~n142 ;
  assign n338 = x1 & ~n337 ;
  assign n339 = x2 & ~n338 ;
  assign n340 = x2 & ~n339 ;
  assign n346 = n340 & x25 ;
  assign n341 = ~x1 & ~n123 ;
  assign n342 = ~x1 & ~n341 ;
  assign n343 = ~x2 & ~n342 ;
  assign n344 = ~x2 & ~n343 ;
  assign n347 = ~n344 & ~x25 ;
  assign n348 = ~n346 & ~n347 ;
  assign n349 = x2 & ~n47 ;
  assign n350 = x2 & ~n349 ;
  assign n354 = n350 & x26 ;
  assign n351 = ~x2 & ~n60 ;
  assign n352 = ~x2 & ~n351 ;
  assign n355 = ~n352 & ~x26 ;
  assign n356 = ~n354 & ~n355 ;
  assign n357 = x0 & x1 ;
  assign n358 = ~n115 & n357 ;
  assign n359 = n8 & ~n70 ;
  assign n360 = ~x2 & ~n359 ;
  assign n361 = ~n358 & n360 ;
  assign n362 = x1 & ~n40 ;
  assign n363 = ~n167 & ~n362 ;
  assign n364 = x2 & ~n363 ;
  assign n365 = ~n361 & ~n364 ;
  assign n376 = n365 & x27 ;
  assign n366 = ~x0 & ~x1 ;
  assign n367 = ~n134 & n366 ;
  assign n368 = n23 & ~n77 ;
  assign n369 = x2 & ~n368 ;
  assign n370 = ~n367 & n369 ;
  assign n371 = ~x1 & ~n53 ;
  assign n372 = ~n178 & ~n371 ;
  assign n373 = ~x2 & ~n372 ;
  assign n374 = ~n370 & ~n373 ;
  assign n377 = ~n374 & ~x27 ;
  assign n378 = ~n376 & ~n377 ;
  assign n379 = x5 & n9 ;
  assign n380 = ~x6 & ~n379 ;
  assign n381 = ~x6 & ~n380 ;
  assign n382 = x0 & ~n381 ;
  assign n383 = x0 & ~n382 ;
  assign n384 = x1 & ~n383 ;
  assign n385 = ~n216 & ~n384 ;
  assign n386 = ~x2 & ~n385 ;
  assign n387 = ~x2 & ~n386 ;
  assign n398 = n387 & x28 ;
  assign n388 = ~x5 & n17 ;
  assign n389 = x6 & ~n388 ;
  assign n390 = x6 & ~n389 ;
  assign n391 = ~x0 & ~n390 ;
  assign n392 = ~x0 & ~n391 ;
  assign n393 = ~x1 & ~n392 ;
  assign n394 = ~n210 & ~n393 ;
  assign n395 = x2 & ~n394 ;
  assign n396 = x2 & ~n395 ;
  assign n399 = ~n396 & ~x28 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = ~n117 & n357 ;
  assign n402 = ~x2 & ~n401 ;
  assign n403 = ~n364 & ~n402 ;
  assign n408 = n403 & x29 ;
  assign n404 = ~n136 & n366 ;
  assign n405 = x2 & ~n404 ;
  assign n406 = ~n373 & ~n405 ;
  assign n409 = ~n406 & ~x29 ;
  assign n410 = ~n408 & ~n409 ;
  assign n412 = ~n307 & ~n329 ;
  assign n413 = ~x2 & ~n412 ;
  assign n414 = ~x2 & ~n413 ;
  assign n419 = n414 & x31 ;
  assign n415 = ~n303 & ~n325 ;
  assign n416 = x2 & ~n415 ;
  assign n417 = x2 & ~n416 ;
  assign n420 = ~n417 & ~x31 ;
  assign n421 = ~n419 & ~n420 ;
  assign n423 = n344 & x32 ;
  assign n424 = ~n340 & ~x32 ;
  assign n425 = ~n423 & ~n424 ;
  assign y0 = ~n38 ;
  assign y1 = ~n68 ;
  assign y2 = ~n86 ;
  assign y3 = ~n106 ;
  assign y4 = ~n148 ;
  assign y5 = ~n166 ;
  assign y6 = ~n192 ;
  assign y7 = ~n208 ;
  assign y8 = ~n224 ;
  assign y9 = ~n234 ;
  assign y10 = ~n248 ;
  assign y11 = ~n264 ;
  assign y12 = ~n284 ;
  assign y13 = ~n294 ;
  assign y14 = ~n302 ;
  assign y15 = ~n314 ;
  assign y16 = ~n324 ;
  assign y17 = ~n336 ;
  assign y18 = ~n348 ;
  assign y19 = ~n356 ;
  assign y20 = ~n378 ;
  assign y21 = ~n400 ;
  assign y22 = ~n410 ;
  assign y23 = x30 ;
  assign y24 = ~n421 ;
  assign y25 = ~n425 ;
endmodule
