module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 , y23806 , y23807 , y23808 , y23809 , y23810 , y23811 , y23812 , y23813 , y23814 , y23815 , y23816 , y23817 , y23818 , y23819 , y23820 , y23821 , y23822 , y23823 , y23824 , y23825 , y23826 , y23827 , y23828 , y23829 , y23830 , y23831 , y23832 , y23833 , y23834 , y23835 , y23836 , y23837 , y23838 , y23839 , y23840 , y23841 , y23842 , y23843 , y23844 , y23845 , y23846 , y23847 , y23848 , y23849 , y23850 , y23851 , y23852 , y23853 , y23854 , y23855 , y23856 , y23857 , y23858 , y23859 , y23860 , y23861 , y23862 , y23863 , y23864 , y23865 , y23866 , y23867 , y23868 , y23869 , y23870 , y23871 , y23872 , y23873 , y23874 , y23875 , y23876 , y23877 , y23878 , y23879 , y23880 , y23881 , y23882 , y23883 , y23884 , y23885 , y23886 , y23887 , y23888 , y23889 , y23890 , y23891 , y23892 , y23893 , y23894 , y23895 , y23896 , y23897 , y23898 , y23899 , y23900 , y23901 , y23902 , y23903 , y23904 , y23905 , y23906 , y23907 , y23908 , y23909 , y23910 , y23911 , y23912 , y23913 , y23914 , y23915 , y23916 , y23917 , y23918 , y23919 , y23920 , y23921 , y23922 , y23923 , y23924 , y23925 , y23926 , y23927 , y23928 , y23929 , y23930 , y23931 , y23932 , y23933 , y23934 , y23935 , y23936 , y23937 , y23938 , y23939 , y23940 , y23941 , y23942 , y23943 , y23944 , y23945 , y23946 , y23947 , y23948 , y23949 , y23950 , y23951 , y23952 , y23953 , y23954 , y23955 , y23956 , y23957 , y23958 , y23959 , y23960 , y23961 , y23962 , y23963 , y23964 , y23965 , y23966 , y23967 , y23968 , y23969 , y23970 , y23971 , y23972 , y23973 , y23974 , y23975 , y23976 , y23977 , y23978 , y23979 , y23980 , y23981 , y23982 , y23983 , y23984 , y23985 , y23986 , y23987 , y23988 , y23989 , y23990 , y23991 , y23992 , y23993 , y23994 , y23995 , y23996 , y23997 , y23998 , y23999 , y24000 , y24001 , y24002 , y24003 , y24004 , y24005 , y24006 , y24007 , y24008 , y24009 , y24010 , y24011 , y24012 , y24013 , y24014 , y24015 , y24016 , y24017 , y24018 , y24019 , y24020 , y24021 , y24022 , y24023 , y24024 , y24025 , y24026 , y24027 , y24028 , y24029 , y24030 , y24031 , y24032 , y24033 , y24034 , y24035 , y24036 , y24037 , y24038 , y24039 , y24040 , y24041 , y24042 , y24043 , y24044 , y24045 , y24046 , y24047 , y24048 , y24049 , y24050 , y24051 , y24052 , y24053 , y24054 , y24055 , y24056 , y24057 , y24058 , y24059 , y24060 , y24061 , y24062 , y24063 , y24064 , y24065 , y24066 , y24067 , y24068 , y24069 , y24070 , y24071 , y24072 , y24073 , y24074 , y24075 , y24076 , y24077 , y24078 , y24079 , y24080 , y24081 , y24082 , y24083 , y24084 , y24085 , y24086 , y24087 , y24088 , y24089 , y24090 , y24091 , y24092 , y24093 , y24094 , y24095 , y24096 , y24097 , y24098 , y24099 , y24100 , y24101 , y24102 , y24103 , y24104 , y24105 , y24106 , y24107 , y24108 , y24109 , y24110 , y24111 , y24112 , y24113 , y24114 , y24115 , y24116 , y24117 , y24118 , y24119 , y24120 , y24121 , y24122 , y24123 , y24124 , y24125 , y24126 , y24127 , y24128 , y24129 , y24130 , y24131 , y24132 , y24133 , y24134 , y24135 , y24136 , y24137 , y24138 , y24139 , y24140 , y24141 , y24142 , y24143 , y24144 , y24145 , y24146 , y24147 , y24148 , y24149 , y24150 , y24151 , y24152 , y24153 , y24154 , y24155 , y24156 , y24157 , y24158 , y24159 , y24160 , y24161 , y24162 , y24163 , y24164 , y24165 , y24166 , y24167 , y24168 , y24169 , y24170 , y24171 , y24172 , y24173 , y24174 , y24175 , y24176 , y24177 , y24178 , y24179 , y24180 , y24181 , y24182 , y24183 , y24184 , y24185 , y24186 , y24187 , y24188 , y24189 , y24190 , y24191 , y24192 , y24193 , y24194 , y24195 , y24196 , y24197 , y24198 , y24199 , y24200 , y24201 , y24202 , y24203 , y24204 , y24205 , y24206 , y24207 , y24208 , y24209 , y24210 , y24211 , y24212 , y24213 , y24214 , y24215 , y24216 , y24217 , y24218 , y24219 , y24220 , y24221 , y24222 , y24223 , y24224 , y24225 , y24226 , y24227 , y24228 , y24229 , y24230 , y24231 , y24232 , y24233 , y24234 , y24235 , y24236 , y24237 , y24238 , y24239 , y24240 , y24241 , y24242 , y24243 , y24244 , y24245 , y24246 , y24247 , y24248 , y24249 , y24250 , y24251 , y24252 , y24253 , y24254 , y24255 , y24256 , y24257 , y24258 , y24259 , y24260 , y24261 , y24262 , y24263 , y24264 , y24265 , y24266 , y24267 , y24268 , y24269 , y24270 , y24271 , y24272 , y24273 , y24274 , y24275 , y24276 , y24277 , y24278 , y24279 , y24280 , y24281 , y24282 , y24283 , y24284 , y24285 , y24286 , y24287 , y24288 , y24289 , y24290 , y24291 , y24292 , y24293 , y24294 , y24295 , y24296 , y24297 , y24298 , y24299 , y24300 , y24301 , y24302 , y24303 , y24304 , y24305 , y24306 , y24307 , y24308 , y24309 , y24310 , y24311 , y24312 , y24313 , y24314 , y24315 , y24316 , y24317 , y24318 , y24319 , y24320 , y24321 , y24322 , y24323 , y24324 , y24325 , y24326 , y24327 , y24328 , y24329 , y24330 , y24331 , y24332 , y24333 , y24334 , y24335 , y24336 , y24337 , y24338 , y24339 , y24340 , y24341 , y24342 , y24343 , y24344 , y24345 , y24346 , y24347 , y24348 , y24349 , y24350 , y24351 , y24352 , y24353 , y24354 , y24355 , y24356 , y24357 , y24358 , y24359 , y24360 , y24361 , y24362 , y24363 , y24364 , y24365 , y24366 , y24367 , y24368 , y24369 , y24370 , y24371 , y24372 , y24373 , y24374 , y24375 , y24376 , y24377 , y24378 , y24379 , y24380 , y24381 , y24382 , y24383 , y24384 , y24385 , y24386 , y24387 , y24388 , y24389 , y24390 , y24391 , y24392 , y24393 , y24394 , y24395 , y24396 , y24397 , y24398 , y24399 , y24400 , y24401 , y24402 , y24403 , y24404 , y24405 , y24406 , y24407 , y24408 , y24409 , y24410 , y24411 , y24412 , y24413 , y24414 , y24415 , y24416 , y24417 , y24418 , y24419 , y24420 , y24421 , y24422 , y24423 , y24424 , y24425 , y24426 , y24427 , y24428 , y24429 , y24430 , y24431 , y24432 , y24433 , y24434 , y24435 , y24436 , y24437 , y24438 , y24439 , y24440 , y24441 , y24442 , y24443 , y24444 , y24445 , y24446 , y24447 , y24448 , y24449 , y24450 , y24451 , y24452 , y24453 , y24454 , y24455 , y24456 , y24457 , y24458 , y24459 , y24460 , y24461 , y24462 , y24463 , y24464 , y24465 , y24466 , y24467 , y24468 , y24469 , y24470 , y24471 , y24472 , y24473 , y24474 , y24475 , y24476 , y24477 , y24478 , y24479 , y24480 , y24481 , y24482 , y24483 , y24484 , y24485 , y24486 , y24487 , y24488 , y24489 , y24490 , y24491 , y24492 , y24493 , y24494 , y24495 , y24496 , y24497 , y24498 , y24499 , y24500 , y24501 , y24502 , y24503 , y24504 , y24505 , y24506 , y24507 , y24508 , y24509 , y24510 , y24511 , y24512 , y24513 , y24514 , y24515 , y24516 , y24517 , y24518 , y24519 , y24520 , y24521 , y24522 , y24523 , y24524 , y24525 , y24526 , y24527 , y24528 , y24529 , y24530 , y24531 , y24532 , y24533 , y24534 , y24535 , y24536 , y24537 , y24538 , y24539 , y24540 , y24541 , y24542 , y24543 , y24544 , y24545 , y24546 , y24547 , y24548 , y24549 , y24550 , y24551 , y24552 , y24553 , y24554 , y24555 , y24556 , y24557 , y24558 , y24559 , y24560 , y24561 , y24562 , y24563 , y24564 , y24565 , y24566 , y24567 , y24568 , y24569 , y24570 , y24571 , y24572 , y24573 , y24574 , y24575 , y24576 , y24577 , y24578 , y24579 , y24580 , y24581 , y24582 , y24583 , y24584 , y24585 , y24586 , y24587 , y24588 , y24589 , y24590 , y24591 , y24592 , y24593 , y24594 , y24595 , y24596 , y24597 , y24598 , y24599 , y24600 , y24601 , y24602 , y24603 , y24604 , y24605 , y24606 , y24607 , y24608 , y24609 , y24610 , y24611 , y24612 , y24613 , y24614 , y24615 , y24616 , y24617 , y24618 , y24619 , y24620 , y24621 , y24622 , y24623 , y24624 , y24625 , y24626 , y24627 , y24628 , y24629 , y24630 , y24631 , y24632 , y24633 , y24634 , y24635 , y24636 , y24637 , y24638 , y24639 , y24640 , y24641 , y24642 , y24643 , y24644 , y24645 , y24646 , y24647 , y24648 , y24649 , y24650 , y24651 , y24652 , y24653 , y24654 , y24655 , y24656 , y24657 , y24658 , y24659 , y24660 , y24661 , y24662 , y24663 , y24664 , y24665 , y24666 , y24667 , y24668 , y24669 , y24670 , y24671 , y24672 , y24673 , y24674 , y24675 , y24676 , y24677 , y24678 , y24679 , y24680 , y24681 , y24682 , y24683 , y24684 , y24685 , y24686 , y24687 , y24688 , y24689 , y24690 , y24691 , y24692 , y24693 , y24694 , y24695 , y24696 , y24697 , y24698 , y24699 , y24700 , y24701 , y24702 , y24703 , y24704 , y24705 , y24706 , y24707 , y24708 , y24709 , y24710 , y24711 , y24712 , y24713 , y24714 , y24715 , y24716 , y24717 , y24718 , y24719 , y24720 , y24721 , y24722 , y24723 , y24724 , y24725 , y24726 , y24727 , y24728 , y24729 , y24730 , y24731 , y24732 , y24733 , y24734 , y24735 , y24736 , y24737 , y24738 , y24739 , y24740 , y24741 , y24742 , y24743 , y24744 , y24745 , y24746 , y24747 , y24748 , y24749 , y24750 , y24751 , y24752 , y24753 , y24754 , y24755 , y24756 , y24757 , y24758 , y24759 , y24760 , y24761 , y24762 , y24763 , y24764 , y24765 , y24766 , y24767 , y24768 , y24769 , y24770 , y24771 , y24772 , y24773 , y24774 , y24775 , y24776 , y24777 , y24778 , y24779 , y24780 , y24781 , y24782 , y24783 , y24784 , y24785 , y24786 , y24787 , y24788 , y24789 , y24790 , y24791 , y24792 , y24793 , y24794 , y24795 , y24796 , y24797 , y24798 , y24799 , y24800 , y24801 , y24802 , y24803 , y24804 , y24805 , y24806 , y24807 , y24808 , y24809 , y24810 , y24811 , y24812 , y24813 , y24814 , y24815 , y24816 , y24817 , y24818 , y24819 , y24820 , y24821 , y24822 , y24823 , y24824 , y24825 , y24826 , y24827 , y24828 , y24829 , y24830 , y24831 , y24832 , y24833 , y24834 , y24835 , y24836 , y24837 , y24838 , y24839 , y24840 , y24841 , y24842 , y24843 , y24844 , y24845 , y24846 , y24847 , y24848 , y24849 , y24850 , y24851 , y24852 , y24853 , y24854 , y24855 , y24856 , y24857 , y24858 , y24859 , y24860 , y24861 , y24862 , y24863 , y24864 , y24865 , y24866 , y24867 , y24868 , y24869 , y24870 , y24871 , y24872 , y24873 , y24874 , y24875 , y24876 , y24877 , y24878 , y24879 , y24880 , y24881 , y24882 , y24883 , y24884 , y24885 , y24886 , y24887 , y24888 , y24889 , y24890 , y24891 , y24892 , y24893 , y24894 , y24895 , y24896 , y24897 , y24898 , y24899 , y24900 , y24901 , y24902 , y24903 , y24904 , y24905 , y24906 , y24907 , y24908 , y24909 , y24910 , y24911 , y24912 , y24913 , y24914 , y24915 , y24916 , y24917 , y24918 , y24919 , y24920 , y24921 , y24922 , y24923 , y24924 , y24925 , y24926 , y24927 , y24928 , y24929 , y24930 , y24931 , y24932 , y24933 , y24934 , y24935 , y24936 , y24937 , y24938 , y24939 , y24940 , y24941 , y24942 , y24943 , y24944 , y24945 , y24946 , y24947 , y24948 , y24949 , y24950 , y24951 , y24952 , y24953 , y24954 , y24955 , y24956 , y24957 , y24958 , y24959 , y24960 , y24961 , y24962 , y24963 , y24964 , y24965 , y24966 , y24967 , y24968 , y24969 , y24970 , y24971 , y24972 , y24973 , y24974 , y24975 , y24976 , y24977 , y24978 , y24979 , y24980 , y24981 , y24982 , y24983 , y24984 , y24985 , y24986 , y24987 , y24988 , y24989 , y24990 , y24991 , y24992 , y24993 , y24994 , y24995 , y24996 , y24997 , y24998 , y24999 , y25000 , y25001 , y25002 , y25003 , y25004 , y25005 , y25006 , y25007 , y25008 , y25009 , y25010 , y25011 , y25012 , y25013 , y25014 , y25015 , y25016 , y25017 , y25018 , y25019 , y25020 , y25021 , y25022 , y25023 , y25024 , y25025 , y25026 , y25027 , y25028 , y25029 , y25030 , y25031 , y25032 , y25033 , y25034 , y25035 , y25036 , y25037 , y25038 , y25039 , y25040 , y25041 , y25042 , y25043 , y25044 , y25045 , y25046 , y25047 , y25048 , y25049 , y25050 , y25051 , y25052 , y25053 , y25054 , y25055 , y25056 , y25057 , y25058 , y25059 , y25060 , y25061 , y25062 , y25063 , y25064 , y25065 , y25066 , y25067 , y25068 , y25069 , y25070 , y25071 , y25072 , y25073 , y25074 , y25075 , y25076 , y25077 , y25078 , y25079 , y25080 , y25081 , y25082 , y25083 , y25084 , y25085 , y25086 , y25087 , y25088 , y25089 , y25090 , y25091 , y25092 , y25093 , y25094 , y25095 , y25096 , y25097 , y25098 , y25099 , y25100 , y25101 , y25102 , y25103 , y25104 , y25105 , y25106 , y25107 , y25108 , y25109 , y25110 , y25111 , y25112 , y25113 , y25114 , y25115 , y25116 , y25117 , y25118 , y25119 , y25120 , y25121 , y25122 , y25123 , y25124 , y25125 , y25126 , y25127 , y25128 , y25129 , y25130 , y25131 , y25132 , y25133 , y25134 , y25135 , y25136 , y25137 , y25138 , y25139 , y25140 , y25141 , y25142 , y25143 , y25144 , y25145 , y25146 , y25147 , y25148 , y25149 , y25150 , y25151 , y25152 , y25153 , y25154 , y25155 , y25156 , y25157 , y25158 , y25159 , y25160 , y25161 , y25162 , y25163 , y25164 , y25165 , y25166 , y25167 , y25168 , y25169 , y25170 , y25171 , y25172 , y25173 , y25174 , y25175 , y25176 , y25177 , y25178 , y25179 , y25180 , y25181 , y25182 , y25183 , y25184 , y25185 , y25186 , y25187 , y25188 , y25189 , y25190 , y25191 , y25192 , y25193 , y25194 , y25195 , y25196 , y25197 , y25198 , y25199 , y25200 , y25201 , y25202 , y25203 , y25204 , y25205 , y25206 , y25207 , y25208 , y25209 , y25210 , y25211 , y25212 , y25213 , y25214 , y25215 , y25216 , y25217 , y25218 , y25219 , y25220 , y25221 , y25222 , y25223 , y25224 , y25225 , y25226 , y25227 , y25228 , y25229 , y25230 , y25231 , y25232 , y25233 , y25234 , y25235 , y25236 , y25237 , y25238 , y25239 , y25240 , y25241 , y25242 , y25243 , y25244 , y25245 , y25246 , y25247 , y25248 , y25249 , y25250 , y25251 , y25252 , y25253 , y25254 , y25255 , y25256 , y25257 , y25258 , y25259 , y25260 , y25261 , y25262 , y25263 , y25264 , y25265 , y25266 , y25267 , y25268 , y25269 , y25270 , y25271 , y25272 , y25273 , y25274 , y25275 , y25276 , y25277 , y25278 , y25279 , y25280 , y25281 , y25282 , y25283 , y25284 , y25285 , y25286 , y25287 , y25288 , y25289 , y25290 , y25291 , y25292 , y25293 , y25294 , y25295 , y25296 , y25297 , y25298 , y25299 , y25300 , y25301 , y25302 , y25303 , y25304 , y25305 , y25306 , y25307 , y25308 , y25309 , y25310 , y25311 , y25312 , y25313 , y25314 , y25315 , y25316 , y25317 , y25318 , y25319 , y25320 , y25321 , y25322 , y25323 , y25324 , y25325 , y25326 , y25327 , y25328 , y25329 , y25330 , y25331 , y25332 , y25333 , y25334 , y25335 , y25336 , y25337 , y25338 , y25339 , y25340 , y25341 , y25342 , y25343 , y25344 , y25345 , y25346 , y25347 , y25348 , y25349 , y25350 , y25351 , y25352 , y25353 , y25354 , y25355 , y25356 , y25357 , y25358 , y25359 , y25360 , y25361 , y25362 , y25363 , y25364 , y25365 , y25366 , y25367 , y25368 , y25369 , y25370 , y25371 , y25372 , y25373 , y25374 , y25375 , y25376 , y25377 , y25378 , y25379 , y25380 , y25381 , y25382 , y25383 , y25384 , y25385 , y25386 , y25387 , y25388 , y25389 , y25390 , y25391 , y25392 , y25393 , y25394 , y25395 , y25396 , y25397 , y25398 , y25399 , y25400 , y25401 , y25402 , y25403 , y25404 , y25405 , y25406 , y25407 , y25408 , y25409 , y25410 , y25411 , y25412 , y25413 , y25414 , y25415 , y25416 , y25417 , y25418 , y25419 , y25420 , y25421 , y25422 , y25423 , y25424 , y25425 , y25426 , y25427 , y25428 , y25429 , y25430 , y25431 , y25432 , y25433 , y25434 , y25435 , y25436 , y25437 , y25438 , y25439 , y25440 , y25441 , y25442 , y25443 , y25444 , y25445 , y25446 , y25447 , y25448 , y25449 , y25450 , y25451 , y25452 , y25453 , y25454 , y25455 , y25456 , y25457 , y25458 , y25459 , y25460 , y25461 , y25462 , y25463 , y25464 , y25465 , y25466 , y25467 , y25468 , y25469 , y25470 , y25471 , y25472 , y25473 , y25474 , y25475 , y25476 , y25477 , y25478 , y25479 , y25480 , y25481 , y25482 , y25483 , y25484 , y25485 , y25486 , y25487 , y25488 , y25489 , y25490 , y25491 , y25492 , y25493 , y25494 , y25495 , y25496 , y25497 , y25498 , y25499 , y25500 , y25501 , y25502 , y25503 , y25504 , y25505 , y25506 , y25507 , y25508 , y25509 , y25510 , y25511 , y25512 , y25513 , y25514 , y25515 , y25516 , y25517 , y25518 , y25519 , y25520 , y25521 , y25522 , y25523 , y25524 , y25525 , y25526 , y25527 , y25528 , y25529 , y25530 , y25531 , y25532 , y25533 , y25534 , y25535 , y25536 , y25537 , y25538 , y25539 , y25540 , y25541 , y25542 , y25543 , y25544 , y25545 , y25546 , y25547 , y25548 , y25549 , y25550 , y25551 , y25552 , y25553 , y25554 , y25555 , y25556 , y25557 , y25558 , y25559 , y25560 , y25561 , y25562 , y25563 , y25564 , y25565 , y25566 , y25567 , y25568 , y25569 , y25570 , y25571 , y25572 , y25573 , y25574 , y25575 , y25576 , y25577 , y25578 , y25579 , y25580 , y25581 , y25582 , y25583 , y25584 , y25585 , y25586 , y25587 , y25588 , y25589 , y25590 , y25591 , y25592 , y25593 , y25594 , y25595 , y25596 , y25597 , y25598 , y25599 , y25600 , y25601 , y25602 , y25603 , y25604 , y25605 , y25606 , y25607 , y25608 , y25609 , y25610 , y25611 , y25612 , y25613 , y25614 , y25615 , y25616 , y25617 , y25618 , y25619 , y25620 , y25621 , y25622 , y25623 , y25624 , y25625 , y25626 , y25627 , y25628 , y25629 , y25630 , y25631 , y25632 , y25633 , y25634 , y25635 , y25636 , y25637 , y25638 , y25639 , y25640 , y25641 , y25642 , y25643 , y25644 , y25645 , y25646 , y25647 , y25648 , y25649 , y25650 , y25651 , y25652 , y25653 , y25654 , y25655 , y25656 , y25657 , y25658 , y25659 , y25660 , y25661 , y25662 , y25663 , y25664 , y25665 , y25666 , y25667 , y25668 , y25669 , y25670 , y25671 , y25672 , y25673 , y25674 , y25675 , y25676 , y25677 , y25678 , y25679 , y25680 , y25681 , y25682 , y25683 , y25684 , y25685 , y25686 , y25687 , y25688 , y25689 , y25690 , y25691 , y25692 , y25693 , y25694 , y25695 , y25696 , y25697 , y25698 , y25699 , y25700 , y25701 , y25702 , y25703 , y25704 , y25705 , y25706 , y25707 , y25708 , y25709 , y25710 , y25711 , y25712 , y25713 , y25714 , y25715 , y25716 , y25717 , y25718 , y25719 , y25720 , y25721 , y25722 , y25723 , y25724 , y25725 , y25726 , y25727 , y25728 , y25729 , y25730 , y25731 , y25732 , y25733 , y25734 , y25735 , y25736 , y25737 , y25738 , y25739 , y25740 , y25741 , y25742 , y25743 , y25744 , y25745 , y25746 , y25747 , y25748 , y25749 , y25750 , y25751 , y25752 , y25753 , y25754 , y25755 , y25756 , y25757 , y25758 , y25759 , y25760 , y25761 , y25762 , y25763 , y25764 , y25765 , y25766 , y25767 , y25768 , y25769 , y25770 , y25771 , y25772 , y25773 , y25774 , y25775 , y25776 , y25777 , y25778 , y25779 , y25780 , y25781 , y25782 , y25783 , y25784 , y25785 , y25786 , y25787 , y25788 , y25789 , y25790 , y25791 , y25792 , y25793 , y25794 , y25795 , y25796 , y25797 , y25798 , y25799 , y25800 , y25801 , y25802 , y25803 , y25804 , y25805 , y25806 , y25807 , y25808 , y25809 , y25810 , y25811 , y25812 , y25813 , y25814 , y25815 , y25816 , y25817 , y25818 , y25819 , y25820 , y25821 , y25822 , y25823 , y25824 , y25825 , y25826 , y25827 , y25828 , y25829 , y25830 , y25831 , y25832 , y25833 , y25834 , y25835 , y25836 , y25837 , y25838 , y25839 , y25840 , y25841 , y25842 , y25843 , y25844 , y25845 , y25846 , y25847 , y25848 , y25849 , y25850 , y25851 , y25852 , y25853 , y25854 , y25855 , y25856 , y25857 , y25858 , y25859 , y25860 , y25861 , y25862 , y25863 , y25864 , y25865 , y25866 , y25867 , y25868 , y25869 , y25870 , y25871 , y25872 , y25873 , y25874 , y25875 , y25876 , y25877 , y25878 , y25879 , y25880 , y25881 , y25882 , y25883 , y25884 , y25885 , y25886 , y25887 , y25888 , y25889 , y25890 , y25891 , y25892 , y25893 , y25894 , y25895 , y25896 , y25897 , y25898 , y25899 , y25900 , y25901 , y25902 , y25903 , y25904 , y25905 , y25906 , y25907 , y25908 , y25909 , y25910 , y25911 , y25912 , y25913 , y25914 , y25915 , y25916 , y25917 , y25918 , y25919 , y25920 , y25921 , y25922 , y25923 , y25924 , y25925 , y25926 , y25927 , y25928 , y25929 , y25930 , y25931 , y25932 , y25933 , y25934 , y25935 , y25936 , y25937 , y25938 , y25939 , y25940 , y25941 , y25942 , y25943 , y25944 , y25945 , y25946 , y25947 , y25948 , y25949 , y25950 , y25951 , y25952 , y25953 , y25954 , y25955 , y25956 , y25957 , y25958 , y25959 , y25960 , y25961 , y25962 , y25963 , y25964 , y25965 , y25966 , y25967 , y25968 , y25969 , y25970 , y25971 , y25972 , y25973 , y25974 , y25975 , y25976 , y25977 , y25978 , y25979 , y25980 , y25981 , y25982 , y25983 , y25984 , y25985 , y25986 , y25987 , y25988 , y25989 , y25990 , y25991 , y25992 , y25993 , y25994 , y25995 , y25996 , y25997 , y25998 , y25999 , y26000 , y26001 , y26002 , y26003 , y26004 , y26005 , y26006 , y26007 , y26008 , y26009 , y26010 , y26011 , y26012 , y26013 , y26014 , y26015 , y26016 , y26017 , y26018 , y26019 , y26020 , y26021 , y26022 , y26023 , y26024 , y26025 , y26026 , y26027 , y26028 , y26029 , y26030 , y26031 , y26032 , y26033 , y26034 , y26035 , y26036 , y26037 , y26038 , y26039 , y26040 , y26041 , y26042 , y26043 , y26044 , y26045 , y26046 , y26047 , y26048 , y26049 , y26050 , y26051 , y26052 , y26053 , y26054 , y26055 , y26056 , y26057 , y26058 , y26059 , y26060 , y26061 , y26062 , y26063 , y26064 , y26065 , y26066 , y26067 , y26068 , y26069 , y26070 , y26071 , y26072 , y26073 , y26074 , y26075 , y26076 , y26077 , y26078 , y26079 , y26080 , y26081 , y26082 , y26083 , y26084 , y26085 , y26086 , y26087 , y26088 , y26089 , y26090 , y26091 , y26092 , y26093 , y26094 , y26095 , y26096 , y26097 , y26098 , y26099 , y26100 , y26101 , y26102 , y26103 , y26104 , y26105 , y26106 , y26107 , y26108 , y26109 , y26110 , y26111 , y26112 , y26113 , y26114 , y26115 , y26116 , y26117 , y26118 , y26119 , y26120 , y26121 , y26122 , y26123 , y26124 , y26125 , y26126 , y26127 , y26128 , y26129 , y26130 , y26131 , y26132 , y26133 , y26134 , y26135 , y26136 , y26137 , y26138 , y26139 , y26140 , y26141 , y26142 , y26143 , y26144 , y26145 , y26146 , y26147 , y26148 , y26149 , y26150 , y26151 , y26152 , y26153 , y26154 , y26155 , y26156 , y26157 , y26158 , y26159 , y26160 , y26161 , y26162 , y26163 , y26164 , y26165 , y26166 , y26167 , y26168 , y26169 , y26170 , y26171 , y26172 , y26173 , y26174 , y26175 , y26176 , y26177 , y26178 , y26179 , y26180 , y26181 , y26182 , y26183 , y26184 , y26185 , y26186 , y26187 , y26188 , y26189 , y26190 , y26191 , y26192 , y26193 , y26194 , y26195 , y26196 , y26197 , y26198 , y26199 , y26200 , y26201 , y26202 , y26203 , y26204 , y26205 , y26206 , y26207 , y26208 , y26209 , y26210 , y26211 , y26212 , y26213 , y26214 , y26215 , y26216 , y26217 , y26218 , y26219 , y26220 , y26221 , y26222 , y26223 , y26224 , y26225 , y26226 , y26227 , y26228 , y26229 , y26230 , y26231 , y26232 , y26233 , y26234 , y26235 , y26236 , y26237 , y26238 , y26239 , y26240 , y26241 , y26242 , y26243 , y26244 , y26245 , y26246 , y26247 , y26248 , y26249 , y26250 , y26251 , y26252 , y26253 , y26254 , y26255 , y26256 , y26257 , y26258 , y26259 , y26260 , y26261 , y26262 , y26263 , y26264 , y26265 , y26266 , y26267 , y26268 , y26269 , y26270 , y26271 , y26272 , y26273 , y26274 , y26275 , y26276 , y26277 , y26278 , y26279 , y26280 , y26281 , y26282 , y26283 , y26284 , y26285 , y26286 , y26287 , y26288 , y26289 , y26290 , y26291 , y26292 , y26293 , y26294 , y26295 , y26296 , y26297 , y26298 , y26299 , y26300 , y26301 , y26302 , y26303 , y26304 , y26305 , y26306 , y26307 , y26308 , y26309 , y26310 , y26311 , y26312 , y26313 , y26314 , y26315 , y26316 , y26317 , y26318 , y26319 , y26320 , y26321 , y26322 , y26323 , y26324 , y26325 , y26326 , y26327 , y26328 , y26329 , y26330 , y26331 , y26332 , y26333 , y26334 , y26335 , y26336 , y26337 , y26338 , y26339 , y26340 , y26341 , y26342 , y26343 , y26344 , y26345 , y26346 , y26347 , y26348 , y26349 , y26350 , y26351 , y26352 , y26353 , y26354 , y26355 , y26356 , y26357 , y26358 , y26359 , y26360 , y26361 , y26362 , y26363 , y26364 , y26365 , y26366 , y26367 , y26368 , y26369 , y26370 , y26371 , y26372 , y26373 , y26374 , y26375 , y26376 , y26377 , y26378 , y26379 , y26380 , y26381 , y26382 , y26383 , y26384 , y26385 , y26386 , y26387 , y26388 , y26389 , y26390 , y26391 , y26392 , y26393 , y26394 , y26395 , y26396 , y26397 , y26398 , y26399 , y26400 , y26401 , y26402 , y26403 , y26404 , y26405 , y26406 , y26407 , y26408 , y26409 , y26410 , y26411 , y26412 , y26413 , y26414 , y26415 , y26416 , y26417 , y26418 , y26419 , y26420 , y26421 , y26422 , y26423 , y26424 , y26425 , y26426 , y26427 , y26428 , y26429 , y26430 , y26431 , y26432 , y26433 , y26434 , y26435 , y26436 , y26437 , y26438 , y26439 , y26440 , y26441 , y26442 , y26443 , y26444 , y26445 , y26446 , y26447 , y26448 , y26449 , y26450 , y26451 , y26452 , y26453 , y26454 , y26455 , y26456 , y26457 , y26458 , y26459 , y26460 , y26461 , y26462 , y26463 , y26464 , y26465 , y26466 , y26467 , y26468 , y26469 , y26470 , y26471 , y26472 , y26473 , y26474 , y26475 , y26476 , y26477 , y26478 , y26479 , y26480 , y26481 , y26482 , y26483 , y26484 , y26485 , y26486 , y26487 , y26488 , y26489 , y26490 , y26491 , y26492 , y26493 , y26494 , y26495 , y26496 , y26497 , y26498 , y26499 , y26500 , y26501 , y26502 , y26503 , y26504 , y26505 , y26506 , y26507 , y26508 , y26509 , y26510 , y26511 , y26512 , y26513 , y26514 , y26515 , y26516 , y26517 , y26518 , y26519 , y26520 , y26521 , y26522 , y26523 , y26524 , y26525 , y26526 , y26527 , y26528 , y26529 , y26530 , y26531 , y26532 , y26533 , y26534 , y26535 , y26536 , y26537 , y26538 , y26539 , y26540 , y26541 , y26542 , y26543 , y26544 , y26545 , y26546 , y26547 , y26548 , y26549 , y26550 , y26551 , y26552 , y26553 , y26554 , y26555 , y26556 , y26557 , y26558 , y26559 , y26560 , y26561 , y26562 , y26563 , y26564 , y26565 , y26566 , y26567 , y26568 , y26569 , y26570 , y26571 , y26572 , y26573 , y26574 , y26575 , y26576 , y26577 , y26578 , y26579 , y26580 , y26581 , y26582 , y26583 , y26584 , y26585 , y26586 , y26587 , y26588 , y26589 , y26590 , y26591 , y26592 , y26593 , y26594 , y26595 , y26596 , y26597 , y26598 , y26599 , y26600 , y26601 , y26602 , y26603 , y26604 , y26605 , y26606 , y26607 , y26608 , y26609 , y26610 , y26611 , y26612 , y26613 , y26614 , y26615 , y26616 , y26617 , y26618 , y26619 , y26620 , y26621 , y26622 , y26623 , y26624 , y26625 , y26626 , y26627 , y26628 , y26629 , y26630 , y26631 , y26632 , y26633 , y26634 , y26635 , y26636 , y26637 , y26638 , y26639 , y26640 , y26641 , y26642 , y26643 , y26644 , y26645 , y26646 , y26647 , y26648 , y26649 , y26650 , y26651 , y26652 , y26653 , y26654 , y26655 , y26656 , y26657 , y26658 , y26659 , y26660 , y26661 , y26662 , y26663 , y26664 , y26665 , y26666 , y26667 , y26668 , y26669 , y26670 , y26671 , y26672 , y26673 , y26674 , y26675 , y26676 , y26677 , y26678 , y26679 , y26680 , y26681 , y26682 , y26683 , y26684 , y26685 , y26686 , y26687 , y26688 , y26689 , y26690 , y26691 , y26692 , y26693 , y26694 , y26695 , y26696 , y26697 , y26698 , y26699 , y26700 , y26701 , y26702 , y26703 , y26704 , y26705 , y26706 , y26707 , y26708 , y26709 , y26710 , y26711 , y26712 , y26713 , y26714 , y26715 , y26716 , y26717 , y26718 , y26719 , y26720 , y26721 , y26722 , y26723 , y26724 , y26725 , y26726 , y26727 , y26728 , y26729 , y26730 , y26731 , y26732 , y26733 , y26734 , y26735 , y26736 , y26737 , y26738 , y26739 , y26740 , y26741 , y26742 , y26743 , y26744 , y26745 , y26746 , y26747 , y26748 , y26749 , y26750 , y26751 , y26752 , y26753 , y26754 , y26755 , y26756 , y26757 , y26758 , y26759 , y26760 , y26761 , y26762 , y26763 , y26764 , y26765 , y26766 , y26767 , y26768 , y26769 , y26770 , y26771 , y26772 , y26773 , y26774 , y26775 , y26776 , y26777 , y26778 , y26779 , y26780 , y26781 , y26782 , y26783 , y26784 , y26785 , y26786 , y26787 , y26788 , y26789 , y26790 , y26791 , y26792 , y26793 , y26794 , y26795 , y26796 , y26797 , y26798 , y26799 , y26800 , y26801 , y26802 , y26803 , y26804 , y26805 , y26806 , y26807 , y26808 , y26809 , y26810 , y26811 , y26812 , y26813 , y26814 , y26815 , y26816 , y26817 , y26818 , y26819 , y26820 , y26821 , y26822 , y26823 , y26824 , y26825 , y26826 , y26827 , y26828 , y26829 , y26830 , y26831 , y26832 , y26833 , y26834 , y26835 , y26836 , y26837 , y26838 , y26839 , y26840 , y26841 , y26842 , y26843 , y26844 , y26845 , y26846 , y26847 , y26848 , y26849 , y26850 , y26851 , y26852 , y26853 , y26854 , y26855 , y26856 , y26857 , y26858 , y26859 , y26860 , y26861 , y26862 , y26863 , y26864 , y26865 , y26866 , y26867 , y26868 , y26869 , y26870 , y26871 , y26872 , y26873 , y26874 , y26875 , y26876 , y26877 , y26878 , y26879 , y26880 , y26881 , y26882 , y26883 , y26884 , y26885 , y26886 , y26887 , y26888 , y26889 , y26890 , y26891 , y26892 , y26893 , y26894 , y26895 , y26896 , y26897 , y26898 , y26899 , y26900 , y26901 , y26902 , y26903 , y26904 , y26905 , y26906 , y26907 , y26908 , y26909 , y26910 , y26911 , y26912 , y26913 , y26914 , y26915 , y26916 , y26917 , y26918 , y26919 , y26920 , y26921 , y26922 , y26923 , y26924 , y26925 , y26926 , y26927 , y26928 , y26929 , y26930 , y26931 , y26932 , y26933 , y26934 , y26935 , y26936 , y26937 , y26938 , y26939 , y26940 , y26941 , y26942 , y26943 , y26944 , y26945 , y26946 , y26947 , y26948 , y26949 , y26950 , y26951 , y26952 , y26953 , y26954 , y26955 , y26956 , y26957 , y26958 , y26959 , y26960 , y26961 , y26962 , y26963 , y26964 , y26965 , y26966 , y26967 , y26968 , y26969 , y26970 , y26971 , y26972 , y26973 , y26974 , y26975 , y26976 , y26977 , y26978 , y26979 , y26980 , y26981 , y26982 , y26983 , y26984 , y26985 , y26986 , y26987 , y26988 , y26989 , y26990 , y26991 , y26992 , y26993 , y26994 , y26995 , y26996 , y26997 , y26998 , y26999 , y27000 , y27001 , y27002 , y27003 , y27004 , y27005 , y27006 , y27007 , y27008 , y27009 , y27010 , y27011 , y27012 , y27013 , y27014 , y27015 , y27016 , y27017 , y27018 , y27019 , y27020 , y27021 , y27022 , y27023 , y27024 , y27025 , y27026 , y27027 , y27028 , y27029 , y27030 , y27031 , y27032 , y27033 , y27034 , y27035 , y27036 , y27037 , y27038 , y27039 , y27040 , y27041 , y27042 , y27043 , y27044 , y27045 , y27046 , y27047 , y27048 , y27049 , y27050 , y27051 , y27052 , y27053 , y27054 , y27055 , y27056 , y27057 , y27058 , y27059 , y27060 , y27061 , y27062 , y27063 , y27064 , y27065 , y27066 , y27067 , y27068 , y27069 , y27070 , y27071 , y27072 , y27073 , y27074 , y27075 , y27076 , y27077 , y27078 , y27079 , y27080 , y27081 , y27082 , y27083 , y27084 , y27085 , y27086 , y27087 , y27088 , y27089 , y27090 , y27091 , y27092 , y27093 , y27094 , y27095 , y27096 , y27097 , y27098 , y27099 , y27100 , y27101 , y27102 , y27103 , y27104 , y27105 , y27106 , y27107 , y27108 , y27109 , y27110 , y27111 , y27112 , y27113 , y27114 , y27115 , y27116 , y27117 , y27118 , y27119 , y27120 , y27121 , y27122 , y27123 , y27124 , y27125 , y27126 , y27127 , y27128 , y27129 , y27130 , y27131 , y27132 , y27133 , y27134 , y27135 , y27136 , y27137 , y27138 , y27139 , y27140 , y27141 , y27142 , y27143 , y27144 , y27145 , y27146 , y27147 , y27148 , y27149 , y27150 , y27151 , y27152 , y27153 , y27154 , y27155 , y27156 , y27157 , y27158 , y27159 , y27160 , y27161 , y27162 , y27163 , y27164 , y27165 , y27166 , y27167 , y27168 , y27169 , y27170 , y27171 , y27172 , y27173 , y27174 , y27175 , y27176 , y27177 , y27178 , y27179 , y27180 , y27181 , y27182 , y27183 , y27184 , y27185 , y27186 , y27187 , y27188 , y27189 , y27190 , y27191 , y27192 , y27193 , y27194 , y27195 , y27196 , y27197 , y27198 , y27199 , y27200 , y27201 , y27202 , y27203 , y27204 , y27205 , y27206 , y27207 , y27208 , y27209 , y27210 , y27211 , y27212 , y27213 , y27214 , y27215 , y27216 , y27217 , y27218 , y27219 , y27220 , y27221 , y27222 , y27223 , y27224 , y27225 , y27226 , y27227 , y27228 , y27229 , y27230 , y27231 , y27232 , y27233 , y27234 , y27235 , y27236 , y27237 , y27238 , y27239 , y27240 , y27241 , y27242 , y27243 , y27244 , y27245 , y27246 , y27247 , y27248 , y27249 , y27250 , y27251 , y27252 , y27253 , y27254 , y27255 , y27256 , y27257 , y27258 , y27259 , y27260 , y27261 , y27262 , y27263 , y27264 , y27265 , y27266 , y27267 , y27268 , y27269 , y27270 , y27271 , y27272 , y27273 , y27274 , y27275 , y27276 , y27277 , y27278 , y27279 , y27280 , y27281 , y27282 , y27283 , y27284 , y27285 , y27286 , y27287 , y27288 , y27289 , y27290 , y27291 , y27292 , y27293 , y27294 , y27295 , y27296 , y27297 , y27298 , y27299 , y27300 , y27301 , y27302 , y27303 , y27304 , y27305 , y27306 , y27307 , y27308 , y27309 , y27310 , y27311 , y27312 , y27313 , y27314 , y27315 , y27316 , y27317 , y27318 , y27319 , y27320 , y27321 , y27322 , y27323 , y27324 , y27325 , y27326 , y27327 , y27328 , y27329 , y27330 , y27331 , y27332 , y27333 , y27334 , y27335 , y27336 , y27337 , y27338 , y27339 , y27340 , y27341 , y27342 , y27343 , y27344 , y27345 , y27346 , y27347 , y27348 , y27349 , y27350 , y27351 , y27352 , y27353 , y27354 , y27355 , y27356 , y27357 , y27358 , y27359 , y27360 , y27361 , y27362 , y27363 , y27364 , y27365 , y27366 , y27367 , y27368 , y27369 , y27370 , y27371 , y27372 , y27373 , y27374 , y27375 , y27376 , y27377 , y27378 , y27379 , y27380 , y27381 , y27382 , y27383 , y27384 , y27385 , y27386 , y27387 , y27388 , y27389 , y27390 , y27391 , y27392 , y27393 , y27394 , y27395 , y27396 , y27397 , y27398 , y27399 , y27400 , y27401 , y27402 , y27403 , y27404 , y27405 , y27406 , y27407 , y27408 , y27409 , y27410 , y27411 , y27412 , y27413 , y27414 , y27415 , y27416 , y27417 , y27418 , y27419 , y27420 , y27421 , y27422 , y27423 , y27424 , y27425 , y27426 , y27427 , y27428 , y27429 , y27430 , y27431 , y27432 , y27433 , y27434 , y27435 , y27436 , y27437 , y27438 , y27439 , y27440 , y27441 , y27442 , y27443 , y27444 , y27445 , y27446 , y27447 , y27448 , y27449 , y27450 , y27451 , y27452 , y27453 , y27454 , y27455 , y27456 , y27457 , y27458 , y27459 , y27460 , y27461 , y27462 , y27463 , y27464 , y27465 , y27466 , y27467 , y27468 , y27469 , y27470 , y27471 , y27472 , y27473 , y27474 , y27475 , y27476 , y27477 , y27478 , y27479 , y27480 , y27481 , y27482 , y27483 , y27484 , y27485 , y27486 , y27487 , y27488 , y27489 , y27490 , y27491 , y27492 , y27493 , y27494 , y27495 , y27496 , y27497 , y27498 , y27499 , y27500 , y27501 , y27502 , y27503 , y27504 , y27505 , y27506 , y27507 , y27508 , y27509 , y27510 , y27511 , y27512 , y27513 , y27514 , y27515 , y27516 , y27517 , y27518 , y27519 , y27520 , y27521 , y27522 , y27523 , y27524 , y27525 , y27526 , y27527 , y27528 , y27529 , y27530 , y27531 , y27532 , y27533 , y27534 , y27535 , y27536 , y27537 , y27538 , y27539 , y27540 , y27541 , y27542 , y27543 , y27544 , y27545 , y27546 , y27547 , y27548 , y27549 , y27550 , y27551 , y27552 , y27553 , y27554 , y27555 , y27556 , y27557 , y27558 , y27559 , y27560 , y27561 , y27562 , y27563 , y27564 , y27565 , y27566 , y27567 , y27568 , y27569 , y27570 , y27571 , y27572 , y27573 , y27574 , y27575 , y27576 , y27577 , y27578 , y27579 , y27580 , y27581 , y27582 , y27583 , y27584 , y27585 , y27586 , y27587 , y27588 , y27589 , y27590 , y27591 , y27592 , y27593 , y27594 , y27595 , y27596 , y27597 , y27598 , y27599 , y27600 , y27601 , y27602 , y27603 , y27604 , y27605 , y27606 , y27607 , y27608 , y27609 , y27610 , y27611 , y27612 , y27613 , y27614 , y27615 , y27616 , y27617 , y27618 , y27619 , y27620 , y27621 , y27622 , y27623 , y27624 , y27625 , y27626 , y27627 , y27628 , y27629 , y27630 , y27631 , y27632 , y27633 , y27634 , y27635 , y27636 , y27637 , y27638 , y27639 , y27640 , y27641 , y27642 , y27643 , y27644 , y27645 , y27646 , y27647 , y27648 , y27649 , y27650 , y27651 , y27652 , y27653 , y27654 , y27655 , y27656 , y27657 , y27658 , y27659 , y27660 , y27661 , y27662 , y27663 , y27664 , y27665 , y27666 , y27667 , y27668 , y27669 , y27670 , y27671 , y27672 , y27673 , y27674 , y27675 , y27676 , y27677 , y27678 , y27679 , y27680 , y27681 , y27682 , y27683 , y27684 , y27685 , y27686 , y27687 , y27688 , y27689 , y27690 , y27691 , y27692 , y27693 , y27694 , y27695 , y27696 , y27697 , y27698 , y27699 , y27700 , y27701 , y27702 , y27703 , y27704 , y27705 , y27706 , y27707 , y27708 , y27709 , y27710 , y27711 , y27712 , y27713 , y27714 , y27715 , y27716 , y27717 , y27718 , y27719 , y27720 , y27721 , y27722 , y27723 , y27724 , y27725 , y27726 , y27727 , y27728 , y27729 , y27730 , y27731 , y27732 , y27733 , y27734 , y27735 , y27736 , y27737 , y27738 , y27739 , y27740 , y27741 , y27742 , y27743 , y27744 , y27745 , y27746 , y27747 , y27748 , y27749 , y27750 , y27751 , y27752 , y27753 , y27754 , y27755 , y27756 , y27757 , y27758 , y27759 , y27760 , y27761 , y27762 , y27763 , y27764 , y27765 , y27766 , y27767 , y27768 , y27769 , y27770 , y27771 , y27772 , y27773 , y27774 , y27775 , y27776 , y27777 , y27778 , y27779 , y27780 , y27781 , y27782 , y27783 , y27784 , y27785 , y27786 , y27787 , y27788 , y27789 , y27790 , y27791 , y27792 , y27793 , y27794 , y27795 , y27796 , y27797 , y27798 , y27799 , y27800 , y27801 , y27802 , y27803 , y27804 , y27805 , y27806 , y27807 , y27808 , y27809 , y27810 , y27811 , y27812 , y27813 , y27814 , y27815 , y27816 , y27817 , y27818 , y27819 , y27820 , y27821 , y27822 , y27823 , y27824 , y27825 , y27826 , y27827 , y27828 , y27829 , y27830 , y27831 , y27832 , y27833 , y27834 , y27835 , y27836 , y27837 , y27838 , y27839 , y27840 , y27841 , y27842 , y27843 , y27844 , y27845 , y27846 , y27847 , y27848 , y27849 , y27850 , y27851 , y27852 , y27853 , y27854 , y27855 , y27856 , y27857 , y27858 , y27859 , y27860 , y27861 , y27862 , y27863 , y27864 , y27865 , y27866 , y27867 , y27868 , y27869 , y27870 , y27871 , y27872 , y27873 , y27874 , y27875 , y27876 , y27877 , y27878 , y27879 , y27880 , y27881 , y27882 , y27883 , y27884 , y27885 , y27886 , y27887 , y27888 , y27889 , y27890 , y27891 , y27892 , y27893 , y27894 , y27895 , y27896 , y27897 , y27898 , y27899 , y27900 , y27901 , y27902 , y27903 , y27904 , y27905 , y27906 , y27907 , y27908 , y27909 , y27910 , y27911 , y27912 , y27913 , y27914 , y27915 , y27916 , y27917 , y27918 , y27919 , y27920 , y27921 , y27922 , y27923 , y27924 , y27925 , y27926 , y27927 , y27928 , y27929 , y27930 , y27931 , y27932 , y27933 , y27934 , y27935 , y27936 , y27937 , y27938 , y27939 , y27940 , y27941 , y27942 , y27943 , y27944 , y27945 , y27946 , y27947 , y27948 , y27949 , y27950 , y27951 , y27952 , y27953 , y27954 , y27955 , y27956 , y27957 , y27958 , y27959 , y27960 , y27961 , y27962 , y27963 , y27964 , y27965 , y27966 , y27967 , y27968 , y27969 , y27970 , y27971 , y27972 , y27973 , y27974 , y27975 , y27976 , y27977 , y27978 , y27979 , y27980 , y27981 , y27982 , y27983 , y27984 , y27985 , y27986 , y27987 , y27988 , y27989 , y27990 , y27991 , y27992 , y27993 , y27994 , y27995 , y27996 , y27997 , y27998 , y27999 , y28000 , y28001 , y28002 , y28003 , y28004 , y28005 , y28006 , y28007 , y28008 , y28009 , y28010 , y28011 , y28012 , y28013 , y28014 , y28015 , y28016 , y28017 , y28018 , y28019 , y28020 , y28021 , y28022 , y28023 , y28024 , y28025 , y28026 , y28027 , y28028 , y28029 , y28030 , y28031 , y28032 , y28033 , y28034 , y28035 , y28036 , y28037 , y28038 , y28039 , y28040 , y28041 , y28042 , y28043 , y28044 , y28045 , y28046 , y28047 , y28048 , y28049 , y28050 , y28051 , y28052 , y28053 , y28054 , y28055 , y28056 , y28057 , y28058 , y28059 , y28060 , y28061 , y28062 , y28063 , y28064 , y28065 , y28066 , y28067 , y28068 , y28069 , y28070 , y28071 , y28072 , y28073 , y28074 , y28075 , y28076 , y28077 , y28078 , y28079 , y28080 , y28081 , y28082 , y28083 , y28084 , y28085 , y28086 , y28087 , y28088 , y28089 , y28090 , y28091 , y28092 , y28093 , y28094 , y28095 , y28096 , y28097 , y28098 , y28099 , y28100 , y28101 , y28102 , y28103 , y28104 , y28105 , y28106 , y28107 , y28108 , y28109 , y28110 , y28111 , y28112 , y28113 , y28114 , y28115 , y28116 , y28117 , y28118 , y28119 , y28120 , y28121 , y28122 , y28123 , y28124 , y28125 , y28126 , y28127 , y28128 , y28129 , y28130 , y28131 , y28132 , y28133 , y28134 , y28135 , y28136 , y28137 , y28138 , y28139 , y28140 , y28141 , y28142 , y28143 , y28144 , y28145 , y28146 , y28147 , y28148 , y28149 , y28150 , y28151 , y28152 , y28153 , y28154 , y28155 , y28156 , y28157 , y28158 , y28159 , y28160 , y28161 , y28162 , y28163 , y28164 , y28165 , y28166 , y28167 , y28168 , y28169 , y28170 , y28171 , y28172 , y28173 , y28174 , y28175 , y28176 , y28177 , y28178 , y28179 , y28180 , y28181 , y28182 , y28183 , y28184 , y28185 , y28186 , y28187 , y28188 , y28189 , y28190 , y28191 , y28192 , y28193 , y28194 , y28195 , y28196 , y28197 , y28198 , y28199 , y28200 , y28201 , y28202 , y28203 , y28204 , y28205 , y28206 , y28207 , y28208 , y28209 , y28210 , y28211 , y28212 , y28213 , y28214 , y28215 , y28216 , y28217 , y28218 , y28219 , y28220 , y28221 , y28222 , y28223 , y28224 , y28225 , y28226 , y28227 , y28228 , y28229 , y28230 , y28231 , y28232 , y28233 , y28234 , y28235 , y28236 , y28237 , y28238 , y28239 , y28240 , y28241 , y28242 , y28243 , y28244 , y28245 , y28246 , y28247 , y28248 , y28249 , y28250 , y28251 , y28252 , y28253 , y28254 , y28255 , y28256 , y28257 , y28258 , y28259 , y28260 , y28261 , y28262 , y28263 , y28264 , y28265 , y28266 , y28267 , y28268 , y28269 , y28270 , y28271 , y28272 , y28273 , y28274 , y28275 , y28276 , y28277 , y28278 , y28279 , y28280 , y28281 , y28282 , y28283 , y28284 , y28285 , y28286 , y28287 , y28288 , y28289 , y28290 , y28291 , y28292 , y28293 , y28294 , y28295 , y28296 , y28297 , y28298 , y28299 , y28300 , y28301 , y28302 , y28303 , y28304 , y28305 , y28306 , y28307 , y28308 , y28309 , y28310 , y28311 , y28312 , y28313 , y28314 , y28315 , y28316 , y28317 , y28318 , y28319 , y28320 , y28321 , y28322 , y28323 , y28324 , y28325 , y28326 , y28327 , y28328 , y28329 , y28330 , y28331 , y28332 , y28333 , y28334 , y28335 , y28336 , y28337 , y28338 , y28339 , y28340 , y28341 , y28342 , y28343 , y28344 , y28345 , y28346 , y28347 , y28348 , y28349 , y28350 , y28351 , y28352 , y28353 , y28354 , y28355 , y28356 , y28357 , y28358 , y28359 , y28360 , y28361 , y28362 , y28363 , y28364 , y28365 , y28366 , y28367 , y28368 , y28369 , y28370 , y28371 , y28372 , y28373 , y28374 , y28375 , y28376 , y28377 , y28378 , y28379 , y28380 , y28381 , y28382 , y28383 , y28384 , y28385 , y28386 , y28387 , y28388 , y28389 , y28390 , y28391 , y28392 , y28393 , y28394 , y28395 , y28396 , y28397 , y28398 , y28399 , y28400 , y28401 , y28402 , y28403 , y28404 , y28405 , y28406 , y28407 , y28408 , y28409 , y28410 , y28411 , y28412 , y28413 , y28414 , y28415 , y28416 , y28417 , y28418 , y28419 , y28420 , y28421 , y28422 , y28423 , y28424 , y28425 , y28426 , y28427 , y28428 , y28429 , y28430 , y28431 , y28432 , y28433 , y28434 , y28435 , y28436 , y28437 , y28438 , y28439 , y28440 , y28441 , y28442 , y28443 , y28444 , y28445 , y28446 , y28447 , y28448 , y28449 , y28450 , y28451 , y28452 , y28453 , y28454 , y28455 , y28456 , y28457 , y28458 , y28459 , y28460 , y28461 , y28462 , y28463 , y28464 , y28465 , y28466 , y28467 , y28468 , y28469 , y28470 , y28471 , y28472 , y28473 , y28474 , y28475 , y28476 , y28477 , y28478 , y28479 , y28480 , y28481 , y28482 , y28483 , y28484 , y28485 , y28486 , y28487 , y28488 , y28489 , y28490 , y28491 , y28492 , y28493 , y28494 , y28495 , y28496 , y28497 , y28498 , y28499 , y28500 , y28501 , y28502 , y28503 , y28504 , y28505 , y28506 , y28507 , y28508 , y28509 , y28510 , y28511 , y28512 , y28513 , y28514 , y28515 , y28516 , y28517 , y28518 , y28519 , y28520 , y28521 , y28522 , y28523 , y28524 , y28525 , y28526 , y28527 , y28528 , y28529 , y28530 , y28531 , y28532 , y28533 , y28534 , y28535 , y28536 , y28537 , y28538 , y28539 , y28540 , y28541 , y28542 , y28543 , y28544 , y28545 , y28546 , y28547 , y28548 , y28549 , y28550 , y28551 , y28552 , y28553 , y28554 , y28555 , y28556 , y28557 , y28558 , y28559 , y28560 , y28561 , y28562 , y28563 , y28564 , y28565 , y28566 , y28567 , y28568 , y28569 , y28570 , y28571 , y28572 , y28573 , y28574 , y28575 , y28576 , y28577 , y28578 , y28579 , y28580 , y28581 , y28582 , y28583 , y28584 , y28585 , y28586 , y28587 , y28588 , y28589 , y28590 , y28591 , y28592 , y28593 , y28594 , y28595 , y28596 , y28597 , y28598 , y28599 , y28600 , y28601 , y28602 , y28603 , y28604 , y28605 , y28606 , y28607 , y28608 , y28609 , y28610 , y28611 , y28612 , y28613 , y28614 , y28615 , y28616 , y28617 , y28618 , y28619 , y28620 , y28621 , y28622 , y28623 , y28624 , y28625 , y28626 , y28627 , y28628 , y28629 , y28630 , y28631 , y28632 , y28633 , y28634 , y28635 , y28636 , y28637 , y28638 , y28639 , y28640 , y28641 , y28642 , y28643 , y28644 , y28645 , y28646 , y28647 , y28648 , y28649 , y28650 , y28651 , y28652 , y28653 , y28654 , y28655 , y28656 , y28657 , y28658 , y28659 , y28660 , y28661 , y28662 , y28663 , y28664 , y28665 , y28666 , y28667 , y28668 , y28669 , y28670 , y28671 , y28672 , y28673 , y28674 , y28675 , y28676 , y28677 , y28678 , y28679 , y28680 , y28681 , y28682 , y28683 , y28684 , y28685 , y28686 , y28687 , y28688 , y28689 , y28690 , y28691 , y28692 , y28693 , y28694 , y28695 , y28696 , y28697 , y28698 , y28699 , y28700 , y28701 , y28702 , y28703 , y28704 , y28705 , y28706 , y28707 , y28708 , y28709 , y28710 , y28711 , y28712 , y28713 , y28714 , y28715 , y28716 , y28717 , y28718 , y28719 , y28720 , y28721 , y28722 , y28723 , y28724 , y28725 , y28726 , y28727 , y28728 , y28729 , y28730 , y28731 , y28732 , y28733 , y28734 , y28735 , y28736 , y28737 , y28738 , y28739 , y28740 , y28741 , y28742 , y28743 , y28744 , y28745 , y28746 , y28747 , y28748 , y28749 , y28750 , y28751 , y28752 , y28753 , y28754 , y28755 , y28756 , y28757 , y28758 , y28759 , y28760 , y28761 , y28762 , y28763 , y28764 , y28765 , y28766 , y28767 , y28768 , y28769 , y28770 , y28771 , y28772 , y28773 , y28774 , y28775 , y28776 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 , y23806 , y23807 , y23808 , y23809 , y23810 , y23811 , y23812 , y23813 , y23814 , y23815 , y23816 , y23817 , y23818 , y23819 , y23820 , y23821 , y23822 , y23823 , y23824 , y23825 , y23826 , y23827 , y23828 , y23829 , y23830 , y23831 , y23832 , y23833 , y23834 , y23835 , y23836 , y23837 , y23838 , y23839 , y23840 , y23841 , y23842 , y23843 , y23844 , y23845 , y23846 , y23847 , y23848 , y23849 , y23850 , y23851 , y23852 , y23853 , y23854 , y23855 , y23856 , y23857 , y23858 , y23859 , y23860 , y23861 , y23862 , y23863 , y23864 , y23865 , y23866 , y23867 , y23868 , y23869 , y23870 , y23871 , y23872 , y23873 , y23874 , y23875 , y23876 , y23877 , y23878 , y23879 , y23880 , y23881 , y23882 , y23883 , y23884 , y23885 , y23886 , y23887 , y23888 , y23889 , y23890 , y23891 , y23892 , y23893 , y23894 , y23895 , y23896 , y23897 , y23898 , y23899 , y23900 , y23901 , y23902 , y23903 , y23904 , y23905 , y23906 , y23907 , y23908 , y23909 , y23910 , y23911 , y23912 , y23913 , y23914 , y23915 , y23916 , y23917 , y23918 , y23919 , y23920 , y23921 , y23922 , y23923 , y23924 , y23925 , y23926 , y23927 , y23928 , y23929 , y23930 , y23931 , y23932 , y23933 , y23934 , y23935 , y23936 , y23937 , y23938 , y23939 , y23940 , y23941 , y23942 , y23943 , y23944 , y23945 , y23946 , y23947 , y23948 , y23949 , y23950 , y23951 , y23952 , y23953 , y23954 , y23955 , y23956 , y23957 , y23958 , y23959 , y23960 , y23961 , y23962 , y23963 , y23964 , y23965 , y23966 , y23967 , y23968 , y23969 , y23970 , y23971 , y23972 , y23973 , y23974 , y23975 , y23976 , y23977 , y23978 , y23979 , y23980 , y23981 , y23982 , y23983 , y23984 , y23985 , y23986 , y23987 , y23988 , y23989 , y23990 , y23991 , y23992 , y23993 , y23994 , y23995 , y23996 , y23997 , y23998 , y23999 , y24000 , y24001 , y24002 , y24003 , y24004 , y24005 , y24006 , y24007 , y24008 , y24009 , y24010 , y24011 , y24012 , y24013 , y24014 , y24015 , y24016 , y24017 , y24018 , y24019 , y24020 , y24021 , y24022 , y24023 , y24024 , y24025 , y24026 , y24027 , y24028 , y24029 , y24030 , y24031 , y24032 , y24033 , y24034 , y24035 , y24036 , y24037 , y24038 , y24039 , y24040 , y24041 , y24042 , y24043 , y24044 , y24045 , y24046 , y24047 , y24048 , y24049 , y24050 , y24051 , y24052 , y24053 , y24054 , y24055 , y24056 , y24057 , y24058 , y24059 , y24060 , y24061 , y24062 , y24063 , y24064 , y24065 , y24066 , y24067 , y24068 , y24069 , y24070 , y24071 , y24072 , y24073 , y24074 , y24075 , y24076 , y24077 , y24078 , y24079 , y24080 , y24081 , y24082 , y24083 , y24084 , y24085 , y24086 , y24087 , y24088 , y24089 , y24090 , y24091 , y24092 , y24093 , y24094 , y24095 , y24096 , y24097 , y24098 , y24099 , y24100 , y24101 , y24102 , y24103 , y24104 , y24105 , y24106 , y24107 , y24108 , y24109 , y24110 , y24111 , y24112 , y24113 , y24114 , y24115 , y24116 , y24117 , y24118 , y24119 , y24120 , y24121 , y24122 , y24123 , y24124 , y24125 , y24126 , y24127 , y24128 , y24129 , y24130 , y24131 , y24132 , y24133 , y24134 , y24135 , y24136 , y24137 , y24138 , y24139 , y24140 , y24141 , y24142 , y24143 , y24144 , y24145 , y24146 , y24147 , y24148 , y24149 , y24150 , y24151 , y24152 , y24153 , y24154 , y24155 , y24156 , y24157 , y24158 , y24159 , y24160 , y24161 , y24162 , y24163 , y24164 , y24165 , y24166 , y24167 , y24168 , y24169 , y24170 , y24171 , y24172 , y24173 , y24174 , y24175 , y24176 , y24177 , y24178 , y24179 , y24180 , y24181 , y24182 , y24183 , y24184 , y24185 , y24186 , y24187 , y24188 , y24189 , y24190 , y24191 , y24192 , y24193 , y24194 , y24195 , y24196 , y24197 , y24198 , y24199 , y24200 , y24201 , y24202 , y24203 , y24204 , y24205 , y24206 , y24207 , y24208 , y24209 , y24210 , y24211 , y24212 , y24213 , y24214 , y24215 , y24216 , y24217 , y24218 , y24219 , y24220 , y24221 , y24222 , y24223 , y24224 , y24225 , y24226 , y24227 , y24228 , y24229 , y24230 , y24231 , y24232 , y24233 , y24234 , y24235 , y24236 , y24237 , y24238 , y24239 , y24240 , y24241 , y24242 , y24243 , y24244 , y24245 , y24246 , y24247 , y24248 , y24249 , y24250 , y24251 , y24252 , y24253 , y24254 , y24255 , y24256 , y24257 , y24258 , y24259 , y24260 , y24261 , y24262 , y24263 , y24264 , y24265 , y24266 , y24267 , y24268 , y24269 , y24270 , y24271 , y24272 , y24273 , y24274 , y24275 , y24276 , y24277 , y24278 , y24279 , y24280 , y24281 , y24282 , y24283 , y24284 , y24285 , y24286 , y24287 , y24288 , y24289 , y24290 , y24291 , y24292 , y24293 , y24294 , y24295 , y24296 , y24297 , y24298 , y24299 , y24300 , y24301 , y24302 , y24303 , y24304 , y24305 , y24306 , y24307 , y24308 , y24309 , y24310 , y24311 , y24312 , y24313 , y24314 , y24315 , y24316 , y24317 , y24318 , y24319 , y24320 , y24321 , y24322 , y24323 , y24324 , y24325 , y24326 , y24327 , y24328 , y24329 , y24330 , y24331 , y24332 , y24333 , y24334 , y24335 , y24336 , y24337 , y24338 , y24339 , y24340 , y24341 , y24342 , y24343 , y24344 , y24345 , y24346 , y24347 , y24348 , y24349 , y24350 , y24351 , y24352 , y24353 , y24354 , y24355 , y24356 , y24357 , y24358 , y24359 , y24360 , y24361 , y24362 , y24363 , y24364 , y24365 , y24366 , y24367 , y24368 , y24369 , y24370 , y24371 , y24372 , y24373 , y24374 , y24375 , y24376 , y24377 , y24378 , y24379 , y24380 , y24381 , y24382 , y24383 , y24384 , y24385 , y24386 , y24387 , y24388 , y24389 , y24390 , y24391 , y24392 , y24393 , y24394 , y24395 , y24396 , y24397 , y24398 , y24399 , y24400 , y24401 , y24402 , y24403 , y24404 , y24405 , y24406 , y24407 , y24408 , y24409 , y24410 , y24411 , y24412 , y24413 , y24414 , y24415 , y24416 , y24417 , y24418 , y24419 , y24420 , y24421 , y24422 , y24423 , y24424 , y24425 , y24426 , y24427 , y24428 , y24429 , y24430 , y24431 , y24432 , y24433 , y24434 , y24435 , y24436 , y24437 , y24438 , y24439 , y24440 , y24441 , y24442 , y24443 , y24444 , y24445 , y24446 , y24447 , y24448 , y24449 , y24450 , y24451 , y24452 , y24453 , y24454 , y24455 , y24456 , y24457 , y24458 , y24459 , y24460 , y24461 , y24462 , y24463 , y24464 , y24465 , y24466 , y24467 , y24468 , y24469 , y24470 , y24471 , y24472 , y24473 , y24474 , y24475 , y24476 , y24477 , y24478 , y24479 , y24480 , y24481 , y24482 , y24483 , y24484 , y24485 , y24486 , y24487 , y24488 , y24489 , y24490 , y24491 , y24492 , y24493 , y24494 , y24495 , y24496 , y24497 , y24498 , y24499 , y24500 , y24501 , y24502 , y24503 , y24504 , y24505 , y24506 , y24507 , y24508 , y24509 , y24510 , y24511 , y24512 , y24513 , y24514 , y24515 , y24516 , y24517 , y24518 , y24519 , y24520 , y24521 , y24522 , y24523 , y24524 , y24525 , y24526 , y24527 , y24528 , y24529 , y24530 , y24531 , y24532 , y24533 , y24534 , y24535 , y24536 , y24537 , y24538 , y24539 , y24540 , y24541 , y24542 , y24543 , y24544 , y24545 , y24546 , y24547 , y24548 , y24549 , y24550 , y24551 , y24552 , y24553 , y24554 , y24555 , y24556 , y24557 , y24558 , y24559 , y24560 , y24561 , y24562 , y24563 , y24564 , y24565 , y24566 , y24567 , y24568 , y24569 , y24570 , y24571 , y24572 , y24573 , y24574 , y24575 , y24576 , y24577 , y24578 , y24579 , y24580 , y24581 , y24582 , y24583 , y24584 , y24585 , y24586 , y24587 , y24588 , y24589 , y24590 , y24591 , y24592 , y24593 , y24594 , y24595 , y24596 , y24597 , y24598 , y24599 , y24600 , y24601 , y24602 , y24603 , y24604 , y24605 , y24606 , y24607 , y24608 , y24609 , y24610 , y24611 , y24612 , y24613 , y24614 , y24615 , y24616 , y24617 , y24618 , y24619 , y24620 , y24621 , y24622 , y24623 , y24624 , y24625 , y24626 , y24627 , y24628 , y24629 , y24630 , y24631 , y24632 , y24633 , y24634 , y24635 , y24636 , y24637 , y24638 , y24639 , y24640 , y24641 , y24642 , y24643 , y24644 , y24645 , y24646 , y24647 , y24648 , y24649 , y24650 , y24651 , y24652 , y24653 , y24654 , y24655 , y24656 , y24657 , y24658 , y24659 , y24660 , y24661 , y24662 , y24663 , y24664 , y24665 , y24666 , y24667 , y24668 , y24669 , y24670 , y24671 , y24672 , y24673 , y24674 , y24675 , y24676 , y24677 , y24678 , y24679 , y24680 , y24681 , y24682 , y24683 , y24684 , y24685 , y24686 , y24687 , y24688 , y24689 , y24690 , y24691 , y24692 , y24693 , y24694 , y24695 , y24696 , y24697 , y24698 , y24699 , y24700 , y24701 , y24702 , y24703 , y24704 , y24705 , y24706 , y24707 , y24708 , y24709 , y24710 , y24711 , y24712 , y24713 , y24714 , y24715 , y24716 , y24717 , y24718 , y24719 , y24720 , y24721 , y24722 , y24723 , y24724 , y24725 , y24726 , y24727 , y24728 , y24729 , y24730 , y24731 , y24732 , y24733 , y24734 , y24735 , y24736 , y24737 , y24738 , y24739 , y24740 , y24741 , y24742 , y24743 , y24744 , y24745 , y24746 , y24747 , y24748 , y24749 , y24750 , y24751 , y24752 , y24753 , y24754 , y24755 , y24756 , y24757 , y24758 , y24759 , y24760 , y24761 , y24762 , y24763 , y24764 , y24765 , y24766 , y24767 , y24768 , y24769 , y24770 , y24771 , y24772 , y24773 , y24774 , y24775 , y24776 , y24777 , y24778 , y24779 , y24780 , y24781 , y24782 , y24783 , y24784 , y24785 , y24786 , y24787 , y24788 , y24789 , y24790 , y24791 , y24792 , y24793 , y24794 , y24795 , y24796 , y24797 , y24798 , y24799 , y24800 , y24801 , y24802 , y24803 , y24804 , y24805 , y24806 , y24807 , y24808 , y24809 , y24810 , y24811 , y24812 , y24813 , y24814 , y24815 , y24816 , y24817 , y24818 , y24819 , y24820 , y24821 , y24822 , y24823 , y24824 , y24825 , y24826 , y24827 , y24828 , y24829 , y24830 , y24831 , y24832 , y24833 , y24834 , y24835 , y24836 , y24837 , y24838 , y24839 , y24840 , y24841 , y24842 , y24843 , y24844 , y24845 , y24846 , y24847 , y24848 , y24849 , y24850 , y24851 , y24852 , y24853 , y24854 , y24855 , y24856 , y24857 , y24858 , y24859 , y24860 , y24861 , y24862 , y24863 , y24864 , y24865 , y24866 , y24867 , y24868 , y24869 , y24870 , y24871 , y24872 , y24873 , y24874 , y24875 , y24876 , y24877 , y24878 , y24879 , y24880 , y24881 , y24882 , y24883 , y24884 , y24885 , y24886 , y24887 , y24888 , y24889 , y24890 , y24891 , y24892 , y24893 , y24894 , y24895 , y24896 , y24897 , y24898 , y24899 , y24900 , y24901 , y24902 , y24903 , y24904 , y24905 , y24906 , y24907 , y24908 , y24909 , y24910 , y24911 , y24912 , y24913 , y24914 , y24915 , y24916 , y24917 , y24918 , y24919 , y24920 , y24921 , y24922 , y24923 , y24924 , y24925 , y24926 , y24927 , y24928 , y24929 , y24930 , y24931 , y24932 , y24933 , y24934 , y24935 , y24936 , y24937 , y24938 , y24939 , y24940 , y24941 , y24942 , y24943 , y24944 , y24945 , y24946 , y24947 , y24948 , y24949 , y24950 , y24951 , y24952 , y24953 , y24954 , y24955 , y24956 , y24957 , y24958 , y24959 , y24960 , y24961 , y24962 , y24963 , y24964 , y24965 , y24966 , y24967 , y24968 , y24969 , y24970 , y24971 , y24972 , y24973 , y24974 , y24975 , y24976 , y24977 , y24978 , y24979 , y24980 , y24981 , y24982 , y24983 , y24984 , y24985 , y24986 , y24987 , y24988 , y24989 , y24990 , y24991 , y24992 , y24993 , y24994 , y24995 , y24996 , y24997 , y24998 , y24999 , y25000 , y25001 , y25002 , y25003 , y25004 , y25005 , y25006 , y25007 , y25008 , y25009 , y25010 , y25011 , y25012 , y25013 , y25014 , y25015 , y25016 , y25017 , y25018 , y25019 , y25020 , y25021 , y25022 , y25023 , y25024 , y25025 , y25026 , y25027 , y25028 , y25029 , y25030 , y25031 , y25032 , y25033 , y25034 , y25035 , y25036 , y25037 , y25038 , y25039 , y25040 , y25041 , y25042 , y25043 , y25044 , y25045 , y25046 , y25047 , y25048 , y25049 , y25050 , y25051 , y25052 , y25053 , y25054 , y25055 , y25056 , y25057 , y25058 , y25059 , y25060 , y25061 , y25062 , y25063 , y25064 , y25065 , y25066 , y25067 , y25068 , y25069 , y25070 , y25071 , y25072 , y25073 , y25074 , y25075 , y25076 , y25077 , y25078 , y25079 , y25080 , y25081 , y25082 , y25083 , y25084 , y25085 , y25086 , y25087 , y25088 , y25089 , y25090 , y25091 , y25092 , y25093 , y25094 , y25095 , y25096 , y25097 , y25098 , y25099 , y25100 , y25101 , y25102 , y25103 , y25104 , y25105 , y25106 , y25107 , y25108 , y25109 , y25110 , y25111 , y25112 , y25113 , y25114 , y25115 , y25116 , y25117 , y25118 , y25119 , y25120 , y25121 , y25122 , y25123 , y25124 , y25125 , y25126 , y25127 , y25128 , y25129 , y25130 , y25131 , y25132 , y25133 , y25134 , y25135 , y25136 , y25137 , y25138 , y25139 , y25140 , y25141 , y25142 , y25143 , y25144 , y25145 , y25146 , y25147 , y25148 , y25149 , y25150 , y25151 , y25152 , y25153 , y25154 , y25155 , y25156 , y25157 , y25158 , y25159 , y25160 , y25161 , y25162 , y25163 , y25164 , y25165 , y25166 , y25167 , y25168 , y25169 , y25170 , y25171 , y25172 , y25173 , y25174 , y25175 , y25176 , y25177 , y25178 , y25179 , y25180 , y25181 , y25182 , y25183 , y25184 , y25185 , y25186 , y25187 , y25188 , y25189 , y25190 , y25191 , y25192 , y25193 , y25194 , y25195 , y25196 , y25197 , y25198 , y25199 , y25200 , y25201 , y25202 , y25203 , y25204 , y25205 , y25206 , y25207 , y25208 , y25209 , y25210 , y25211 , y25212 , y25213 , y25214 , y25215 , y25216 , y25217 , y25218 , y25219 , y25220 , y25221 , y25222 , y25223 , y25224 , y25225 , y25226 , y25227 , y25228 , y25229 , y25230 , y25231 , y25232 , y25233 , y25234 , y25235 , y25236 , y25237 , y25238 , y25239 , y25240 , y25241 , y25242 , y25243 , y25244 , y25245 , y25246 , y25247 , y25248 , y25249 , y25250 , y25251 , y25252 , y25253 , y25254 , y25255 , y25256 , y25257 , y25258 , y25259 , y25260 , y25261 , y25262 , y25263 , y25264 , y25265 , y25266 , y25267 , y25268 , y25269 , y25270 , y25271 , y25272 , y25273 , y25274 , y25275 , y25276 , y25277 , y25278 , y25279 , y25280 , y25281 , y25282 , y25283 , y25284 , y25285 , y25286 , y25287 , y25288 , y25289 , y25290 , y25291 , y25292 , y25293 , y25294 , y25295 , y25296 , y25297 , y25298 , y25299 , y25300 , y25301 , y25302 , y25303 , y25304 , y25305 , y25306 , y25307 , y25308 , y25309 , y25310 , y25311 , y25312 , y25313 , y25314 , y25315 , y25316 , y25317 , y25318 , y25319 , y25320 , y25321 , y25322 , y25323 , y25324 , y25325 , y25326 , y25327 , y25328 , y25329 , y25330 , y25331 , y25332 , y25333 , y25334 , y25335 , y25336 , y25337 , y25338 , y25339 , y25340 , y25341 , y25342 , y25343 , y25344 , y25345 , y25346 , y25347 , y25348 , y25349 , y25350 , y25351 , y25352 , y25353 , y25354 , y25355 , y25356 , y25357 , y25358 , y25359 , y25360 , y25361 , y25362 , y25363 , y25364 , y25365 , y25366 , y25367 , y25368 , y25369 , y25370 , y25371 , y25372 , y25373 , y25374 , y25375 , y25376 , y25377 , y25378 , y25379 , y25380 , y25381 , y25382 , y25383 , y25384 , y25385 , y25386 , y25387 , y25388 , y25389 , y25390 , y25391 , y25392 , y25393 , y25394 , y25395 , y25396 , y25397 , y25398 , y25399 , y25400 , y25401 , y25402 , y25403 , y25404 , y25405 , y25406 , y25407 , y25408 , y25409 , y25410 , y25411 , y25412 , y25413 , y25414 , y25415 , y25416 , y25417 , y25418 , y25419 , y25420 , y25421 , y25422 , y25423 , y25424 , y25425 , y25426 , y25427 , y25428 , y25429 , y25430 , y25431 , y25432 , y25433 , y25434 , y25435 , y25436 , y25437 , y25438 , y25439 , y25440 , y25441 , y25442 , y25443 , y25444 , y25445 , y25446 , y25447 , y25448 , y25449 , y25450 , y25451 , y25452 , y25453 , y25454 , y25455 , y25456 , y25457 , y25458 , y25459 , y25460 , y25461 , y25462 , y25463 , y25464 , y25465 , y25466 , y25467 , y25468 , y25469 , y25470 , y25471 , y25472 , y25473 , y25474 , y25475 , y25476 , y25477 , y25478 , y25479 , y25480 , y25481 , y25482 , y25483 , y25484 , y25485 , y25486 , y25487 , y25488 , y25489 , y25490 , y25491 , y25492 , y25493 , y25494 , y25495 , y25496 , y25497 , y25498 , y25499 , y25500 , y25501 , y25502 , y25503 , y25504 , y25505 , y25506 , y25507 , y25508 , y25509 , y25510 , y25511 , y25512 , y25513 , y25514 , y25515 , y25516 , y25517 , y25518 , y25519 , y25520 , y25521 , y25522 , y25523 , y25524 , y25525 , y25526 , y25527 , y25528 , y25529 , y25530 , y25531 , y25532 , y25533 , y25534 , y25535 , y25536 , y25537 , y25538 , y25539 , y25540 , y25541 , y25542 , y25543 , y25544 , y25545 , y25546 , y25547 , y25548 , y25549 , y25550 , y25551 , y25552 , y25553 , y25554 , y25555 , y25556 , y25557 , y25558 , y25559 , y25560 , y25561 , y25562 , y25563 , y25564 , y25565 , y25566 , y25567 , y25568 , y25569 , y25570 , y25571 , y25572 , y25573 , y25574 , y25575 , y25576 , y25577 , y25578 , y25579 , y25580 , y25581 , y25582 , y25583 , y25584 , y25585 , y25586 , y25587 , y25588 , y25589 , y25590 , y25591 , y25592 , y25593 , y25594 , y25595 , y25596 , y25597 , y25598 , y25599 , y25600 , y25601 , y25602 , y25603 , y25604 , y25605 , y25606 , y25607 , y25608 , y25609 , y25610 , y25611 , y25612 , y25613 , y25614 , y25615 , y25616 , y25617 , y25618 , y25619 , y25620 , y25621 , y25622 , y25623 , y25624 , y25625 , y25626 , y25627 , y25628 , y25629 , y25630 , y25631 , y25632 , y25633 , y25634 , y25635 , y25636 , y25637 , y25638 , y25639 , y25640 , y25641 , y25642 , y25643 , y25644 , y25645 , y25646 , y25647 , y25648 , y25649 , y25650 , y25651 , y25652 , y25653 , y25654 , y25655 , y25656 , y25657 , y25658 , y25659 , y25660 , y25661 , y25662 , y25663 , y25664 , y25665 , y25666 , y25667 , y25668 , y25669 , y25670 , y25671 , y25672 , y25673 , y25674 , y25675 , y25676 , y25677 , y25678 , y25679 , y25680 , y25681 , y25682 , y25683 , y25684 , y25685 , y25686 , y25687 , y25688 , y25689 , y25690 , y25691 , y25692 , y25693 , y25694 , y25695 , y25696 , y25697 , y25698 , y25699 , y25700 , y25701 , y25702 , y25703 , y25704 , y25705 , y25706 , y25707 , y25708 , y25709 , y25710 , y25711 , y25712 , y25713 , y25714 , y25715 , y25716 , y25717 , y25718 , y25719 , y25720 , y25721 , y25722 , y25723 , y25724 , y25725 , y25726 , y25727 , y25728 , y25729 , y25730 , y25731 , y25732 , y25733 , y25734 , y25735 , y25736 , y25737 , y25738 , y25739 , y25740 , y25741 , y25742 , y25743 , y25744 , y25745 , y25746 , y25747 , y25748 , y25749 , y25750 , y25751 , y25752 , y25753 , y25754 , y25755 , y25756 , y25757 , y25758 , y25759 , y25760 , y25761 , y25762 , y25763 , y25764 , y25765 , y25766 , y25767 , y25768 , y25769 , y25770 , y25771 , y25772 , y25773 , y25774 , y25775 , y25776 , y25777 , y25778 , y25779 , y25780 , y25781 , y25782 , y25783 , y25784 , y25785 , y25786 , y25787 , y25788 , y25789 , y25790 , y25791 , y25792 , y25793 , y25794 , y25795 , y25796 , y25797 , y25798 , y25799 , y25800 , y25801 , y25802 , y25803 , y25804 , y25805 , y25806 , y25807 , y25808 , y25809 , y25810 , y25811 , y25812 , y25813 , y25814 , y25815 , y25816 , y25817 , y25818 , y25819 , y25820 , y25821 , y25822 , y25823 , y25824 , y25825 , y25826 , y25827 , y25828 , y25829 , y25830 , y25831 , y25832 , y25833 , y25834 , y25835 , y25836 , y25837 , y25838 , y25839 , y25840 , y25841 , y25842 , y25843 , y25844 , y25845 , y25846 , y25847 , y25848 , y25849 , y25850 , y25851 , y25852 , y25853 , y25854 , y25855 , y25856 , y25857 , y25858 , y25859 , y25860 , y25861 , y25862 , y25863 , y25864 , y25865 , y25866 , y25867 , y25868 , y25869 , y25870 , y25871 , y25872 , y25873 , y25874 , y25875 , y25876 , y25877 , y25878 , y25879 , y25880 , y25881 , y25882 , y25883 , y25884 , y25885 , y25886 , y25887 , y25888 , y25889 , y25890 , y25891 , y25892 , y25893 , y25894 , y25895 , y25896 , y25897 , y25898 , y25899 , y25900 , y25901 , y25902 , y25903 , y25904 , y25905 , y25906 , y25907 , y25908 , y25909 , y25910 , y25911 , y25912 , y25913 , y25914 , y25915 , y25916 , y25917 , y25918 , y25919 , y25920 , y25921 , y25922 , y25923 , y25924 , y25925 , y25926 , y25927 , y25928 , y25929 , y25930 , y25931 , y25932 , y25933 , y25934 , y25935 , y25936 , y25937 , y25938 , y25939 , y25940 , y25941 , y25942 , y25943 , y25944 , y25945 , y25946 , y25947 , y25948 , y25949 , y25950 , y25951 , y25952 , y25953 , y25954 , y25955 , y25956 , y25957 , y25958 , y25959 , y25960 , y25961 , y25962 , y25963 , y25964 , y25965 , y25966 , y25967 , y25968 , y25969 , y25970 , y25971 , y25972 , y25973 , y25974 , y25975 , y25976 , y25977 , y25978 , y25979 , y25980 , y25981 , y25982 , y25983 , y25984 , y25985 , y25986 , y25987 , y25988 , y25989 , y25990 , y25991 , y25992 , y25993 , y25994 , y25995 , y25996 , y25997 , y25998 , y25999 , y26000 , y26001 , y26002 , y26003 , y26004 , y26005 , y26006 , y26007 , y26008 , y26009 , y26010 , y26011 , y26012 , y26013 , y26014 , y26015 , y26016 , y26017 , y26018 , y26019 , y26020 , y26021 , y26022 , y26023 , y26024 , y26025 , y26026 , y26027 , y26028 , y26029 , y26030 , y26031 , y26032 , y26033 , y26034 , y26035 , y26036 , y26037 , y26038 , y26039 , y26040 , y26041 , y26042 , y26043 , y26044 , y26045 , y26046 , y26047 , y26048 , y26049 , y26050 , y26051 , y26052 , y26053 , y26054 , y26055 , y26056 , y26057 , y26058 , y26059 , y26060 , y26061 , y26062 , y26063 , y26064 , y26065 , y26066 , y26067 , y26068 , y26069 , y26070 , y26071 , y26072 , y26073 , y26074 , y26075 , y26076 , y26077 , y26078 , y26079 , y26080 , y26081 , y26082 , y26083 , y26084 , y26085 , y26086 , y26087 , y26088 , y26089 , y26090 , y26091 , y26092 , y26093 , y26094 , y26095 , y26096 , y26097 , y26098 , y26099 , y26100 , y26101 , y26102 , y26103 , y26104 , y26105 , y26106 , y26107 , y26108 , y26109 , y26110 , y26111 , y26112 , y26113 , y26114 , y26115 , y26116 , y26117 , y26118 , y26119 , y26120 , y26121 , y26122 , y26123 , y26124 , y26125 , y26126 , y26127 , y26128 , y26129 , y26130 , y26131 , y26132 , y26133 , y26134 , y26135 , y26136 , y26137 , y26138 , y26139 , y26140 , y26141 , y26142 , y26143 , y26144 , y26145 , y26146 , y26147 , y26148 , y26149 , y26150 , y26151 , y26152 , y26153 , y26154 , y26155 , y26156 , y26157 , y26158 , y26159 , y26160 , y26161 , y26162 , y26163 , y26164 , y26165 , y26166 , y26167 , y26168 , y26169 , y26170 , y26171 , y26172 , y26173 , y26174 , y26175 , y26176 , y26177 , y26178 , y26179 , y26180 , y26181 , y26182 , y26183 , y26184 , y26185 , y26186 , y26187 , y26188 , y26189 , y26190 , y26191 , y26192 , y26193 , y26194 , y26195 , y26196 , y26197 , y26198 , y26199 , y26200 , y26201 , y26202 , y26203 , y26204 , y26205 , y26206 , y26207 , y26208 , y26209 , y26210 , y26211 , y26212 , y26213 , y26214 , y26215 , y26216 , y26217 , y26218 , y26219 , y26220 , y26221 , y26222 , y26223 , y26224 , y26225 , y26226 , y26227 , y26228 , y26229 , y26230 , y26231 , y26232 , y26233 , y26234 , y26235 , y26236 , y26237 , y26238 , y26239 , y26240 , y26241 , y26242 , y26243 , y26244 , y26245 , y26246 , y26247 , y26248 , y26249 , y26250 , y26251 , y26252 , y26253 , y26254 , y26255 , y26256 , y26257 , y26258 , y26259 , y26260 , y26261 , y26262 , y26263 , y26264 , y26265 , y26266 , y26267 , y26268 , y26269 , y26270 , y26271 , y26272 , y26273 , y26274 , y26275 , y26276 , y26277 , y26278 , y26279 , y26280 , y26281 , y26282 , y26283 , y26284 , y26285 , y26286 , y26287 , y26288 , y26289 , y26290 , y26291 , y26292 , y26293 , y26294 , y26295 , y26296 , y26297 , y26298 , y26299 , y26300 , y26301 , y26302 , y26303 , y26304 , y26305 , y26306 , y26307 , y26308 , y26309 , y26310 , y26311 , y26312 , y26313 , y26314 , y26315 , y26316 , y26317 , y26318 , y26319 , y26320 , y26321 , y26322 , y26323 , y26324 , y26325 , y26326 , y26327 , y26328 , y26329 , y26330 , y26331 , y26332 , y26333 , y26334 , y26335 , y26336 , y26337 , y26338 , y26339 , y26340 , y26341 , y26342 , y26343 , y26344 , y26345 , y26346 , y26347 , y26348 , y26349 , y26350 , y26351 , y26352 , y26353 , y26354 , y26355 , y26356 , y26357 , y26358 , y26359 , y26360 , y26361 , y26362 , y26363 , y26364 , y26365 , y26366 , y26367 , y26368 , y26369 , y26370 , y26371 , y26372 , y26373 , y26374 , y26375 , y26376 , y26377 , y26378 , y26379 , y26380 , y26381 , y26382 , y26383 , y26384 , y26385 , y26386 , y26387 , y26388 , y26389 , y26390 , y26391 , y26392 , y26393 , y26394 , y26395 , y26396 , y26397 , y26398 , y26399 , y26400 , y26401 , y26402 , y26403 , y26404 , y26405 , y26406 , y26407 , y26408 , y26409 , y26410 , y26411 , y26412 , y26413 , y26414 , y26415 , y26416 , y26417 , y26418 , y26419 , y26420 , y26421 , y26422 , y26423 , y26424 , y26425 , y26426 , y26427 , y26428 , y26429 , y26430 , y26431 , y26432 , y26433 , y26434 , y26435 , y26436 , y26437 , y26438 , y26439 , y26440 , y26441 , y26442 , y26443 , y26444 , y26445 , y26446 , y26447 , y26448 , y26449 , y26450 , y26451 , y26452 , y26453 , y26454 , y26455 , y26456 , y26457 , y26458 , y26459 , y26460 , y26461 , y26462 , y26463 , y26464 , y26465 , y26466 , y26467 , y26468 , y26469 , y26470 , y26471 , y26472 , y26473 , y26474 , y26475 , y26476 , y26477 , y26478 , y26479 , y26480 , y26481 , y26482 , y26483 , y26484 , y26485 , y26486 , y26487 , y26488 , y26489 , y26490 , y26491 , y26492 , y26493 , y26494 , y26495 , y26496 , y26497 , y26498 , y26499 , y26500 , y26501 , y26502 , y26503 , y26504 , y26505 , y26506 , y26507 , y26508 , y26509 , y26510 , y26511 , y26512 , y26513 , y26514 , y26515 , y26516 , y26517 , y26518 , y26519 , y26520 , y26521 , y26522 , y26523 , y26524 , y26525 , y26526 , y26527 , y26528 , y26529 , y26530 , y26531 , y26532 , y26533 , y26534 , y26535 , y26536 , y26537 , y26538 , y26539 , y26540 , y26541 , y26542 , y26543 , y26544 , y26545 , y26546 , y26547 , y26548 , y26549 , y26550 , y26551 , y26552 , y26553 , y26554 , y26555 , y26556 , y26557 , y26558 , y26559 , y26560 , y26561 , y26562 , y26563 , y26564 , y26565 , y26566 , y26567 , y26568 , y26569 , y26570 , y26571 , y26572 , y26573 , y26574 , y26575 , y26576 , y26577 , y26578 , y26579 , y26580 , y26581 , y26582 , y26583 , y26584 , y26585 , y26586 , y26587 , y26588 , y26589 , y26590 , y26591 , y26592 , y26593 , y26594 , y26595 , y26596 , y26597 , y26598 , y26599 , y26600 , y26601 , y26602 , y26603 , y26604 , y26605 , y26606 , y26607 , y26608 , y26609 , y26610 , y26611 , y26612 , y26613 , y26614 , y26615 , y26616 , y26617 , y26618 , y26619 , y26620 , y26621 , y26622 , y26623 , y26624 , y26625 , y26626 , y26627 , y26628 , y26629 , y26630 , y26631 , y26632 , y26633 , y26634 , y26635 , y26636 , y26637 , y26638 , y26639 , y26640 , y26641 , y26642 , y26643 , y26644 , y26645 , y26646 , y26647 , y26648 , y26649 , y26650 , y26651 , y26652 , y26653 , y26654 , y26655 , y26656 , y26657 , y26658 , y26659 , y26660 , y26661 , y26662 , y26663 , y26664 , y26665 , y26666 , y26667 , y26668 , y26669 , y26670 , y26671 , y26672 , y26673 , y26674 , y26675 , y26676 , y26677 , y26678 , y26679 , y26680 , y26681 , y26682 , y26683 , y26684 , y26685 , y26686 , y26687 , y26688 , y26689 , y26690 , y26691 , y26692 , y26693 , y26694 , y26695 , y26696 , y26697 , y26698 , y26699 , y26700 , y26701 , y26702 , y26703 , y26704 , y26705 , y26706 , y26707 , y26708 , y26709 , y26710 , y26711 , y26712 , y26713 , y26714 , y26715 , y26716 , y26717 , y26718 , y26719 , y26720 , y26721 , y26722 , y26723 , y26724 , y26725 , y26726 , y26727 , y26728 , y26729 , y26730 , y26731 , y26732 , y26733 , y26734 , y26735 , y26736 , y26737 , y26738 , y26739 , y26740 , y26741 , y26742 , y26743 , y26744 , y26745 , y26746 , y26747 , y26748 , y26749 , y26750 , y26751 , y26752 , y26753 , y26754 , y26755 , y26756 , y26757 , y26758 , y26759 , y26760 , y26761 , y26762 , y26763 , y26764 , y26765 , y26766 , y26767 , y26768 , y26769 , y26770 , y26771 , y26772 , y26773 , y26774 , y26775 , y26776 , y26777 , y26778 , y26779 , y26780 , y26781 , y26782 , y26783 , y26784 , y26785 , y26786 , y26787 , y26788 , y26789 , y26790 , y26791 , y26792 , y26793 , y26794 , y26795 , y26796 , y26797 , y26798 , y26799 , y26800 , y26801 , y26802 , y26803 , y26804 , y26805 , y26806 , y26807 , y26808 , y26809 , y26810 , y26811 , y26812 , y26813 , y26814 , y26815 , y26816 , y26817 , y26818 , y26819 , y26820 , y26821 , y26822 , y26823 , y26824 , y26825 , y26826 , y26827 , y26828 , y26829 , y26830 , y26831 , y26832 , y26833 , y26834 , y26835 , y26836 , y26837 , y26838 , y26839 , y26840 , y26841 , y26842 , y26843 , y26844 , y26845 , y26846 , y26847 , y26848 , y26849 , y26850 , y26851 , y26852 , y26853 , y26854 , y26855 , y26856 , y26857 , y26858 , y26859 , y26860 , y26861 , y26862 , y26863 , y26864 , y26865 , y26866 , y26867 , y26868 , y26869 , y26870 , y26871 , y26872 , y26873 , y26874 , y26875 , y26876 , y26877 , y26878 , y26879 , y26880 , y26881 , y26882 , y26883 , y26884 , y26885 , y26886 , y26887 , y26888 , y26889 , y26890 , y26891 , y26892 , y26893 , y26894 , y26895 , y26896 , y26897 , y26898 , y26899 , y26900 , y26901 , y26902 , y26903 , y26904 , y26905 , y26906 , y26907 , y26908 , y26909 , y26910 , y26911 , y26912 , y26913 , y26914 , y26915 , y26916 , y26917 , y26918 , y26919 , y26920 , y26921 , y26922 , y26923 , y26924 , y26925 , y26926 , y26927 , y26928 , y26929 , y26930 , y26931 , y26932 , y26933 , y26934 , y26935 , y26936 , y26937 , y26938 , y26939 , y26940 , y26941 , y26942 , y26943 , y26944 , y26945 , y26946 , y26947 , y26948 , y26949 , y26950 , y26951 , y26952 , y26953 , y26954 , y26955 , y26956 , y26957 , y26958 , y26959 , y26960 , y26961 , y26962 , y26963 , y26964 , y26965 , y26966 , y26967 , y26968 , y26969 , y26970 , y26971 , y26972 , y26973 , y26974 , y26975 , y26976 , y26977 , y26978 , y26979 , y26980 , y26981 , y26982 , y26983 , y26984 , y26985 , y26986 , y26987 , y26988 , y26989 , y26990 , y26991 , y26992 , y26993 , y26994 , y26995 , y26996 , y26997 , y26998 , y26999 , y27000 , y27001 , y27002 , y27003 , y27004 , y27005 , y27006 , y27007 , y27008 , y27009 , y27010 , y27011 , y27012 , y27013 , y27014 , y27015 , y27016 , y27017 , y27018 , y27019 , y27020 , y27021 , y27022 , y27023 , y27024 , y27025 , y27026 , y27027 , y27028 , y27029 , y27030 , y27031 , y27032 , y27033 , y27034 , y27035 , y27036 , y27037 , y27038 , y27039 , y27040 , y27041 , y27042 , y27043 , y27044 , y27045 , y27046 , y27047 , y27048 , y27049 , y27050 , y27051 , y27052 , y27053 , y27054 , y27055 , y27056 , y27057 , y27058 , y27059 , y27060 , y27061 , y27062 , y27063 , y27064 , y27065 , y27066 , y27067 , y27068 , y27069 , y27070 , y27071 , y27072 , y27073 , y27074 , y27075 , y27076 , y27077 , y27078 , y27079 , y27080 , y27081 , y27082 , y27083 , y27084 , y27085 , y27086 , y27087 , y27088 , y27089 , y27090 , y27091 , y27092 , y27093 , y27094 , y27095 , y27096 , y27097 , y27098 , y27099 , y27100 , y27101 , y27102 , y27103 , y27104 , y27105 , y27106 , y27107 , y27108 , y27109 , y27110 , y27111 , y27112 , y27113 , y27114 , y27115 , y27116 , y27117 , y27118 , y27119 , y27120 , y27121 , y27122 , y27123 , y27124 , y27125 , y27126 , y27127 , y27128 , y27129 , y27130 , y27131 , y27132 , y27133 , y27134 , y27135 , y27136 , y27137 , y27138 , y27139 , y27140 , y27141 , y27142 , y27143 , y27144 , y27145 , y27146 , y27147 , y27148 , y27149 , y27150 , y27151 , y27152 , y27153 , y27154 , y27155 , y27156 , y27157 , y27158 , y27159 , y27160 , y27161 , y27162 , y27163 , y27164 , y27165 , y27166 , y27167 , y27168 , y27169 , y27170 , y27171 , y27172 , y27173 , y27174 , y27175 , y27176 , y27177 , y27178 , y27179 , y27180 , y27181 , y27182 , y27183 , y27184 , y27185 , y27186 , y27187 , y27188 , y27189 , y27190 , y27191 , y27192 , y27193 , y27194 , y27195 , y27196 , y27197 , y27198 , y27199 , y27200 , y27201 , y27202 , y27203 , y27204 , y27205 , y27206 , y27207 , y27208 , y27209 , y27210 , y27211 , y27212 , y27213 , y27214 , y27215 , y27216 , y27217 , y27218 , y27219 , y27220 , y27221 , y27222 , y27223 , y27224 , y27225 , y27226 , y27227 , y27228 , y27229 , y27230 , y27231 , y27232 , y27233 , y27234 , y27235 , y27236 , y27237 , y27238 , y27239 , y27240 , y27241 , y27242 , y27243 , y27244 , y27245 , y27246 , y27247 , y27248 , y27249 , y27250 , y27251 , y27252 , y27253 , y27254 , y27255 , y27256 , y27257 , y27258 , y27259 , y27260 , y27261 , y27262 , y27263 , y27264 , y27265 , y27266 , y27267 , y27268 , y27269 , y27270 , y27271 , y27272 , y27273 , y27274 , y27275 , y27276 , y27277 , y27278 , y27279 , y27280 , y27281 , y27282 , y27283 , y27284 , y27285 , y27286 , y27287 , y27288 , y27289 , y27290 , y27291 , y27292 , y27293 , y27294 , y27295 , y27296 , y27297 , y27298 , y27299 , y27300 , y27301 , y27302 , y27303 , y27304 , y27305 , y27306 , y27307 , y27308 , y27309 , y27310 , y27311 , y27312 , y27313 , y27314 , y27315 , y27316 , y27317 , y27318 , y27319 , y27320 , y27321 , y27322 , y27323 , y27324 , y27325 , y27326 , y27327 , y27328 , y27329 , y27330 , y27331 , y27332 , y27333 , y27334 , y27335 , y27336 , y27337 , y27338 , y27339 , y27340 , y27341 , y27342 , y27343 , y27344 , y27345 , y27346 , y27347 , y27348 , y27349 , y27350 , y27351 , y27352 , y27353 , y27354 , y27355 , y27356 , y27357 , y27358 , y27359 , y27360 , y27361 , y27362 , y27363 , y27364 , y27365 , y27366 , y27367 , y27368 , y27369 , y27370 , y27371 , y27372 , y27373 , y27374 , y27375 , y27376 , y27377 , y27378 , y27379 , y27380 , y27381 , y27382 , y27383 , y27384 , y27385 , y27386 , y27387 , y27388 , y27389 , y27390 , y27391 , y27392 , y27393 , y27394 , y27395 , y27396 , y27397 , y27398 , y27399 , y27400 , y27401 , y27402 , y27403 , y27404 , y27405 , y27406 , y27407 , y27408 , y27409 , y27410 , y27411 , y27412 , y27413 , y27414 , y27415 , y27416 , y27417 , y27418 , y27419 , y27420 , y27421 , y27422 , y27423 , y27424 , y27425 , y27426 , y27427 , y27428 , y27429 , y27430 , y27431 , y27432 , y27433 , y27434 , y27435 , y27436 , y27437 , y27438 , y27439 , y27440 , y27441 , y27442 , y27443 , y27444 , y27445 , y27446 , y27447 , y27448 , y27449 , y27450 , y27451 , y27452 , y27453 , y27454 , y27455 , y27456 , y27457 , y27458 , y27459 , y27460 , y27461 , y27462 , y27463 , y27464 , y27465 , y27466 , y27467 , y27468 , y27469 , y27470 , y27471 , y27472 , y27473 , y27474 , y27475 , y27476 , y27477 , y27478 , y27479 , y27480 , y27481 , y27482 , y27483 , y27484 , y27485 , y27486 , y27487 , y27488 , y27489 , y27490 , y27491 , y27492 , y27493 , y27494 , y27495 , y27496 , y27497 , y27498 , y27499 , y27500 , y27501 , y27502 , y27503 , y27504 , y27505 , y27506 , y27507 , y27508 , y27509 , y27510 , y27511 , y27512 , y27513 , y27514 , y27515 , y27516 , y27517 , y27518 , y27519 , y27520 , y27521 , y27522 , y27523 , y27524 , y27525 , y27526 , y27527 , y27528 , y27529 , y27530 , y27531 , y27532 , y27533 , y27534 , y27535 , y27536 , y27537 , y27538 , y27539 , y27540 , y27541 , y27542 , y27543 , y27544 , y27545 , y27546 , y27547 , y27548 , y27549 , y27550 , y27551 , y27552 , y27553 , y27554 , y27555 , y27556 , y27557 , y27558 , y27559 , y27560 , y27561 , y27562 , y27563 , y27564 , y27565 , y27566 , y27567 , y27568 , y27569 , y27570 , y27571 , y27572 , y27573 , y27574 , y27575 , y27576 , y27577 , y27578 , y27579 , y27580 , y27581 , y27582 , y27583 , y27584 , y27585 , y27586 , y27587 , y27588 , y27589 , y27590 , y27591 , y27592 , y27593 , y27594 , y27595 , y27596 , y27597 , y27598 , y27599 , y27600 , y27601 , y27602 , y27603 , y27604 , y27605 , y27606 , y27607 , y27608 , y27609 , y27610 , y27611 , y27612 , y27613 , y27614 , y27615 , y27616 , y27617 , y27618 , y27619 , y27620 , y27621 , y27622 , y27623 , y27624 , y27625 , y27626 , y27627 , y27628 , y27629 , y27630 , y27631 , y27632 , y27633 , y27634 , y27635 , y27636 , y27637 , y27638 , y27639 , y27640 , y27641 , y27642 , y27643 , y27644 , y27645 , y27646 , y27647 , y27648 , y27649 , y27650 , y27651 , y27652 , y27653 , y27654 , y27655 , y27656 , y27657 , y27658 , y27659 , y27660 , y27661 , y27662 , y27663 , y27664 , y27665 , y27666 , y27667 , y27668 , y27669 , y27670 , y27671 , y27672 , y27673 , y27674 , y27675 , y27676 , y27677 , y27678 , y27679 , y27680 , y27681 , y27682 , y27683 , y27684 , y27685 , y27686 , y27687 , y27688 , y27689 , y27690 , y27691 , y27692 , y27693 , y27694 , y27695 , y27696 , y27697 , y27698 , y27699 , y27700 , y27701 , y27702 , y27703 , y27704 , y27705 , y27706 , y27707 , y27708 , y27709 , y27710 , y27711 , y27712 , y27713 , y27714 , y27715 , y27716 , y27717 , y27718 , y27719 , y27720 , y27721 , y27722 , y27723 , y27724 , y27725 , y27726 , y27727 , y27728 , y27729 , y27730 , y27731 , y27732 , y27733 , y27734 , y27735 , y27736 , y27737 , y27738 , y27739 , y27740 , y27741 , y27742 , y27743 , y27744 , y27745 , y27746 , y27747 , y27748 , y27749 , y27750 , y27751 , y27752 , y27753 , y27754 , y27755 , y27756 , y27757 , y27758 , y27759 , y27760 , y27761 , y27762 , y27763 , y27764 , y27765 , y27766 , y27767 , y27768 , y27769 , y27770 , y27771 , y27772 , y27773 , y27774 , y27775 , y27776 , y27777 , y27778 , y27779 , y27780 , y27781 , y27782 , y27783 , y27784 , y27785 , y27786 , y27787 , y27788 , y27789 , y27790 , y27791 , y27792 , y27793 , y27794 , y27795 , y27796 , y27797 , y27798 , y27799 , y27800 , y27801 , y27802 , y27803 , y27804 , y27805 , y27806 , y27807 , y27808 , y27809 , y27810 , y27811 , y27812 , y27813 , y27814 , y27815 , y27816 , y27817 , y27818 , y27819 , y27820 , y27821 , y27822 , y27823 , y27824 , y27825 , y27826 , y27827 , y27828 , y27829 , y27830 , y27831 , y27832 , y27833 , y27834 , y27835 , y27836 , y27837 , y27838 , y27839 , y27840 , y27841 , y27842 , y27843 , y27844 , y27845 , y27846 , y27847 , y27848 , y27849 , y27850 , y27851 , y27852 , y27853 , y27854 , y27855 , y27856 , y27857 , y27858 , y27859 , y27860 , y27861 , y27862 , y27863 , y27864 , y27865 , y27866 , y27867 , y27868 , y27869 , y27870 , y27871 , y27872 , y27873 , y27874 , y27875 , y27876 , y27877 , y27878 , y27879 , y27880 , y27881 , y27882 , y27883 , y27884 , y27885 , y27886 , y27887 , y27888 , y27889 , y27890 , y27891 , y27892 , y27893 , y27894 , y27895 , y27896 , y27897 , y27898 , y27899 , y27900 , y27901 , y27902 , y27903 , y27904 , y27905 , y27906 , y27907 , y27908 , y27909 , y27910 , y27911 , y27912 , y27913 , y27914 , y27915 , y27916 , y27917 , y27918 , y27919 , y27920 , y27921 , y27922 , y27923 , y27924 , y27925 , y27926 , y27927 , y27928 , y27929 , y27930 , y27931 , y27932 , y27933 , y27934 , y27935 , y27936 , y27937 , y27938 , y27939 , y27940 , y27941 , y27942 , y27943 , y27944 , y27945 , y27946 , y27947 , y27948 , y27949 , y27950 , y27951 , y27952 , y27953 , y27954 , y27955 , y27956 , y27957 , y27958 , y27959 , y27960 , y27961 , y27962 , y27963 , y27964 , y27965 , y27966 , y27967 , y27968 , y27969 , y27970 , y27971 , y27972 , y27973 , y27974 , y27975 , y27976 , y27977 , y27978 , y27979 , y27980 , y27981 , y27982 , y27983 , y27984 , y27985 , y27986 , y27987 , y27988 , y27989 , y27990 , y27991 , y27992 , y27993 , y27994 , y27995 , y27996 , y27997 , y27998 , y27999 , y28000 , y28001 , y28002 , y28003 , y28004 , y28005 , y28006 , y28007 , y28008 , y28009 , y28010 , y28011 , y28012 , y28013 , y28014 , y28015 , y28016 , y28017 , y28018 , y28019 , y28020 , y28021 , y28022 , y28023 , y28024 , y28025 , y28026 , y28027 , y28028 , y28029 , y28030 , y28031 , y28032 , y28033 , y28034 , y28035 , y28036 , y28037 , y28038 , y28039 , y28040 , y28041 , y28042 , y28043 , y28044 , y28045 , y28046 , y28047 , y28048 , y28049 , y28050 , y28051 , y28052 , y28053 , y28054 , y28055 , y28056 , y28057 , y28058 , y28059 , y28060 , y28061 , y28062 , y28063 , y28064 , y28065 , y28066 , y28067 , y28068 , y28069 , y28070 , y28071 , y28072 , y28073 , y28074 , y28075 , y28076 , y28077 , y28078 , y28079 , y28080 , y28081 , y28082 , y28083 , y28084 , y28085 , y28086 , y28087 , y28088 , y28089 , y28090 , y28091 , y28092 , y28093 , y28094 , y28095 , y28096 , y28097 , y28098 , y28099 , y28100 , y28101 , y28102 , y28103 , y28104 , y28105 , y28106 , y28107 , y28108 , y28109 , y28110 , y28111 , y28112 , y28113 , y28114 , y28115 , y28116 , y28117 , y28118 , y28119 , y28120 , y28121 , y28122 , y28123 , y28124 , y28125 , y28126 , y28127 , y28128 , y28129 , y28130 , y28131 , y28132 , y28133 , y28134 , y28135 , y28136 , y28137 , y28138 , y28139 , y28140 , y28141 , y28142 , y28143 , y28144 , y28145 , y28146 , y28147 , y28148 , y28149 , y28150 , y28151 , y28152 , y28153 , y28154 , y28155 , y28156 , y28157 , y28158 , y28159 , y28160 , y28161 , y28162 , y28163 , y28164 , y28165 , y28166 , y28167 , y28168 , y28169 , y28170 , y28171 , y28172 , y28173 , y28174 , y28175 , y28176 , y28177 , y28178 , y28179 , y28180 , y28181 , y28182 , y28183 , y28184 , y28185 , y28186 , y28187 , y28188 , y28189 , y28190 , y28191 , y28192 , y28193 , y28194 , y28195 , y28196 , y28197 , y28198 , y28199 , y28200 , y28201 , y28202 , y28203 , y28204 , y28205 , y28206 , y28207 , y28208 , y28209 , y28210 , y28211 , y28212 , y28213 , y28214 , y28215 , y28216 , y28217 , y28218 , y28219 , y28220 , y28221 , y28222 , y28223 , y28224 , y28225 , y28226 , y28227 , y28228 , y28229 , y28230 , y28231 , y28232 , y28233 , y28234 , y28235 , y28236 , y28237 , y28238 , y28239 , y28240 , y28241 , y28242 , y28243 , y28244 , y28245 , y28246 , y28247 , y28248 , y28249 , y28250 , y28251 , y28252 , y28253 , y28254 , y28255 , y28256 , y28257 , y28258 , y28259 , y28260 , y28261 , y28262 , y28263 , y28264 , y28265 , y28266 , y28267 , y28268 , y28269 , y28270 , y28271 , y28272 , y28273 , y28274 , y28275 , y28276 , y28277 , y28278 , y28279 , y28280 , y28281 , y28282 , y28283 , y28284 , y28285 , y28286 , y28287 , y28288 , y28289 , y28290 , y28291 , y28292 , y28293 , y28294 , y28295 , y28296 , y28297 , y28298 , y28299 , y28300 , y28301 , y28302 , y28303 , y28304 , y28305 , y28306 , y28307 , y28308 , y28309 , y28310 , y28311 , y28312 , y28313 , y28314 , y28315 , y28316 , y28317 , y28318 , y28319 , y28320 , y28321 , y28322 , y28323 , y28324 , y28325 , y28326 , y28327 , y28328 , y28329 , y28330 , y28331 , y28332 , y28333 , y28334 , y28335 , y28336 , y28337 , y28338 , y28339 , y28340 , y28341 , y28342 , y28343 , y28344 , y28345 , y28346 , y28347 , y28348 , y28349 , y28350 , y28351 , y28352 , y28353 , y28354 , y28355 , y28356 , y28357 , y28358 , y28359 , y28360 , y28361 , y28362 , y28363 , y28364 , y28365 , y28366 , y28367 , y28368 , y28369 , y28370 , y28371 , y28372 , y28373 , y28374 , y28375 , y28376 , y28377 , y28378 , y28379 , y28380 , y28381 , y28382 , y28383 , y28384 , y28385 , y28386 , y28387 , y28388 , y28389 , y28390 , y28391 , y28392 , y28393 , y28394 , y28395 , y28396 , y28397 , y28398 , y28399 , y28400 , y28401 , y28402 , y28403 , y28404 , y28405 , y28406 , y28407 , y28408 , y28409 , y28410 , y28411 , y28412 , y28413 , y28414 , y28415 , y28416 , y28417 , y28418 , y28419 , y28420 , y28421 , y28422 , y28423 , y28424 , y28425 , y28426 , y28427 , y28428 , y28429 , y28430 , y28431 , y28432 , y28433 , y28434 , y28435 , y28436 , y28437 , y28438 , y28439 , y28440 , y28441 , y28442 , y28443 , y28444 , y28445 , y28446 , y28447 , y28448 , y28449 , y28450 , y28451 , y28452 , y28453 , y28454 , y28455 , y28456 , y28457 , y28458 , y28459 , y28460 , y28461 , y28462 , y28463 , y28464 , y28465 , y28466 , y28467 , y28468 , y28469 , y28470 , y28471 , y28472 , y28473 , y28474 , y28475 , y28476 , y28477 , y28478 , y28479 , y28480 , y28481 , y28482 , y28483 , y28484 , y28485 , y28486 , y28487 , y28488 , y28489 , y28490 , y28491 , y28492 , y28493 , y28494 , y28495 , y28496 , y28497 , y28498 , y28499 , y28500 , y28501 , y28502 , y28503 , y28504 , y28505 , y28506 , y28507 , y28508 , y28509 , y28510 , y28511 , y28512 , y28513 , y28514 , y28515 , y28516 , y28517 , y28518 , y28519 , y28520 , y28521 , y28522 , y28523 , y28524 , y28525 , y28526 , y28527 , y28528 , y28529 , y28530 , y28531 , y28532 , y28533 , y28534 , y28535 , y28536 , y28537 , y28538 , y28539 , y28540 , y28541 , y28542 , y28543 , y28544 , y28545 , y28546 , y28547 , y28548 , y28549 , y28550 , y28551 , y28552 , y28553 , y28554 , y28555 , y28556 , y28557 , y28558 , y28559 , y28560 , y28561 , y28562 , y28563 , y28564 , y28565 , y28566 , y28567 , y28568 , y28569 , y28570 , y28571 , y28572 , y28573 , y28574 , y28575 , y28576 , y28577 , y28578 , y28579 , y28580 , y28581 , y28582 , y28583 , y28584 , y28585 , y28586 , y28587 , y28588 , y28589 , y28590 , y28591 , y28592 , y28593 , y28594 , y28595 , y28596 , y28597 , y28598 , y28599 , y28600 , y28601 , y28602 , y28603 , y28604 , y28605 , y28606 , y28607 , y28608 , y28609 , y28610 , y28611 , y28612 , y28613 , y28614 , y28615 , y28616 , y28617 , y28618 , y28619 , y28620 , y28621 , y28622 , y28623 , y28624 , y28625 , y28626 , y28627 , y28628 , y28629 , y28630 , y28631 , y28632 , y28633 , y28634 , y28635 , y28636 , y28637 , y28638 , y28639 , y28640 , y28641 , y28642 , y28643 , y28644 , y28645 , y28646 , y28647 , y28648 , y28649 , y28650 , y28651 , y28652 , y28653 , y28654 , y28655 , y28656 , y28657 , y28658 , y28659 , y28660 , y28661 , y28662 , y28663 , y28664 , y28665 , y28666 , y28667 , y28668 , y28669 , y28670 , y28671 , y28672 , y28673 , y28674 , y28675 , y28676 , y28677 , y28678 , y28679 , y28680 , y28681 , y28682 , y28683 , y28684 , y28685 , y28686 , y28687 , y28688 , y28689 , y28690 , y28691 , y28692 , y28693 , y28694 , y28695 , y28696 , y28697 , y28698 , y28699 , y28700 , y28701 , y28702 , y28703 , y28704 , y28705 , y28706 , y28707 , y28708 , y28709 , y28710 , y28711 , y28712 , y28713 , y28714 , y28715 , y28716 , y28717 , y28718 , y28719 , y28720 , y28721 , y28722 , y28723 , y28724 , y28725 , y28726 , y28727 , y28728 , y28729 , y28730 , y28731 , y28732 , y28733 , y28734 , y28735 , y28736 , y28737 , y28738 , y28739 , y28740 , y28741 , y28742 , y28743 , y28744 , y28745 , y28746 , y28747 , y28748 , y28749 , y28750 , y28751 , y28752 , y28753 , y28754 , y28755 , y28756 , y28757 , y28758 , y28759 , y28760 , y28761 , y28762 , y28763 , y28764 , y28765 , y28766 , y28767 , y28768 , y28769 , y28770 , y28771 , y28772 , y28773 , y28774 , y28775 , y28776 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 ;
  assign n13 = ( x1 & ~x4 ) | ( x1 & x8 ) | ( ~x4 & x8 ) ;
  assign n14 = n13 ^ x0 ^ 1'b0 ;
  assign n15 = x1 & n14 ;
  assign n16 = ( x4 & x7 ) | ( x4 & ~x11 ) | ( x7 & ~x11 ) ;
  assign n19 = x3 & n15 ;
  assign n20 = n19 ^ n13 ^ 1'b0 ;
  assign n17 = x9 ^ x6 ^ 1'b0 ;
  assign n18 = x6 & n17 ;
  assign n21 = n20 ^ n18 ^ 1'b0 ;
  assign n22 = n16 & ~n21 ;
  assign n23 = ~x3 & x11 ;
  assign n32 = ( x6 & ~x10 ) | ( x6 & x11 ) | ( ~x10 & x11 ) ;
  assign n24 = x0 & x3 ;
  assign n25 = ~n18 & n24 ;
  assign n26 = n25 ^ n18 ^ n15 ;
  assign n27 = x11 & n18 ;
  assign n28 = n27 ^ x9 ^ 1'b0 ;
  assign n29 = n16 & ~n28 ;
  assign n30 = ~n26 & n29 ;
  assign n31 = x3 & ~n30 ;
  assign n33 = n32 ^ n31 ^ 1'b0 ;
  assign n35 = ( ~x2 & x3 ) | ( ~x2 & x5 ) | ( x3 & x5 ) ;
  assign n36 = x10 | n28 ;
  assign n37 = ( ~n22 & n35 ) | ( ~n22 & n36 ) | ( n35 & n36 ) ;
  assign n34 = x3 & n26 ;
  assign n38 = n37 ^ n34 ^ 1'b0 ;
  assign n39 = n37 ^ n20 ^ 1'b0 ;
  assign n40 = n25 ^ x4 ^ x2 ;
  assign n41 = n25 & n40 ;
  assign n42 = n41 ^ x6 ^ x0 ;
  assign n43 = n35 ^ x4 ^ 1'b0 ;
  assign n44 = n43 ^ x10 ^ x1 ;
  assign n45 = ~x7 & n41 ;
  assign n46 = ( x8 & n25 ) | ( x8 & ~n45 ) | ( n25 & ~n45 ) ;
  assign n47 = n37 & ~n45 ;
  assign n48 = n47 ^ n42 ^ 1'b0 ;
  assign n49 = n15 ^ x10 ^ x5 ;
  assign n50 = x5 & x9 ;
  assign n51 = n49 & n50 ;
  assign n52 = x5 & n47 ;
  assign n53 = n52 ^ n42 ^ 1'b0 ;
  assign n54 = n42 ^ n22 ^ x6 ;
  assign n55 = x3 & ~x10 ;
  assign n56 = n35 ^ x3 ^ 1'b0 ;
  assign n57 = x0 & n56 ;
  assign n58 = n18 & n57 ;
  assign n59 = ~n26 & n58 ;
  assign n60 = x10 & ~n59 ;
  assign n61 = ~n16 & n60 ;
  assign n62 = n20 ^ x11 ^ 1'b0 ;
  assign n63 = n49 ^ n33 ^ x6 ;
  assign n64 = n26 & n44 ;
  assign n65 = ~x9 & n64 ;
  assign n66 = n45 | n65 ;
  assign n67 = n66 ^ n43 ^ 1'b0 ;
  assign n68 = n67 ^ x5 ^ 1'b0 ;
  assign n69 = x8 & x9 ;
  assign n70 = n69 ^ n42 ^ 1'b0 ;
  assign n71 = x1 & n70 ;
  assign n72 = n28 & n71 ;
  assign n73 = n72 ^ n26 ^ 1'b0 ;
  assign n74 = n73 ^ n59 ^ n44 ;
  assign n75 = n63 ^ n22 ^ 1'b0 ;
  assign n76 = x11 & n51 ;
  assign n77 = x0 & n76 ;
  assign n78 = ~n16 & n77 ;
  assign n79 = n38 ^ x0 ^ 1'b0 ;
  assign n80 = n43 ^ n41 ^ x6 ;
  assign n81 = ~n23 & n80 ;
  assign n82 = n81 ^ n38 ^ 1'b0 ;
  assign n84 = n20 | n25 ;
  assign n83 = x0 & ~n42 ;
  assign n85 = n84 ^ n83 ^ 1'b0 ;
  assign n86 = n16 & ~n23 ;
  assign n87 = ~n37 & n86 ;
  assign n88 = n87 ^ n18 ^ 1'b0 ;
  assign n89 = n22 & ~n88 ;
  assign n90 = n18 & ~n49 ;
  assign n91 = n90 ^ n62 ^ 1'b0 ;
  assign n92 = ~n25 & n68 ;
  assign n93 = n36 & n92 ;
  assign n94 = n33 | n51 ;
  assign n95 = n94 ^ n28 ^ 1'b0 ;
  assign n96 = n95 ^ n93 ^ n63 ;
  assign n97 = ( x10 & n93 ) | ( x10 & ~n96 ) | ( n93 & ~n96 ) ;
  assign n98 = ~x10 & n35 ;
  assign n99 = n32 & ~n98 ;
  assign n100 = n59 ^ x7 ^ x6 ;
  assign n101 = n100 ^ x7 ^ 1'b0 ;
  assign n102 = ( ~x3 & n99 ) | ( ~x3 & n101 ) | ( n99 & n101 ) ;
  assign n104 = x0 | n20 ;
  assign n103 = ~n20 & n54 ;
  assign n105 = n104 ^ n103 ^ 1'b0 ;
  assign n106 = n65 ^ n55 ^ 1'b0 ;
  assign n107 = ~n42 & n106 ;
  assign n108 = ( x3 & n76 ) | ( x3 & n107 ) | ( n76 & n107 ) ;
  assign n109 = n63 ^ n41 ^ 1'b0 ;
  assign n110 = ( x6 & x8 ) | ( x6 & n32 ) | ( x8 & n32 ) ;
  assign n111 = n110 ^ n85 ^ 1'b0 ;
  assign n112 = n111 ^ n44 ^ 1'b0 ;
  assign n113 = n22 & n72 ;
  assign n114 = n57 & ~n93 ;
  assign n115 = ~n113 & n114 ;
  assign n116 = n115 ^ x3 ^ 1'b0 ;
  assign n117 = n75 | n116 ;
  assign n118 = n99 & n100 ;
  assign n119 = n96 | n112 ;
  assign n120 = x4 ^ x3 ^ 1'b0 ;
  assign n121 = x6 & n120 ;
  assign n122 = n121 ^ n55 ^ 1'b0 ;
  assign n123 = ~n61 & n122 ;
  assign n124 = ~n40 & n123 ;
  assign n125 = n124 ^ n96 ^ n95 ;
  assign n126 = n65 & n70 ;
  assign n127 = n32 ^ n16 ^ 1'b0 ;
  assign n128 = x10 & n127 ;
  assign n129 = n128 ^ n44 ^ 1'b0 ;
  assign n130 = ( n67 & ~n126 ) | ( n67 & n129 ) | ( ~n126 & n129 ) ;
  assign n131 = n51 | n59 ;
  assign n132 = ( n51 & n89 ) | ( n51 & ~n131 ) | ( n89 & ~n131 ) ;
  assign n133 = ~n25 & n46 ;
  assign n134 = n133 ^ n55 ^ 1'b0 ;
  assign n135 = ~x9 & n134 ;
  assign n136 = n45 ^ n25 ^ 1'b0 ;
  assign n137 = n38 & ~n104 ;
  assign n138 = n32 & n137 ;
  assign n139 = ~x9 & n138 ;
  assign n140 = n32 ^ x3 ^ 1'b0 ;
  assign n141 = x11 & n140 ;
  assign n142 = ( x6 & n112 ) | ( x6 & ~n141 ) | ( n112 & ~n141 ) ;
  assign n143 = n23 & ~n84 ;
  assign n144 = n143 ^ n33 ^ 1'b0 ;
  assign n145 = ~n124 & n144 ;
  assign n146 = n137 & n145 ;
  assign n147 = n43 & n146 ;
  assign n148 = x5 & n46 ;
  assign n149 = n148 ^ n93 ^ 1'b0 ;
  assign n150 = ( n55 & ~n135 ) | ( n55 & n149 ) | ( ~n135 & n149 ) ;
  assign n151 = ( n37 & n59 ) | ( n37 & ~n150 ) | ( n59 & ~n150 ) ;
  assign n152 = ( ~n20 & n63 ) | ( ~n20 & n89 ) | ( n63 & n89 ) ;
  assign n153 = n68 ^ n41 ^ 1'b0 ;
  assign n154 = n124 ^ n67 ^ 1'b0 ;
  assign n155 = ~n101 & n154 ;
  assign n156 = n155 ^ x10 ^ 1'b0 ;
  assign n157 = n43 ^ x7 ^ 1'b0 ;
  assign n158 = ( n111 & n121 ) | ( n111 & n157 ) | ( n121 & n157 ) ;
  assign n159 = n37 & ~n158 ;
  assign n160 = n16 & ~n45 ;
  assign n161 = n63 | n93 ;
  assign n162 = n161 ^ n143 ^ 1'b0 ;
  assign n163 = n162 ^ n79 ^ 1'b0 ;
  assign n164 = n160 & ~n163 ;
  assign n165 = n119 & n164 ;
  assign n166 = ~x4 & x8 ;
  assign n167 = n166 ^ n137 ^ 1'b0 ;
  assign n168 = ~n73 & n167 ;
  assign n169 = ( ~x4 & n108 ) | ( ~x4 & n168 ) | ( n108 & n168 ) ;
  assign n170 = n169 ^ n75 ^ 1'b0 ;
  assign n171 = ~n124 & n170 ;
  assign n172 = n171 ^ n43 ^ 1'b0 ;
  assign n173 = n142 ^ n43 ^ 1'b0 ;
  assign n174 = n141 & n173 ;
  assign n175 = n89 & ~n126 ;
  assign n176 = ~n82 & n175 ;
  assign n177 = n59 ^ x10 ^ 1'b0 ;
  assign n178 = n109 | n117 ;
  assign n179 = n178 ^ n102 ^ n44 ;
  assign n180 = ( x0 & n154 ) | ( x0 & n162 ) | ( n154 & n162 ) ;
  assign n181 = n101 & ~n180 ;
  assign n182 = n181 ^ n23 ^ 1'b0 ;
  assign n183 = n51 | n182 ;
  assign n184 = n61 ^ n32 ^ 1'b0 ;
  assign n185 = n101 | n184 ;
  assign n186 = n42 | n157 ;
  assign n187 = ~x3 & n186 ;
  assign n188 = ( n41 & n59 ) | ( n41 & n98 ) | ( n59 & n98 ) ;
  assign n189 = n125 | n188 ;
  assign n190 = n187 & ~n189 ;
  assign n191 = ( x2 & n62 ) | ( x2 & ~n186 ) | ( n62 & ~n186 ) ;
  assign n192 = n191 ^ n152 ^ 1'b0 ;
  assign n193 = n124 ^ n59 ^ 1'b0 ;
  assign n194 = n121 ^ n18 ^ x6 ;
  assign n195 = n193 & n194 ;
  assign n196 = n147 ^ x9 ^ 1'b0 ;
  assign n197 = n195 & ~n196 ;
  assign n204 = ~n150 & n164 ;
  assign n199 = n26 & ~n28 ;
  assign n200 = n67 & n199 ;
  assign n201 = n16 & n36 ;
  assign n202 = n200 | n201 ;
  assign n198 = n47 & n145 ;
  assign n203 = n202 ^ n198 ^ 1'b0 ;
  assign n205 = n204 ^ n203 ^ 1'b0 ;
  assign n206 = ~n99 & n127 ;
  assign n207 = n181 & ~n206 ;
  assign n208 = ~x1 & n207 ;
  assign n209 = n77 | n143 ;
  assign n210 = n209 ^ x8 ^ 1'b0 ;
  assign n211 = n204 ^ n98 ^ n47 ;
  assign n212 = n59 | n211 ;
  assign n213 = n169 | n212 ;
  assign n214 = n125 ^ n59 ^ 1'b0 ;
  assign n215 = n75 | n142 ;
  assign n216 = n147 & ~n215 ;
  assign n217 = ~n49 & n216 ;
  assign n218 = x9 | n95 ;
  assign n219 = n201 ^ n65 ^ 1'b0 ;
  assign n220 = n210 | n219 ;
  assign n221 = n101 ^ n53 ^ 1'b0 ;
  assign n222 = n221 ^ n112 ^ 1'b0 ;
  assign n223 = ~n97 & n115 ;
  assign n224 = ( n41 & n55 ) | ( n41 & n223 ) | ( n55 & n223 ) ;
  assign n225 = n119 ^ n33 ^ 1'b0 ;
  assign n226 = n141 ^ n44 ^ 1'b0 ;
  assign n227 = n226 ^ n41 ^ 1'b0 ;
  assign n228 = n47 & ~n227 ;
  assign n229 = n228 ^ n208 ^ 1'b0 ;
  assign n230 = ~n159 & n229 ;
  assign n231 = n51 ^ x10 ^ 1'b0 ;
  assign n233 = n187 ^ n108 ^ 1'b0 ;
  assign n234 = n141 & ~n233 ;
  assign n235 = ( x10 & n45 ) | ( x10 & ~n162 ) | ( n45 & ~n162 ) ;
  assign n236 = n234 & ~n235 ;
  assign n232 = n44 | n84 ;
  assign n237 = n236 ^ n232 ^ 1'b0 ;
  assign n238 = n231 & n237 ;
  assign n239 = ~n32 & n119 ;
  assign n240 = n239 ^ n13 ^ 1'b0 ;
  assign n241 = n240 ^ n190 ^ n40 ;
  assign n242 = n44 & ~n87 ;
  assign n243 = ( x3 & ~n13 ) | ( x3 & n132 ) | ( ~n13 & n132 ) ;
  assign n244 = n143 ^ n57 ^ 1'b0 ;
  assign n245 = n107 & ~n244 ;
  assign n246 = ( n44 & n100 ) | ( n44 & n245 ) | ( n100 & n245 ) ;
  assign n247 = n131 | n246 ;
  assign n248 = n82 & n247 ;
  assign n249 = n248 ^ n46 ^ 1'b0 ;
  assign n250 = n249 ^ n77 ^ 1'b0 ;
  assign n251 = x10 | n65 ;
  assign n252 = n37 | n251 ;
  assign n253 = n122 & n130 ;
  assign n254 = n253 ^ n159 ^ 1'b0 ;
  assign n255 = n119 & n147 ;
  assign n256 = n179 ^ n78 ^ n62 ;
  assign n257 = n89 & ~n246 ;
  assign n258 = n257 ^ n170 ^ 1'b0 ;
  assign n259 = n256 & n258 ;
  assign n260 = n16 ^ x5 ^ x4 ;
  assign n261 = n60 & n78 ;
  assign n262 = n98 | n101 ;
  assign n263 = n261 & ~n262 ;
  assign n264 = n263 ^ n250 ^ 1'b0 ;
  assign n265 = n131 | n264 ;
  assign n266 = n245 ^ n40 ^ 1'b0 ;
  assign n267 = n119 & n266 ;
  assign n268 = ~n226 & n259 ;
  assign n269 = ~n267 & n268 ;
  assign n270 = ~n36 & n194 ;
  assign n271 = n152 | n270 ;
  assign n272 = n271 ^ n129 ^ n102 ;
  assign n274 = n23 & ~n62 ;
  assign n275 = n191 & n274 ;
  assign n273 = n75 | n206 ;
  assign n276 = n275 ^ n273 ^ 1'b0 ;
  assign n277 = n39 | n87 ;
  assign n278 = n41 | n277 ;
  assign n279 = n154 & ~n278 ;
  assign n280 = n279 ^ n124 ^ x7 ;
  assign n281 = ~n276 & n280 ;
  assign n282 = n272 ^ n51 ^ 1'b0 ;
  assign n283 = ~n112 & n282 ;
  assign n286 = n49 | n63 ;
  assign n287 = n39 & ~n286 ;
  assign n284 = n111 ^ n108 ^ 1'b0 ;
  assign n285 = n72 | n284 ;
  assign n288 = n287 ^ n285 ^ 1'b0 ;
  assign n289 = ~n115 & n288 ;
  assign n290 = x11 & ~n183 ;
  assign n291 = n290 ^ n48 ^ 1'b0 ;
  assign n292 = n78 | n156 ;
  assign n293 = n59 & ~n292 ;
  assign n294 = ( n62 & n63 ) | ( n62 & n149 ) | ( n63 & n149 ) ;
  assign n303 = ~n23 & n38 ;
  assign n295 = n26 & n157 ;
  assign n296 = ~n246 & n295 ;
  assign n297 = n150 ^ n100 ^ 1'b0 ;
  assign n298 = x7 & n297 ;
  assign n299 = n298 ^ n181 ^ n53 ;
  assign n300 = n22 & ~n299 ;
  assign n301 = n300 ^ n263 ^ 1'b0 ;
  assign n302 = ~n296 & n301 ;
  assign n304 = n303 ^ n302 ^ 1'b0 ;
  assign n305 = ( n99 & n294 ) | ( n99 & n304 ) | ( n294 & n304 ) ;
  assign n306 = n294 ^ n98 ^ n59 ;
  assign n308 = n54 ^ n26 ^ 1'b0 ;
  assign n307 = n40 | n218 ;
  assign n309 = n308 ^ n307 ^ 1'b0 ;
  assign n310 = n270 ^ n67 ^ 1'b0 ;
  assign n311 = n174 ^ n77 ^ 1'b0 ;
  assign n312 = n310 & n311 ;
  assign n313 = x0 & ~n157 ;
  assign n314 = x10 & ~n275 ;
  assign n315 = n314 ^ n150 ^ 1'b0 ;
  assign n316 = ( x0 & n313 ) | ( x0 & n315 ) | ( n313 & n315 ) ;
  assign n317 = n127 & n316 ;
  assign n318 = n278 ^ n126 ^ n55 ;
  assign n319 = ~n177 & n318 ;
  assign n320 = n246 ^ n35 ^ 1'b0 ;
  assign n321 = n320 ^ n143 ^ 1'b0 ;
  assign n322 = x5 & n67 ;
  assign n323 = n49 | n87 ;
  assign n324 = n23 | n323 ;
  assign n325 = n119 & n324 ;
  assign n326 = n325 ^ n63 ^ 1'b0 ;
  assign n327 = n326 ^ x0 ^ 1'b0 ;
  assign n328 = n132 & n327 ;
  assign n329 = n38 | n328 ;
  assign n330 = n57 & ~n188 ;
  assign n331 = n285 & n330 ;
  assign n332 = n331 ^ n251 ^ 1'b0 ;
  assign n333 = n147 | n183 ;
  assign n334 = n333 ^ n164 ^ 1'b0 ;
  assign n335 = ~n177 & n334 ;
  assign n336 = n335 ^ n139 ^ 1'b0 ;
  assign n337 = n336 ^ n283 ^ 1'b0 ;
  assign n338 = n283 & n337 ;
  assign n339 = n254 ^ n95 ^ 1'b0 ;
  assign n340 = n256 & ~n339 ;
  assign n341 = n340 ^ n322 ^ 1'b0 ;
  assign n342 = n48 ^ n47 ^ n33 ;
  assign n343 = n225 ^ n44 ^ 1'b0 ;
  assign n344 = n36 & ~n343 ;
  assign n345 = n342 & n344 ;
  assign n346 = ( n15 & n180 ) | ( n15 & ~n324 ) | ( n180 & ~n324 ) ;
  assign n351 = n143 ^ n125 ^ 1'b0 ;
  assign n348 = n168 ^ n23 ^ 1'b0 ;
  assign n349 = n95 | n348 ;
  assign n347 = ~n126 & n256 ;
  assign n350 = n349 ^ n347 ^ 1'b0 ;
  assign n352 = n351 ^ n350 ^ 1'b0 ;
  assign n353 = ( n220 & n346 ) | ( n220 & n352 ) | ( n346 & n352 ) ;
  assign n354 = n150 ^ n48 ^ 1'b0 ;
  assign n355 = n354 ^ n51 ^ n38 ;
  assign n356 = n296 ^ n134 ^ 1'b0 ;
  assign n357 = n356 ^ n206 ^ 1'b0 ;
  assign n358 = x1 & ~n357 ;
  assign n372 = n110 ^ n23 ^ x3 ;
  assign n369 = x0 & n74 ;
  assign n370 = n22 & n165 ;
  assign n371 = n369 & n370 ;
  assign n361 = ( n48 & ~n206 ) | ( n48 & n231 ) | ( ~n206 & n231 ) ;
  assign n362 = n361 ^ n115 ^ 1'b0 ;
  assign n363 = n26 & ~n362 ;
  assign n364 = n231 & n363 ;
  assign n365 = n188 ^ n156 ^ 1'b0 ;
  assign n366 = ~n364 & n365 ;
  assign n359 = n166 ^ n26 ^ 1'b0 ;
  assign n360 = n79 & n359 ;
  assign n367 = n366 ^ n360 ^ 1'b0 ;
  assign n368 = n318 & n367 ;
  assign n373 = n372 ^ n371 ^ n368 ;
  assign n374 = n174 & ~n346 ;
  assign n375 = n179 ^ n80 ^ 1'b0 ;
  assign n376 = n375 ^ n214 ^ 1'b0 ;
  assign n377 = n169 & n304 ;
  assign n378 = ~n350 & n377 ;
  assign n379 = ( ~n303 & n376 ) | ( ~n303 & n378 ) | ( n376 & n378 ) ;
  assign n380 = n188 ^ n48 ^ 1'b0 ;
  assign n381 = ~n231 & n380 ;
  assign n382 = n381 ^ n111 ^ 1'b0 ;
  assign n383 = n263 | n382 ;
  assign n384 = n221 ^ n217 ^ x4 ;
  assign n385 = n383 | n384 ;
  assign n386 = n385 ^ x0 ^ 1'b0 ;
  assign n387 = n344 ^ x9 ^ 1'b0 ;
  assign n388 = ~n222 & n387 ;
  assign n389 = n328 ^ n159 ^ 1'b0 ;
  assign n390 = n13 & ~n389 ;
  assign n391 = n226 ^ n197 ^ 1'b0 ;
  assign n392 = n55 | n391 ;
  assign n393 = n304 & ~n355 ;
  assign n394 = n393 ^ n115 ^ 1'b0 ;
  assign n395 = x1 & ~n59 ;
  assign n396 = ~n145 & n395 ;
  assign n397 = n396 ^ n283 ^ 1'b0 ;
  assign n398 = n246 & ~n397 ;
  assign n399 = ~n111 & n246 ;
  assign n400 = n398 & n399 ;
  assign n401 = n340 | n400 ;
  assign n402 = n231 ^ n183 ^ 1'b0 ;
  assign n403 = n100 & n402 ;
  assign n404 = n285 ^ n23 ^ 1'b0 ;
  assign n405 = n169 & ~n404 ;
  assign n406 = n405 ^ x4 ^ 1'b0 ;
  assign n407 = n137 ^ n107 ^ 1'b0 ;
  assign n408 = ~n95 & n407 ;
  assign n409 = n408 ^ n324 ^ n91 ;
  assign n414 = ( ~n97 & n102 ) | ( ~n97 & n188 ) | ( n102 & n188 ) ;
  assign n410 = n74 | n315 ;
  assign n411 = n125 & ~n410 ;
  assign n412 = n240 & ~n411 ;
  assign n413 = ~n275 & n412 ;
  assign n415 = n414 ^ n413 ^ 1'b0 ;
  assign n416 = x10 | n44 ;
  assign n417 = n204 ^ n201 ^ x1 ;
  assign n418 = n91 & n313 ;
  assign n419 = n203 ^ n158 ^ 1'b0 ;
  assign n420 = n418 & n419 ;
  assign n421 = ( n33 & n412 ) | ( n33 & ~n420 ) | ( n412 & ~n420 ) ;
  assign n422 = n254 & ~n272 ;
  assign n423 = ~n301 & n422 ;
  assign n424 = n179 & ~n238 ;
  assign n425 = n49 ^ n45 ^ 1'b0 ;
  assign n426 = ~n28 & n425 ;
  assign n427 = n228 & n426 ;
  assign n428 = n427 ^ n23 ^ 1'b0 ;
  assign n429 = n74 | n204 ;
  assign n430 = n429 ^ n145 ^ 1'b0 ;
  assign n431 = n430 ^ n326 ^ 1'b0 ;
  assign n432 = n154 ^ n61 ^ 1'b0 ;
  assign n433 = n224 & n432 ;
  assign n434 = n433 ^ n194 ^ 1'b0 ;
  assign n435 = n434 ^ n241 ^ n55 ;
  assign n436 = n44 & n178 ;
  assign n437 = n289 ^ n91 ^ 1'b0 ;
  assign n438 = x6 & n369 ;
  assign n439 = n139 | n185 ;
  assign n442 = n41 & ~n77 ;
  assign n443 = n97 ^ n53 ^ x8 ;
  assign n444 = n443 ^ n313 ^ 1'b0 ;
  assign n445 = n442 & ~n444 ;
  assign n440 = n107 ^ x3 ^ 1'b0 ;
  assign n441 = n440 ^ n77 ^ 1'b0 ;
  assign n446 = n445 ^ n441 ^ 1'b0 ;
  assign n447 = ~n51 & n177 ;
  assign n448 = n226 ^ n37 ^ 1'b0 ;
  assign n449 = n237 & n448 ;
  assign n450 = n449 ^ n261 ^ 1'b0 ;
  assign n451 = n450 ^ n220 ^ 1'b0 ;
  assign n452 = n451 ^ n113 ^ 1'b0 ;
  assign n453 = n320 ^ n51 ^ 1'b0 ;
  assign n454 = x10 & ~n95 ;
  assign n455 = n454 ^ x0 ^ 1'b0 ;
  assign n456 = n102 | n112 ;
  assign n457 = n455 & ~n456 ;
  assign n458 = n457 ^ n179 ^ 1'b0 ;
  assign n459 = n458 ^ x3 ^ 1'b0 ;
  assign n462 = n32 & n164 ;
  assign n460 = n287 ^ n15 ^ 1'b0 ;
  assign n461 = n217 | n460 ;
  assign n463 = n462 ^ n461 ^ n80 ;
  assign n464 = n74 | n283 ;
  assign n465 = n185 ^ n135 ^ n105 ;
  assign n466 = n465 ^ n63 ^ 1'b0 ;
  assign n467 = n102 ^ n51 ^ 1'b0 ;
  assign n468 = n32 & ~n51 ;
  assign n469 = n468 ^ n36 ^ 1'b0 ;
  assign n470 = n440 ^ n234 ^ 1'b0 ;
  assign n471 = n190 | n470 ;
  assign n472 = n44 & ~n122 ;
  assign n473 = n472 ^ n75 ^ 1'b0 ;
  assign n474 = ~n471 & n473 ;
  assign n475 = n474 ^ n202 ^ 1'b0 ;
  assign n476 = n96 ^ x5 ^ 1'b0 ;
  assign n477 = n475 & n476 ;
  assign n478 = n417 & ~n477 ;
  assign n479 = n158 & ~n383 ;
  assign n480 = n479 ^ x1 ^ 1'b0 ;
  assign n481 = n350 & n480 ;
  assign n483 = n283 ^ n63 ^ 1'b0 ;
  assign n482 = n141 & n352 ;
  assign n484 = n483 ^ n482 ^ 1'b0 ;
  assign n485 = ~x0 & n340 ;
  assign n486 = ( ~x4 & n256 ) | ( ~x4 & n351 ) | ( n256 & n351 ) ;
  assign n489 = ~n185 & n237 ;
  assign n490 = n489 ^ n59 ^ 1'b0 ;
  assign n491 = ( n72 & n224 ) | ( n72 & n490 ) | ( n224 & n490 ) ;
  assign n487 = ~n63 & n306 ;
  assign n488 = n45 & n487 ;
  assign n492 = n491 ^ n488 ^ 1'b0 ;
  assign n493 = ( x9 & n191 ) | ( x9 & ~n492 ) | ( n191 & ~n492 ) ;
  assign n494 = n486 & ~n493 ;
  assign n495 = ~n112 & n195 ;
  assign n496 = n495 ^ n53 ^ 1'b0 ;
  assign n497 = n496 ^ n184 ^ 1'b0 ;
  assign n498 = ~n492 & n497 ;
  assign n499 = n149 ^ n107 ^ 1'b0 ;
  assign n500 = x9 & n319 ;
  assign n501 = n76 ^ n57 ^ 1'b0 ;
  assign n502 = n37 & ~n501 ;
  assign n503 = n57 ^ x10 ^ 1'b0 ;
  assign n504 = n41 & n503 ;
  assign n505 = n504 ^ n231 ^ 1'b0 ;
  assign n509 = n218 ^ n55 ^ 1'b0 ;
  assign n510 = n109 & n509 ;
  assign n506 = n102 ^ n26 ^ 1'b0 ;
  assign n507 = n152 & n506 ;
  assign n508 = ~n40 & n507 ;
  assign n511 = n510 ^ n508 ^ n91 ;
  assign n512 = n505 & ~n511 ;
  assign n513 = n218 & n512 ;
  assign n514 = n252 ^ n251 ^ n119 ;
  assign n515 = n23 & n514 ;
  assign n516 = n35 & ~n74 ;
  assign n517 = n184 & n516 ;
  assign n518 = n265 | n517 ;
  assign n519 = ( n241 & n488 ) | ( n241 & ~n518 ) | ( n488 & ~n518 ) ;
  assign n520 = n38 & n157 ;
  assign n521 = ~n432 & n520 ;
  assign n522 = n130 & ~n521 ;
  assign n523 = ~n464 & n522 ;
  assign n524 = n210 ^ n33 ^ 1'b0 ;
  assign n525 = n350 & ~n524 ;
  assign n526 = x11 & ~n471 ;
  assign n527 = n526 ^ n36 ^ 1'b0 ;
  assign n528 = ~n93 & n527 ;
  assign n529 = ~n525 & n528 ;
  assign n530 = n129 & ~n484 ;
  assign n531 = n206 ^ n102 ^ 1'b0 ;
  assign n532 = n44 & n531 ;
  assign n533 = ( n321 & ~n332 ) | ( n321 & n443 ) | ( ~n332 & n443 ) ;
  assign n534 = n40 & n462 ;
  assign n535 = ~n355 & n534 ;
  assign n536 = n535 ^ n149 ^ 1'b0 ;
  assign n537 = n105 & ~n536 ;
  assign n538 = n537 ^ n450 ^ 1'b0 ;
  assign n539 = n139 ^ x9 ^ 1'b0 ;
  assign n540 = n539 ^ n272 ^ 1'b0 ;
  assign n541 = ~n231 & n540 ;
  assign n542 = n541 ^ n536 ^ 1'b0 ;
  assign n543 = n224 ^ n23 ^ n15 ;
  assign n544 = n543 ^ n486 ^ 1'b0 ;
  assign n545 = ~n55 & n318 ;
  assign n546 = n344 ^ n65 ^ 1'b0 ;
  assign n547 = n141 | n546 ;
  assign n548 = n188 ^ n23 ^ 1'b0 ;
  assign n549 = n441 ^ n426 ^ 1'b0 ;
  assign n550 = ~n548 & n549 ;
  assign n551 = n550 ^ n334 ^ n22 ;
  assign n552 = n536 ^ n127 ^ 1'b0 ;
  assign n553 = n551 | n552 ;
  assign n554 = ( n236 & n430 ) | ( n236 & ~n462 ) | ( n430 & ~n462 ) ;
  assign n555 = n41 & ~n222 ;
  assign n556 = ~n186 & n555 ;
  assign n557 = n372 ^ n36 ^ 1'b0 ;
  assign n558 = n46 & n225 ;
  assign n559 = n558 ^ n283 ^ 1'b0 ;
  assign n560 = n341 & ~n559 ;
  assign n561 = n547 ^ n263 ^ n201 ;
  assign n562 = n298 ^ n15 ^ 1'b0 ;
  assign n563 = ~n294 & n562 ;
  assign n564 = n411 ^ n129 ^ n118 ;
  assign n565 = n168 & ~n272 ;
  assign n566 = n565 ^ n192 ^ 1'b0 ;
  assign n567 = ( n202 & n564 ) | ( n202 & ~n566 ) | ( n564 & ~n566 ) ;
  assign n568 = n16 & n567 ;
  assign n569 = n568 ^ n164 ^ 1'b0 ;
  assign n570 = x6 & n364 ;
  assign n571 = ~n181 & n570 ;
  assign n572 = n480 | n485 ;
  assign n573 = n572 ^ n415 ^ 1'b0 ;
  assign n574 = n571 & n573 ;
  assign n577 = ( n40 & ~n70 ) | ( n40 & n234 ) | ( ~n70 & n234 ) ;
  assign n576 = n375 ^ x10 ^ 1'b0 ;
  assign n575 = n119 ^ x3 ^ 1'b0 ;
  assign n578 = n577 ^ n576 ^ n575 ;
  assign n579 = n278 & n532 ;
  assign n580 = n579 ^ n177 ^ 1'b0 ;
  assign n581 = n200 ^ n107 ^ 1'b0 ;
  assign n582 = n53 | n581 ;
  assign n583 = n341 ^ n242 ^ 1'b0 ;
  assign n584 = n443 & n583 ;
  assign n585 = ~n582 & n584 ;
  assign n586 = x0 & ~n548 ;
  assign n587 = ( n539 & n585 ) | ( n539 & n586 ) | ( n585 & n586 ) ;
  assign n588 = ( n177 & ~n279 ) | ( n177 & n346 ) | ( ~n279 & n346 ) ;
  assign n589 = n254 & ~n396 ;
  assign n590 = n589 ^ n44 ^ 1'b0 ;
  assign n591 = n424 ^ n336 ^ 1'b0 ;
  assign n592 = ~n61 & n591 ;
  assign n593 = n592 ^ n78 ^ 1'b0 ;
  assign n594 = n499 ^ x3 ^ 1'b0 ;
  assign n595 = n415 ^ n101 ^ 1'b0 ;
  assign n596 = ~n423 & n595 ;
  assign n597 = ~n46 & n596 ;
  assign n599 = n77 & ~n411 ;
  assign n600 = n599 ^ n331 ^ 1'b0 ;
  assign n598 = n350 ^ n91 ^ n74 ;
  assign n601 = n600 ^ n598 ^ 1'b0 ;
  assign n602 = x10 & n192 ;
  assign n603 = ~n197 & n602 ;
  assign n604 = ~n597 & n603 ;
  assign n605 = n142 & ~n435 ;
  assign n606 = n372 | n513 ;
  assign n607 = n324 | n606 ;
  assign n608 = ~n149 & n607 ;
  assign n609 = n183 | n534 ;
  assign n610 = n37 & n609 ;
  assign n611 = n610 ^ n230 ^ 1'b0 ;
  assign n612 = n143 | n450 ;
  assign n613 = n195 & ~n211 ;
  assign n614 = n613 ^ n205 ^ 1'b0 ;
  assign n615 = ( n32 & n242 ) | ( n32 & n308 ) | ( n242 & n308 ) ;
  assign n616 = n614 & ~n615 ;
  assign n617 = n517 & n616 ;
  assign n618 = n46 & n57 ;
  assign n619 = n618 ^ n98 ^ 1'b0 ;
  assign n620 = n213 | n349 ;
  assign n621 = n620 ^ n201 ^ 1'b0 ;
  assign n622 = n67 | n435 ;
  assign n623 = ~n621 & n622 ;
  assign n624 = n623 ^ n209 ^ 1'b0 ;
  assign n625 = n624 ^ n45 ^ 1'b0 ;
  assign n626 = n619 & n625 ;
  assign n627 = n626 ^ n588 ^ n319 ;
  assign n628 = n566 ^ n39 ^ 1'b0 ;
  assign n629 = n588 ^ n132 ^ n40 ;
  assign n630 = n236 | n362 ;
  assign n631 = n156 | n160 ;
  assign n632 = n91 | n631 ;
  assign n633 = n630 | n632 ;
  assign n634 = ~n398 & n622 ;
  assign n635 = n634 ^ n577 ^ 1'b0 ;
  assign n636 = n427 & ~n635 ;
  assign n637 = n261 & ~n263 ;
  assign n638 = n313 | n637 ;
  assign n639 = n638 ^ n319 ^ 1'b0 ;
  assign n640 = ~n466 & n639 ;
  assign n641 = n147 ^ n68 ^ 1'b0 ;
  assign n643 = n457 ^ n152 ^ 1'b0 ;
  assign n644 = n234 & ~n643 ;
  assign n642 = n384 | n621 ;
  assign n645 = n644 ^ n642 ^ 1'b0 ;
  assign n646 = ( x10 & n40 ) | ( x10 & n490 ) | ( n40 & n490 ) ;
  assign n647 = ~n453 & n646 ;
  assign n648 = n93 & n334 ;
  assign n649 = ( n381 & ~n469 ) | ( n381 & n648 ) | ( ~n469 & n648 ) ;
  assign n650 = ~n596 & n649 ;
  assign n654 = n68 | n112 ;
  assign n651 = n503 ^ n152 ^ 1'b0 ;
  assign n652 = ~n59 & n651 ;
  assign n653 = n37 & n652 ;
  assign n655 = n654 ^ n653 ^ 1'b0 ;
  assign n656 = n655 ^ n312 ^ 1'b0 ;
  assign n657 = n33 & n77 ;
  assign n658 = n168 & ~n657 ;
  assign n659 = n658 ^ n112 ^ 1'b0 ;
  assign n660 = n659 ^ n469 ^ 1'b0 ;
  assign n661 = n532 & n660 ;
  assign n665 = n143 ^ n68 ^ 1'b0 ;
  assign n662 = n181 ^ n44 ^ 1'b0 ;
  assign n663 = n201 ^ n44 ^ 1'b0 ;
  assign n664 = ( n44 & n662 ) | ( n44 & n663 ) | ( n662 & n663 ) ;
  assign n666 = n665 ^ n664 ^ 1'b0 ;
  assign n667 = n105 & ~n397 ;
  assign n668 = ( n281 & ~n532 ) | ( n281 & n667 ) | ( ~n532 & n667 ) ;
  assign n669 = ~n513 & n527 ;
  assign n670 = ~x10 & n669 ;
  assign n681 = n217 ^ x3 ^ 1'b0 ;
  assign n682 = n313 | n681 ;
  assign n683 = n132 | n682 ;
  assign n684 = n683 ^ n548 ^ 1'b0 ;
  assign n677 = ~n421 & n486 ;
  assign n678 = n677 ^ n220 ^ 1'b0 ;
  assign n679 = n678 ^ n278 ^ 1'b0 ;
  assign n680 = ~n272 & n679 ;
  assign n671 = ~n162 & n381 ;
  assign n672 = ~n194 & n671 ;
  assign n673 = n417 & ~n672 ;
  assign n674 = n275 & n673 ;
  assign n675 = n139 | n674 ;
  assign n676 = n675 ^ n361 ^ 1'b0 ;
  assign n685 = n684 ^ n680 ^ n676 ;
  assign n686 = n61 & n203 ;
  assign n687 = n448 ^ n151 ^ 1'b0 ;
  assign n688 = n686 | n687 ;
  assign n689 = n506 & n545 ;
  assign n690 = n689 ^ n63 ^ 1'b0 ;
  assign n691 = n75 | n164 ;
  assign n692 = n220 ^ n154 ^ 1'b0 ;
  assign n693 = n91 & ~n147 ;
  assign n694 = n693 ^ n152 ^ 1'b0 ;
  assign n695 = n576 & ~n694 ;
  assign n696 = n318 & n695 ;
  assign n697 = n696 ^ n659 ^ n260 ;
  assign n698 = n245 ^ n179 ^ 1'b0 ;
  assign n699 = ~n226 & n503 ;
  assign n700 = n414 & n699 ;
  assign n701 = n700 ^ n247 ^ 1'b0 ;
  assign n702 = n109 & ~n701 ;
  assign n703 = n113 & n534 ;
  assign n704 = ~x7 & n703 ;
  assign n705 = ( n306 & ~n473 ) | ( n306 & n694 ) | ( ~n473 & n694 ) ;
  assign n706 = ( n524 & n704 ) | ( n524 & n705 ) | ( n704 & n705 ) ;
  assign n707 = n251 ^ x9 ^ 1'b0 ;
  assign n708 = ( n169 & n306 ) | ( n169 & n707 ) | ( n306 & n707 ) ;
  assign n709 = n646 ^ n269 ^ n36 ;
  assign n710 = n46 & ~n709 ;
  assign n711 = n291 ^ n112 ^ x0 ;
  assign n712 = n63 & n525 ;
  assign n713 = ( n355 & ~n711 ) | ( n355 & n712 ) | ( ~n711 & n712 ) ;
  assign n714 = x8 & n713 ;
  assign n715 = ~n30 & n99 ;
  assign n716 = n715 ^ n285 ^ 1'b0 ;
  assign n717 = n493 ^ n231 ^ 1'b0 ;
  assign n718 = n688 & ~n717 ;
  assign n719 = ( n368 & ~n716 ) | ( n368 & n718 ) | ( ~n716 & n718 ) ;
  assign n720 = n477 ^ n68 ^ 1'b0 ;
  assign n721 = n686 ^ n526 ^ 1'b0 ;
  assign n722 = n228 | n721 ;
  assign n723 = n567 & n722 ;
  assign n724 = n532 & ~n576 ;
  assign n725 = n724 ^ n74 ^ 1'b0 ;
  assign n726 = ( n102 & n723 ) | ( n102 & n725 ) | ( n723 & n725 ) ;
  assign n728 = n177 ^ n121 ^ 1'b0 ;
  assign n727 = n446 & n583 ;
  assign n729 = n728 ^ n727 ^ n139 ;
  assign n730 = n666 ^ n601 ^ 1'b0 ;
  assign n731 = n115 & n519 ;
  assign n732 = n731 ^ n153 ^ 1'b0 ;
  assign n733 = n360 & ~n732 ;
  assign n734 = n42 & ~n139 ;
  assign n735 = n688 & ~n734 ;
  assign n736 = n448 ^ n102 ^ 1'b0 ;
  assign n737 = n37 & ~n315 ;
  assign n738 = n737 ^ n170 ^ 1'b0 ;
  assign n739 = n738 ^ x10 ^ 1'b0 ;
  assign n740 = ~n131 & n142 ;
  assign n741 = n467 | n672 ;
  assign n742 = n741 ^ n223 ^ n40 ;
  assign n743 = n177 | n200 ;
  assign n744 = n743 ^ n548 ^ 1'b0 ;
  assign n745 = n396 & ~n744 ;
  assign n746 = n745 ^ n255 ^ 1'b0 ;
  assign n747 = n197 & n746 ;
  assign n748 = n493 & n747 ;
  assign n749 = n748 ^ n318 ^ 1'b0 ;
  assign n750 = n108 & ~n641 ;
  assign n751 = n432 & n727 ;
  assign n752 = n147 & n751 ;
  assign n753 = n469 ^ n436 ^ 1'b0 ;
  assign n754 = n589 & n753 ;
  assign n755 = ( n403 & ~n431 ) | ( n403 & n754 ) | ( ~n431 & n754 ) ;
  assign n756 = n63 ^ n37 ^ 1'b0 ;
  assign n758 = n35 & ~n548 ;
  assign n759 = n758 ^ n57 ^ 1'b0 ;
  assign n757 = x6 & n178 ;
  assign n760 = n759 ^ n757 ^ 1'b0 ;
  assign n761 = n760 ^ n548 ^ x10 ;
  assign n765 = n33 | n190 ;
  assign n762 = n318 ^ n102 ^ 1'b0 ;
  assign n763 = n384 ^ n202 ^ x0 ;
  assign n764 = n762 | n763 ;
  assign n766 = n765 ^ n764 ^ n181 ;
  assign n767 = n178 ^ n93 ^ x6 ;
  assign n768 = ~n44 & n767 ;
  assign n769 = n768 ^ n127 ^ 1'b0 ;
  assign n770 = n527 ^ n25 ^ 1'b0 ;
  assign n771 = n431 & ~n770 ;
  assign n772 = n345 & n368 ;
  assign n773 = n772 ^ n655 ^ 1'b0 ;
  assign n774 = n42 & ~n349 ;
  assign n775 = ~n608 & n774 ;
  assign n776 = n773 & n775 ;
  assign n777 = n680 & ~n755 ;
  assign n778 = n344 ^ n168 ^ 1'b0 ;
  assign n779 = n57 & n778 ;
  assign n780 = ( ~n100 & n435 ) | ( ~n100 & n779 ) | ( n435 & n779 ) ;
  assign n781 = n37 & n432 ;
  assign n782 = n781 ^ n299 ^ 1'b0 ;
  assign n783 = n782 ^ n156 ^ 1'b0 ;
  assign n784 = n352 & ~n783 ;
  assign n785 = n784 ^ n63 ^ 1'b0 ;
  assign n786 = n636 | n785 ;
  assign n787 = n786 ^ n435 ^ n72 ;
  assign n791 = n135 ^ n87 ^ 1'b0 ;
  assign n792 = ( n36 & ~n63 ) | ( n36 & n791 ) | ( ~n63 & n791 ) ;
  assign n788 = n145 & n306 ;
  assign n789 = n788 ^ n682 ^ 1'b0 ;
  assign n790 = n426 | n789 ;
  assign n793 = n792 ^ n790 ^ 1'b0 ;
  assign n794 = n77 & ~n793 ;
  assign n798 = ~n62 & n728 ;
  assign n799 = n798 ^ n534 ^ 1'b0 ;
  assign n795 = n299 ^ x10 ^ 1'b0 ;
  assign n796 = n381 & ~n795 ;
  assign n797 = n796 ^ n392 ^ 1'b0 ;
  assign n800 = n799 ^ n797 ^ n313 ;
  assign n801 = n415 ^ n310 ^ n209 ;
  assign n802 = ~n716 & n801 ;
  assign n803 = ~n211 & n416 ;
  assign n804 = n506 & ~n524 ;
  assign n805 = n312 | n320 ;
  assign n806 = n805 ^ n195 ^ 1'b0 ;
  assign n807 = n383 ^ n345 ^ 1'b0 ;
  assign n808 = n806 & n807 ;
  assign n809 = ( ~n165 & n426 ) | ( ~n165 & n589 ) | ( n426 & n589 ) ;
  assign n810 = n82 | n809 ;
  assign n811 = n810 ^ n105 ^ 1'b0 ;
  assign n812 = n139 | n332 ;
  assign n813 = n165 | n812 ;
  assign n814 = n263 | n813 ;
  assign n815 = ~n28 & n644 ;
  assign n816 = n48 & n815 ;
  assign n817 = n627 | n816 ;
  assign n818 = ~x10 & n178 ;
  assign n819 = n818 ^ n678 ^ 1'b0 ;
  assign n821 = n614 & n648 ;
  assign n822 = n821 ^ n525 ^ 1'b0 ;
  assign n820 = n577 & ~n593 ;
  assign n823 = n822 ^ n820 ^ 1'b0 ;
  assign n824 = n440 & n823 ;
  assign n825 = ( n246 & n439 ) | ( n246 & ~n637 ) | ( n439 & ~n637 ) ;
  assign n826 = n825 ^ n188 ^ n168 ;
  assign n827 = n180 & ~n826 ;
  assign n828 = n283 & ~n379 ;
  assign n829 = ~n827 & n828 ;
  assign n830 = n829 ^ n324 ^ 1'b0 ;
  assign n832 = n46 & ~n440 ;
  assign n833 = ~n241 & n832 ;
  assign n834 = n833 ^ n646 ^ 1'b0 ;
  assign n831 = ~n98 & n105 ;
  assign n835 = n834 ^ n831 ^ 1'b0 ;
  assign n836 = ~n830 & n835 ;
  assign n837 = n110 & n587 ;
  assign n838 = ( n241 & n496 ) | ( n241 & ~n704 ) | ( n496 & ~n704 ) ;
  assign n839 = ( n513 & ~n649 ) | ( n513 & n838 ) | ( ~n649 & n838 ) ;
  assign n840 = n839 ^ n174 ^ 1'b0 ;
  assign n841 = n283 & ~n840 ;
  assign n842 = ~n65 & n200 ;
  assign n843 = n842 ^ n641 ^ 1'b0 ;
  assign n844 = n320 | n843 ;
  assign n845 = n346 ^ n122 ^ 1'b0 ;
  assign n846 = n667 ^ n453 ^ n276 ;
  assign n847 = n63 | n299 ;
  assign n848 = n442 | n847 ;
  assign n849 = n848 ^ n459 ^ n341 ;
  assign n850 = n37 & ~n849 ;
  assign n851 = n738 & n850 ;
  assign n852 = ~n725 & n851 ;
  assign n853 = n99 & ~n170 ;
  assign n854 = ~n375 & n853 ;
  assign n858 = n445 & n614 ;
  assign n859 = n858 ^ n127 ^ 1'b0 ;
  assign n855 = n250 & ~n426 ;
  assign n856 = n26 & n255 ;
  assign n857 = n855 & n856 ;
  assign n860 = n859 ^ n857 ^ 1'b0 ;
  assign n861 = n356 ^ x11 ^ 1'b0 ;
  assign n862 = n587 ^ n350 ^ 1'b0 ;
  assign n863 = n388 & ~n862 ;
  assign n865 = n168 ^ n39 ^ 1'b0 ;
  assign n864 = n166 ^ n153 ^ 1'b0 ;
  assign n866 = n865 ^ n864 ^ 1'b0 ;
  assign n867 = n213 ^ n115 ^ 1'b0 ;
  assign n868 = n496 | n867 ;
  assign n869 = n484 ^ n73 ^ 1'b0 ;
  assign n870 = x0 & n869 ;
  assign n871 = ~n790 & n870 ;
  assign n872 = n154 & ~n435 ;
  assign n873 = n872 ^ n430 ^ 1'b0 ;
  assign n874 = n263 | n451 ;
  assign n875 = n873 & ~n874 ;
  assign n876 = ( ~n186 & n203 ) | ( ~n186 & n269 ) | ( n203 & n269 ) ;
  assign n877 = n245 | n876 ;
  assign n878 = n600 ^ n125 ^ 1'b0 ;
  assign n879 = n304 & n878 ;
  assign n880 = n41 & ~n276 ;
  assign n881 = n880 ^ n466 ^ 1'b0 ;
  assign n882 = n478 ^ n428 ^ n59 ;
  assign n883 = n882 ^ n825 ^ 1'b0 ;
  assign n884 = n186 | n883 ;
  assign n887 = n127 ^ n113 ^ 1'b0 ;
  assign n888 = n575 & ~n887 ;
  assign n885 = n585 ^ n475 ^ n350 ;
  assign n886 = n885 ^ n835 ^ x1 ;
  assign n889 = n888 ^ n886 ^ n51 ;
  assign n890 = n491 ^ n353 ^ n41 ;
  assign n891 = n184 & ~n211 ;
  assign n893 = n159 | n598 ;
  assign n894 = ~n369 & n664 ;
  assign n895 = ~n169 & n894 ;
  assign n896 = x2 & ~n895 ;
  assign n897 = ~n420 & n896 ;
  assign n898 = n893 | n897 ;
  assign n899 = n898 ^ n141 ^ 1'b0 ;
  assign n892 = ~x10 & n118 ;
  assign n900 = n899 ^ n892 ^ 1'b0 ;
  assign n901 = n51 | n829 ;
  assign n902 = n901 ^ n126 ^ 1'b0 ;
  assign n903 = n355 | n397 ;
  assign n904 = n118 & ~n797 ;
  assign n905 = ~n44 & n904 ;
  assign n906 = ~n214 & n270 ;
  assign n907 = n47 & ~n183 ;
  assign n908 = n694 & n907 ;
  assign n909 = n908 ^ n773 ^ n713 ;
  assign n910 = n506 ^ n412 ^ 1'b0 ;
  assign n911 = n181 & ~n190 ;
  assign n912 = n525 & n911 ;
  assign n913 = n912 ^ n23 ^ 1'b0 ;
  assign n914 = ~n461 & n913 ;
  assign n915 = ~n910 & n914 ;
  assign n917 = n96 & ~n156 ;
  assign n918 = ~n767 & n917 ;
  assign n916 = n855 ^ n412 ^ n298 ;
  assign n919 = n918 ^ n916 ^ 1'b0 ;
  assign n920 = n728 & ~n919 ;
  assign n921 = ~n712 & n920 ;
  assign n922 = n91 | n496 ;
  assign n923 = n543 ^ n494 ^ 1'b0 ;
  assign n924 = n923 ^ n349 ^ 1'b0 ;
  assign n925 = n840 & n924 ;
  assign n926 = n61 & n481 ;
  assign n927 = n441 & n514 ;
  assign n928 = ( n160 & ~n763 ) | ( n160 & n927 ) | ( ~n763 & n927 ) ;
  assign n929 = n928 ^ n338 ^ 1'b0 ;
  assign n930 = n152 & ~n705 ;
  assign n931 = n930 ^ n257 ^ 1'b0 ;
  assign n933 = n744 ^ n601 ^ 1'b0 ;
  assign n932 = n252 | n631 ;
  assign n934 = n933 ^ n932 ^ 1'b0 ;
  assign n935 = n475 | n511 ;
  assign n936 = n935 ^ n532 ^ 1'b0 ;
  assign n937 = ~n686 & n936 ;
  assign n938 = ~n506 & n937 ;
  assign n939 = n126 ^ n33 ^ 1'b0 ;
  assign n940 = ~n59 & n939 ;
  assign n941 = ( ~n130 & n221 ) | ( ~n130 & n940 ) | ( n221 & n940 ) ;
  assign n942 = n637 | n941 ;
  assign n943 = n544 & ~n548 ;
  assign n944 = n942 & n943 ;
  assign n945 = ~n388 & n443 ;
  assign n946 = n578 ^ n405 ^ 1'b0 ;
  assign n947 = n841 ^ n648 ^ n309 ;
  assign n948 = n139 & ~n345 ;
  assign n949 = n948 ^ n416 ^ n397 ;
  assign n953 = ( n42 & n401 ) | ( n42 & ~n471 ) | ( n401 & ~n471 ) ;
  assign n951 = n418 ^ n267 ^ 1'b0 ;
  assign n952 = n918 | n951 ;
  assign n954 = n953 ^ n952 ^ 1'b0 ;
  assign n950 = n38 | n269 ;
  assign n955 = n954 ^ n950 ^ 1'b0 ;
  assign n956 = n955 ^ n137 ^ 1'b0 ;
  assign n957 = n876 | n956 ;
  assign n958 = n791 ^ n690 ^ n372 ;
  assign n959 = n33 & n928 ;
  assign n961 = ( n28 & n272 ) | ( n28 & n334 ) | ( n272 & n334 ) ;
  assign n960 = n41 & ~n374 ;
  assign n962 = n961 ^ n960 ^ n209 ;
  assign n963 = n962 ^ n833 ^ n650 ;
  assign n964 = n63 & n395 ;
  assign n965 = n255 & n964 ;
  assign n966 = n965 ^ n38 ^ 1'b0 ;
  assign n967 = n716 & n761 ;
  assign n968 = n967 ^ n329 ^ 1'b0 ;
  assign n969 = n166 & n411 ;
  assign n970 = n85 & ~n895 ;
  assign n971 = n970 ^ n124 ^ 1'b0 ;
  assign n972 = n928 & n938 ;
  assign n973 = n971 & n972 ;
  assign n974 = n861 & n892 ;
  assign n975 = ~x0 & n644 ;
  assign n976 = n164 | n961 ;
  assign n983 = n665 ^ n183 ^ 1'b0 ;
  assign n981 = n469 ^ n280 ^ 1'b0 ;
  assign n982 = ~n51 & n981 ;
  assign n984 = n983 ^ n982 ^ 1'b0 ;
  assign n977 = n82 & n760 ;
  assign n978 = n977 ^ n876 ^ n510 ;
  assign n979 = n63 & ~n978 ;
  assign n980 = n566 & n979 ;
  assign n985 = n984 ^ n982 ^ n980 ;
  assign n986 = n166 & ~n816 ;
  assign n987 = n986 ^ n539 ^ 1'b0 ;
  assign n988 = n260 | n830 ;
  assign n989 = n542 & ~n988 ;
  assign n990 = ( ~n469 & n987 ) | ( ~n469 & n989 ) | ( n987 & n989 ) ;
  assign n991 = n63 | n176 ;
  assign n992 = n873 ^ n23 ^ 1'b0 ;
  assign n993 = ~n249 & n992 ;
  assign n994 = n465 ^ n48 ^ 1'b0 ;
  assign n995 = ~n663 & n680 ;
  assign n996 = n690 & ~n995 ;
  assign n997 = n415 ^ n51 ^ 1'b0 ;
  assign n998 = n668 | n839 ;
  assign n1000 = n524 & ~n918 ;
  assign n1001 = ( ~n44 & n767 ) | ( ~n44 & n1000 ) | ( n767 & n1000 ) ;
  assign n999 = n281 ^ n223 ^ n35 ;
  assign n1002 = n1001 ^ n999 ^ 1'b0 ;
  assign n1003 = n885 & n1002 ;
  assign n1004 = n864 ^ n446 ^ 1'b0 ;
  assign n1005 = n303 ^ n157 ^ 1'b0 ;
  assign n1006 = n51 | n1005 ;
  assign n1007 = n1006 ^ n441 ^ n126 ;
  assign n1008 = x10 & ~n1007 ;
  assign n1009 = n1008 ^ n406 ^ 1'b0 ;
  assign n1010 = n648 ^ n39 ^ 1'b0 ;
  assign n1011 = n1010 ^ n63 ^ 1'b0 ;
  assign n1012 = n117 ^ n46 ^ 1'b0 ;
  assign n1013 = n42 | n1012 ;
  assign n1014 = n1013 ^ n279 ^ 1'b0 ;
  assign n1015 = n1011 & ~n1014 ;
  assign n1016 = n867 ^ n269 ^ 1'b0 ;
  assign n1017 = ~n1001 & n1016 ;
  assign n1018 = ( n111 & n191 ) | ( n111 & n1017 ) | ( n191 & n1017 ) ;
  assign n1020 = ~n74 & n346 ;
  assign n1021 = ~n1017 & n1020 ;
  assign n1022 = ~n51 & n1021 ;
  assign n1019 = n953 ^ n464 ^ 1'b0 ;
  assign n1023 = n1022 ^ n1019 ^ 1'b0 ;
  assign n1024 = n739 ^ n563 ^ 1'b0 ;
  assign n1025 = n818 ^ n124 ^ 1'b0 ;
  assign n1026 = ~n352 & n649 ;
  assign n1027 = ~n484 & n1026 ;
  assign n1028 = n1027 ^ n28 ^ 1'b0 ;
  assign n1029 = n762 ^ n521 ^ 1'b0 ;
  assign n1030 = n806 ^ n666 ^ 1'b0 ;
  assign n1031 = n955 ^ n20 ^ 1'b0 ;
  assign n1032 = n1031 ^ n421 ^ 1'b0 ;
  assign n1033 = ~n533 & n578 ;
  assign n1034 = n224 & n491 ;
  assign n1035 = n1034 ^ n36 ^ 1'b0 ;
  assign n1036 = n541 ^ n437 ^ 1'b0 ;
  assign n1037 = n1035 | n1036 ;
  assign n1038 = n432 ^ n80 ^ n59 ;
  assign n1039 = n270 & n1038 ;
  assign n1040 = ( n313 & n637 ) | ( n313 & n762 ) | ( n637 & n762 ) ;
  assign n1041 = ~n867 & n1040 ;
  assign n1042 = n250 & ~n1041 ;
  assign n1043 = n627 & n1042 ;
  assign n1044 = n376 | n1043 ;
  assign n1045 = n1044 ^ n686 ^ 1'b0 ;
  assign n1046 = ~n1039 & n1045 ;
  assign n1047 = ( n241 & ~n395 ) | ( n241 & n502 ) | ( ~n395 & n502 ) ;
  assign n1048 = n1047 ^ n324 ^ 1'b0 ;
  assign n1049 = n756 & ~n819 ;
  assign n1050 = n548 ^ n356 ^ 1'b0 ;
  assign n1051 = n628 ^ x3 ^ 1'b0 ;
  assign n1052 = ~n20 & n668 ;
  assign n1053 = n320 ^ n200 ^ 1'b0 ;
  assign n1054 = ~n850 & n1053 ;
  assign n1055 = n525 & ~n1054 ;
  assign n1056 = ~n82 & n711 ;
  assign n1057 = n328 & n1056 ;
  assign n1058 = n1057 ^ n834 ^ 1'b0 ;
  assign n1059 = n842 & n1058 ;
  assign n1060 = ~n1055 & n1059 ;
  assign n1061 = n216 & n590 ;
  assign n1062 = n1061 ^ n824 ^ 1'b0 ;
  assign n1063 = n1026 ^ n462 ^ n39 ;
  assign n1064 = n1063 ^ n977 ^ n374 ;
  assign n1065 = n118 & ~n265 ;
  assign n1066 = n1065 ^ n503 ^ 1'b0 ;
  assign n1067 = n463 & ~n1066 ;
  assign n1068 = ~n483 & n1067 ;
  assign n1069 = n864 ^ n259 ^ 1'b0 ;
  assign n1070 = n249 & n1069 ;
  assign n1071 = n1070 ^ n756 ^ 1'b0 ;
  assign n1072 = ~n275 & n711 ;
  assign n1073 = ( n63 & n139 ) | ( n63 & ~n371 ) | ( n139 & ~n371 ) ;
  assign n1074 = n1073 ^ n816 ^ 1'b0 ;
  assign n1075 = n644 & n1074 ;
  assign n1076 = ~n181 & n589 ;
  assign n1077 = n22 & ~n1076 ;
  assign n1078 = n478 & n1077 ;
  assign n1079 = ( n923 & n1075 ) | ( n923 & n1078 ) | ( n1075 & n1078 ) ;
  assign n1082 = n609 ^ n500 ^ 1'b0 ;
  assign n1080 = n30 & n132 ;
  assign n1081 = n1080 ^ n1035 ^ 1'b0 ;
  assign n1083 = n1082 ^ n1081 ^ 1'b0 ;
  assign n1084 = n220 & n250 ;
  assign n1085 = ( n46 & n201 ) | ( n46 & ~n390 ) | ( n201 & ~n390 ) ;
  assign n1086 = n884 ^ n469 ^ 1'b0 ;
  assign n1087 = n1085 & ~n1086 ;
  assign n1088 = n213 & n324 ;
  assign n1089 = x2 & n1088 ;
  assign n1090 = ( n794 & n874 ) | ( n794 & n918 ) | ( n874 & n918 ) ;
  assign n1091 = ~n398 & n728 ;
  assign n1092 = ~n435 & n1091 ;
  assign n1093 = ( n542 & n614 ) | ( n542 & ~n1092 ) | ( n614 & ~n1092 ) ;
  assign n1094 = n596 | n686 ;
  assign n1095 = n1094 ^ n121 ^ 1'b0 ;
  assign n1096 = ~n210 & n1095 ;
  assign n1097 = n1096 ^ n741 ^ 1'b0 ;
  assign n1103 = n147 | n563 ;
  assign n1098 = ~n217 & n532 ;
  assign n1099 = n1098 ^ n75 ^ 1'b0 ;
  assign n1100 = n329 & ~n1099 ;
  assign n1101 = n1100 ^ n104 ^ 1'b0 ;
  assign n1102 = ~n112 & n1101 ;
  assign n1104 = n1103 ^ n1102 ^ n51 ;
  assign n1105 = ~n734 & n969 ;
  assign n1106 = ~n187 & n903 ;
  assign n1107 = n1106 ^ n271 ^ 1'b0 ;
  assign n1108 = n37 & ~n604 ;
  assign n1109 = n194 | n601 ;
  assign n1110 = n511 & n1109 ;
  assign n1111 = n329 & ~n890 ;
  assign n1112 = n1111 ^ n570 ^ 1'b0 ;
  assign n1113 = n688 & ~n1112 ;
  assign n1114 = ~n417 & n1113 ;
  assign n1115 = ( ~n762 & n1110 ) | ( ~n762 & n1114 ) | ( n1110 & n1114 ) ;
  assign n1116 = ~n358 & n644 ;
  assign n1117 = ~n115 & n409 ;
  assign n1118 = n427 & n1117 ;
  assign n1119 = n1118 ^ n177 ^ 1'b0 ;
  assign n1120 = n929 & ~n1119 ;
  assign n1121 = n131 ^ n63 ^ 1'b0 ;
  assign n1122 = n940 & n1121 ;
  assign n1123 = n694 ^ n209 ^ 1'b0 ;
  assign n1124 = n1017 & ~n1123 ;
  assign n1125 = ~n457 & n855 ;
  assign n1126 = n1125 ^ n48 ^ 1'b0 ;
  assign n1127 = ( n445 & ~n1124 ) | ( n445 & n1126 ) | ( ~n1124 & n1126 ) ;
  assign n1128 = n238 | n635 ;
  assign n1129 = n1128 ^ n637 ^ 1'b0 ;
  assign n1130 = n955 | n1129 ;
  assign n1131 = n1130 ^ n678 ^ 1'b0 ;
  assign n1132 = n55 & ~n293 ;
  assign n1133 = ~n570 & n1132 ;
  assign n1134 = n1133 ^ n550 ^ n226 ;
  assign n1135 = n717 & n1134 ;
  assign n1136 = n108 & ~n954 ;
  assign n1137 = ~x9 & n1136 ;
  assign n1138 = ( ~n572 & n709 ) | ( ~n572 & n1137 ) | ( n709 & n1137 ) ;
  assign n1139 = n451 & ~n472 ;
  assign n1140 = n1139 ^ n672 ^ 1'b0 ;
  assign n1141 = n685 ^ n654 ^ 1'b0 ;
  assign n1142 = n1140 | n1141 ;
  assign n1143 = n231 & ~n759 ;
  assign n1144 = n1143 ^ n204 ^ 1'b0 ;
  assign n1145 = ~n667 & n1144 ;
  assign n1146 = n220 | n769 ;
  assign n1147 = n464 | n1146 ;
  assign n1148 = n640 & n645 ;
  assign n1149 = ( n441 & n841 ) | ( n441 & ~n1148 ) | ( n841 & ~n1148 ) ;
  assign n1150 = n676 ^ n551 ^ n490 ;
  assign n1151 = ( n283 & n650 ) | ( n283 & n888 ) | ( n650 & n888 ) ;
  assign n1152 = n1151 ^ n384 ^ 1'b0 ;
  assign n1153 = n589 & ~n1152 ;
  assign n1154 = n688 ^ n371 ^ n362 ;
  assign n1155 = ~n1114 & n1154 ;
  assign n1156 = n1155 ^ n332 ^ 1'b0 ;
  assign n1157 = n784 & ~n795 ;
  assign n1158 = n263 | n461 ;
  assign n1159 = n80 | n1158 ;
  assign n1160 = n1159 ^ n646 ^ 1'b0 ;
  assign n1161 = ~n1157 & n1160 ;
  assign n1162 = ~n842 & n1161 ;
  assign n1163 = n80 & n806 ;
  assign n1164 = ~n1153 & n1163 ;
  assign n1165 = n41 & n105 ;
  assign n1166 = n1165 ^ n782 ^ 1'b0 ;
  assign n1167 = n833 & ~n1166 ;
  assign n1168 = n1167 ^ n826 ^ n747 ;
  assign n1169 = n791 & ~n1168 ;
  assign n1170 = n459 & n1169 ;
  assign n1171 = n445 ^ n408 ^ 1'b0 ;
  assign n1172 = n238 | n384 ;
  assign n1173 = n1058 & ~n1172 ;
  assign n1174 = n154 ^ n51 ^ 1'b0 ;
  assign n1175 = n42 | n1174 ;
  assign n1176 = n1175 ^ n206 ^ n110 ;
  assign n1177 = ~n688 & n835 ;
  assign n1178 = ( ~x0 & n41 ) | ( ~x0 & n223 ) | ( n41 & n223 ) ;
  assign n1179 = n1178 ^ n593 ^ n334 ;
  assign n1180 = n839 & n1179 ;
  assign n1181 = ( n1176 & n1177 ) | ( n1176 & ~n1180 ) | ( n1177 & ~n1180 ) ;
  assign n1182 = n63 & n477 ;
  assign n1183 = n626 & n1082 ;
  assign n1184 = ~n508 & n865 ;
  assign n1185 = n1184 ^ n709 ^ n596 ;
  assign n1186 = ( n403 & ~n816 ) | ( n403 & n1185 ) | ( ~n816 & n1185 ) ;
  assign n1187 = n1186 ^ n829 ^ 1'b0 ;
  assign n1188 = n37 & ~n1187 ;
  assign n1189 = n1013 ^ n209 ^ n23 ;
  assign n1190 = ~n935 & n1189 ;
  assign n1191 = n1190 ^ n870 ^ 1'b0 ;
  assign n1192 = n561 | n1191 ;
  assign n1193 = n1192 ^ n844 ^ x8 ;
  assign n1194 = n32 & n1109 ;
  assign n1195 = ~n550 & n1194 ;
  assign n1196 = n710 ^ n676 ^ 1'b0 ;
  assign n1197 = ( n97 & n941 ) | ( n97 & ~n1196 ) | ( n941 & ~n1196 ) ;
  assign n1198 = ( n310 & n1195 ) | ( n310 & n1197 ) | ( n1195 & n1197 ) ;
  assign n1199 = n181 ^ n77 ^ 1'b0 ;
  assign n1200 = ~n1073 & n1199 ;
  assign n1201 = ( n865 & n868 ) | ( n865 & n1200 ) | ( n868 & n1200 ) ;
  assign n1202 = n1201 ^ n1177 ^ n287 ;
  assign n1203 = n267 & n922 ;
  assign n1204 = n1203 ^ n926 ^ 1'b0 ;
  assign n1205 = n121 & ~n502 ;
  assign n1206 = n1205 ^ n130 ^ 1'b0 ;
  assign n1207 = ~n684 & n1206 ;
  assign n1208 = n1207 ^ n309 ^ 1'b0 ;
  assign n1209 = x0 & ~n1208 ;
  assign n1210 = n844 ^ n332 ^ 1'b0 ;
  assign n1212 = n259 & ~n849 ;
  assign n1213 = n1212 ^ n1088 ^ 1'b0 ;
  assign n1211 = n666 & ~n1167 ;
  assign n1214 = n1213 ^ n1211 ^ 1'b0 ;
  assign n1215 = n1214 ^ n518 ^ 1'b0 ;
  assign n1216 = ~n1000 & n1215 ;
  assign n1217 = n301 & n1216 ;
  assign n1218 = n1217 ^ n208 ^ 1'b0 ;
  assign n1220 = n57 | n720 ;
  assign n1219 = n353 & ~n607 ;
  assign n1221 = n1220 ^ n1219 ^ 1'b0 ;
  assign n1222 = n1218 & ~n1221 ;
  assign n1223 = n822 & n1222 ;
  assign n1224 = n152 & ~n226 ;
  assign n1225 = n895 & n1224 ;
  assign n1226 = n1225 ^ n263 ^ 1'b0 ;
  assign n1227 = ~n665 & n794 ;
  assign n1228 = n1227 ^ n1019 ^ 1'b0 ;
  assign n1229 = n1228 ^ n209 ^ 1'b0 ;
  assign n1230 = ~n822 & n1229 ;
  assign n1231 = n726 | n1124 ;
  assign n1232 = n1231 ^ n975 ^ 1'b0 ;
  assign n1233 = n834 | n1088 ;
  assign n1234 = n310 & ~n445 ;
  assign n1235 = n1234 ^ n1050 ^ 1'b0 ;
  assign n1236 = n93 | n416 ;
  assign n1237 = n1236 ^ n160 ^ 1'b0 ;
  assign n1238 = n1237 ^ n384 ^ 1'b0 ;
  assign n1239 = n397 & ~n1133 ;
  assign n1240 = n299 & n1239 ;
  assign n1241 = n317 & ~n1240 ;
  assign n1242 = n918 & n1241 ;
  assign n1243 = ~n711 & n1242 ;
  assign n1244 = n369 | n1243 ;
  assign n1245 = n1103 ^ n334 ^ 1'b0 ;
  assign n1246 = n592 ^ n411 ^ 1'b0 ;
  assign n1247 = n1063 ^ n379 ^ n371 ;
  assign n1248 = x10 | n1247 ;
  assign n1249 = n941 ^ n855 ^ n596 ;
  assign n1250 = n1248 & ~n1249 ;
  assign n1251 = ( n408 & ~n1246 ) | ( n408 & n1250 ) | ( ~n1246 & n1250 ) ;
  assign n1252 = n32 | n44 ;
  assign n1253 = n100 | n1252 ;
  assign n1254 = n344 & n1253 ;
  assign n1255 = ~n875 & n1254 ;
  assign n1256 = n174 ^ n23 ^ 1'b0 ;
  assign n1257 = n633 & ~n1256 ;
  assign n1258 = n1257 ^ n551 ^ 1'b0 ;
  assign n1259 = ~n755 & n772 ;
  assign n1260 = n1259 ^ n414 ^ 1'b0 ;
  assign n1261 = n1221 & n1260 ;
  assign n1262 = n263 | n577 ;
  assign n1263 = n742 ^ n299 ^ 1'b0 ;
  assign n1264 = n581 ^ n364 ^ n33 ;
  assign n1265 = n469 ^ n97 ^ 1'b0 ;
  assign n1266 = n524 & ~n1265 ;
  assign n1267 = ~n1264 & n1266 ;
  assign n1268 = n1183 | n1267 ;
  assign n1269 = n376 & ~n1268 ;
  assign n1270 = n1263 & ~n1269 ;
  assign n1275 = n321 ^ n59 ^ 1'b0 ;
  assign n1276 = ~n654 & n1275 ;
  assign n1271 = n356 ^ n54 ^ 1'b0 ;
  assign n1272 = ~n373 & n1271 ;
  assign n1273 = n1272 ^ n586 ^ 1'b0 ;
  assign n1274 = n600 & n1273 ;
  assign n1277 = n1276 ^ n1274 ^ n303 ;
  assign n1278 = n349 ^ n230 ^ 1'b0 ;
  assign n1279 = ( n442 & n1256 ) | ( n442 & ~n1278 ) | ( n1256 & ~n1278 ) ;
  assign n1280 = ( n160 & n517 ) | ( n160 & ~n637 ) | ( n517 & ~n637 ) ;
  assign n1281 = n1280 ^ n788 ^ n210 ;
  assign n1282 = n1281 ^ n1189 ^ 1'b0 ;
  assign n1283 = ( n183 & n769 ) | ( n183 & ~n1282 ) | ( n769 & ~n1282 ) ;
  assign n1284 = n1274 & ~n1283 ;
  assign n1285 = n1284 ^ n728 ^ 1'b0 ;
  assign n1286 = ~n527 & n1237 ;
  assign n1290 = ~n500 & n722 ;
  assign n1287 = n445 ^ n315 ^ n61 ;
  assign n1288 = ( n67 & ~n183 ) | ( n67 & n473 ) | ( ~n183 & n473 ) ;
  assign n1289 = ( ~n222 & n1287 ) | ( ~n222 & n1288 ) | ( n1287 & n1288 ) ;
  assign n1291 = n1290 ^ n1289 ^ 1'b0 ;
  assign n1292 = n1286 | n1291 ;
  assign n1293 = n1292 ^ n710 ^ 1'b0 ;
  assign n1297 = n801 | n965 ;
  assign n1298 = n1297 ^ n293 ^ 1'b0 ;
  assign n1299 = n1298 ^ n324 ^ 1'b0 ;
  assign n1300 = n341 & ~n1299 ;
  assign n1294 = n906 ^ n893 ^ n473 ;
  assign n1295 = ~n576 & n1076 ;
  assign n1296 = ~n1294 & n1295 ;
  assign n1301 = n1300 ^ n1296 ^ 1'b0 ;
  assign n1302 = ~n214 & n1301 ;
  assign n1303 = n37 & ~n729 ;
  assign n1304 = ~n319 & n1303 ;
  assign n1305 = n1304 ^ n159 ^ 1'b0 ;
  assign n1306 = n440 | n711 ;
  assign n1307 = n1305 | n1306 ;
  assign n1308 = n344 & ~n1153 ;
  assign n1309 = n1195 ^ n752 ^ 1'b0 ;
  assign n1310 = n624 & ~n890 ;
  assign n1311 = ( x10 & ~n80 ) | ( x10 & n672 ) | ( ~n80 & n672 ) ;
  assign n1312 = n1311 ^ n467 ^ n234 ;
  assign n1313 = ~n1310 & n1312 ;
  assign n1314 = n603 & n1313 ;
  assign n1315 = n164 & ~n624 ;
  assign n1316 = n221 | n1315 ;
  assign n1317 = n885 ^ n686 ^ 1'b0 ;
  assign n1318 = n1198 ^ n991 ^ 1'b0 ;
  assign n1319 = ~n374 & n604 ;
  assign n1320 = n585 & ~n1319 ;
  assign n1321 = n1320 ^ n733 ^ 1'b0 ;
  assign n1322 = n1318 | n1321 ;
  assign n1323 = ~n102 & n356 ;
  assign n1324 = n772 & n1323 ;
  assign n1325 = n1324 ^ n192 ^ 1'b0 ;
  assign n1326 = n1154 | n1325 ;
  assign n1327 = n556 | n1326 ;
  assign n1328 = ~n667 & n1243 ;
  assign n1329 = n162 ^ n156 ^ 1'b0 ;
  assign n1330 = n1329 ^ x8 ^ 1'b0 ;
  assign n1331 = n637 ^ n162 ^ 1'b0 ;
  assign n1332 = n1094 & n1331 ;
  assign n1334 = n40 | n152 ;
  assign n1333 = n53 & ~n1175 ;
  assign n1335 = n1334 ^ n1333 ^ 1'b0 ;
  assign n1336 = n1335 ^ n1195 ^ 1'b0 ;
  assign n1337 = n344 ^ n322 ^ 1'b0 ;
  assign n1338 = ~n1177 & n1288 ;
  assign n1339 = ~n368 & n1338 ;
  assign n1340 = n224 ^ n113 ^ 1'b0 ;
  assign n1341 = n1037 & n1340 ;
  assign n1342 = n126 | n819 ;
  assign n1343 = n1342 ^ n298 ^ 1'b0 ;
  assign n1344 = n1159 ^ n89 ^ 1'b0 ;
  assign n1345 = n1344 ^ n859 ^ n183 ;
  assign n1346 = n1345 ^ n846 ^ 1'b0 ;
  assign n1347 = n791 ^ n437 ^ 1'b0 ;
  assign n1348 = n428 & ~n1347 ;
  assign n1351 = n44 | n135 ;
  assign n1352 = n805 & ~n1351 ;
  assign n1353 = n587 & n1352 ;
  assign n1349 = n23 | n87 ;
  assign n1350 = x7 | n1349 ;
  assign n1354 = n1353 ^ n1350 ^ 1'b0 ;
  assign n1355 = n1348 & ~n1354 ;
  assign n1358 = n13 & ~n753 ;
  assign n1359 = n1358 ^ n842 ^ 1'b0 ;
  assign n1360 = n414 & ~n1359 ;
  assign n1357 = n137 & ~n431 ;
  assign n1361 = n1360 ^ n1357 ^ 1'b0 ;
  assign n1356 = n250 & n848 ;
  assign n1362 = n1361 ^ n1356 ^ 1'b0 ;
  assign n1363 = ( n619 & n1287 ) | ( n619 & n1362 ) | ( n1287 & n1362 ) ;
  assign n1364 = ~n276 & n972 ;
  assign n1365 = n1364 ^ n308 ^ 1'b0 ;
  assign n1366 = n513 | n893 ;
  assign n1367 = n257 & ~n1366 ;
  assign n1368 = ~n1359 & n1367 ;
  assign n1369 = n141 | n190 ;
  assign n1370 = n1369 ^ n1139 ^ 1'b0 ;
  assign n1371 = n1370 ^ n764 ^ 1'b0 ;
  assign n1372 = n897 ^ n63 ^ 1'b0 ;
  assign n1373 = n432 & ~n1372 ;
  assign n1374 = ~n575 & n1373 ;
  assign n1375 = n674 | n686 ;
  assign n1376 = n1375 ^ n355 ^ 1'b0 ;
  assign n1377 = n874 ^ n534 ^ 1'b0 ;
  assign n1378 = n63 | n1377 ;
  assign n1379 = n1376 | n1378 ;
  assign n1380 = n1379 ^ x10 ^ 1'b0 ;
  assign n1381 = n1374 | n1380 ;
  assign n1382 = n521 & ~n1381 ;
  assign n1383 = ( n711 & n1080 ) | ( n711 & ~n1196 ) | ( n1080 & ~n1196 ) ;
  assign n1384 = n172 & n228 ;
  assign n1385 = n1384 ^ n276 ^ 1'b0 ;
  assign n1386 = x4 & ~n1385 ;
  assign n1387 = ( n39 & n612 ) | ( n39 & ~n1386 ) | ( n612 & ~n1386 ) ;
  assign n1388 = n428 & ~n1387 ;
  assign n1389 = ~n55 & n1388 ;
  assign n1390 = n1278 & ~n1389 ;
  assign n1391 = n745 & n1390 ;
  assign n1392 = n791 & n947 ;
  assign n1393 = n1290 & n1392 ;
  assign n1394 = ~n211 & n301 ;
  assign n1395 = n1394 ^ n115 ^ 1'b0 ;
  assign n1396 = n478 | n1395 ;
  assign n1397 = n1393 & ~n1396 ;
  assign n1398 = n241 & n409 ;
  assign n1399 = n1398 ^ n100 ^ 1'b0 ;
  assign n1400 = ( ~n706 & n998 ) | ( ~n706 & n1399 ) | ( n998 & n1399 ) ;
  assign n1401 = x3 & ~n837 ;
  assign n1402 = n289 ^ n20 ^ 1'b0 ;
  assign n1403 = n508 ^ n503 ^ 1'b0 ;
  assign n1404 = n426 ^ n225 ^ 1'b0 ;
  assign n1405 = n1011 & ~n1404 ;
  assign n1406 = n1405 ^ n922 ^ n682 ;
  assign n1407 = ( n35 & ~n523 ) | ( n35 & n829 ) | ( ~n523 & n829 ) ;
  assign n1408 = n358 ^ n328 ^ 1'b0 ;
  assign n1409 = n1407 & ~n1408 ;
  assign n1410 = n1409 ^ n808 ^ n39 ;
  assign n1411 = n1410 ^ n1389 ^ n749 ;
  assign n1412 = n1411 ^ n82 ^ 1'b0 ;
  assign n1413 = n1336 & ~n1412 ;
  assign n1414 = n1104 & n1413 ;
  assign n1415 = n136 & ~n176 ;
  assign n1416 = n521 & n1415 ;
  assign n1417 = n1402 ^ n445 ^ 1'b0 ;
  assign n1418 = n1151 & ~n1417 ;
  assign n1419 = n408 & ~n1213 ;
  assign n1420 = n738 & n1419 ;
  assign n1421 = ~n659 & n1420 ;
  assign n1422 = n720 | n884 ;
  assign n1423 = n523 & ~n1422 ;
  assign n1424 = ( ~n698 & n1110 ) | ( ~n698 & n1168 ) | ( n1110 & n1168 ) ;
  assign n1425 = n1424 ^ n283 ^ 1'b0 ;
  assign n1426 = n1121 ^ n884 ^ 1'b0 ;
  assign n1427 = ( n371 & n628 ) | ( n371 & n1056 ) | ( n628 & n1056 ) ;
  assign n1428 = n36 & n762 ;
  assign n1429 = ( n911 & n999 ) | ( n911 & n1428 ) | ( n999 & n1428 ) ;
  assign n1430 = n1429 ^ n903 ^ 1'b0 ;
  assign n1431 = ~n1427 & n1430 ;
  assign n1432 = n803 & ~n1133 ;
  assign n1433 = n109 & n1432 ;
  assign n1434 = n525 & n1433 ;
  assign n1435 = ~n910 & n1434 ;
  assign n1436 = ( n165 & n1294 ) | ( n165 & ~n1311 ) | ( n1294 & ~n1311 ) ;
  assign n1437 = ~n298 & n1436 ;
  assign n1438 = n1094 ^ n54 ^ 1'b0 ;
  assign n1439 = ~n65 & n1438 ;
  assign n1440 = n1439 ^ n1272 ^ 1'b0 ;
  assign n1441 = n572 & n1440 ;
  assign n1442 = n529 & n1441 ;
  assign n1443 = n1442 ^ n1309 ^ 1'b0 ;
  assign n1452 = n132 & ~n392 ;
  assign n1453 = n1452 ^ n1214 ^ 1'b0 ;
  assign n1451 = n206 | n615 ;
  assign n1454 = n1453 ^ n1451 ^ 1'b0 ;
  assign n1444 = n121 & n283 ;
  assign n1445 = n316 ^ n57 ^ 1'b0 ;
  assign n1446 = n291 & ~n1445 ;
  assign n1447 = ( ~n296 & n888 ) | ( ~n296 & n1446 ) | ( n888 & n1446 ) ;
  assign n1448 = n1447 ^ n411 ^ 1'b0 ;
  assign n1449 = n676 | n1448 ;
  assign n1450 = n1444 | n1449 ;
  assign n1455 = n1454 ^ n1450 ^ n830 ;
  assign n1456 = n281 & ~n813 ;
  assign n1457 = n1131 ^ n764 ^ 1'b0 ;
  assign n1461 = n131 | n893 ;
  assign n1458 = n98 | n514 ;
  assign n1459 = x10 | n1458 ;
  assign n1460 = ~n408 & n1459 ;
  assign n1462 = n1461 ^ n1460 ^ n1426 ;
  assign n1463 = n803 ^ n499 ^ n211 ;
  assign n1464 = n1463 ^ n379 ^ 1'b0 ;
  assign n1465 = n383 & n457 ;
  assign n1466 = n356 & n445 ;
  assign n1467 = n1465 & n1466 ;
  assign n1468 = n361 ^ n153 ^ 1'b0 ;
  assign n1469 = ~n1467 & n1468 ;
  assign n1470 = n1469 ^ n502 ^ 1'b0 ;
  assign n1471 = ~n1464 & n1470 ;
  assign n1472 = n191 | n650 ;
  assign n1473 = n411 | n714 ;
  assign n1474 = n1094 | n1473 ;
  assign n1475 = ( ~n856 & n1472 ) | ( ~n856 & n1474 ) | ( n1472 & n1474 ) ;
  assign n1476 = n644 ^ n519 ^ n59 ;
  assign n1477 = n1475 & n1476 ;
  assign n1478 = ~n57 & n1477 ;
  assign n1479 = n1172 ^ n427 ^ 1'b0 ;
  assign n1480 = ~n553 & n1479 ;
  assign n1481 = ( n941 & n1378 ) | ( n941 & n1480 ) | ( n1378 & n1480 ) ;
  assign n1482 = ~n78 & n374 ;
  assign n1483 = ~n191 & n1482 ;
  assign n1484 = n1169 ^ n588 ^ n543 ;
  assign n1485 = n519 & ~n903 ;
  assign n1486 = n200 | n434 ;
  assign n1487 = n548 & ~n1486 ;
  assign n1488 = ~n1116 & n1487 ;
  assign n1489 = n1052 ^ n551 ^ 1'b0 ;
  assign n1490 = n816 ^ n305 ^ 1'b0 ;
  assign n1492 = n228 & n593 ;
  assign n1491 = ( n43 & ~n242 ) | ( n43 & n865 ) | ( ~n242 & n865 ) ;
  assign n1493 = n1492 ^ n1491 ^ n1178 ;
  assign n1494 = n554 ^ n211 ^ 1'b0 ;
  assign n1495 = n40 & ~n1494 ;
  assign n1496 = ( ~n1050 & n1493 ) | ( ~n1050 & n1495 ) | ( n1493 & n1495 ) ;
  assign n1501 = n916 ^ n213 ^ 1'b0 ;
  assign n1502 = n427 | n1501 ;
  assign n1498 = n435 | n508 ;
  assign n1499 = n37 | n1498 ;
  assign n1497 = n16 & n1085 ;
  assign n1500 = n1499 ^ n1497 ^ 1'b0 ;
  assign n1503 = n1502 ^ n1500 ^ n911 ;
  assign n1504 = n234 & ~n954 ;
  assign n1505 = n1504 ^ n310 ^ 1'b0 ;
  assign n1506 = n1000 ^ n237 ^ 1'b0 ;
  assign n1507 = n647 | n1035 ;
  assign n1508 = n1018 ^ n177 ^ 1'b0 ;
  assign n1509 = n231 | n1508 ;
  assign n1510 = n1507 & ~n1509 ;
  assign n1511 = n1510 ^ n186 ^ 1'b0 ;
  assign n1512 = ( n305 & n830 ) | ( n305 & n1080 ) | ( n830 & n1080 ) ;
  assign n1513 = n20 | n44 ;
  assign n1514 = n1171 ^ n1037 ^ 1'b0 ;
  assign n1515 = n1513 | n1514 ;
  assign n1516 = n383 ^ n121 ^ 1'b0 ;
  assign n1517 = n494 & n717 ;
  assign n1518 = ~n1516 & n1517 ;
  assign n1519 = n1035 ^ n801 ^ 1'b0 ;
  assign n1520 = n99 & n1519 ;
  assign n1521 = n583 ^ n59 ^ 1'b0 ;
  assign n1522 = n98 | n1521 ;
  assign n1523 = ( n73 & n766 ) | ( n73 & ~n1522 ) | ( n766 & ~n1522 ) ;
  assign n1524 = n130 & ~n398 ;
  assign n1525 = n67 & n1524 ;
  assign n1527 = ( n201 & n756 ) | ( n201 & n938 ) | ( n756 & n938 ) ;
  assign n1528 = n1527 ^ n1218 ^ 1'b0 ;
  assign n1529 = n1160 & ~n1528 ;
  assign n1526 = n109 & n1278 ;
  assign n1530 = n1529 ^ n1526 ^ 1'b0 ;
  assign n1531 = n772 & n1530 ;
  assign n1532 = n1525 | n1531 ;
  assign n1533 = ~n177 & n1465 ;
  assign n1534 = n533 & ~n818 ;
  assign n1535 = n320 & n1534 ;
  assign n1536 = n79 & ~n1535 ;
  assign n1537 = n1536 ^ n1156 ^ 1'b0 ;
  assign n1538 = ~n108 & n1226 ;
  assign n1539 = n53 & ~n1234 ;
  assign n1540 = n572 ^ x10 ^ 1'b0 ;
  assign n1542 = n23 | n1245 ;
  assign n1541 = n180 & n1334 ;
  assign n1543 = n1542 ^ n1541 ^ 1'b0 ;
  assign n1544 = ~n59 & n688 ;
  assign n1545 = n251 & n1544 ;
  assign n1546 = n169 & n558 ;
  assign n1547 = n639 ^ n576 ^ n62 ;
  assign n1548 = n260 & n881 ;
  assign n1549 = ( ~n294 & n1547 ) | ( ~n294 & n1548 ) | ( n1547 & n1548 ) ;
  assign n1550 = n498 ^ n41 ^ 1'b0 ;
  assign n1551 = n153 & n1055 ;
  assign n1552 = n1551 ^ n177 ^ 1'b0 ;
  assign n1553 = ~n55 & n814 ;
  assign n1554 = ~n919 & n1178 ;
  assign n1555 = n334 & n863 ;
  assign n1556 = ~n1554 & n1555 ;
  assign n1557 = n44 & ~n1427 ;
  assign n1558 = n1557 ^ n804 ^ 1'b0 ;
  assign n1559 = n763 ^ n40 ^ 1'b0 ;
  assign n1560 = n586 & ~n1559 ;
  assign n1561 = ~n1558 & n1560 ;
  assign n1562 = n722 & ~n1561 ;
  assign n1563 = ~n1237 & n1562 ;
  assign n1564 = n151 ^ x10 ^ 1'b0 ;
  assign n1565 = ~n1135 & n1564 ;
  assign n1566 = n466 & ~n1516 ;
  assign n1567 = n1566 ^ n1476 ^ 1'b0 ;
  assign n1568 = n427 | n1567 ;
  assign n1569 = n77 & n886 ;
  assign n1570 = n350 & n991 ;
  assign n1571 = n684 & n1570 ;
  assign n1572 = ( n1041 & ~n1569 ) | ( n1041 & n1571 ) | ( ~n1569 & n1571 ) ;
  assign n1573 = n1572 ^ n1515 ^ 1'b0 ;
  assign n1574 = ~n245 & n612 ;
  assign n1575 = ~n150 & n577 ;
  assign n1576 = n1196 | n1335 ;
  assign n1577 = n1575 | n1576 ;
  assign n1578 = n209 & n728 ;
  assign n1579 = x1 & ~n190 ;
  assign n1580 = n281 & n1579 ;
  assign n1581 = n548 & n1580 ;
  assign n1582 = n840 ^ n554 ^ 1'b0 ;
  assign n1583 = ~x1 & n1582 ;
  assign n1584 = n37 & n1302 ;
  assign n1585 = ~n885 & n1584 ;
  assign n1586 = n381 ^ x10 ^ 1'b0 ;
  assign n1587 = ~n318 & n1087 ;
  assign n1588 = ~n439 & n644 ;
  assign n1589 = ~n1587 & n1588 ;
  assign n1591 = n711 ^ n38 ^ 1'b0 ;
  assign n1590 = ( n30 & ~n576 ) | ( n30 & n1063 ) | ( ~n576 & n1063 ) ;
  assign n1592 = n1591 ^ n1590 ^ 1'b0 ;
  assign n1593 = n774 & ~n1509 ;
  assign n1594 = ~n1241 & n1593 ;
  assign n1595 = n427 | n747 ;
  assign n1596 = n1595 ^ n1105 ^ 1'b0 ;
  assign n1597 = n1192 ^ n230 ^ x3 ;
  assign n1598 = n525 & n645 ;
  assign n1599 = n1598 ^ n1024 ^ 1'b0 ;
  assign n1600 = ~n1456 & n1599 ;
  assign n1601 = ~n723 & n1600 ;
  assign n1602 = ~n1597 & n1601 ;
  assign n1603 = n874 ^ n356 ^ 1'b0 ;
  assign n1604 = ~n423 & n1603 ;
  assign n1605 = ( ~n1341 & n1599 ) | ( ~n1341 & n1604 ) | ( n1599 & n1604 ) ;
  assign n1606 = n1605 ^ n982 ^ 1'b0 ;
  assign n1607 = n905 ^ n101 ^ 1'b0 ;
  assign n1608 = ~n426 & n1607 ;
  assign n1609 = ~n647 & n1608 ;
  assign n1610 = n923 | n1189 ;
  assign n1611 = n269 & n526 ;
  assign n1612 = n1611 ^ n428 ^ 1'b0 ;
  assign n1613 = n1610 & ~n1612 ;
  assign n1614 = n107 & n192 ;
  assign n1615 = n205 ^ n150 ^ 1'b0 ;
  assign n1616 = x0 & ~n1615 ;
  assign n1617 = n350 & n1175 ;
  assign n1618 = n1616 & ~n1617 ;
  assign n1619 = n637 & n1618 ;
  assign n1620 = n1066 ^ n550 ^ 1'b0 ;
  assign n1621 = n974 & ~n1620 ;
  assign n1622 = ( n100 & n1619 ) | ( n100 & n1621 ) | ( n1619 & n1621 ) ;
  assign n1623 = ( ~n166 & n1614 ) | ( ~n166 & n1622 ) | ( n1614 & n1622 ) ;
  assign n1624 = x0 & n725 ;
  assign n1625 = n1624 ^ n53 ^ 1'b0 ;
  assign n1626 = ~n1045 & n1614 ;
  assign n1627 = n1626 ^ n361 ^ 1'b0 ;
  assign n1628 = n1506 | n1627 ;
  assign n1629 = n360 & ~n441 ;
  assign n1630 = n1629 ^ n1573 ^ 1'b0 ;
  assign n1632 = n607 ^ n91 ^ 1'b0 ;
  assign n1633 = n1260 & ~n1632 ;
  assign n1631 = n716 & n1457 ;
  assign n1634 = n1633 ^ n1631 ^ 1'b0 ;
  assign n1635 = ~n265 & n1147 ;
  assign n1636 = ~n519 & n1058 ;
  assign n1637 = n498 ^ n37 ^ 1'b0 ;
  assign n1638 = n1636 | n1637 ;
  assign n1639 = n471 & n1241 ;
  assign n1640 = ( n346 & n684 ) | ( n346 & ~n1639 ) | ( n684 & ~n1639 ) ;
  assign n1641 = n1640 ^ n1048 ^ 1'b0 ;
  assign n1642 = ( n890 & ~n942 ) | ( n890 & n1180 ) | ( ~n942 & n1180 ) ;
  assign n1643 = n498 | n953 ;
  assign n1644 = n842 ^ n108 ^ 1'b0 ;
  assign n1645 = n436 & n1644 ;
  assign n1649 = n458 & ~n1095 ;
  assign n1646 = n547 ^ n115 ^ 1'b0 ;
  assign n1647 = n218 | n1646 ;
  assign n1648 = n74 | n1647 ;
  assign n1650 = n1649 ^ n1648 ^ 1'b0 ;
  assign n1651 = n1062 & n1418 ;
  assign n1652 = n1651 ^ n533 ^ 1'b0 ;
  assign n1653 = n1531 ^ n315 ^ 1'b0 ;
  assign n1654 = n1387 ^ n1142 ^ 1'b0 ;
  assign n1655 = ~n707 & n953 ;
  assign n1656 = n1655 ^ n720 ^ 1'b0 ;
  assign n1657 = n1407 ^ n1048 ^ 1'b0 ;
  assign n1658 = n1656 | n1657 ;
  assign n1659 = n994 & n1210 ;
  assign n1660 = ~n860 & n1659 ;
  assign n1662 = ( ~n955 & n972 ) | ( ~n955 & n1095 ) | ( n972 & n1095 ) ;
  assign n1661 = n1395 ^ n256 ^ 1'b0 ;
  assign n1663 = n1662 ^ n1661 ^ 1'b0 ;
  assign n1664 = n550 & ~n1663 ;
  assign n1665 = n1664 ^ n1149 ^ n77 ;
  assign n1666 = n722 ^ n324 ^ 1'b0 ;
  assign n1667 = n980 | n1666 ;
  assign n1668 = n1667 ^ n73 ^ 1'b0 ;
  assign n1669 = n800 & n1159 ;
  assign n1670 = ~n16 & n1669 ;
  assign n1671 = n151 | n321 ;
  assign n1672 = n192 | n1671 ;
  assign n1673 = n791 & n823 ;
  assign n1674 = n1673 ^ n682 ^ 1'b0 ;
  assign n1675 = n1672 & n1674 ;
  assign n1676 = ~n735 & n1675 ;
  assign n1677 = n1138 ^ n431 ^ 1'b0 ;
  assign n1678 = n1566 ^ n205 ^ 1'b0 ;
  assign n1679 = x11 & n1678 ;
  assign n1681 = n885 ^ n299 ^ 1'b0 ;
  assign n1682 = n569 | n1021 ;
  assign n1683 = n1682 ^ n135 ^ 1'b0 ;
  assign n1684 = ~n1681 & n1683 ;
  assign n1680 = ~x11 & n486 ;
  assign n1685 = n1684 ^ n1680 ^ 1'b0 ;
  assign n1686 = n1679 & ~n1685 ;
  assign n1687 = n532 & n1686 ;
  assign n1688 = n1687 ^ n541 ^ 1'b0 ;
  assign n1689 = n1677 | n1688 ;
  assign n1690 = n1676 | n1689 ;
  assign n1691 = n1167 | n1619 ;
  assign n1692 = n102 | n455 ;
  assign n1693 = n230 & ~n1692 ;
  assign n1694 = n738 & n1693 ;
  assign n1695 = n225 ^ n93 ^ 1'b0 ;
  assign n1696 = n42 | n1695 ;
  assign n1697 = n1696 ^ n334 ^ 1'b0 ;
  assign n1698 = n420 & ~n1697 ;
  assign n1699 = n973 & ~n1698 ;
  assign n1708 = n747 & n791 ;
  assign n1709 = n1708 ^ n174 ^ 1'b0 ;
  assign n1700 = ~n111 & n153 ;
  assign n1701 = n521 ^ n364 ^ n228 ;
  assign n1702 = n698 | n1701 ;
  assign n1703 = n922 & n1702 ;
  assign n1704 = n1703 ^ n752 ^ 1'b0 ;
  assign n1705 = n1138 ^ n554 ^ 1'b0 ;
  assign n1706 = n1704 & ~n1705 ;
  assign n1707 = ~n1700 & n1706 ;
  assign n1710 = n1709 ^ n1707 ^ 1'b0 ;
  assign n1711 = n539 | n951 ;
  assign n1712 = n1711 ^ n1680 ^ 1'b0 ;
  assign n1713 = n408 ^ n121 ^ 1'b0 ;
  assign n1714 = ~n238 & n1061 ;
  assign n1715 = ~n1713 & n1714 ;
  assign n1716 = n432 & n1715 ;
  assign n1717 = ( ~n136 & n570 ) | ( ~n136 & n1200 ) | ( n570 & n1200 ) ;
  assign n1718 = n63 & n705 ;
  assign n1719 = n1717 & ~n1718 ;
  assign n1720 = ~n1094 & n1719 ;
  assign n1721 = n494 & ~n1720 ;
  assign n1722 = n750 ^ n201 ^ 1'b0 ;
  assign n1723 = ( x1 & ~n195 ) | ( x1 & n816 ) | ( ~n195 & n816 ) ;
  assign n1724 = n1723 ^ n43 ^ 1'b0 ;
  assign n1725 = n1335 ^ n925 ^ 1'b0 ;
  assign n1726 = n846 & ~n1725 ;
  assign n1727 = ~n691 & n860 ;
  assign n1728 = n1200 ^ n214 ^ 1'b0 ;
  assign n1729 = ~n381 & n1728 ;
  assign n1730 = n792 & n1729 ;
  assign n1731 = n1730 ^ n905 ^ 1'b0 ;
  assign n1732 = n1640 ^ n1258 ^ 1'b0 ;
  assign n1733 = n147 | n1732 ;
  assign n1734 = n990 & ~n1733 ;
  assign n1735 = n745 ^ n250 ^ 1'b0 ;
  assign n1736 = ~n1426 & n1735 ;
  assign n1737 = n174 & ~n1112 ;
  assign n1743 = n67 | n865 ;
  assign n1744 = n1743 ^ n428 ^ 1'b0 ;
  assign n1739 = n254 ^ n179 ^ 1'b0 ;
  assign n1740 = n396 | n1739 ;
  assign n1738 = ~n132 & n283 ;
  assign n1741 = n1740 ^ n1738 ^ 1'b0 ;
  assign n1742 = n1741 ^ n563 ^ 1'b0 ;
  assign n1745 = n1744 ^ n1742 ^ n1155 ;
  assign n1746 = ( n158 & n830 ) | ( n158 & ~n1439 ) | ( n830 & ~n1439 ) ;
  assign n1747 = ~n639 & n782 ;
  assign n1748 = n125 & n1747 ;
  assign n1749 = n322 ^ n44 ^ 1'b0 ;
  assign n1750 = n923 | n1749 ;
  assign n1751 = n1748 & ~n1750 ;
  assign n1752 = n918 ^ n334 ^ 1'b0 ;
  assign n1753 = n561 | n1752 ;
  assign n1754 = n1753 ^ n316 ^ 1'b0 ;
  assign n1755 = n716 & ~n916 ;
  assign n1756 = n1754 & n1755 ;
  assign n1757 = n1243 | n1756 ;
  assign n1758 = n353 | n1757 ;
  assign n1759 = n1566 ^ n126 ^ 1'b0 ;
  assign n1760 = n431 & ~n1759 ;
  assign n1761 = n1287 ^ n990 ^ 1'b0 ;
  assign n1762 = n129 & ~n440 ;
  assign n1763 = n1741 ^ n1153 ^ 1'b0 ;
  assign n1764 = n1762 & n1763 ;
  assign n1765 = n324 & n1764 ;
  assign n1766 = ~n309 & n1765 ;
  assign n1767 = n132 ^ n102 ^ n36 ;
  assign n1768 = n1767 ^ n886 ^ 1'b0 ;
  assign n1769 = n1189 ^ n607 ^ 1'b0 ;
  assign n1770 = n223 & ~n1769 ;
  assign n1771 = ~n250 & n1770 ;
  assign n1773 = n527 & ~n532 ;
  assign n1774 = n174 & ~n457 ;
  assign n1775 = n1351 & n1774 ;
  assign n1776 = n210 | n1775 ;
  assign n1777 = n1776 ^ n1247 ^ 1'b0 ;
  assign n1778 = n514 | n1777 ;
  assign n1779 = n1778 ^ n48 ^ 1'b0 ;
  assign n1780 = n1779 ^ n464 ^ 1'b0 ;
  assign n1781 = n1773 & ~n1780 ;
  assign n1782 = n1334 & n1781 ;
  assign n1783 = ~n1472 & n1782 ;
  assign n1784 = n1783 ^ n766 ^ n79 ;
  assign n1772 = n332 & n1698 ;
  assign n1785 = n1784 ^ n1772 ^ 1'b0 ;
  assign n1786 = n23 | n1785 ;
  assign n1787 = n887 ^ n313 ^ 1'b0 ;
  assign n1788 = n32 & n55 ;
  assign n1789 = ~n85 & n1788 ;
  assign n1790 = n1789 ^ n224 ^ 1'b0 ;
  assign n1791 = n99 & ~n1790 ;
  assign n1792 = n842 & n1791 ;
  assign n1793 = n955 & n1792 ;
  assign n1794 = ~n243 & n1072 ;
  assign n1795 = n695 & n1794 ;
  assign n1796 = n1795 ^ n448 ^ 1'b0 ;
  assign n1797 = ~n93 & n564 ;
  assign n1798 = n1797 ^ n475 ^ 1'b0 ;
  assign n1799 = n1196 ^ n895 ^ 1'b0 ;
  assign n1800 = ~n1798 & n1799 ;
  assign n1801 = ( ~n150 & n1495 ) | ( ~n150 & n1800 ) | ( n1495 & n1800 ) ;
  assign n1802 = n1796 & n1801 ;
  assign n1803 = n1802 ^ n63 ^ 1'b0 ;
  assign n1804 = n154 & ~n1596 ;
  assign n1805 = ~n160 & n1804 ;
  assign n1806 = n1594 | n1805 ;
  assign n1807 = n1153 | n1806 ;
  assign n1808 = n426 & ~n435 ;
  assign n1809 = n1509 ^ n589 ^ n136 ;
  assign n1810 = n405 | n694 ;
  assign n1811 = n916 & ~n1682 ;
  assign n1812 = n633 ^ n237 ^ 1'b0 ;
  assign n1813 = n462 ^ n63 ^ 1'b0 ;
  assign n1814 = n1813 ^ n1103 ^ 1'b0 ;
  assign n1815 = n779 & ~n1814 ;
  assign n1816 = n354 | n1815 ;
  assign n1817 = n947 ^ n408 ^ 1'b0 ;
  assign n1818 = ~n1816 & n1817 ;
  assign n1819 = ~n637 & n838 ;
  assign n1820 = ~n22 & n1819 ;
  assign n1821 = n846 & ~n1820 ;
  assign n1822 = n1821 ^ n1362 ^ 1'b0 ;
  assign n1823 = ~n51 & n238 ;
  assign n1824 = n503 ^ n44 ^ n22 ;
  assign n1825 = n1188 ^ n115 ^ 1'b0 ;
  assign n1826 = n556 & ~n672 ;
  assign n1827 = n916 ^ n816 ^ 1'b0 ;
  assign n1828 = n263 | n1827 ;
  assign n1829 = n510 & n962 ;
  assign n1830 = ~n1418 & n1829 ;
  assign n1834 = n46 & n583 ;
  assign n1835 = n1834 ^ n336 ^ 1'b0 ;
  assign n1836 = ~n48 & n1835 ;
  assign n1831 = n918 ^ n756 ^ 1'b0 ;
  assign n1832 = n475 & ~n1831 ;
  assign n1833 = ~n1397 & n1832 ;
  assign n1837 = n1836 ^ n1833 ^ 1'b0 ;
  assign n1838 = n1073 & n1837 ;
  assign n1839 = n760 & ~n811 ;
  assign n1840 = n1839 ^ n1197 ^ 1'b0 ;
  assign n1841 = ~n1370 & n1374 ;
  assign n1842 = n649 ^ n176 ^ 1'b0 ;
  assign n1843 = n1842 ^ n977 ^ 1'b0 ;
  assign n1845 = n210 & n811 ;
  assign n1844 = x11 & ~n641 ;
  assign n1846 = n1845 ^ n1844 ^ 1'b0 ;
  assign n1847 = n947 ^ n922 ^ 1'b0 ;
  assign n1848 = x6 & n1847 ;
  assign n1849 = n1848 ^ n1046 ^ n438 ;
  assign n1850 = n955 | n1849 ;
  assign n1851 = n332 & ~n1850 ;
  assign n1852 = n1094 & n1527 ;
  assign n1859 = n1444 ^ n1035 ^ n261 ;
  assign n1856 = n431 ^ n319 ^ 1'b0 ;
  assign n1857 = ~n951 & n1856 ;
  assign n1853 = n483 & ~n903 ;
  assign n1854 = n1853 ^ n47 ^ 1'b0 ;
  assign n1855 = n1744 & n1854 ;
  assign n1858 = n1857 ^ n1855 ^ 1'b0 ;
  assign n1860 = n1859 ^ n1858 ^ 1'b0 ;
  assign n1861 = n524 & ~n1860 ;
  assign n1862 = n1666 ^ n263 ^ 1'b0 ;
  assign n1863 = n1861 & n1862 ;
  assign n1864 = ~n1169 & n1863 ;
  assign n1865 = n790 ^ n216 ^ 1'b0 ;
  assign n1866 = ( n376 & n1731 ) | ( n376 & n1865 ) | ( n1731 & n1865 ) ;
  assign n1867 = n619 ^ n361 ^ 1'b0 ;
  assign n1868 = n1221 | n1867 ;
  assign n1873 = n91 ^ n20 ^ 1'b0 ;
  assign n1874 = n1633 & n1873 ;
  assign n1875 = n228 | n230 ;
  assign n1876 = ( n1316 & ~n1563 ) | ( n1316 & n1875 ) | ( ~n1563 & n1875 ) ;
  assign n1877 = ( n97 & n1874 ) | ( n97 & n1876 ) | ( n1874 & n1876 ) ;
  assign n1869 = ~n352 & n1334 ;
  assign n1870 = n806 & ~n1869 ;
  assign n1871 = n1870 ^ n397 ^ 1'b0 ;
  assign n1872 = n78 | n1871 ;
  assign n1878 = n1877 ^ n1872 ^ 1'b0 ;
  assign n1879 = n580 & n1607 ;
  assign n1880 = n1879 ^ n1491 ^ 1'b0 ;
  assign n1881 = n1609 | n1880 ;
  assign n1882 = n153 & ~n361 ;
  assign n1883 = n963 | n1636 ;
  assign n1884 = n853 & ~n1871 ;
  assign n1885 = ~n134 & n1884 ;
  assign n1886 = n506 & ~n1885 ;
  assign n1887 = n1817 ^ n766 ^ 1'b0 ;
  assign n1888 = n1886 & n1887 ;
  assign n1889 = n30 ^ n13 ^ 1'b0 ;
  assign n1890 = n1889 ^ n1157 ^ 1'b0 ;
  assign n1891 = n263 | n326 ;
  assign n1892 = n169 & n177 ;
  assign n1893 = ~x10 & n1892 ;
  assign n1894 = n1573 & n1726 ;
  assign n1895 = n941 & ~n1167 ;
  assign n1896 = n1078 | n1895 ;
  assign n1897 = n1896 ^ n285 ^ 1'b0 ;
  assign n1898 = ( n576 & n830 ) | ( n576 & n1897 ) | ( n830 & n1897 ) ;
  assign n1899 = n361 | n1898 ;
  assign n1900 = n1272 | n1899 ;
  assign n1901 = ~n176 & n1575 ;
  assign n1902 = n1901 ^ n51 ^ 1'b0 ;
  assign n1903 = n1902 ^ n306 ^ 1'b0 ;
  assign n1904 = n1903 ^ n1770 ^ n1489 ;
  assign n1905 = n1871 ^ n619 ^ 1'b0 ;
  assign n1910 = ~n98 & n226 ;
  assign n1911 = n77 & n350 ;
  assign n1912 = n1910 & n1911 ;
  assign n1907 = ~n592 & n983 ;
  assign n1908 = n563 ^ n362 ^ 1'b0 ;
  assign n1909 = n1907 & ~n1908 ;
  assign n1906 = n252 ^ n57 ^ 1'b0 ;
  assign n1913 = n1912 ^ n1909 ^ n1906 ;
  assign n1918 = n624 ^ n44 ^ 1'b0 ;
  assign n1914 = n364 | n1121 ;
  assign n1915 = n1914 ^ n272 ^ 1'b0 ;
  assign n1916 = n1138 | n1915 ;
  assign n1917 = n1207 & ~n1916 ;
  assign n1919 = n1918 ^ n1917 ^ 1'b0 ;
  assign n1920 = ~n478 & n1919 ;
  assign n1921 = ~n22 & n1920 ;
  assign n1926 = n1495 ^ n933 ^ 1'b0 ;
  assign n1922 = n1777 ^ n619 ^ 1'b0 ;
  assign n1923 = n417 & ~n1922 ;
  assign n1924 = n1403 & n1923 ;
  assign n1925 = n654 | n1924 ;
  assign n1927 = n1926 ^ n1925 ^ 1'b0 ;
  assign n1928 = ~x3 & n1062 ;
  assign n1929 = ( n527 & n794 ) | ( n527 & ~n1061 ) | ( n794 & ~n1061 ) ;
  assign n1930 = n1929 ^ n1280 ^ 1'b0 ;
  assign n1931 = n1930 ^ n1419 ^ 1'b0 ;
  assign n1932 = n1871 ^ n604 ^ 1'b0 ;
  assign n1933 = n1886 & ~n1932 ;
  assign n1934 = n415 & ~n1029 ;
  assign n1935 = n68 & n164 ;
  assign n1936 = n184 & n1935 ;
  assign n1937 = n1936 ^ n109 ^ 1'b0 ;
  assign n1938 = n1859 ^ n767 ^ n612 ;
  assign n1939 = n1938 ^ n1190 ^ 1'b0 ;
  assign n1940 = n1937 | n1939 ;
  assign n1941 = ~n961 & n1400 ;
  assign n1942 = n1941 ^ n1909 ^ 1'b0 ;
  assign n1943 = n1942 ^ n508 ^ 1'b0 ;
  assign n1944 = n334 & ~n541 ;
  assign n1945 = n1876 & n1944 ;
  assign n1946 = n251 ^ n136 ^ 1'b0 ;
  assign n1947 = n558 | n1946 ;
  assign n1948 = n1947 ^ x3 ^ 1'b0 ;
  assign n1949 = n1041 | n1367 ;
  assign n1950 = n908 & ~n1949 ;
  assign n1951 = n918 & n1950 ;
  assign n1952 = n1629 & n1951 ;
  assign n1955 = n178 & n1262 ;
  assign n1956 = ~n283 & n1955 ;
  assign n1953 = n63 & n1273 ;
  assign n1954 = n756 | n1953 ;
  assign n1957 = n1956 ^ n1954 ^ 1'b0 ;
  assign n1958 = ( ~n102 & n210 ) | ( ~n102 & n1682 ) | ( n210 & n1682 ) ;
  assign n1959 = ~n79 & n203 ;
  assign n1960 = n1959 ^ n1818 ^ 1'b0 ;
  assign n1961 = n739 ^ n542 ^ 1'b0 ;
  assign n1962 = n590 & ~n1961 ;
  assign n1963 = n1339 ^ n309 ^ 1'b0 ;
  assign n1964 = n1922 | n1963 ;
  assign n1965 = n231 | n1538 ;
  assign n1966 = n1964 | n1965 ;
  assign n1967 = n1846 | n1966 ;
  assign n1968 = n437 | n494 ;
  assign n1969 = n1968 ^ n1699 ^ 1'b0 ;
  assign n1970 = ~n1784 & n1969 ;
  assign n1971 = n1956 | n1970 ;
  assign n1972 = n1971 ^ n218 ^ 1'b0 ;
  assign n1973 = n26 & ~n61 ;
  assign n1974 = n969 & n1973 ;
  assign n1975 = n875 & n1131 ;
  assign n1976 = n1974 & n1975 ;
  assign n1977 = n877 | n1748 ;
  assign n1978 = ~n1871 & n1977 ;
  assign n1979 = n354 & n1978 ;
  assign n1980 = n401 & ~n641 ;
  assign n1981 = n1980 ^ n1699 ^ 1'b0 ;
  assign n1982 = n1979 | n1981 ;
  assign n1983 = ( n484 & n1096 ) | ( n484 & n1164 ) | ( n1096 & n1164 ) ;
  assign n1984 = n914 & ~n1983 ;
  assign n1985 = n169 & ~n1958 ;
  assign n1986 = ~n263 & n1985 ;
  assign n1987 = n1357 ^ n989 ^ 1'b0 ;
  assign n1988 = n1318 | n1987 ;
  assign n1993 = n1813 ^ n738 ^ x6 ;
  assign n1989 = n612 ^ n126 ^ 1'b0 ;
  assign n1990 = n46 & n1989 ;
  assign n1991 = n922 & n1990 ;
  assign n1992 = n767 & ~n1991 ;
  assign n1994 = n1993 ^ n1992 ^ 1'b0 ;
  assign n1995 = ~n332 & n1994 ;
  assign n1996 = ( n40 & n187 ) | ( n40 & n760 ) | ( n187 & n760 ) ;
  assign n1997 = n1996 ^ n1915 ^ 1'b0 ;
  assign n1998 = n704 | n1996 ;
  assign n1999 = n1998 ^ n1670 ^ 1'b0 ;
  assign n2000 = n1511 ^ n108 ^ 1'b0 ;
  assign n2001 = n594 & ~n2000 ;
  assign n2002 = ( ~n360 & n1942 ) | ( ~n360 & n2001 ) | ( n1942 & n2001 ) ;
  assign n2003 = ~n217 & n1419 ;
  assign n2004 = ~n341 & n2003 ;
  assign n2005 = n130 & ~n321 ;
  assign n2006 = n2004 & ~n2005 ;
  assign n2007 = ~n886 & n1169 ;
  assign n2008 = n686 & n2007 ;
  assign n2009 = n340 & ~n1990 ;
  assign n2010 = n2009 ^ n592 ^ 1'b0 ;
  assign n2011 = n2008 | n2010 ;
  assign n2013 = n1134 ^ n773 ^ 1'b0 ;
  assign n2014 = n892 & n2013 ;
  assign n2012 = n893 | n1340 ;
  assign n2015 = n2014 ^ n2012 ^ 1'b0 ;
  assign n2016 = n811 | n1653 ;
  assign n2017 = n1720 & ~n2016 ;
  assign n2018 = n249 | n355 ;
  assign n2019 = n608 & ~n2018 ;
  assign n2020 = n567 & ~n2019 ;
  assign n2021 = n948 ^ n583 ^ 1'b0 ;
  assign n2022 = n2020 & ~n2021 ;
  assign n2023 = n356 ^ n203 ^ 1'b0 ;
  assign n2024 = n1977 & ~n2023 ;
  assign n2025 = n332 & n2024 ;
  assign n2026 = n269 ^ n55 ^ 1'b0 ;
  assign n2027 = n2025 | n2026 ;
  assign n2028 = n1153 ^ n951 ^ n59 ;
  assign n2029 = n2008 ^ n1647 ^ n67 ;
  assign n2030 = n1772 ^ n1425 ^ n321 ;
  assign n2031 = n322 | n345 ;
  assign n2032 = n2031 ^ n792 ^ 1'b0 ;
  assign n2033 = ~n63 & n2032 ;
  assign n2034 = n2033 ^ n172 ^ 1'b0 ;
  assign n2035 = n166 & ~n2034 ;
  assign n2036 = n1041 & n2035 ;
  assign n2037 = n2036 ^ n505 ^ 1'b0 ;
  assign n2038 = n563 & n708 ;
  assign n2039 = n378 & n2038 ;
  assign n2040 = n63 | n1441 ;
  assign n2041 = n101 & ~n2040 ;
  assign n2043 = n59 | n908 ;
  assign n2044 = n763 & ~n2043 ;
  assign n2045 = n1246 ^ n154 ^ n108 ;
  assign n2046 = ~n2044 & n2045 ;
  assign n2047 = n376 & n2046 ;
  assign n2042 = n1672 & n1791 ;
  assign n2048 = n2047 ^ n2042 ^ 1'b0 ;
  assign n2049 = ( n304 & n2041 ) | ( n304 & ~n2048 ) | ( n2041 & ~n2048 ) ;
  assign n2050 = n1526 ^ n1180 ^ 1'b0 ;
  assign n2051 = n740 ^ n458 ^ 1'b0 ;
  assign n2052 = n2051 ^ n774 ^ 1'b0 ;
  assign n2053 = n2050 & n2052 ;
  assign n2054 = n603 ^ n48 ^ 1'b0 ;
  assign n2055 = n1636 ^ n694 ^ 1'b0 ;
  assign n2056 = ~n2054 & n2055 ;
  assign n2057 = n2056 ^ n57 ^ 1'b0 ;
  assign n2058 = n1980 | n2057 ;
  assign n2059 = n2058 ^ n757 ^ 1'b0 ;
  assign n2060 = n1450 & n1991 ;
  assign n2061 = n30 | n2060 ;
  assign n2062 = n2061 ^ n35 ^ 1'b0 ;
  assign n2063 = x10 & ~n1427 ;
  assign n2064 = ~n1109 & n2063 ;
  assign n2065 = n2064 ^ n1910 ^ n1460 ;
  assign n2066 = n2065 ^ n1277 ^ 1'b0 ;
  assign n2067 = n40 | n2066 ;
  assign n2068 = n596 | n629 ;
  assign n2069 = n230 & n1320 ;
  assign n2070 = n2069 ^ n1279 ^ 1'b0 ;
  assign n2071 = n2070 ^ n1262 ^ 1'b0 ;
  assign n2072 = ~n210 & n859 ;
  assign n2073 = n289 ^ n118 ^ 1'b0 ;
  assign n2074 = n2073 ^ n313 ^ 1'b0 ;
  assign n2075 = n183 ^ n162 ^ 1'b0 ;
  assign n2076 = n2074 & n2075 ;
  assign n2089 = n861 ^ n315 ^ 1'b0 ;
  assign n2084 = n346 & n400 ;
  assign n2085 = n863 & ~n2084 ;
  assign n2086 = n2085 ^ n905 ^ 1'b0 ;
  assign n2087 = n827 & ~n1779 ;
  assign n2088 = ~n2086 & n2087 ;
  assign n2090 = n2089 ^ n2088 ^ 1'b0 ;
  assign n2077 = n36 & ~n685 ;
  assign n2078 = n53 & ~n2077 ;
  assign n2079 = x7 & ~n1709 ;
  assign n2080 = n2079 ^ n501 ^ 1'b0 ;
  assign n2081 = n214 & ~n2080 ;
  assign n2082 = n2081 ^ n1591 ^ 1'b0 ;
  assign n2083 = ( n450 & ~n2078 ) | ( n450 & n2082 ) | ( ~n2078 & n2082 ) ;
  assign n2091 = n2090 ^ n2083 ^ 1'b0 ;
  assign n2092 = n842 & n2091 ;
  assign n2093 = n1329 ^ n548 ^ 1'b0 ;
  assign n2094 = n152 & ~n2093 ;
  assign n2095 = n837 & n2094 ;
  assign n2096 = n1761 ^ n1401 ^ 1'b0 ;
  assign n2097 = ~n2095 & n2096 ;
  assign n2098 = n37 & n1326 ;
  assign n2099 = ~n57 & n2098 ;
  assign n2100 = ~n2059 & n2099 ;
  assign n2101 = n246 & n730 ;
  assign n2102 = ~n1940 & n2101 ;
  assign n2108 = n197 & ~n747 ;
  assign n2109 = n2108 ^ n1619 ^ 1'b0 ;
  assign n2110 = n381 & n2109 ;
  assign n2106 = ~n461 & n691 ;
  assign n2107 = n2106 ^ n893 ^ 1'b0 ;
  assign n2103 = n655 & n887 ;
  assign n2104 = n726 & n2103 ;
  assign n2105 = n1010 & ~n2104 ;
  assign n2111 = n2110 ^ n2107 ^ n2105 ;
  assign n2112 = n774 ^ n717 ^ 1'b0 ;
  assign n2113 = n649 & n2112 ;
  assign n2114 = n641 ^ n607 ^ 1'b0 ;
  assign n2115 = n2114 ^ n472 ^ n458 ;
  assign n2118 = ~n569 & n838 ;
  assign n2116 = n216 | n1133 ;
  assign n2117 = n263 & ~n2116 ;
  assign n2119 = n2118 ^ n2117 ^ n1893 ;
  assign n2120 = n1091 ^ n752 ^ n742 ;
  assign n2121 = n1320 ^ n98 ^ 1'b0 ;
  assign n2122 = n2120 & ~n2121 ;
  assign n2123 = n809 ^ x8 ^ 1'b0 ;
  assign n2124 = n2123 ^ n1075 ^ n358 ;
  assign n2125 = n2124 ^ n545 ^ 1'b0 ;
  assign n2127 = n1112 ^ n884 ^ 1'b0 ;
  assign n2128 = ~n875 & n2127 ;
  assign n2126 = n684 & n800 ;
  assign n2129 = n2128 ^ n2126 ^ 1'b0 ;
  assign n2130 = n159 | n656 ;
  assign n2131 = n121 & n1168 ;
  assign n2132 = n2131 ^ n801 ^ 1'b0 ;
  assign n2133 = n1865 ^ n997 ^ 1'b0 ;
  assign n2134 = n411 | n2133 ;
  assign n2135 = n1170 | n1885 ;
  assign n2136 = ~n890 & n1125 ;
  assign n2137 = ~n2135 & n2136 ;
  assign n2138 = n1167 & n2137 ;
  assign n2139 = ( ~n517 & n1617 ) | ( ~n517 & n2138 ) | ( n1617 & n2138 ) ;
  assign n2140 = n13 & n1716 ;
  assign n2141 = n2140 ^ n854 ^ 1'b0 ;
  assign n2142 = n1506 | n2141 ;
  assign n2143 = n447 ^ n272 ^ 1'b0 ;
  assign n2144 = n1371 ^ n557 ^ 1'b0 ;
  assign n2145 = n2143 | n2144 ;
  assign n2146 = n510 | n1148 ;
  assign n2147 = n2146 ^ n1389 ^ n401 ;
  assign n2148 = ( n121 & n411 ) | ( n121 & ~n1177 ) | ( n411 & ~n1177 ) ;
  assign n2149 = ( n523 & ~n2019 ) | ( n523 & n2148 ) | ( ~n2019 & n2148 ) ;
  assign n2150 = n2149 ^ n1401 ^ 1'b0 ;
  assign n2151 = n318 & ~n1856 ;
  assign n2152 = n1542 & n2151 ;
  assign n2153 = n1488 & ~n2152 ;
  assign n2154 = n2153 ^ n1752 ^ 1'b0 ;
  assign n2155 = n57 & ~n923 ;
  assign n2156 = n2155 ^ n577 ^ 1'b0 ;
  assign n2157 = n2156 ^ n836 ^ 1'b0 ;
  assign n2158 = n2157 ^ n779 ^ n686 ;
  assign n2159 = n1676 ^ n1370 ^ 1'b0 ;
  assign n2160 = n1527 ^ n298 ^ 1'b0 ;
  assign n2161 = ( ~n401 & n2159 ) | ( ~n401 & n2160 ) | ( n2159 & n2160 ) ;
  assign n2167 = n608 | n1001 ;
  assign n2168 = n441 | n2167 ;
  assign n2162 = n1225 ^ n576 ^ 1'b0 ;
  assign n2163 = n2162 ^ n23 ^ 1'b0 ;
  assign n2164 = n1052 ^ n394 ^ n259 ;
  assign n2165 = n2163 & ~n2164 ;
  assign n2166 = n572 | n2165 ;
  assign n2169 = n2168 ^ n2166 ^ 1'b0 ;
  assign n2170 = n353 ^ n20 ^ 1'b0 ;
  assign n2171 = ~n383 & n2118 ;
  assign n2172 = n2170 & n2171 ;
  assign n2173 = n1591 | n2045 ;
  assign n2174 = n2173 ^ n899 ^ n126 ;
  assign n2175 = n179 | n523 ;
  assign n2176 = n2175 ^ x3 ^ 1'b0 ;
  assign n2177 = n1946 & n2176 ;
  assign n2178 = n1167 ^ n890 ^ 1'b0 ;
  assign n2179 = n93 & n1334 ;
  assign n2180 = ( ~n73 & n719 ) | ( ~n73 & n2179 ) | ( n719 & n2179 ) ;
  assign n2181 = n534 | n1930 ;
  assign n2182 = ( ~n82 & n249 ) | ( ~n82 & n684 ) | ( n249 & n684 ) ;
  assign n2183 = n1839 ^ n842 ^ 1'b0 ;
  assign n2184 = ~n2182 & n2183 ;
  assign n2185 = ~n1283 & n2184 ;
  assign n2186 = n692 & n2185 ;
  assign n2187 = n2186 ^ n1542 ^ 1'b0 ;
  assign n2188 = n1197 & ~n1225 ;
  assign n2189 = n1045 ^ n481 ^ 1'b0 ;
  assign n2190 = n1095 & n2189 ;
  assign n2191 = n1320 & n2190 ;
  assign n2192 = ~n1746 & n2191 ;
  assign n2193 = n127 & ~n2192 ;
  assign n2194 = n217 & n2193 ;
  assign n2195 = n435 | n517 ;
  assign n2196 = n1889 & n2195 ;
  assign n2197 = n125 ^ x10 ^ 1'b0 ;
  assign n2198 = ~n1166 & n2197 ;
  assign n2199 = n2196 & n2198 ;
  assign n2201 = n85 & n695 ;
  assign n2200 = ~n918 & n1178 ;
  assign n2202 = n2201 ^ n2200 ^ 1'b0 ;
  assign n2203 = n954 ^ n833 ^ n127 ;
  assign n2204 = n2086 & ~n2203 ;
  assign n2205 = n2204 ^ n1554 ^ 1'b0 ;
  assign n2206 = n650 ^ n85 ^ 1'b0 ;
  assign n2207 = n51 & ~n2143 ;
  assign n2208 = n2207 ^ n607 ^ n496 ;
  assign n2209 = n16 & ~n1758 ;
  assign n2210 = n1084 | n2209 ;
  assign n2211 = n1368 | n2210 ;
  assign n2212 = ~n876 & n1889 ;
  assign n2213 = ~n797 & n2212 ;
  assign n2217 = n436 ^ n383 ^ n350 ;
  assign n2218 = n249 ^ n37 ^ 1'b0 ;
  assign n2219 = n2217 & ~n2218 ;
  assign n2220 = ~n1679 & n2219 ;
  assign n2221 = n2220 ^ n969 ^ n151 ;
  assign n2215 = n1380 ^ n572 ^ 1'b0 ;
  assign n2216 = n767 & ~n2215 ;
  assign n2222 = n2221 ^ n2216 ^ x3 ;
  assign n2214 = ~n147 & n995 ;
  assign n2223 = n2222 ^ n2214 ^ n897 ;
  assign n2224 = ~n1553 & n1558 ;
  assign n2225 = ~n1264 & n2224 ;
  assign n2226 = ~n941 & n1156 ;
  assign n2230 = ( n622 & n639 ) | ( n622 & n1190 ) | ( n639 & n1190 ) ;
  assign n2227 = n188 | n1311 ;
  assign n2228 = n913 | n2227 ;
  assign n2229 = n2228 ^ n346 ^ 1'b0 ;
  assign n2231 = n2230 ^ n2229 ^ n55 ;
  assign n2232 = ~n498 & n1621 ;
  assign n2233 = n502 & ~n893 ;
  assign n2234 = n2017 | n2233 ;
  assign n2235 = ~n2232 & n2234 ;
  assign n2236 = n2231 & n2235 ;
  assign n2237 = n1184 ^ n875 ^ 1'b0 ;
  assign n2238 = n2237 ^ n916 ^ 1'b0 ;
  assign n2239 = n1435 | n2238 ;
  assign n2240 = n2239 ^ n874 ^ 1'b0 ;
  assign n2241 = ~n1410 & n2240 ;
  assign n2242 = n1453 ^ n91 ^ 1'b0 ;
  assign n2243 = n74 & ~n755 ;
  assign n2244 = n1874 & n2243 ;
  assign n2245 = ~n1109 & n2244 ;
  assign n2246 = ( ~n1295 & n2242 ) | ( ~n1295 & n2245 ) | ( n2242 & n2245 ) ;
  assign n2247 = ( ~n214 & n1539 ) | ( ~n214 & n2246 ) | ( n1539 & n2246 ) ;
  assign n2248 = n98 & ~n676 ;
  assign n2249 = ~n40 & n2248 ;
  assign n2250 = n98 & ~n285 ;
  assign n2251 = n993 | n2250 ;
  assign n2252 = n82 & ~n1171 ;
  assign n2253 = n2252 ^ n1890 ^ 1'b0 ;
  assign n2254 = n1120 ^ n491 ^ 1'b0 ;
  assign n2255 = n2158 ^ n2068 ^ 1'b0 ;
  assign n2256 = n2254 | n2255 ;
  assign n2257 = ~n548 & n1238 ;
  assign n2258 = n2257 ^ n1402 ^ 1'b0 ;
  assign n2259 = n1182 ^ n890 ^ 1'b0 ;
  assign n2260 = n649 & n1037 ;
  assign n2261 = n2260 ^ n1031 ^ 1'b0 ;
  assign n2262 = n1859 ^ n374 ^ 1'b0 ;
  assign n2263 = n2261 & n2262 ;
  assign n2264 = ~n2259 & n2263 ;
  assign n2265 = n1322 ^ n617 ^ 1'b0 ;
  assign n2266 = ~n802 & n2265 ;
  assign n2267 = n1484 & n2266 ;
  assign n2268 = n2267 ^ n836 ^ 1'b0 ;
  assign n2269 = n466 | n2143 ;
  assign n2270 = n1431 | n2269 ;
  assign n2276 = ( n132 & n217 ) | ( n132 & n532 ) | ( n217 & n532 ) ;
  assign n2273 = n1022 & n1164 ;
  assign n2271 = n2218 ^ n1055 ^ 1'b0 ;
  assign n2272 = n2242 & n2271 ;
  assign n2274 = n2273 ^ n2272 ^ 1'b0 ;
  assign n2275 = n1656 | n2274 ;
  assign n2277 = n2276 ^ n2275 ^ 1'b0 ;
  assign n2278 = n2084 & n2216 ;
  assign n2279 = n124 ^ n63 ^ 1'b0 ;
  assign n2280 = ~n184 & n2279 ;
  assign n2281 = n2280 ^ n957 ^ 1'b0 ;
  assign n2282 = n1245 ^ n74 ^ 1'b0 ;
  assign n2283 = n2282 ^ n411 ^ 1'b0 ;
  assign n2284 = n1875 ^ n126 ^ n55 ;
  assign n2285 = n1230 & ~n2284 ;
  assign n2286 = n2285 ^ n1599 ^ 1'b0 ;
  assign n2288 = n53 | n1912 ;
  assign n2287 = n177 & ~n782 ;
  assign n2289 = n2288 ^ n2287 ^ n1535 ;
  assign n2290 = n687 & n1482 ;
  assign n2291 = n218 & n2290 ;
  assign n2292 = n648 ^ n493 ^ 1'b0 ;
  assign n2293 = n2291 | n2292 ;
  assign n2294 = n2293 ^ n1433 ^ 1'b0 ;
  assign n2296 = ~n118 & n1178 ;
  assign n2295 = n360 & ~n1090 ;
  assign n2297 = n2296 ^ n2295 ^ 1'b0 ;
  assign n2298 = n97 | n2297 ;
  assign n2299 = n53 & n816 ;
  assign n2300 = n2299 ^ n1071 ^ 1'b0 ;
  assign n2301 = n195 & n791 ;
  assign n2302 = n2301 ^ x10 ^ 1'b0 ;
  assign n2303 = x6 & ~n332 ;
  assign n2304 = n2302 | n2303 ;
  assign n2305 = n1213 ^ n1017 ^ 1'b0 ;
  assign n2306 = ~n628 & n636 ;
  assign n2307 = ~n2305 & n2306 ;
  assign n2308 = n612 & ~n2307 ;
  assign n2309 = n2304 & n2308 ;
  assign n2310 = ~n131 & n1822 ;
  assign n2311 = ~n108 & n2310 ;
  assign n2312 = n2058 ^ n272 ^ 1'b0 ;
  assign n2313 = n1848 ^ n508 ^ n228 ;
  assign n2314 = ( n755 & n2217 ) | ( n755 & ~n2313 ) | ( n2217 & ~n2313 ) ;
  assign n2315 = n1701 ^ n1343 ^ 1'b0 ;
  assign n2316 = ~n2314 & n2315 ;
  assign n2317 = ( n795 & n1021 ) | ( n795 & n2316 ) | ( n1021 & n2316 ) ;
  assign n2318 = ~n32 & n1439 ;
  assign n2319 = n2318 ^ n1573 ^ 1'b0 ;
  assign n2320 = n187 ^ n78 ^ n49 ;
  assign n2321 = ~n1575 & n2320 ;
  assign n2322 = n2321 ^ n960 ^ n411 ;
  assign n2323 = ~n42 & n1410 ;
  assign n2324 = n2323 ^ x10 ^ 1'b0 ;
  assign n2325 = n1026 & ~n1249 ;
  assign n2326 = n2325 ^ n102 ^ 1'b0 ;
  assign n2327 = n406 & n525 ;
  assign n2328 = n119 & n908 ;
  assign n2329 = n2327 & ~n2328 ;
  assign n2330 = n2172 & n2329 ;
  assign n2331 = n345 ^ n271 ^ 1'b0 ;
  assign n2332 = ~n733 & n2331 ;
  assign n2333 = n838 & n2332 ;
  assign n2334 = ( n799 & ~n1139 ) | ( n799 & n2333 ) | ( ~n1139 & n2333 ) ;
  assign n2335 = n1416 ^ n461 ^ n142 ;
  assign n2336 = ~n203 & n780 ;
  assign n2337 = n2336 ^ n447 ^ 1'b0 ;
  assign n2338 = n1532 & ~n2337 ;
  assign n2339 = n2328 ^ n1389 ^ n426 ;
  assign n2340 = ~n401 & n2339 ;
  assign n2341 = n2340 ^ n887 ^ 1'b0 ;
  assign n2342 = n96 & n687 ;
  assign n2343 = n2342 ^ n349 ^ 1'b0 ;
  assign n2344 = n866 & n2343 ;
  assign n2345 = n928 ^ n125 ^ 1'b0 ;
  assign n2346 = n2344 | n2345 ;
  assign n2347 = n318 ^ n156 ^ 1'b0 ;
  assign n2348 = ~n98 & n1210 ;
  assign n2349 = ~n2025 & n2348 ;
  assign n2350 = ~n2179 & n2349 ;
  assign n2351 = n698 ^ n247 ^ 1'b0 ;
  assign n2352 = n1741 & n2351 ;
  assign n2353 = n871 ^ x5 ^ 1'b0 ;
  assign n2354 = n2328 & ~n2353 ;
  assign n2355 = n2354 ^ n726 ^ 1'b0 ;
  assign n2356 = n2355 ^ n567 ^ 1'b0 ;
  assign n2357 = n524 & n639 ;
  assign n2358 = n1061 | n2143 ;
  assign n2359 = n2358 ^ n605 ^ 1'b0 ;
  assign n2360 = n2359 ^ n908 ^ 1'b0 ;
  assign n2361 = n730 | n1798 ;
  assign n2362 = n2361 ^ n57 ^ 1'b0 ;
  assign n2363 = n1019 ^ n162 ^ n55 ;
  assign n2364 = n2362 & n2363 ;
  assign n2365 = ~n2014 & n2364 ;
  assign n2366 = ~n285 & n877 ;
  assign n2367 = n2365 & n2366 ;
  assign n2368 = ( n397 & ~n911 ) | ( n397 & n1632 ) | ( ~n911 & n1632 ) ;
  assign n2369 = n2368 ^ n1110 ^ 1'b0 ;
  assign n2370 = n876 & n2369 ;
  assign n2371 = n711 & ~n756 ;
  assign n2372 = n2371 ^ n1124 ^ 1'b0 ;
  assign n2373 = ( ~n441 & n1332 ) | ( ~n441 & n1499 ) | ( n1332 & n1499 ) ;
  assign n2374 = n124 & n1722 ;
  assign n2375 = ~n2373 & n2374 ;
  assign n2376 = n1339 & ~n2253 ;
  assign n2377 = n2376 ^ n1010 ^ 1'b0 ;
  assign n2378 = ( n493 & n922 ) | ( n493 & n1061 ) | ( n922 & n1061 ) ;
  assign n2379 = ~n104 & n855 ;
  assign n2380 = n2379 ^ n38 ^ 1'b0 ;
  assign n2381 = n1052 | n2380 ;
  assign n2382 = n965 & ~n2381 ;
  assign n2383 = n621 ^ n458 ^ 1'b0 ;
  assign n2384 = n586 & ~n2383 ;
  assign n2385 = ( n728 & n1115 ) | ( n728 & ~n2384 ) | ( n1115 & ~n2384 ) ;
  assign n2386 = n2382 | n2385 ;
  assign n2387 = n686 & ~n2386 ;
  assign n2388 = n2378 & ~n2387 ;
  assign n2389 = n2388 ^ n524 ^ 1'b0 ;
  assign n2390 = ~n1896 & n2236 ;
  assign n2391 = n95 & n1038 ;
  assign n2392 = n630 & n2391 ;
  assign n2393 = n1464 & n2392 ;
  assign n2394 = n2250 ^ n572 ^ 1'b0 ;
  assign n2395 = n1278 & ~n2394 ;
  assign n2396 = n799 ^ n121 ^ 1'b0 ;
  assign n2397 = n2328 & ~n2396 ;
  assign n2398 = n35 & n2397 ;
  assign n2399 = ~n2395 & n2398 ;
  assign n2402 = n67 & n101 ;
  assign n2400 = n159 | n700 ;
  assign n2401 = n2400 ^ n1343 ^ 1'b0 ;
  assign n2403 = n2402 ^ n2401 ^ n101 ;
  assign n2404 = n126 | n383 ;
  assign n2405 = n2404 ^ n1361 ^ 1'b0 ;
  assign n2407 = n108 & n1436 ;
  assign n2408 = n2407 ^ n973 ^ 1'b0 ;
  assign n2406 = n230 | n2307 ;
  assign n2409 = n2408 ^ n2406 ^ 1'b0 ;
  assign n2410 = n2131 ^ n617 ^ 1'b0 ;
  assign n2411 = n1642 & n2410 ;
  assign n2412 = ( n761 & ~n808 ) | ( n761 & n1253 ) | ( ~n808 & n1253 ) ;
  assign n2413 = ( n230 & n918 ) | ( n230 & n2412 ) | ( n918 & n2412 ) ;
  assign n2414 = n1406 & ~n1956 ;
  assign n2418 = ~n838 & n892 ;
  assign n2415 = n517 | n1859 ;
  assign n2416 = n1281 | n2415 ;
  assign n2417 = ~n1917 & n2416 ;
  assign n2419 = n2418 ^ n2417 ^ 1'b0 ;
  assign n2420 = n2419 ^ n77 ^ 1'b0 ;
  assign n2421 = n708 & n2420 ;
  assign n2422 = n471 & n2373 ;
  assign n2423 = n53 & ~n735 ;
  assign n2424 = n2337 ^ n1041 ^ 1'b0 ;
  assign n2425 = n459 & n2424 ;
  assign n2426 = ~n2423 & n2425 ;
  assign n2427 = n620 & n2426 ;
  assign n2428 = ~n670 & n2427 ;
  assign n2429 = n1686 ^ n1647 ^ n744 ;
  assign n2430 = n2075 ^ n400 ^ 1'b0 ;
  assign n2431 = ~n124 & n2430 ;
  assign n2432 = n657 & n1058 ;
  assign n2433 = ( n1120 & n2431 ) | ( n1120 & n2432 ) | ( n2431 & n2432 ) ;
  assign n2435 = n1315 ^ n792 ^ n484 ;
  assign n2434 = n1777 ^ n823 ^ n191 ;
  assign n2436 = n2435 ^ n2434 ^ n234 ;
  assign n2437 = n1245 ^ n230 ^ 1'b0 ;
  assign n2438 = n16 & n2437 ;
  assign n2439 = n129 & ~n485 ;
  assign n2440 = n2439 ^ n493 ^ 1'b0 ;
  assign n2441 = n1134 & ~n2440 ;
  assign n2442 = n2441 ^ n210 ^ 1'b0 ;
  assign n2443 = n2438 & ~n2442 ;
  assign n2444 = n2436 & n2443 ;
  assign n2445 = n411 & n2444 ;
  assign n2446 = ~n131 & n834 ;
  assign n2447 = ( ~n786 & n925 ) | ( ~n786 & n2337 ) | ( n925 & n2337 ) ;
  assign n2448 = n2447 ^ n982 ^ 1'b0 ;
  assign n2449 = ~n2446 & n2448 ;
  assign n2450 = n2449 ^ n59 ^ 1'b0 ;
  assign n2451 = n852 | n2450 ;
  assign n2452 = ( n729 & n759 ) | ( n729 & ~n1959 ) | ( n759 & ~n1959 ) ;
  assign n2453 = n1848 ^ n1594 ^ 1'b0 ;
  assign n2454 = n356 & n2225 ;
  assign n2455 = n1085 ^ n209 ^ 1'b0 ;
  assign n2456 = ~n414 & n2455 ;
  assign n2457 = n2456 ^ n571 ^ 1'b0 ;
  assign n2458 = n230 & ~n1945 ;
  assign n2459 = n2458 ^ n984 ^ 1'b0 ;
  assign n2460 = ( n57 & n1756 ) | ( n57 & ~n2459 ) | ( n1756 & ~n2459 ) ;
  assign n2461 = ~n205 & n662 ;
  assign n2462 = n1272 ^ n1225 ^ 1'b0 ;
  assign n2463 = n2461 & ~n2462 ;
  assign n2464 = n2463 ^ n1049 ^ 1'b0 ;
  assign n2465 = ~n1081 & n2464 ;
  assign n2466 = ~n1418 & n2465 ;
  assign n2468 = n154 & n1439 ;
  assign n2469 = n221 & n2468 ;
  assign n2467 = n1262 & ~n1921 ;
  assign n2470 = n2469 ^ n2467 ^ 1'b0 ;
  assign n2471 = n178 & ~n633 ;
  assign n2472 = n1365 | n2471 ;
  assign n2474 = n471 & ~n946 ;
  assign n2473 = n259 & n661 ;
  assign n2475 = n2474 ^ n2473 ^ 1'b0 ;
  assign n2476 = n2475 ^ n704 ^ 1'b0 ;
  assign n2477 = ( ~n501 & n578 ) | ( ~n501 & n990 ) | ( n578 & n990 ) ;
  assign n2478 = n2477 ^ n191 ^ 1'b0 ;
  assign n2479 = n1842 & n2478 ;
  assign n2480 = n1513 ^ n141 ^ 1'b0 ;
  assign n2481 = n525 & n2480 ;
  assign n2482 = n1525 | n2481 ;
  assign n2483 = ( n309 & n486 ) | ( n309 & ~n1706 ) | ( n486 & ~n1706 ) ;
  assign n2484 = n1917 ^ n341 ^ x1 ;
  assign n2485 = ~n951 & n2484 ;
  assign n2486 = n1307 ^ n1250 ^ 1'b0 ;
  assign n2487 = n2486 ^ n498 ^ 1'b0 ;
  assign n2488 = ~n1777 & n2487 ;
  assign n2489 = ( ~x3 & n1328 ) | ( ~x3 & n2266 ) | ( n1328 & n2266 ) ;
  assign n2490 = ~n54 & n358 ;
  assign n2492 = n686 ^ n183 ^ 1'b0 ;
  assign n2491 = n98 | n2359 ;
  assign n2493 = n2492 ^ n2491 ^ 1'b0 ;
  assign n2494 = ( n115 & ~n2179 ) | ( n115 & n2493 ) | ( ~n2179 & n2493 ) ;
  assign n2495 = ~n51 & n1917 ;
  assign n2496 = n448 & ~n767 ;
  assign n2497 = n2496 ^ n434 ^ 1'b0 ;
  assign n2498 = n241 & n1022 ;
  assign n2499 = ~n993 & n2498 ;
  assign n2500 = n2499 ^ n41 ^ n36 ;
  assign n2501 = n524 & ~n1589 ;
  assign n2502 = n1594 & n2501 ;
  assign n2503 = ( ~n1932 & n2320 ) | ( ~n1932 & n2502 ) | ( n2320 & n2502 ) ;
  assign n2504 = n2379 ^ n2198 ^ 1'b0 ;
  assign n2505 = n213 & ~n2504 ;
  assign n2506 = n2163 ^ n1131 ^ 1'b0 ;
  assign n2507 = n2168 & n2506 ;
  assign n2508 = ( n1475 & n2414 ) | ( n1475 & ~n2507 ) | ( n2414 & ~n2507 ) ;
  assign n2509 = n285 | n1549 ;
  assign n2510 = n1909 ^ n78 ^ 1'b0 ;
  assign n2511 = n2510 ^ n1133 ^ n259 ;
  assign n2512 = n1433 & n2511 ;
  assign n2513 = n2512 ^ n561 ^ 1'b0 ;
  assign n2514 = n2509 & n2513 ;
  assign n2515 = n2379 ^ n2237 ^ n2070 ;
  assign n2516 = n2515 ^ n762 ^ 1'b0 ;
  assign n2517 = n753 & ~n1082 ;
  assign n2518 = ~n801 & n825 ;
  assign n2519 = ~n1959 & n2518 ;
  assign n2520 = ~n736 & n1762 ;
  assign n2521 = n2148 & n2520 ;
  assign n2522 = n135 ^ n102 ^ 1'b0 ;
  assign n2523 = ~n2423 & n2522 ;
  assign n2524 = n41 ^ n23 ^ 1'b0 ;
  assign n2525 = n2524 ^ n1437 ^ 1'b0 ;
  assign n2526 = n1487 | n2525 ;
  assign n2529 = n941 | n1200 ;
  assign n2527 = n285 | n609 ;
  assign n2528 = n2527 ^ n1736 ^ 1'b0 ;
  assign n2530 = n2529 ^ n2528 ^ 1'b0 ;
  assign n2531 = ~n2526 & n2530 ;
  assign n2533 = n394 & ~n957 ;
  assign n2534 = n2533 ^ n1400 ^ 1'b0 ;
  assign n2532 = ( n973 & n1052 ) | ( n973 & n2250 ) | ( n1052 & n2250 ) ;
  assign n2535 = n2534 ^ n2532 ^ n607 ;
  assign n2536 = ~n1409 & n2535 ;
  assign n2537 = n2278 & n2536 ;
  assign n2538 = ( n68 & ~n1441 ) | ( n68 & n1464 ) | ( ~n1441 & n1464 ) ;
  assign n2539 = n2538 ^ n1527 ^ n1485 ;
  assign n2543 = ~n890 & n1245 ;
  assign n2544 = n2543 ^ n135 ^ 1'b0 ;
  assign n2540 = n1210 ^ n78 ^ 1'b0 ;
  assign n2541 = n1026 & ~n2540 ;
  assign n2542 = n469 & ~n2541 ;
  assign n2545 = n2544 ^ n2542 ^ n1339 ;
  assign n2546 = n2432 ^ n784 ^ 1'b0 ;
  assign n2547 = n465 ^ n174 ^ 1'b0 ;
  assign n2548 = n1231 & ~n2547 ;
  assign n2549 = n2548 ^ n1468 ^ 1'b0 ;
  assign n2550 = n852 | n2549 ;
  assign n2551 = n1459 | n2550 ;
  assign n2552 = ( n1076 & n1962 ) | ( n1076 & n2551 ) | ( n1962 & n2551 ) ;
  assign n2553 = n186 & n923 ;
  assign n2554 = n1481 ^ n371 ^ 1'b0 ;
  assign n2555 = ~n2553 & n2554 ;
  assign n2556 = n164 & n1238 ;
  assign n2557 = ~n511 & n2556 ;
  assign n2558 = n879 & ~n1992 ;
  assign n2559 = n1959 ^ n717 ^ 1'b0 ;
  assign n2560 = n1547 & n2559 ;
  assign n2561 = n91 & ~n1456 ;
  assign n2562 = n65 | n961 ;
  assign n2563 = n2562 ^ n2314 ^ 1'b0 ;
  assign n2564 = n1276 ^ n249 ^ 1'b0 ;
  assign n2565 = n759 | n2564 ;
  assign n2566 = n2565 ^ n1368 ^ 1'b0 ;
  assign n2567 = n1609 & n2566 ;
  assign n2568 = n2567 ^ n174 ^ 1'b0 ;
  assign n2569 = ~n170 & n1371 ;
  assign n2570 = n1527 & n2569 ;
  assign n2571 = n2570 ^ n1553 ^ 1'b0 ;
  assign n2572 = n652 ^ n151 ^ 1'b0 ;
  assign n2573 = n544 & ~n2572 ;
  assign n2574 = n2573 ^ n2002 ^ 1'b0 ;
  assign n2575 = n2571 & ~n2574 ;
  assign n2576 = n41 & ~n344 ;
  assign n2577 = n247 & n2576 ;
  assign n2579 = n1061 & n1491 ;
  assign n2578 = n112 | n1895 ;
  assign n2580 = n2579 ^ n2578 ^ 1'b0 ;
  assign n2581 = n2134 ^ n1302 ^ 1'b0 ;
  assign n2582 = n2374 & n2581 ;
  assign n2583 = n1017 ^ n436 ^ x3 ;
  assign n2584 = n26 | n1630 ;
  assign n2585 = n2583 | n2584 ;
  assign n2586 = n2585 ^ n1120 ^ 1'b0 ;
  assign n2587 = ~n168 & n2118 ;
  assign n2588 = n654 ^ n249 ^ 1'b0 ;
  assign n2589 = ( ~n190 & n1853 ) | ( ~n190 & n2588 ) | ( n1853 & n2588 ) ;
  assign n2595 = n1575 ^ n999 ^ 1'b0 ;
  assign n2596 = n187 & n2595 ;
  assign n2590 = n521 ^ n48 ^ 1'b0 ;
  assign n2591 = n35 & n2590 ;
  assign n2592 = n2591 ^ n567 ^ 1'b0 ;
  assign n2593 = ~n313 & n695 ;
  assign n2594 = ~n2592 & n2593 ;
  assign n2597 = n2596 ^ n2594 ^ 1'b0 ;
  assign n2598 = ~n1682 & n2597 ;
  assign n2599 = n2598 ^ n583 ^ 1'b0 ;
  assign n2600 = n54 & ~n515 ;
  assign n2601 = n598 & n2600 ;
  assign n2602 = n2601 ^ n2149 ^ 1'b0 ;
  assign n2604 = n1521 ^ n484 ^ 1'b0 ;
  assign n2605 = n2604 ^ n567 ^ 1'b0 ;
  assign n2603 = ~n772 & n2333 ;
  assign n2606 = n2605 ^ n2603 ^ n1032 ;
  assign n2607 = ~n2597 & n2606 ;
  assign n2608 = n57 & ~n1353 ;
  assign n2609 = ~n2510 & n2608 ;
  assign n2610 = n2609 ^ n1647 ^ n1453 ;
  assign n2611 = n324 & ~n627 ;
  assign n2612 = ~n448 & n2611 ;
  assign n2613 = n1623 | n2612 ;
  assign n2614 = n2613 ^ n1589 ^ n1175 ;
  assign n2615 = n2111 ^ n588 ^ 1'b0 ;
  assign n2616 = n2615 ^ n2160 ^ 1'b0 ;
  assign n2617 = ( ~n755 & n1296 ) | ( ~n755 & n1569 ) | ( n1296 & n1569 ) ;
  assign n2618 = ( n431 & n829 ) | ( n431 & n1063 ) | ( n829 & n1063 ) ;
  assign n2619 = n44 & n2618 ;
  assign n2620 = n2617 & ~n2619 ;
  assign n2621 = ~n1061 & n2276 ;
  assign n2622 = n2621 ^ n23 ^ 1'b0 ;
  assign n2623 = n2101 ^ n645 ^ 1'b0 ;
  assign n2624 = n1096 ^ n299 ^ 1'b0 ;
  assign n2625 = n1078 & ~n2624 ;
  assign n2626 = ~n1021 & n2370 ;
  assign n2627 = n2626 ^ n1056 ^ 1'b0 ;
  assign n2628 = ( x4 & n408 ) | ( x4 & ~n1436 ) | ( n408 & ~n1436 ) ;
  assign n2629 = n1381 | n2628 ;
  assign n2630 = n30 & ~n2629 ;
  assign n2643 = n2095 ^ n259 ^ 1'b0 ;
  assign n2644 = n2073 & ~n2643 ;
  assign n2635 = n435 ^ n431 ^ n152 ;
  assign n2634 = n441 & ~n1682 ;
  assign n2636 = n2635 ^ n2634 ^ 1'b0 ;
  assign n2637 = n2636 ^ n2198 ^ 1'b0 ;
  assign n2638 = n1938 & n2637 ;
  assign n2639 = n1110 ^ n1073 ^ 1'b0 ;
  assign n2640 = n1079 | n2639 ;
  assign n2641 = n2640 ^ n2601 ^ 1'b0 ;
  assign n2642 = n2638 & n2641 ;
  assign n2631 = n30 | n513 ;
  assign n2632 = n169 & ~n2631 ;
  assign n2633 = n2632 ^ n1255 ^ 1'b0 ;
  assign n2645 = n2644 ^ n2642 ^ n2633 ;
  assign n2646 = n18 & n2645 ;
  assign n2647 = n1022 ^ n953 ^ 1'b0 ;
  assign n2648 = n246 & ~n2647 ;
  assign n2649 = n2648 ^ n1729 ^ n714 ;
  assign n2650 = n2305 ^ n1153 ^ n1090 ;
  assign n2651 = ~n1317 & n2615 ;
  assign n2652 = ~n63 & n2651 ;
  assign n2653 = ( n1842 & n2145 ) | ( n1842 & ~n2652 ) | ( n2145 & ~n2652 ) ;
  assign n2654 = n1554 & n1932 ;
  assign n2655 = n2654 ^ n394 ^ 1'b0 ;
  assign n2656 = n2655 ^ n2128 ^ 1'b0 ;
  assign n2657 = n1515 | n2656 ;
  assign n2658 = ~n96 & n655 ;
  assign n2659 = n293 | n2658 ;
  assign n2660 = n2523 | n2659 ;
  assign n2661 = ( n583 & n1107 ) | ( n583 & n1282 ) | ( n1107 & n1282 ) ;
  assign n2662 = n2661 ^ n1241 ^ 1'b0 ;
  assign n2663 = ~n536 & n1085 ;
  assign n2664 = n2454 & n2663 ;
  assign n2665 = n1693 ^ n1355 ^ n664 ;
  assign n2666 = n89 & n448 ;
  assign n2667 = ( n1862 & n2665 ) | ( n1862 & ~n2666 ) | ( n2665 & ~n2666 ) ;
  assign n2668 = ~n1049 & n2658 ;
  assign n2670 = n351 & n1932 ;
  assign n2671 = n667 & n2670 ;
  assign n2669 = ~n859 & n1110 ;
  assign n2672 = n2671 ^ n2669 ^ 1'b0 ;
  assign n2673 = n1345 ^ n1267 ^ 1'b0 ;
  assign n2677 = n1460 | n1485 ;
  assign n2674 = n493 & ~n2477 ;
  assign n2675 = n2513 & n2674 ;
  assign n2676 = ~n2405 & n2675 ;
  assign n2678 = n2677 ^ n2676 ^ 1'b0 ;
  assign n2679 = n1527 ^ n1084 ^ n368 ;
  assign n2681 = n818 ^ n706 ^ 1'b0 ;
  assign n2682 = n1839 & n2681 ;
  assign n2680 = n1049 ^ n75 ^ 1'b0 ;
  assign n2683 = n2682 ^ n2680 ^ 1'b0 ;
  assign n2684 = n1959 & ~n2683 ;
  assign n2685 = n251 ^ n126 ^ 1'b0 ;
  assign n2686 = ~n139 & n2685 ;
  assign n2687 = ~n426 & n2606 ;
  assign n2688 = n2373 & ~n2687 ;
  assign n2689 = n2688 ^ n1680 ^ 1'b0 ;
  assign n2690 = n2243 & n2474 ;
  assign n2691 = ~n1309 & n2690 ;
  assign n2692 = n2691 ^ n467 ^ n400 ;
  assign n2693 = n2177 ^ n1037 ^ n415 ;
  assign n2694 = n2693 ^ n202 ^ 1'b0 ;
  assign n2698 = n2601 ^ n521 ^ 1'b0 ;
  assign n2699 = ( n440 & ~n704 ) | ( n440 & n2698 ) | ( ~n704 & n2698 ) ;
  assign n2695 = n1554 ^ n368 ^ 1'b0 ;
  assign n2696 = n1319 | n2695 ;
  assign n2697 = ( n569 & n1216 ) | ( n569 & n2696 ) | ( n1216 & n2696 ) ;
  assign n2700 = n2699 ^ n2697 ^ 1'b0 ;
  assign n2701 = n1052 | n2700 ;
  assign n2702 = n2694 & n2701 ;
  assign n2703 = n940 & n1099 ;
  assign n2704 = ~n126 & n2703 ;
  assign n2705 = ( n338 & n1903 ) | ( n338 & ~n2704 ) | ( n1903 & ~n2704 ) ;
  assign n2706 = n569 & n1793 ;
  assign n2709 = n2583 ^ n730 ^ 1'b0 ;
  assign n2710 = ~n809 & n2709 ;
  assign n2707 = n1945 ^ n1722 ^ 1'b0 ;
  assign n2708 = n811 | n2707 ;
  assign n2711 = n2710 ^ n2708 ^ 1'b0 ;
  assign n2712 = n2489 | n2711 ;
  assign n2713 = n1133 ^ n870 ^ 1'b0 ;
  assign n2714 = n119 & n963 ;
  assign n2715 = n2714 ^ n1642 ^ 1'b0 ;
  assign n2716 = n1506 & ~n2715 ;
  assign n2717 = n305 & n2716 ;
  assign n2718 = ~n2217 & n2717 ;
  assign n2719 = n1184 | n1882 ;
  assign n2720 = ~n16 & n2719 ;
  assign n2721 = n360 & ~n1139 ;
  assign n2722 = n2186 ^ n1185 ^ 1'b0 ;
  assign n2723 = ( ~n581 & n2721 ) | ( ~n581 & n2722 ) | ( n2721 & n2722 ) ;
  assign n2724 = n1169 & n1587 ;
  assign n2725 = n2724 ^ n1185 ^ 1'b0 ;
  assign n2726 = n141 & ~n1912 ;
  assign n2727 = n780 & ~n2726 ;
  assign n2728 = n922 | n1353 ;
  assign n2729 = ~n276 & n2728 ;
  assign n2730 = n164 & n1061 ;
  assign n2731 = n2730 ^ n1395 ^ 1'b0 ;
  assign n2732 = n2731 ^ n1357 ^ n1058 ;
  assign n2733 = n2732 ^ n698 ^ 1'b0 ;
  assign n2734 = n985 & n2471 ;
  assign n2735 = n2734 ^ n2291 ^ 1'b0 ;
  assign n2736 = n1801 ^ n564 ^ 1'b0 ;
  assign n2737 = n345 ^ n78 ^ 1'b0 ;
  assign n2738 = ~n1866 & n2737 ;
  assign n2739 = ~n957 & n2030 ;
  assign n2740 = ~n777 & n2739 ;
  assign n2741 = n1882 ^ n570 ^ 1'b0 ;
  assign n2742 = n1364 ^ n750 ^ 1'b0 ;
  assign n2743 = n464 & n2742 ;
  assign n2744 = n686 | n1247 ;
  assign n2745 = n2744 ^ n178 ^ 1'b0 ;
  assign n2746 = ( n1699 & ~n2111 ) | ( n1699 & n2745 ) | ( ~n2111 & n2745 ) ;
  assign n2747 = n172 & ~n2405 ;
  assign n2748 = ~n263 & n1813 ;
  assign n2749 = n2748 ^ n2220 ^ 1'b0 ;
  assign n2750 = ( n776 & ~n842 ) | ( n776 & n1153 ) | ( ~n842 & n1153 ) ;
  assign n2751 = n2750 ^ n2642 ^ n2258 ;
  assign n2755 = n354 ^ n352 ^ 1'b0 ;
  assign n2756 = n241 & ~n2755 ;
  assign n2752 = n320 & ~n1046 ;
  assign n2753 = n1256 | n2752 ;
  assign n2754 = n1341 | n2753 ;
  assign n2757 = n2756 ^ n2754 ^ 1'b0 ;
  assign n2758 = n1465 ^ n698 ^ 1'b0 ;
  assign n2759 = ( n694 & ~n808 ) | ( n694 & n1468 ) | ( ~n808 & n1468 ) ;
  assign n2760 = n2759 ^ n395 ^ 1'b0 ;
  assign n2761 = n2758 | n2760 ;
  assign n2762 = n230 & n1105 ;
  assign n2763 = n2762 ^ n188 ^ 1'b0 ;
  assign n2764 = n1874 & n2494 ;
  assign n2765 = ( n44 & n272 ) | ( n44 & n1253 ) | ( n272 & n1253 ) ;
  assign n2766 = n1483 ^ n875 ^ n408 ;
  assign n2767 = n37 & n630 ;
  assign n2768 = ~n2261 & n2767 ;
  assign n2769 = n1835 ^ n1791 ^ n331 ;
  assign n2770 = n1684 & n2769 ;
  assign n2771 = n1652 ^ n51 ^ 1'b0 ;
  assign n2772 = ~n2770 & n2771 ;
  assign n2773 = ~n263 & n836 ;
  assign n2774 = n2773 ^ n995 ^ 1'b0 ;
  assign n2775 = n1280 & n2774 ;
  assign n2776 = n1062 & ~n2775 ;
  assign n2777 = n2108 ^ n1083 ^ 1'b0 ;
  assign n2778 = n2776 | n2777 ;
  assign n2779 = x0 & n2778 ;
  assign n2780 = n37 & ~n2779 ;
  assign n2781 = n2780 ^ n684 ^ 1'b0 ;
  assign n2782 = n1001 & n2053 ;
  assign n2783 = n2561 & n2782 ;
  assign n2784 = n400 ^ n313 ^ 1'b0 ;
  assign n2785 = n2784 ^ n260 ^ n217 ;
  assign n2786 = ~n328 & n1429 ;
  assign n2787 = n794 ^ n532 ^ n184 ;
  assign n2788 = n991 & n2787 ;
  assign n2789 = n2788 ^ n105 ^ 1'b0 ;
  assign n2790 = n2789 ^ n1363 ^ 1'b0 ;
  assign n2791 = n2790 ^ n2352 ^ 1'b0 ;
  assign n2792 = n2786 & n2791 ;
  assign n2793 = ~n2785 & n2792 ;
  assign n2794 = n2161 & ~n2793 ;
  assign n2795 = n1095 ^ n1001 ^ n192 ;
  assign n2797 = n1938 ^ n889 ^ n839 ;
  assign n2798 = n2797 ^ x3 ^ 1'b0 ;
  assign n2796 = n1075 & ~n2005 ;
  assign n2799 = n2798 ^ n2796 ^ 1'b0 ;
  assign n2800 = n2799 ^ n2384 ^ 1'b0 ;
  assign n2801 = n1990 & n2800 ;
  assign n2802 = n2795 & n2801 ;
  assign n2803 = n1718 ^ n101 ^ 1'b0 ;
  assign n2804 = ~n548 & n2803 ;
  assign n2805 = n2804 ^ n1234 ^ 1'b0 ;
  assign n2806 = ( n101 & n257 ) | ( n101 & n472 ) | ( n257 & n472 ) ;
  assign n2807 = n2357 | n2806 ;
  assign n2811 = n238 | n2307 ;
  assign n2808 = n772 ^ n508 ^ 1'b0 ;
  assign n2809 = n868 ^ x10 ^ 1'b0 ;
  assign n2810 = n2808 | n2809 ;
  assign n2812 = n2811 ^ n2810 ^ 1'b0 ;
  assign n2813 = n2395 & n2812 ;
  assign n2814 = n2813 ^ n1308 ^ 1'b0 ;
  assign n2815 = n145 & n2814 ;
  assign n2816 = n324 & n951 ;
  assign n2817 = n2048 ^ n949 ^ 1'b0 ;
  assign n2818 = n1455 ^ n814 ^ 1'b0 ;
  assign n2819 = n496 | n2818 ;
  assign n2820 = n1463 ^ n740 ^ 1'b0 ;
  assign n2821 = ~n886 & n2232 ;
  assign n2822 = n744 | n2821 ;
  assign n2823 = n2198 | n2822 ;
  assign n2824 = n2823 ^ n2054 ^ 1'b0 ;
  assign n2825 = n2824 ^ n1957 ^ 1'b0 ;
  assign n2826 = n1013 ^ n381 ^ 1'b0 ;
  assign n2827 = n888 & n2826 ;
  assign n2828 = ( n1168 & n2241 ) | ( n1168 & n2804 ) | ( n2241 & n2804 ) ;
  assign n2829 = n1025 & n2828 ;
  assign n2830 = n2829 ^ n1190 ^ 1'b0 ;
  assign n2831 = n2827 & n2830 ;
  assign n2832 = ~n505 & n2456 ;
  assign n2833 = n1529 & ~n2832 ;
  assign n2834 = n2695 ^ n1216 ^ 1'b0 ;
  assign n2835 = n657 | n2834 ;
  assign n2836 = n102 | n2835 ;
  assign n2837 = n401 & n1125 ;
  assign n2838 = n2837 ^ n1878 ^ 1'b0 ;
  assign n2839 = n430 & ~n2838 ;
  assign n2840 = n1302 ^ n180 ^ 1'b0 ;
  assign n2841 = n451 & ~n1749 ;
  assign n2842 = n2619 ^ n2075 ^ 1'b0 ;
  assign n2843 = n2841 | n2842 ;
  assign n2844 = n2196 ^ n524 ^ n272 ;
  assign n2845 = n882 | n2844 ;
  assign n2846 = n1210 ^ n26 ^ 1'b0 ;
  assign n2847 = n2846 ^ n1212 ^ 1'b0 ;
  assign n2848 = n587 | n2847 ;
  assign n2849 = n2217 ^ n1287 ^ n41 ;
  assign n2850 = n186 & ~n539 ;
  assign n2851 = ~n2849 & n2850 ;
  assign n2852 = n1849 ^ n1274 ^ 1'b0 ;
  assign n2853 = n2851 | n2852 ;
  assign n2854 = n1810 ^ n1133 ^ n799 ;
  assign n2855 = ~n2114 & n2854 ;
  assign n2856 = n631 | n1319 ;
  assign n2857 = n2856 ^ n480 ^ 1'b0 ;
  assign n2858 = n966 ^ n37 ^ 1'b0 ;
  assign n2859 = ~n2857 & n2858 ;
  assign n2860 = n360 & n1745 ;
  assign n2861 = ( n1075 & n1292 ) | ( n1075 & n2860 ) | ( n1292 & n2860 ) ;
  assign n2862 = n2861 ^ n2736 ^ 1'b0 ;
  assign n2863 = n1465 | n2862 ;
  assign n2864 = n2176 | n2502 ;
  assign n2865 = n1172 | n2864 ;
  assign n2866 = n2220 & ~n2865 ;
  assign n2867 = n2535 ^ n1157 ^ 1'b0 ;
  assign n2868 = n465 ^ n401 ^ 1'b0 ;
  assign n2869 = n276 & ~n2088 ;
  assign n2870 = ( ~n147 & n855 ) | ( ~n147 & n2869 ) | ( n855 & n2869 ) ;
  assign n2871 = n511 & n2870 ;
  assign n2872 = n1857 & n2828 ;
  assign n2873 = n2320 ^ n827 ^ n554 ;
  assign n2874 = ( ~n38 & n414 ) | ( ~n38 & n2873 ) | ( n414 & n2873 ) ;
  assign n2875 = n2874 ^ n961 ^ 1'b0 ;
  assign n2876 = ~n1129 & n2875 ;
  assign n2877 = n2876 ^ n2623 ^ n448 ;
  assign n2878 = ( n710 & n848 ) | ( n710 & ~n2259 ) | ( n848 & ~n2259 ) ;
  assign n2879 = n2058 & n2878 ;
  assign n2880 = n1858 & ~n2374 ;
  assign n2881 = ~n250 & n2880 ;
  assign n2882 = n809 & n2881 ;
  assign n2884 = n1095 ^ n1056 ^ 1'b0 ;
  assign n2883 = n1491 & ~n2306 ;
  assign n2885 = n2884 ^ n2883 ^ 1'b0 ;
  assign n2886 = ~n205 & n1339 ;
  assign n2887 = n2363 ^ n2021 ^ 1'b0 ;
  assign n2888 = n705 | n2887 ;
  assign n2889 = ( n511 & n923 ) | ( n511 & n2150 ) | ( n923 & n2150 ) ;
  assign n2890 = n861 ^ x6 ^ 1'b0 ;
  assign n2891 = n2174 & n2890 ;
  assign n2892 = n2889 & n2891 ;
  assign n2893 = ( n1045 & ~n1545 ) | ( n1045 & n2576 ) | ( ~n1545 & n2576 ) ;
  assign n2894 = n2581 ^ n2180 ^ 1'b0 ;
  assign n2895 = ~n656 & n2894 ;
  assign n2898 = n2217 ^ n99 ^ 1'b0 ;
  assign n2896 = n1355 ^ n867 ^ 1'b0 ;
  assign n2897 = n2896 ^ n2869 ^ 1'b0 ;
  assign n2899 = n2898 ^ n2897 ^ 1'b0 ;
  assign n2900 = n2387 ^ x0 ^ 1'b0 ;
  assign n2901 = n2899 & ~n2900 ;
  assign n2902 = n1260 ^ n214 ^ 1'b0 ;
  assign n2903 = n2901 & n2902 ;
  assign n2904 = n2903 ^ n100 ^ 1'b0 ;
  assign n2905 = n2034 & n2524 ;
  assign n2906 = n554 ^ n142 ^ 1'b0 ;
  assign n2907 = n2906 ^ n2452 ^ 1'b0 ;
  assign n2908 = n2589 ^ n1078 ^ 1'b0 ;
  assign n2909 = ~n2367 & n2908 ;
  assign n2910 = n1110 ^ n650 ^ 1'b0 ;
  assign n2911 = ( n1491 & n2184 ) | ( n1491 & ~n2910 ) | ( n2184 & ~n2910 ) ;
  assign n2912 = n312 & ~n890 ;
  assign n2913 = ~n318 & n2912 ;
  assign n2914 = n1909 & ~n2913 ;
  assign n2915 = n2914 ^ n1226 ^ 1'b0 ;
  assign n2916 = n46 & n2915 ;
  assign n2917 = n2887 ^ n1662 ^ 1'b0 ;
  assign n2918 = ~n797 & n856 ;
  assign n2919 = n925 ^ n590 ^ x6 ;
  assign n2920 = n2919 ^ n1418 ^ 1'b0 ;
  assign n2921 = n1026 & n1897 ;
  assign n2922 = n2921 ^ n834 ^ 1'b0 ;
  assign n2923 = ~n2920 & n2922 ;
  assign n2924 = n2846 ^ n664 ^ 1'b0 ;
  assign n2925 = n2384 & ~n2924 ;
  assign n2926 = n360 | n1636 ;
  assign n2927 = ~n95 & n2352 ;
  assign n2928 = n231 & n2927 ;
  assign n2929 = n2411 ^ n1467 ^ 1'b0 ;
  assign n2930 = n2435 & ~n2929 ;
  assign n2931 = n2930 ^ n1623 ^ 1'b0 ;
  assign n2932 = ~n2928 & n2931 ;
  assign n2933 = n2806 ^ n889 ^ 1'b0 ;
  assign n2934 = n2323 & ~n2693 ;
  assign n2935 = n2045 ^ n686 ^ 1'b0 ;
  assign n2936 = n89 & n855 ;
  assign n2937 = n2936 ^ n2550 ^ 1'b0 ;
  assign n2938 = n2192 ^ n1664 ^ 1'b0 ;
  assign n2939 = n2025 | n2938 ;
  assign n2941 = n395 & n1664 ;
  assign n2942 = n2941 ^ n2603 ^ 1'b0 ;
  assign n2940 = n826 & ~n2627 ;
  assign n2943 = n2942 ^ n2940 ^ n2251 ;
  assign n2948 = n1861 ^ n427 ^ 1'b0 ;
  assign n2949 = n2304 | n2948 ;
  assign n2950 = n1813 & ~n2949 ;
  assign n2951 = n170 & n2950 ;
  assign n2944 = ~n1357 & n1428 ;
  assign n2945 = ( n1727 & n1768 ) | ( n1727 & ~n2944 ) | ( n1768 & ~n2944 ) ;
  assign n2946 = ( n852 & n2134 ) | ( n852 & n2945 ) | ( n2134 & n2945 ) ;
  assign n2947 = n1811 & ~n2946 ;
  assign n2952 = n2951 ^ n2947 ^ 1'b0 ;
  assign n2953 = n1200 ^ n201 ^ 1'b0 ;
  assign n2954 = n2953 ^ n2251 ^ n313 ;
  assign n2955 = n2535 ^ n934 ^ n849 ;
  assign n2956 = n532 ^ n484 ^ 1'b0 ;
  assign n2957 = n2939 ^ n1990 ^ 1'b0 ;
  assign n2958 = ~n2956 & n2957 ;
  assign n2959 = n124 | n744 ;
  assign n2960 = n865 & ~n2959 ;
  assign n2961 = n893 & n2960 ;
  assign n2962 = ~n299 & n2876 ;
  assign n2963 = n1150 & n2962 ;
  assign n2964 = n1220 & ~n1832 ;
  assign n2965 = ~n2963 & n2964 ;
  assign n2966 = n2965 ^ n1506 ^ 1'b0 ;
  assign n2967 = ( n1076 & n1415 ) | ( n1076 & n2966 ) | ( n1415 & n2966 ) ;
  assign n2968 = n1841 ^ n1362 ^ 1'b0 ;
  assign n2969 = ~n1351 & n2968 ;
  assign n2970 = n96 & n411 ;
  assign n2971 = n87 & n2970 ;
  assign n2972 = n2971 ^ n57 ^ 1'b0 ;
  assign n2973 = n192 & n887 ;
  assign n2974 = n2973 ^ x4 ^ 1'b0 ;
  assign n2975 = n1062 ^ n418 ^ 1'b0 ;
  assign n2976 = ~n1553 & n2975 ;
  assign n2977 = ( n191 & ~n890 ) | ( n191 & n2976 ) | ( ~n890 & n2976 ) ;
  assign n2978 = n755 ^ n214 ^ 1'b0 ;
  assign n2979 = n690 & n2978 ;
  assign n2980 = n2977 & ~n2979 ;
  assign n2981 = n760 & n1436 ;
  assign n2982 = n829 & n2981 ;
  assign n2983 = ~n1081 & n1724 ;
  assign n2984 = ( ~n1886 & n2333 ) | ( ~n1886 & n2983 ) | ( n2333 & n2983 ) ;
  assign n2985 = n2984 ^ n1547 ^ n1460 ;
  assign n2986 = ~n384 & n897 ;
  assign n2987 = ~n2925 & n2986 ;
  assign n2988 = n2987 ^ n2735 ^ 1'b0 ;
  assign n2989 = n2029 & n2988 ;
  assign n2990 = n145 | n156 ;
  assign n2991 = n823 ^ n461 ^ n304 ;
  assign n2992 = n2991 ^ n2893 ^ n1319 ;
  assign n2993 = n105 & n159 ;
  assign n2994 = n2992 & n2993 ;
  assign n2995 = n411 | n1311 ;
  assign n2996 = n1610 & n2995 ;
  assign n2997 = ~n463 & n2996 ;
  assign n2998 = n1395 | n2986 ;
  assign n2999 = n2998 ^ n1244 ^ 1'b0 ;
  assign n3000 = n1118 & ~n1246 ;
  assign n3001 = n3000 ^ n2176 ^ n2048 ;
  assign n3002 = ( n760 & n1243 ) | ( n760 & ~n2631 ) | ( n1243 & ~n2631 ) ;
  assign n3003 = n1078 & n3002 ;
  assign n3004 = ( n390 & n1339 ) | ( n390 & n1805 ) | ( n1339 & n1805 ) ;
  assign n3005 = n3003 & ~n3004 ;
  assign n3006 = n41 & ~n3005 ;
  assign n3007 = n765 ^ n676 ^ 1'b0 ;
  assign n3008 = ~n142 & n2888 ;
  assign n3009 = ( n688 & ~n1018 ) | ( n688 & n1634 ) | ( ~n1018 & n1634 ) ;
  assign n3010 = n1866 ^ n711 ^ n28 ;
  assign n3011 = n1661 ^ n32 ^ 1'b0 ;
  assign n3012 = n54 & ~n401 ;
  assign n3013 = n3012 ^ n1467 ^ 1'b0 ;
  assign n3014 = ( n641 & ~n993 ) | ( n641 & n1017 ) | ( ~n993 & n1017 ) ;
  assign n3015 = n3014 ^ n308 ^ 1'b0 ;
  assign n3016 = n3013 & ~n3015 ;
  assign n3017 = n1226 ^ n197 ^ 1'b0 ;
  assign n3018 = n3016 & n3017 ;
  assign n3027 = n1263 ^ n469 ^ 1'b0 ;
  assign n3028 = n503 & ~n3027 ;
  assign n3029 = n824 & n3028 ;
  assign n3019 = n2381 ^ n909 ^ n656 ;
  assign n3020 = n331 & ~n607 ;
  assign n3021 = n1733 ^ n1151 ^ 1'b0 ;
  assign n3022 = n3020 & ~n3021 ;
  assign n3023 = n3022 ^ n1929 ^ 1'b0 ;
  assign n3024 = n3019 & n3023 ;
  assign n3025 = ( n87 & ~n2622 ) | ( n87 & n3024 ) | ( ~n2622 & n3024 ) ;
  assign n3026 = ~n2951 & n3025 ;
  assign n3030 = n3029 ^ n3026 ^ 1'b0 ;
  assign n3031 = n1483 ^ n1296 ^ n1184 ;
  assign n3032 = n3031 ^ n1996 ^ 1'b0 ;
  assign n3033 = n564 & ~n3032 ;
  assign n3034 = ~n43 & n1274 ;
  assign n3035 = n1565 & ~n3034 ;
  assign n3036 = ~n364 & n850 ;
  assign n3037 = n49 & n3036 ;
  assign n3038 = n3037 ^ n2995 ^ 1'b0 ;
  assign n3039 = n2077 ^ n585 ^ 1'b0 ;
  assign n3040 = n445 & n782 ;
  assign n3041 = ~n1348 & n3040 ;
  assign n3042 = n1752 | n3041 ;
  assign n3043 = n1367 & ~n3042 ;
  assign n3044 = ( n48 & n578 ) | ( n48 & n1118 ) | ( n578 & n1118 ) ;
  assign n3045 = n328 & n3044 ;
  assign n3046 = ~n250 & n1293 ;
  assign n3047 = n1327 | n3046 ;
  assign n3048 = n3047 ^ n1628 ^ 1'b0 ;
  assign n3049 = n1386 ^ n994 ^ 1'b0 ;
  assign n3050 = ~n3048 & n3049 ;
  assign n3051 = ~n96 & n3050 ;
  assign n3052 = n502 | n3051 ;
  assign n3053 = n3045 & ~n3052 ;
  assign n3054 = ( n26 & n3043 ) | ( n26 & ~n3053 ) | ( n3043 & ~n3053 ) ;
  assign n3056 = n308 & n1039 ;
  assign n3055 = n420 & ~n1298 ;
  assign n3057 = n3056 ^ n3055 ^ 1'b0 ;
  assign n3058 = ~n1591 & n3057 ;
  assign n3059 = n1122 & n3058 ;
  assign n3060 = ( n32 & n279 ) | ( n32 & n2108 ) | ( n279 & n2108 ) ;
  assign n3061 = n3059 | n3060 ;
  assign n3062 = ( n82 & n2886 ) | ( n82 & ~n3061 ) | ( n2886 & ~n3061 ) ;
  assign n3063 = n3062 ^ n2312 ^ 1'b0 ;
  assign n3064 = n3054 & ~n3063 ;
  assign n3067 = n184 ^ n48 ^ 1'b0 ;
  assign n3068 = n28 | n551 ;
  assign n3069 = n1324 & ~n3068 ;
  assign n3070 = n3067 | n3069 ;
  assign n3065 = n957 ^ n63 ^ 1'b0 ;
  assign n3066 = n240 | n3065 ;
  assign n3071 = n3070 ^ n3066 ^ 1'b0 ;
  assign n3072 = ~n1082 & n1815 ;
  assign n3073 = ~n1296 & n3072 ;
  assign n3074 = n3073 ^ n929 ^ 1'b0 ;
  assign n3075 = n473 & ~n3074 ;
  assign n3076 = n561 & n3075 ;
  assign n3077 = ( ~n51 & n1009 ) | ( ~n51 & n2346 ) | ( n1009 & n2346 ) ;
  assign n3078 = n1233 | n2538 ;
  assign n3079 = n1907 | n3078 ;
  assign n3080 = n1029 ^ n168 ^ 1'b0 ;
  assign n3081 = ~n502 & n1918 ;
  assign n3082 = n369 ^ n154 ^ n126 ;
  assign n3083 = n2676 ^ n1969 ^ 1'b0 ;
  assign n3084 = n732 & ~n3083 ;
  assign n3085 = ( n2443 & n3082 ) | ( n2443 & ~n3084 ) | ( n3082 & ~n3084 ) ;
  assign n3086 = n1355 & ~n3085 ;
  assign n3087 = n3081 & n3086 ;
  assign n3088 = n962 ^ n801 ^ n278 ;
  assign n3089 = n2022 & n3088 ;
  assign n3091 = n2499 ^ n1455 ^ 1'b0 ;
  assign n3092 = n2237 | n3091 ;
  assign n3093 = n203 & ~n1000 ;
  assign n3094 = ~n3092 & n3093 ;
  assign n3090 = ( n1613 & n1977 ) | ( n1613 & n2440 ) | ( n1977 & n2440 ) ;
  assign n3095 = n3094 ^ n3090 ^ 1'b0 ;
  assign n3096 = n166 & ~n3095 ;
  assign n3097 = ~x3 & n1476 ;
  assign n3098 = n1432 ^ n1089 ^ n102 ;
  assign n3099 = n1097 ^ x7 ^ 1'b0 ;
  assign n3100 = n130 & n3099 ;
  assign n3101 = ( n1073 & n3098 ) | ( n1073 & n3100 ) | ( n3098 & n3100 ) ;
  assign n3102 = n3101 ^ n1793 ^ 1'b0 ;
  assign n3103 = ~n42 & n1890 ;
  assign n3104 = n3103 ^ n2416 ^ 1'b0 ;
  assign n3105 = n735 & n1225 ;
  assign n3106 = ( ~n1322 & n2500 ) | ( ~n1322 & n3105 ) | ( n2500 & n3105 ) ;
  assign n3107 = n1940 ^ n1653 ^ n82 ;
  assign n3108 = n1322 ^ n1120 ^ 1'b0 ;
  assign n3109 = n3108 ^ n1999 ^ 1'b0 ;
  assign n3110 = n723 ^ n108 ^ 1'b0 ;
  assign n3111 = n1355 & ~n3110 ;
  assign n3112 = n1502 ^ n511 ^ 1'b0 ;
  assign n3113 = n3112 ^ n1204 ^ n30 ;
  assign n3114 = ~n2440 & n2789 ;
  assign n3115 = n57 & ~n1859 ;
  assign n3116 = n3115 ^ n362 ^ 1'b0 ;
  assign n3118 = n41 & ~n1010 ;
  assign n3119 = n3118 ^ n1922 ^ 1'b0 ;
  assign n3117 = n2550 | n2926 ;
  assign n3120 = n3119 ^ n3117 ^ 1'b0 ;
  assign n3121 = n1741 ^ n63 ^ 1'b0 ;
  assign n3122 = n868 | n2547 ;
  assign n3123 = n1922 ^ n526 ^ 1'b0 ;
  assign n3124 = n2220 | n3123 ;
  assign n3126 = ~n1138 & n1650 ;
  assign n3127 = n371 & n3126 ;
  assign n3125 = ( n344 & n1140 ) | ( n344 & n1611 ) | ( n1140 & n1611 ) ;
  assign n3128 = n3127 ^ n3125 ^ 1'b0 ;
  assign n3129 = n53 & ~n548 ;
  assign n3130 = n3129 ^ n1748 ^ 1'b0 ;
  assign n3131 = ( n238 & ~n2583 ) | ( n238 & n3130 ) | ( ~n2583 & n3130 ) ;
  assign n3132 = n149 & n209 ;
  assign n3133 = n3132 ^ n45 ^ 1'b0 ;
  assign n3134 = ~n3131 & n3133 ;
  assign n3135 = ( n652 & n867 ) | ( n652 & ~n2508 ) | ( n867 & ~n2508 ) ;
  assign n3136 = n1209 & n1213 ;
  assign n3137 = n3135 & n3136 ;
  assign n3138 = n3134 | n3137 ;
  assign n3139 = n478 | n704 ;
  assign n3140 = n1153 | n3139 ;
  assign n3141 = n3140 ^ n2403 ^ 1'b0 ;
  assign n3143 = n687 & n1977 ;
  assign n3144 = n132 & n3143 ;
  assign n3142 = n1912 ^ n680 ^ 1'b0 ;
  assign n3145 = n3144 ^ n3142 ^ n2477 ;
  assign n3146 = n3145 ^ n890 ^ 1'b0 ;
  assign n3148 = n1226 ^ n194 ^ 1'b0 ;
  assign n3147 = n186 & n1431 ;
  assign n3149 = n3148 ^ n3147 ^ 1'b0 ;
  assign n3150 = n3149 ^ n2110 ^ 1'b0 ;
  assign n3151 = n3146 & ~n3150 ;
  assign n3152 = n3151 ^ n515 ^ 1'b0 ;
  assign n3153 = n1145 & ~n3152 ;
  assign n3154 = ~n55 & n437 ;
  assign n3155 = ~n376 & n1079 ;
  assign n3156 = ~n1073 & n2524 ;
  assign n3157 = ~n772 & n2350 ;
  assign n3158 = ~n929 & n3157 ;
  assign n3159 = n79 & ~n2886 ;
  assign n3160 = n698 ^ n498 ^ 1'b0 ;
  assign n3161 = n813 & n3160 ;
  assign n3162 = ~n2906 & n3161 ;
  assign n3163 = n1397 | n3162 ;
  assign n3165 = ~n1148 & n1472 ;
  assign n3166 = n3165 ^ n1386 ^ 1'b0 ;
  assign n3164 = n366 & n1461 ;
  assign n3167 = n3166 ^ n3164 ^ 1'b0 ;
  assign n3172 = ~n220 & n1773 ;
  assign n3173 = n1944 & n3172 ;
  assign n3169 = n101 & n1431 ;
  assign n3170 = ~n108 & n3169 ;
  assign n3168 = ( ~n435 & n1245 ) | ( ~n435 & n1279 ) | ( n1245 & n1279 ) ;
  assign n3171 = n3170 ^ n3168 ^ 1'b0 ;
  assign n3174 = n3173 ^ n3171 ^ 1'b0 ;
  assign n3175 = ( n406 & n656 ) | ( n406 & n1000 ) | ( n656 & n1000 ) ;
  assign n3176 = n3175 ^ n2257 ^ n1893 ;
  assign n3177 = n1344 ^ n1281 ^ n711 ;
  assign n3178 = n469 & ~n3177 ;
  assign n3179 = n3178 ^ n2961 ^ 1'b0 ;
  assign n3180 = n809 ^ n650 ^ n97 ;
  assign n3181 = ~n1006 & n3180 ;
  assign n3182 = n3181 ^ n1260 ^ 1'b0 ;
  assign n3183 = ~n177 & n3182 ;
  assign n3184 = n2162 ^ n1009 ^ 1'b0 ;
  assign n3185 = ( n1746 & n2355 ) | ( n1746 & ~n3184 ) | ( n2355 & ~n3184 ) ;
  assign n3186 = n665 ^ n411 ^ 1'b0 ;
  assign n3187 = n2665 & n3186 ;
  assign n3188 = n55 | n1970 ;
  assign n3189 = n3188 ^ n3184 ^ n2081 ;
  assign n3190 = ( n105 & ~n3187 ) | ( n105 & n3189 ) | ( ~n3187 & n3189 ) ;
  assign n3191 = n3190 ^ n1677 ^ n1360 ;
  assign n3192 = n808 ^ n156 ^ 1'b0 ;
  assign n3193 = n3192 ^ n2592 ^ 1'b0 ;
  assign n3194 = ~n2635 & n3193 ;
  assign n3195 = n3194 ^ n1950 ^ 1'b0 ;
  assign n3196 = n3195 ^ n1629 ^ 1'b0 ;
  assign n3197 = ~n882 & n1088 ;
  assign n3198 = ~n1405 & n3197 ;
  assign n3201 = n428 ^ n293 ^ 1'b0 ;
  assign n3199 = n2054 ^ n1280 ^ n846 ;
  assign n3200 = ~n396 & n3199 ;
  assign n3202 = n3201 ^ n3200 ^ 1'b0 ;
  assign n3203 = n3198 | n3202 ;
  assign n3204 = n3203 ^ n1052 ^ 1'b0 ;
  assign n3205 = n2229 & ~n3204 ;
  assign n3206 = n767 & ~n2303 ;
  assign n3207 = n3206 ^ n36 ^ 1'b0 ;
  assign n3208 = ~n287 & n3207 ;
  assign n3209 = n3208 ^ n2140 ^ 1'b0 ;
  assign n3210 = n366 & n3025 ;
  assign n3211 = ~n3209 & n3210 ;
  assign n3212 = n861 | n2203 ;
  assign n3213 = ~n2145 & n3212 ;
  assign n3214 = n3211 & n3213 ;
  assign n3215 = n1286 | n1502 ;
  assign n3216 = n437 & ~n3215 ;
  assign n3217 = n57 & ~n644 ;
  assign n3220 = n80 & n501 ;
  assign n3221 = n3220 ^ x10 ^ 1'b0 ;
  assign n3218 = n597 | n794 ;
  assign n3219 = n259 & ~n3218 ;
  assign n3222 = n3221 ^ n3219 ^ 1'b0 ;
  assign n3223 = ~n3217 & n3222 ;
  assign n3224 = ( n2902 & n3216 ) | ( n2902 & n3223 ) | ( n3216 & n3223 ) ;
  assign n3225 = n1542 ^ n440 ^ n176 ;
  assign n3226 = n889 & n1853 ;
  assign n3227 = n3225 & n3226 ;
  assign n3232 = n1956 ^ n1258 ^ 1'b0 ;
  assign n3228 = ~n45 & n875 ;
  assign n3229 = n871 & n3228 ;
  assign n3230 = n3229 ^ n1265 ^ 1'b0 ;
  assign n3231 = n1810 & n3230 ;
  assign n3233 = n3232 ^ n3231 ^ 1'b0 ;
  assign n3234 = n3227 | n3233 ;
  assign n3235 = n450 & n3234 ;
  assign n3236 = n41 & n700 ;
  assign n3237 = n2130 ^ n769 ^ 1'b0 ;
  assign n3238 = n598 | n833 ;
  assign n3239 = n3238 ^ n35 ^ 1'b0 ;
  assign n3240 = n2337 | n3239 ;
  assign n3241 = n3240 ^ n1771 ^ n84 ;
  assign n3242 = n3168 | n3241 ;
  assign n3243 = n1105 & n2374 ;
  assign n3244 = n1599 & ~n2696 ;
  assign n3245 = n3244 ^ n1051 ^ n953 ;
  assign n3246 = n3245 ^ n2059 ^ 1'b0 ;
  assign n3247 = n1272 & n2505 ;
  assign n3248 = n3247 ^ n1561 ^ 1'b0 ;
  assign n3249 = n1798 | n2161 ;
  assign n3250 = n3249 ^ n102 ^ 1'b0 ;
  assign n3251 = ~n1715 & n1717 ;
  assign n3252 = ~n3250 & n3251 ;
  assign n3253 = n1312 ^ n15 ^ 1'b0 ;
  assign n3254 = ~n139 & n3253 ;
  assign n3255 = ( n289 & n303 ) | ( n289 & ~n777 ) | ( n303 & ~n777 ) ;
  assign n3256 = n2776 ^ n2538 ^ n1255 ;
  assign n3257 = ~n3255 & n3256 ;
  assign n3258 = ~n2664 & n3257 ;
  assign n3259 = n3258 ^ n727 ^ 1'b0 ;
  assign n3264 = n1015 ^ n326 ^ 1'b0 ;
  assign n3260 = ~n398 & n2425 ;
  assign n3261 = ( n448 & n1594 ) | ( n448 & n3260 ) | ( n1594 & n3260 ) ;
  assign n3262 = n3261 ^ n762 ^ 1'b0 ;
  assign n3263 = ~n3229 & n3262 ;
  assign n3265 = n3264 ^ n3263 ^ 1'b0 ;
  assign n3266 = ~n1583 & n3265 ;
  assign n3267 = n661 ^ n590 ^ 1'b0 ;
  assign n3268 = n3266 & n3267 ;
  assign n3269 = n378 ^ n280 ^ 1'b0 ;
  assign n3270 = ~n494 & n3269 ;
  assign n3271 = ~n132 & n1605 ;
  assign n3272 = ~n859 & n1564 ;
  assign n3273 = n2337 & n3272 ;
  assign n3274 = ( n664 & ~n3271 ) | ( n664 & n3273 ) | ( ~n3271 & n3273 ) ;
  assign n3275 = n3274 ^ n1957 ^ 1'b0 ;
  assign n3276 = n366 ^ n194 ^ n36 ;
  assign n3277 = n1084 ^ n973 ^ n426 ;
  assign n3278 = ~n2846 & n3277 ;
  assign n3279 = n3278 ^ n1571 ^ 1'b0 ;
  assign n3280 = n976 ^ n279 ^ 1'b0 ;
  assign n3281 = n1078 | n3280 ;
  assign n3282 = n3281 ^ n1243 ^ 1'b0 ;
  assign n3283 = n220 | n2181 ;
  assign n3284 = n3283 ^ n250 ^ 1'b0 ;
  assign n3285 = n2940 ^ n1139 ^ 1'b0 ;
  assign n3286 = n1697 & ~n3285 ;
  assign n3287 = ~n763 & n1072 ;
  assign n3288 = n3287 ^ n2811 ^ 1'b0 ;
  assign n3289 = ~n1568 & n2702 ;
  assign n3290 = ~n3288 & n3289 ;
  assign n3291 = ~n704 & n3025 ;
  assign n3292 = n3290 & n3291 ;
  assign n3293 = ~n126 & n1532 ;
  assign n3294 = n1089 & n1115 ;
  assign n3295 = n3294 ^ n2074 ^ n1405 ;
  assign n3296 = n2034 ^ n1085 ^ 1'b0 ;
  assign n3297 = n3295 | n3296 ;
  assign n3298 = n3293 & ~n3297 ;
  assign n3299 = n543 ^ n36 ^ 1'b0 ;
  assign n3300 = n2427 ^ n185 ^ 1'b0 ;
  assign n3301 = ~n1311 & n3300 ;
  assign n3302 = n1272 & ~n3301 ;
  assign n3303 = n3302 ^ n2356 ^ 1'b0 ;
  assign n3304 = n3299 | n3303 ;
  assign n3306 = n1611 & ~n2964 ;
  assign n3307 = n3306 ^ n2960 ^ n1817 ;
  assign n3308 = n3307 ^ n3293 ^ 1'b0 ;
  assign n3305 = n1289 ^ n714 ^ 1'b0 ;
  assign n3309 = n3308 ^ n3305 ^ n676 ;
  assign n3310 = n1013 ^ n326 ^ 1'b0 ;
  assign n3311 = ~n515 & n1595 ;
  assign n3312 = n3310 & n3311 ;
  assign n3313 = n1418 ^ n1260 ^ 1'b0 ;
  assign n3314 = n3312 & ~n3313 ;
  assign n3316 = n2960 ^ n864 ^ 1'b0 ;
  assign n3317 = n2694 & n3316 ;
  assign n3315 = ~n941 & n1861 ;
  assign n3318 = n3317 ^ n3315 ^ 1'b0 ;
  assign n3319 = n2017 ^ n1474 ^ 1'b0 ;
  assign n3320 = n3319 ^ n1200 ^ 1'b0 ;
  assign n3321 = ~n3318 & n3320 ;
  assign n3326 = ( n889 & ~n1178 ) | ( n889 & n1418 ) | ( ~n1178 & n1418 ) ;
  assign n3322 = n1110 & ~n1640 ;
  assign n3323 = ~n183 & n3322 ;
  assign n3324 = ~n2098 & n3323 ;
  assign n3325 = n855 & ~n3324 ;
  assign n3327 = n3326 ^ n3325 ^ 1'b0 ;
  assign n3328 = n1775 ^ n1097 ^ 1'b0 ;
  assign n3329 = n23 | n3328 ;
  assign n3330 = n3329 ^ n2049 ^ 1'b0 ;
  assign n3331 = ~n1927 & n3330 ;
  assign n3332 = n3331 ^ n2181 ^ 1'b0 ;
  assign n3333 = n710 | n2729 ;
  assign n3334 = n201 & ~n2120 ;
  assign n3335 = n621 | n1629 ;
  assign n3336 = n3334 & ~n3335 ;
  assign n3337 = n1912 ^ n1656 ^ 1'b0 ;
  assign n3338 = n1832 & ~n3337 ;
  assign n3339 = n3338 ^ n467 ^ 1'b0 ;
  assign n3340 = n3085 ^ n1959 ^ 1'b0 ;
  assign n3341 = n3339 | n3340 ;
  assign n3342 = n3176 ^ n1926 ^ 1'b0 ;
  assign n3343 = n1894 ^ n1439 ^ n349 ;
  assign n3344 = n3343 ^ n2763 ^ 1'b0 ;
  assign n3345 = n2826 & ~n3344 ;
  assign n3346 = n3345 ^ n3173 ^ 1'b0 ;
  assign n3347 = n1483 ^ n195 ^ 1'b0 ;
  assign n3348 = ~n1040 & n3347 ;
  assign n3349 = n532 & ~n1314 ;
  assign n3350 = ~n3348 & n3349 ;
  assign n3351 = n3335 ^ n1206 ^ n331 ;
  assign n3352 = n3351 ^ n267 ^ 1'b0 ;
  assign n3353 = n589 & n3352 ;
  assign n3354 = n3353 ^ n2939 ^ n2381 ;
  assign n3355 = n2262 ^ n590 ^ 1'b0 ;
  assign n3356 = n3253 ^ n1915 ^ 1'b0 ;
  assign n3357 = n929 & ~n3356 ;
  assign n3358 = n3357 ^ n2989 ^ 1'b0 ;
  assign n3360 = n280 ^ n118 ^ 1'b0 ;
  assign n3361 = n38 & n3360 ;
  assign n3359 = ( n611 & ~n1180 ) | ( n611 & n1357 ) | ( ~n1180 & n1357 ) ;
  assign n3362 = n3361 ^ n3359 ^ n960 ;
  assign n3363 = n1875 & ~n3362 ;
  assign n3364 = n1143 ^ n772 ^ 1'b0 ;
  assign n3365 = ( n1223 & ~n1647 ) | ( n1223 & n3364 ) | ( ~n1647 & n3364 ) ;
  assign n3366 = n3175 & n3240 ;
  assign n3367 = n3366 ^ n294 ^ 1'b0 ;
  assign n3368 = ( ~n678 & n2373 ) | ( ~n678 & n3367 ) | ( n2373 & n3367 ) ;
  assign n3369 = n1579 ^ n381 ^ 1'b0 ;
  assign n3370 = n2020 & n3369 ;
  assign n3371 = n654 ^ n139 ^ 1'b0 ;
  assign n3372 = ~n2913 & n3371 ;
  assign n3373 = n1444 & ~n3372 ;
  assign n3374 = n1465 | n2182 ;
  assign n3375 = n3374 ^ n822 ^ 1'b0 ;
  assign n3376 = ( ~n1693 & n3373 ) | ( ~n1693 & n3375 ) | ( n3373 & n3375 ) ;
  assign n3377 = n1461 & ~n2147 ;
  assign n3378 = ~n93 & n1666 ;
  assign n3379 = n3378 ^ n620 ^ 1'b0 ;
  assign n3380 = n3064 & n3379 ;
  assign n3381 = ~n590 & n3380 ;
  assign n3382 = n1039 & ~n3381 ;
  assign n3383 = ( n563 & n1922 ) | ( n563 & ~n2283 ) | ( n1922 & ~n2283 ) ;
  assign n3384 = n1610 & ~n3383 ;
  assign n3385 = n44 & ~n1172 ;
  assign n3386 = n1547 ^ n368 ^ 1'b0 ;
  assign n3387 = n2668 ^ n1218 ^ 1'b0 ;
  assign n3388 = n2555 & n3330 ;
  assign n3389 = n3387 & n3388 ;
  assign n3391 = n201 & n1995 ;
  assign n3392 = ~n887 & n3391 ;
  assign n3390 = ~n139 & n2332 ;
  assign n3393 = n3392 ^ n3390 ^ 1'b0 ;
  assign n3394 = n2758 | n3393 ;
  assign n3395 = n2596 & ~n3394 ;
  assign n3396 = n827 & n994 ;
  assign n3397 = n78 & n3396 ;
  assign n3398 = n2094 | n3397 ;
  assign n3399 = n1149 & ~n3294 ;
  assign n3400 = n3362 ^ n670 ^ 1'b0 ;
  assign n3401 = ~n3399 & n3400 ;
  assign n3402 = n3401 ^ n3101 ^ n400 ;
  assign n3403 = n63 & ~n2655 ;
  assign n3404 = ~n3402 & n3403 ;
  assign n3405 = n234 & ~n3404 ;
  assign n3406 = ~n3398 & n3405 ;
  assign n3407 = n1408 ^ n1095 ^ n63 ;
  assign n3408 = n2419 ^ n910 ^ n878 ;
  assign n3409 = n3408 ^ n1153 ^ n1124 ;
  assign n3410 = ( ~n3299 & n3407 ) | ( ~n3299 & n3409 ) | ( n3407 & n3409 ) ;
  assign n3411 = n2264 ^ n545 ^ 1'b0 ;
  assign n3412 = n868 | n3411 ;
  assign n3413 = n1853 ^ n1681 ^ 1'b0 ;
  assign n3414 = n1641 & n3413 ;
  assign n3415 = n1255 | n3414 ;
  assign n3416 = n3415 ^ n607 ^ 1'b0 ;
  assign n3417 = n2379 & n3057 ;
  assign n3418 = n3417 ^ n2732 ^ 1'b0 ;
  assign n3419 = ~n20 & n1175 ;
  assign n3420 = n3419 ^ n383 ^ 1'b0 ;
  assign n3421 = ( n544 & n1201 ) | ( n544 & ~n3420 ) | ( n1201 & ~n3420 ) ;
  assign n3422 = ( n26 & n185 ) | ( n26 & ~n1553 ) | ( n185 & ~n1553 ) ;
  assign n3423 = n1945 | n3422 ;
  assign n3424 = n1344 & n2470 ;
  assign n3425 = n3424 ^ n1091 ^ 1'b0 ;
  assign n3430 = ( n1307 & n1353 ) | ( n1307 & ~n1762 ) | ( n1353 & ~n1762 ) ;
  assign n3431 = n3430 ^ n1521 ^ 1'b0 ;
  assign n3432 = n589 & n3431 ;
  assign n3428 = n2176 ^ n1387 ^ 1'b0 ;
  assign n3426 = n866 & ~n1668 ;
  assign n3427 = n563 & ~n3426 ;
  assign n3429 = n3428 ^ n3427 ^ 1'b0 ;
  assign n3433 = n3432 ^ n3429 ^ n1816 ;
  assign n3434 = n2156 ^ n306 ^ 1'b0 ;
  assign n3435 = n156 | n3434 ;
  assign n3436 = n729 & n3371 ;
  assign n3437 = n217 & n3436 ;
  assign n3438 = n1395 | n3437 ;
  assign n3439 = n3438 ^ n1682 ^ 1'b0 ;
  assign n3440 = n1490 & n1883 ;
  assign n3441 = ~n2601 & n3440 ;
  assign n3442 = n3439 & n3441 ;
  assign n3443 = ( n966 & n3224 ) | ( n966 & ~n3442 ) | ( n3224 & ~n3442 ) ;
  assign n3447 = n739 ^ n467 ^ 1'b0 ;
  assign n3448 = n3447 ^ n2164 ^ 1'b0 ;
  assign n3449 = n383 | n3448 ;
  assign n3444 = ~n597 & n1212 ;
  assign n3445 = n260 & n3444 ;
  assign n3446 = n3445 ^ n1116 ^ 1'b0 ;
  assign n3450 = n3449 ^ n3446 ^ 1'b0 ;
  assign n3451 = n2418 | n3282 ;
  assign n3452 = n3451 ^ n2665 ^ 1'b0 ;
  assign n3453 = n1234 & ~n2432 ;
  assign n3454 = n3453 ^ n511 ^ 1'b0 ;
  assign n3455 = n1032 ^ n1017 ^ 1'b0 ;
  assign n3457 = n1054 ^ n36 ^ 1'b0 ;
  assign n3458 = ~n1185 & n3457 ;
  assign n3459 = n3458 ^ n1340 ^ 1'b0 ;
  assign n3456 = n577 & n1402 ;
  assign n3460 = n3459 ^ n3456 ^ n1997 ;
  assign n3461 = n949 & n1099 ;
  assign n3462 = n3027 | n3461 ;
  assign n3463 = n3462 ^ n954 ^ 1'b0 ;
  assign n3464 = n3463 ^ n834 ^ 1'b0 ;
  assign n3465 = n3273 ^ n2534 ^ 1'b0 ;
  assign n3466 = n3465 ^ n324 ^ 1'b0 ;
  assign n3467 = n37 & n3466 ;
  assign n3468 = n13 & ~n636 ;
  assign n3469 = n3468 ^ n334 ^ 1'b0 ;
  assign n3470 = n702 | n3469 ;
  assign n3471 = n2710 | n3470 ;
  assign n3472 = n1368 ^ n435 ^ 1'b0 ;
  assign n3473 = n3471 | n3472 ;
  assign n3476 = ~n435 & n823 ;
  assign n3477 = n3476 ^ n639 ^ 1'b0 ;
  assign n3474 = n1118 ^ n37 ^ 1'b0 ;
  assign n3475 = n1157 | n3474 ;
  assign n3478 = n3477 ^ n3475 ^ 1'b0 ;
  assign n3479 = n23 | n38 ;
  assign n3480 = n2334 & ~n3479 ;
  assign n3481 = n3480 ^ n1537 ^ 1'b0 ;
  assign n3482 = n2078 & n3481 ;
  assign n3483 = n1770 & n1927 ;
  assign n3484 = n1235 & ~n1953 ;
  assign n3487 = ~n75 & n784 ;
  assign n3488 = ~n648 & n3487 ;
  assign n3485 = n765 ^ x10 ^ 1'b0 ;
  assign n3486 = n3221 & ~n3485 ;
  assign n3489 = n3488 ^ n3486 ^ n980 ;
  assign n3490 = n2870 & ~n3446 ;
  assign n3491 = n25 & n3490 ;
  assign n3492 = x10 | n3491 ;
  assign n3493 = n3489 & ~n3492 ;
  assign n3495 = ~n427 & n853 ;
  assign n3494 = n25 | n859 ;
  assign n3496 = n3495 ^ n3494 ^ 1'b0 ;
  assign n3497 = n3496 ^ n557 ^ 1'b0 ;
  assign n3498 = n597 | n3497 ;
  assign n3499 = n1591 ^ n922 ^ 1'b0 ;
  assign n3500 = n797 | n3499 ;
  assign n3501 = n3500 ^ n883 ^ 1'b0 ;
  assign n3502 = n379 | n3501 ;
  assign n3503 = n3502 ^ n45 ^ 1'b0 ;
  assign n3504 = n1665 ^ n782 ^ 1'b0 ;
  assign n3505 = n2373 & ~n3504 ;
  assign n3506 = ( ~n105 & n811 ) | ( ~n105 & n1038 ) | ( n811 & n1038 ) ;
  assign n3507 = n2971 ^ n2245 ^ 1'b0 ;
  assign n3508 = ~n214 & n3507 ;
  assign n3509 = n592 & ~n1871 ;
  assign n3510 = n3509 ^ n1255 ^ 1'b0 ;
  assign n3511 = n846 & n3510 ;
  assign n3512 = ~n3508 & n3511 ;
  assign n3513 = n360 | n3512 ;
  assign n3514 = n586 | n3513 ;
  assign n3515 = n3301 ^ n1744 ^ 1'b0 ;
  assign n3516 = n2036 ^ n611 ^ 1'b0 ;
  assign n3517 = n2422 | n3516 ;
  assign n3518 = n710 & ~n2811 ;
  assign n3519 = n711 & ~n1804 ;
  assign n3520 = ~n631 & n1907 ;
  assign n3521 = n218 & n3520 ;
  assign n3522 = n3521 ^ n1089 ^ 1'b0 ;
  assign n3523 = ( ~n137 & n147 ) | ( ~n137 & n3522 ) | ( n147 & n3522 ) ;
  assign n3524 = n1145 ^ n965 ^ 1'b0 ;
  assign n3525 = ~n694 & n1315 ;
  assign n3526 = ~n3524 & n3525 ;
  assign n3527 = n3526 ^ n971 ^ 1'b0 ;
  assign n3528 = n3523 | n3527 ;
  assign n3529 = n2206 & ~n3528 ;
  assign n3530 = n3529 ^ n1360 ^ 1'b0 ;
  assign n3536 = n2425 & ~n2971 ;
  assign n3537 = n3536 ^ n1523 ^ 1'b0 ;
  assign n3538 = n3537 ^ n572 ^ 1'b0 ;
  assign n3539 = ~n2381 & n3538 ;
  assign n3531 = n1339 ^ n1302 ^ n529 ;
  assign n3532 = n1395 & n1822 ;
  assign n3533 = n1348 ^ n1084 ^ n645 ;
  assign n3534 = ( ~n3531 & n3532 ) | ( ~n3531 & n3533 ) | ( n3532 & n3533 ) ;
  assign n3535 = n1862 & ~n3534 ;
  assign n3540 = n3539 ^ n3535 ^ 1'b0 ;
  assign n3543 = n51 | n3027 ;
  assign n3541 = n406 ^ n115 ^ 1'b0 ;
  assign n3542 = n3541 ^ n22 ^ 1'b0 ;
  assign n3544 = n3543 ^ n3542 ^ 1'b0 ;
  assign n3545 = ~n211 & n3544 ;
  assign n3546 = ~n1017 & n3545 ;
  assign n3547 = n942 ^ n394 ^ 1'b0 ;
  assign n3548 = n940 & ~n3547 ;
  assign n3549 = ~n322 & n3231 ;
  assign n3550 = ~n3548 & n3549 ;
  assign n3551 = n572 | n1581 ;
  assign n3552 = n1521 ^ n764 ^ x10 ;
  assign n3553 = n3552 ^ n2471 ^ 1'b0 ;
  assign n3554 = n95 | n3553 ;
  assign n3555 = n3551 & n3554 ;
  assign n3557 = n3253 ^ n2510 ^ n1532 ;
  assign n3556 = n1332 & ~n2640 ;
  assign n3558 = n3557 ^ n3556 ^ 1'b0 ;
  assign n3572 = n462 & n3361 ;
  assign n3573 = ~n1406 & n3572 ;
  assign n3561 = n1582 ^ n79 ^ 1'b0 ;
  assign n3562 = n1365 | n3561 ;
  assign n3563 = n3562 ^ n154 ^ 1'b0 ;
  assign n3560 = n652 & ~n3044 ;
  assign n3564 = n3563 ^ n3560 ^ 1'b0 ;
  assign n3565 = n2002 & ~n3564 ;
  assign n3559 = n788 & ~n2159 ;
  assign n3566 = n3565 ^ n3559 ^ 1'b0 ;
  assign n3568 = n1332 ^ n437 ^ 1'b0 ;
  assign n3567 = n702 & ~n1114 ;
  assign n3569 = n3568 ^ n3567 ^ 1'b0 ;
  assign n3570 = n447 & ~n3569 ;
  assign n3571 = ~n3566 & n3570 ;
  assign n3574 = n3573 ^ n3571 ^ n3040 ;
  assign n3577 = n891 & ~n1848 ;
  assign n3575 = n3364 ^ n3144 ^ n279 ;
  assign n3576 = n899 & ~n3575 ;
  assign n3578 = n3577 ^ n3576 ^ 1'b0 ;
  assign n3580 = ( n636 & n674 ) | ( n636 & n2094 ) | ( n674 & n2094 ) ;
  assign n3579 = ( n726 & n1340 ) | ( n726 & ~n2397 ) | ( n1340 & ~n2397 ) ;
  assign n3581 = n3580 ^ n3579 ^ 1'b0 ;
  assign n3582 = n895 ^ n131 ^ 1'b0 ;
  assign n3583 = n3232 | n3582 ;
  assign n3584 = n3583 ^ n1456 ^ 1'b0 ;
  assign n3585 = ~n2051 & n3584 ;
  assign n3586 = n2756 ^ n1185 ^ 1'b0 ;
  assign n3587 = ~n1164 & n3586 ;
  assign n3588 = n2445 & n3587 ;
  assign n3589 = n2791 ^ n2201 ^ 1'b0 ;
  assign n3590 = n791 & n3589 ;
  assign n3591 = ( n130 & n322 ) | ( n130 & ~n328 ) | ( n322 & ~n328 ) ;
  assign n3592 = n3591 ^ n2528 ^ n2461 ;
  assign n3593 = n55 & ~n544 ;
  assign n3594 = n836 ^ n725 ^ 1'b0 ;
  assign n3595 = ~n3593 & n3594 ;
  assign n3596 = n3592 & n3595 ;
  assign n3597 = ~n3590 & n3596 ;
  assign n3598 = ~n569 & n2483 ;
  assign n3599 = ~n37 & n3598 ;
  assign n3600 = n2837 ^ n1305 ^ 1'b0 ;
  assign n3601 = n358 & n424 ;
  assign n3602 = ~n572 & n3601 ;
  assign n3603 = n3602 ^ n2499 ^ 1'b0 ;
  assign n3604 = n392 ^ x0 ^ 1'b0 ;
  assign n3605 = n3604 ^ n369 ^ 1'b0 ;
  assign n3606 = n420 & n3605 ;
  assign n3607 = ( n2056 & n3603 ) | ( n2056 & n3606 ) | ( n3603 & n3606 ) ;
  assign n3608 = ( n998 & n2089 ) | ( n998 & n3144 ) | ( n2089 & n3144 ) ;
  assign n3609 = n661 & n839 ;
  assign n3610 = ~n3127 & n3609 ;
  assign n3617 = n373 | n902 ;
  assign n3618 = n405 | n3617 ;
  assign n3611 = n322 | n759 ;
  assign n3612 = n583 | n3611 ;
  assign n3614 = n1674 & n2128 ;
  assign n3613 = n492 | n2609 ;
  assign n3615 = n3614 ^ n3613 ^ 1'b0 ;
  assign n3616 = n3612 & n3615 ;
  assign n3619 = n3618 ^ n3616 ^ 1'b0 ;
  assign n3620 = n3619 ^ n33 ^ 1'b0 ;
  assign n3621 = n1849 ^ n344 ^ 1'b0 ;
  assign n3622 = n203 & ~n3621 ;
  assign n3623 = n732 & ~n2044 ;
  assign n3624 = ~n2791 & n3623 ;
  assign n3625 = ( n1874 & ~n2173 ) | ( n1874 & n2231 ) | ( ~n2173 & n2231 ) ;
  assign n3626 = ~n3624 & n3625 ;
  assign n3627 = n467 & n1336 ;
  assign n3628 = n3627 ^ n3041 ^ 1'b0 ;
  assign n3629 = n448 & n1713 ;
  assign n3630 = ~n3628 & n3629 ;
  assign n3631 = n390 ^ n249 ^ 1'b0 ;
  assign n3632 = n3299 | n3631 ;
  assign n3633 = n3632 ^ n1269 ^ 1'b0 ;
  assign n3634 = n2591 | n3633 ;
  assign n3635 = n431 & ~n2535 ;
  assign n3636 = ( n674 & ~n1365 ) | ( n674 & n3375 ) | ( ~n1365 & n3375 ) ;
  assign n3637 = n2837 ^ n1563 ^ 1'b0 ;
  assign n3638 = n1791 ^ n974 ^ n886 ;
  assign n3639 = n3638 ^ n2570 ^ 1'b0 ;
  assign n3640 = n1389 | n3046 ;
  assign n3641 = n2732 & ~n3293 ;
  assign n3642 = n1468 ^ n1207 ^ 1'b0 ;
  assign n3643 = n1126 | n3642 ;
  assign n3644 = n3336 | n3643 ;
  assign n3654 = ~n132 & n1231 ;
  assign n3650 = n1619 ^ n977 ^ n686 ;
  assign n3651 = n3650 ^ n626 ^ 1'b0 ;
  assign n3647 = n30 & n1262 ;
  assign n3645 = n814 | n1048 ;
  assign n3646 = ~n478 & n3645 ;
  assign n3648 = n3647 ^ n3646 ^ 1'b0 ;
  assign n3649 = n550 & n3648 ;
  assign n3652 = n3651 ^ n3649 ^ 1'b0 ;
  assign n3653 = ~n1796 & n3652 ;
  assign n3655 = n3654 ^ n3653 ^ 1'b0 ;
  assign n3656 = n2761 ^ n32 ^ 1'b0 ;
  assign n3657 = n1300 & ~n2023 ;
  assign n3658 = n3657 ^ n526 ^ 1'b0 ;
  assign n3659 = ( ~n561 & n935 ) | ( ~n561 & n3658 ) | ( n935 & n3658 ) ;
  assign n3660 = ~n1032 & n3659 ;
  assign n3661 = n42 & ~n1846 ;
  assign n3662 = ( n2289 & ~n3660 ) | ( n2289 & n3661 ) | ( ~n3660 & n3661 ) ;
  assign n3663 = ~n63 & n753 ;
  assign n3664 = n686 ^ n578 ^ 1'b0 ;
  assign n3665 = n702 & ~n3664 ;
  assign n3666 = n3212 & n3665 ;
  assign n3667 = ( n322 & n564 ) | ( n322 & ~n3666 ) | ( n564 & ~n3666 ) ;
  assign n3668 = n2925 & ~n3667 ;
  assign n3669 = n202 & n3668 ;
  assign n3675 = n1041 ^ n1028 ^ 1'b0 ;
  assign n3676 = n3579 | n3675 ;
  assign n3670 = n648 & ~n2044 ;
  assign n3671 = n2102 & n3670 ;
  assign n3672 = n977 | n3671 ;
  assign n3673 = n1324 & ~n3672 ;
  assign n3674 = n3635 & ~n3673 ;
  assign n3677 = n3676 ^ n3674 ^ 1'b0 ;
  assign n3678 = n1589 | n1945 ;
  assign n3679 = n181 | n3678 ;
  assign n3680 = n3190 | n3679 ;
  assign n3681 = n756 ^ n23 ^ 1'b0 ;
  assign n3682 = n2095 ^ n23 ^ 1'b0 ;
  assign n3683 = n3682 ^ n1680 ^ 1'b0 ;
  assign n3684 = n1793 & ~n3683 ;
  assign n3685 = ( n1789 & n3681 ) | ( n1789 & ~n3684 ) | ( n3681 & ~n3684 ) ;
  assign n3687 = n51 | n2320 ;
  assign n3688 = ~n842 & n3687 ;
  assign n3689 = n2839 | n3688 ;
  assign n3690 = n3001 & ~n3689 ;
  assign n3686 = n371 ^ n303 ^ 1'b0 ;
  assign n3691 = n3690 ^ n3686 ^ 1'b0 ;
  assign n3692 = n3685 & ~n3691 ;
  assign n3693 = n2828 ^ n916 ^ 1'b0 ;
  assign n3694 = n3418 ^ n2481 ^ 1'b0 ;
  assign n3695 = n1856 & n2666 ;
  assign n3696 = n2078 & n3695 ;
  assign n3697 = n168 & ~n1157 ;
  assign n3698 = ~n567 & n3697 ;
  assign n3699 = n1828 | n3698 ;
  assign n3700 = n3699 ^ n82 ^ 1'b0 ;
  assign n3701 = n2097 & ~n3700 ;
  assign n3702 = n1642 & n3701 ;
  assign n3703 = ( n234 & ~n1383 ) | ( n234 & n3569 ) | ( ~n1383 & n3569 ) ;
  assign n3704 = n2108 | n3703 ;
  assign n3705 = n3704 ^ n1186 ^ 1'b0 ;
  assign n3706 = n3702 | n3705 ;
  assign n3707 = n313 | n863 ;
  assign n3708 = ~n1339 & n3166 ;
  assign n3709 = n755 ^ n299 ^ 1'b0 ;
  assign n3710 = ( n1582 & n1805 ) | ( n1582 & n3709 ) | ( n1805 & n3709 ) ;
  assign n3711 = ~n3407 & n3710 ;
  assign n3712 = ( n481 & n3708 ) | ( n481 & n3711 ) | ( n3708 & n3711 ) ;
  assign n3713 = x3 | n2054 ;
  assign n3714 = n2216 & ~n3713 ;
  assign n3715 = n1214 & n2849 ;
  assign n3716 = n1454 & n3715 ;
  assign n3717 = ~n2179 & n3716 ;
  assign n3718 = n965 | n3717 ;
  assign n3719 = n3718 ^ n3408 ^ 1'b0 ;
  assign n3720 = n544 ^ x10 ^ 1'b0 ;
  assign n3721 = n234 & n2362 ;
  assign n3722 = ~n3720 & n3721 ;
  assign n3723 = n467 & n3357 ;
  assign n3724 = n177 | n1127 ;
  assign n3725 = n3723 | n3724 ;
  assign n3726 = n1399 ^ n1127 ^ n621 ;
  assign n3727 = ( n371 & n926 ) | ( n371 & n3726 ) | ( n926 & n3726 ) ;
  assign n3728 = n108 & n2273 ;
  assign n3729 = n3728 ^ n491 ^ 1'b0 ;
  assign n3730 = n3195 & n3729 ;
  assign n3731 = n1731 & n3730 ;
  assign n3732 = n1944 ^ n855 ^ 1'b0 ;
  assign n3733 = n1318 ^ n1235 ^ 1'b0 ;
  assign n3734 = n3732 & n3733 ;
  assign n3735 = n415 & ~n672 ;
  assign n3736 = ~n3734 & n3735 ;
  assign n3737 = n596 & n2665 ;
  assign n3738 = ( ~n510 & n1083 ) | ( ~n510 & n3737 ) | ( n1083 & n3737 ) ;
  assign n3739 = n3738 ^ n1192 ^ n40 ;
  assign n3740 = n3739 ^ n1470 ^ 1'b0 ;
  assign n3741 = n3740 ^ n2505 ^ n1063 ;
  assign n3742 = ( n570 & ~n1447 ) | ( n570 & n2689 ) | ( ~n1447 & n2689 ) ;
  assign n3743 = n1368 & n3742 ;
  assign n3744 = n3743 ^ n3187 ^ 1'b0 ;
  assign n3745 = n1179 ^ n803 ^ 1'b0 ;
  assign n3746 = n2844 & ~n3745 ;
  assign n3747 = n3744 & n3746 ;
  assign n3753 = ~n529 & n2068 ;
  assign n3748 = n1178 ^ n666 ^ 1'b0 ;
  assign n3749 = ~n2143 & n3748 ;
  assign n3750 = ~n214 & n2157 ;
  assign n3751 = n1314 | n3750 ;
  assign n3752 = n3749 & ~n3751 ;
  assign n3754 = n3753 ^ n3752 ^ 1'b0 ;
  assign n3758 = n1820 ^ x8 ^ 1'b0 ;
  assign n3759 = n3758 ^ n1921 ^ 1'b0 ;
  assign n3755 = n1979 & ~n2453 ;
  assign n3756 = n117 | n3755 ;
  assign n3757 = n261 | n3756 ;
  assign n3760 = n3759 ^ n3757 ^ 1'b0 ;
  assign n3766 = n1237 ^ n434 ^ 1'b0 ;
  assign n3767 = n2459 | n3766 ;
  assign n3764 = n91 & ~n272 ;
  assign n3765 = n3764 ^ n1943 ^ 1'b0 ;
  assign n3762 = n1493 ^ n533 ^ n211 ;
  assign n3761 = ( n63 & n1052 ) | ( n63 & ~n1552 ) | ( n1052 & ~n1552 ) ;
  assign n3763 = n3762 ^ n3761 ^ 1'b0 ;
  assign n3768 = n3767 ^ n3765 ^ n3763 ;
  assign n3769 = ( n772 & n2281 ) | ( n772 & n3336 ) | ( n2281 & n3336 ) ;
  assign n3770 = n2359 ^ n826 ^ 1'b0 ;
  assign n3771 = n761 & ~n1464 ;
  assign n3772 = n3771 ^ n1456 ^ 1'b0 ;
  assign n3774 = n1004 ^ n795 ^ 1'b0 ;
  assign n3775 = n3774 ^ n1238 ^ 1'b0 ;
  assign n3773 = ~n1081 & n3123 ;
  assign n3776 = n3775 ^ n3773 ^ n2913 ;
  assign n3777 = ( n313 & ~n3772 ) | ( n313 & n3776 ) | ( ~n3772 & n3776 ) ;
  assign n3778 = n3567 ^ n3263 ^ 1'b0 ;
  assign n3779 = n358 & ~n2844 ;
  assign n3780 = ~n1290 & n2261 ;
  assign n3781 = n3779 & n3780 ;
  assign n3782 = n3781 ^ n2379 ^ 1'b0 ;
  assign n3783 = n1411 & n3740 ;
  assign n3784 = ~n3782 & n3783 ;
  assign n3785 = n1444 & ~n2493 ;
  assign n3786 = n1043 & n3785 ;
  assign n3787 = n1200 & n1300 ;
  assign n3788 = n3787 ^ n583 ^ 1'b0 ;
  assign n3789 = n3786 & ~n3788 ;
  assign n3790 = n84 | n2302 ;
  assign n3791 = ( ~n496 & n563 ) | ( ~n496 & n3790 ) | ( n563 & n3790 ) ;
  assign n3792 = n1848 & ~n3791 ;
  assign n3793 = n2638 ^ n1092 ^ 1'b0 ;
  assign n3794 = n2048 ^ n70 ^ 1'b0 ;
  assign n3795 = ~n3793 & n3794 ;
  assign n3796 = n226 ^ n181 ^ 1'b0 ;
  assign n3797 = n2239 | n3796 ;
  assign n3798 = n51 & ~n3797 ;
  assign n3799 = n2306 ^ n879 ^ 1'b0 ;
  assign n3800 = n131 & ~n2060 ;
  assign n3801 = n121 & ~n3044 ;
  assign n3802 = n3800 & ~n3801 ;
  assign n3803 = ( n717 & n3799 ) | ( n717 & ~n3802 ) | ( n3799 & ~n3802 ) ;
  assign n3804 = ( n1175 & ~n1437 ) | ( n1175 & n3803 ) | ( ~n1437 & n3803 ) ;
  assign n3805 = n2137 ^ n96 ^ 1'b0 ;
  assign n3809 = n1184 | n1190 ;
  assign n3810 = n3809 ^ n1175 ^ 1'b0 ;
  assign n3808 = n947 & ~n1638 ;
  assign n3811 = n3810 ^ n3808 ^ 1'b0 ;
  assign n3806 = n448 & n1096 ;
  assign n3807 = n3806 ^ n1025 ^ 1'b0 ;
  assign n3812 = n3811 ^ n3807 ^ 1'b0 ;
  assign n3813 = n1200 & n3628 ;
  assign n3814 = n1121 & n3813 ;
  assign n3815 = x4 & n583 ;
  assign n3816 = n2956 & n3815 ;
  assign n3817 = ( n457 & ~n1988 ) | ( n457 & n2105 ) | ( ~n1988 & n2105 ) ;
  assign n3818 = ( n186 & n1752 ) | ( n186 & n2360 ) | ( n1752 & n2360 ) ;
  assign n3819 = ( n2273 & ~n2595 ) | ( n2273 & n3818 ) | ( ~n2595 & n3818 ) ;
  assign n3820 = n1278 & n3130 ;
  assign n3821 = ~n2514 & n3820 ;
  assign n3822 = n3774 ^ n503 ^ 1'b0 ;
  assign n3823 = n272 | n3822 ;
  assign n3824 = ~n177 & n3823 ;
  assign n3825 = n3824 ^ n1196 ^ 1'b0 ;
  assign n3826 = n1843 & n2077 ;
  assign n3827 = n3825 & n3826 ;
  assign n3828 = n3821 & n3827 ;
  assign n3829 = n1355 & ~n3828 ;
  assign n3830 = ~n962 & n3829 ;
  assign n3831 = n965 & ~n1024 ;
  assign n3832 = ~n3577 & n3831 ;
  assign n3833 = n1176 ^ n922 ^ 1'b0 ;
  assign n3834 = n2872 ^ n1537 ^ 1'b0 ;
  assign n3835 = ~n3833 & n3834 ;
  assign n3836 = n2391 ^ n1474 ^ 1'b0 ;
  assign n3837 = ~n859 & n3836 ;
  assign n3838 = n3837 ^ n3699 ^ n963 ;
  assign n3839 = n598 | n883 ;
  assign n3840 = n3839 ^ n350 ^ 1'b0 ;
  assign n3841 = n3840 ^ n1287 ^ 1'b0 ;
  assign n3842 = n813 & ~n3841 ;
  assign n3843 = n3842 ^ n2270 ^ n838 ;
  assign n3844 = n3843 ^ n2118 ^ 1'b0 ;
  assign n3845 = n3838 & ~n3844 ;
  assign n3846 = n3845 ^ n3081 ^ 1'b0 ;
  assign n3847 = n1281 ^ n1221 ^ n440 ;
  assign n3848 = ( n1182 & n1389 ) | ( n1182 & n1851 ) | ( n1389 & n1851 ) ;
  assign n3849 = x10 & n2416 ;
  assign n3850 = n3849 ^ n3000 ^ 1'b0 ;
  assign n3851 = n951 | n1060 ;
  assign n3852 = ~n44 & n1918 ;
  assign n3853 = ~n318 & n3852 ;
  assign n3854 = n1026 & ~n3853 ;
  assign n3855 = ~n876 & n3854 ;
  assign n3856 = n1047 ^ n691 ^ n580 ;
  assign n3857 = n234 & ~n3856 ;
  assign n3858 = n3857 ^ n593 ^ 1'b0 ;
  assign n3859 = n3858 ^ n842 ^ 1'b0 ;
  assign n3860 = n1684 & n3859 ;
  assign n3861 = n1951 ^ n1922 ^ n532 ;
  assign n3862 = n1365 | n3861 ;
  assign n3863 = n13 | n3862 ;
  assign n3864 = n483 & n3863 ;
  assign n3865 = ~n1049 & n2648 ;
  assign n3866 = n2302 & n3865 ;
  assign n3867 = n569 & ~n1135 ;
  assign n3868 = n635 ^ n445 ^ n369 ;
  assign n3869 = n2810 ^ n1875 ^ 1'b0 ;
  assign n3870 = n3868 & n3869 ;
  assign n3871 = n55 & n3870 ;
  assign n3872 = n2280 ^ n1051 ^ 1'b0 ;
  assign n3873 = n506 & n3872 ;
  assign n3874 = n3873 ^ n1818 ^ 1'b0 ;
  assign n3875 = n3615 ^ n2653 ^ 1'b0 ;
  assign n3876 = n2493 & ~n3875 ;
  assign n3877 = n854 & n3218 ;
  assign n3878 = n1636 ^ n486 ^ 1'b0 ;
  assign n3879 = n352 ^ n228 ^ 1'b0 ;
  assign n3880 = n1592 & ~n3879 ;
  assign n3881 = ~n1679 & n2694 ;
  assign n3882 = n41 & ~n3779 ;
  assign n3883 = n3882 ^ n3080 ^ n78 ;
  assign n3884 = n3582 ^ n2655 ^ 1'b0 ;
  assign n3885 = n3884 ^ n3301 ^ 1'b0 ;
  assign n3886 = x10 & ~n1454 ;
  assign n3887 = n1959 ^ n129 ^ 1'b0 ;
  assign n3888 = n1490 & n3887 ;
  assign n3889 = n2150 & n3888 ;
  assign n3890 = n3889 ^ n1032 ^ 1'b0 ;
  assign n3891 = ( n865 & n3886 ) | ( n865 & n3890 ) | ( n3886 & n3890 ) ;
  assign n3892 = n1849 ^ n96 ^ 1'b0 ;
  assign n3893 = n3892 ^ n289 ^ 1'b0 ;
  assign n3894 = n1330 & n3466 ;
  assign n3896 = n289 & n564 ;
  assign n3895 = n879 | n1221 ;
  assign n3897 = n3896 ^ n3895 ^ 1'b0 ;
  assign n3898 = n3897 ^ n3019 ^ 1'b0 ;
  assign n3899 = n2668 & ~n3658 ;
  assign n3900 = n3899 ^ n3119 ^ 1'b0 ;
  assign n3901 = ~n3898 & n3900 ;
  assign n3902 = ~n2425 & n3128 ;
  assign n3903 = n2434 ^ n863 ^ 1'b0 ;
  assign n3904 = n945 & ~n3903 ;
  assign n3905 = n1550 & ~n3904 ;
  assign n3906 = n317 & n3832 ;
  assign n3907 = n3082 ^ n991 ^ 1'b0 ;
  assign n3908 = ~n769 & n3907 ;
  assign n3909 = n698 ^ n204 ^ 1'b0 ;
  assign n3910 = ~n1265 & n3909 ;
  assign n3911 = ~n958 & n3910 ;
  assign n3912 = x3 & ~n3911 ;
  assign n3913 = ~n1666 & n3912 ;
  assign n3914 = n2971 & n3913 ;
  assign n3915 = n35 & n2305 ;
  assign n3916 = n3915 ^ n3522 ^ 1'b0 ;
  assign n3917 = n503 & n1125 ;
  assign n3918 = n3917 ^ n2601 ^ 1'b0 ;
  assign n3919 = n3918 ^ n1837 ^ n1204 ;
  assign n3920 = n3919 ^ n2211 ^ n2195 ;
  assign n3921 = n2289 & n3897 ;
  assign n3922 = n3921 ^ n54 ^ 1'b0 ;
  assign n3924 = ~n55 & n664 ;
  assign n3925 = n131 & n3924 ;
  assign n3926 = n3671 | n3925 ;
  assign n3927 = n2343 & ~n3046 ;
  assign n3928 = ~n3926 & n3927 ;
  assign n3929 = n3928 ^ n2199 ^ 1'b0 ;
  assign n3923 = ~n874 & n1679 ;
  assign n3930 = n3929 ^ n3923 ^ 1'b0 ;
  assign n3931 = n523 & n918 ;
  assign n3932 = n132 & ~n1056 ;
  assign n3933 = ~n67 & n3932 ;
  assign n3934 = n3933 ^ n3406 ^ 1'b0 ;
  assign n3935 = ~n921 & n2370 ;
  assign n3936 = ~n3156 & n3935 ;
  assign n3937 = n1881 & n2083 ;
  assign n3938 = n3856 & n3937 ;
  assign n3939 = ( n2615 & n3512 ) | ( n2615 & n3938 ) | ( n3512 & n3938 ) ;
  assign n3940 = n3939 ^ n3902 ^ 1'b0 ;
  assign n3941 = n1480 & n3566 ;
  assign n3942 = n1744 ^ n395 ^ 1'b0 ;
  assign n3943 = ~n570 & n3942 ;
  assign n3944 = n875 & n3943 ;
  assign n3945 = n694 & n3944 ;
  assign n3946 = n2640 ^ n864 ^ 1'b0 ;
  assign n3947 = n1737 & n3628 ;
  assign n3948 = n3946 & n3947 ;
  assign n3949 = ~x5 & n2196 ;
  assign n3950 = n3770 ^ n2701 ^ n2068 ;
  assign n3951 = n3216 ^ n1912 ^ 1'b0 ;
  assign n3952 = ~n1126 & n1380 ;
  assign n3953 = n1591 & n3952 ;
  assign n3954 = n944 ^ n691 ^ 1'b0 ;
  assign n3955 = ~n694 & n3954 ;
  assign n3956 = n3614 & n3955 ;
  assign n3957 = n3956 ^ n2190 ^ 1'b0 ;
  assign n3958 = n41 & n690 ;
  assign n3959 = n3198 & n3958 ;
  assign n3960 = n3959 ^ n3308 ^ 1'b0 ;
  assign n3961 = ~n2864 & n3960 ;
  assign n3962 = n63 & ~n230 ;
  assign n3963 = n3229 ^ n3179 ^ 1'b0 ;
  assign n3964 = n3962 & n3963 ;
  assign n3965 = n41 & ~n342 ;
  assign n3966 = n3965 ^ n674 ^ 1'b0 ;
  assign n3967 = n3359 ^ n2440 ^ 1'b0 ;
  assign n3968 = n1525 | n3967 ;
  assign n3969 = ~n3966 & n3968 ;
  assign n3970 = n403 | n946 ;
  assign n3971 = ~n3969 & n3970 ;
  assign n3972 = n778 ^ n536 ^ 1'b0 ;
  assign n3973 = n517 | n3972 ;
  assign n3974 = n1551 ^ n1213 ^ 1'b0 ;
  assign n3975 = ~n3973 & n3974 ;
  assign n3976 = n1718 ^ n383 ^ 1'b0 ;
  assign n3977 = n3976 ^ n3123 ^ n2284 ;
  assign n3978 = n3977 ^ n2312 ^ 1'b0 ;
  assign n3979 = n1003 | n3978 ;
  assign n3980 = n3975 & ~n3979 ;
  assign n3981 = n3980 ^ n3600 ^ 1'b0 ;
  assign n3982 = n3981 ^ n2494 ^ 1'b0 ;
  assign n3983 = n704 & n1380 ;
  assign n3984 = n3983 ^ n180 ^ n113 ;
  assign n3985 = ( n1807 & ~n2844 ) | ( n1807 & n3034 ) | ( ~n2844 & n3034 ) ;
  assign n3986 = n3985 ^ n1210 ^ 1'b0 ;
  assign n3987 = n334 & n3986 ;
  assign n3988 = n709 ^ n132 ^ 1'b0 ;
  assign n3989 = n3988 ^ n684 ^ 1'b0 ;
  assign n3990 = n2330 ^ n2156 ^ 1'b0 ;
  assign n3991 = n3989 & n3990 ;
  assign n3992 = n1520 & ~n3599 ;
  assign n3993 = ~n3991 & n3992 ;
  assign n3994 = n384 | n2086 ;
  assign n3995 = n722 & n3966 ;
  assign n3996 = n3995 ^ n839 ^ 1'b0 ;
  assign n3997 = n3634 & n3996 ;
  assign n3998 = n65 & ~n1010 ;
  assign n3999 = n3998 ^ n2324 ^ 1'b0 ;
  assign n4000 = n1220 & ~n3999 ;
  assign n4001 = n511 | n2377 ;
  assign n4002 = n4001 ^ n2257 ^ 1'b0 ;
  assign n4003 = n980 | n2078 ;
  assign n4004 = n4003 ^ n1251 ^ 1'b0 ;
  assign n4005 = ( n183 & n462 ) | ( n183 & n1069 ) | ( n462 & n1069 ) ;
  assign n4006 = n3993 | n4005 ;
  assign n4007 = n2731 ^ n1145 ^ 1'b0 ;
  assign n4008 = n63 & n4007 ;
  assign n4009 = n4008 ^ n2423 ^ n448 ;
  assign n4010 = n652 & ~n4009 ;
  assign n4011 = ~n3211 & n4010 ;
  assign n4012 = n2828 ^ n1546 ^ n1273 ;
  assign n4013 = n2858 | n4012 ;
  assign n4014 = n1037 | n4013 ;
  assign n4015 = n1365 ^ n1105 ^ 1'b0 ;
  assign n4016 = x2 & ~n4015 ;
  assign n4017 = n4016 ^ n2944 ^ 1'b0 ;
  assign n4018 = n645 | n4017 ;
  assign n4019 = ~n883 & n4018 ;
  assign n4020 = n237 & n4019 ;
  assign n4021 = ~n4014 & n4020 ;
  assign n4022 = n43 | n2181 ;
  assign n4023 = n1518 & ~n4022 ;
  assign n4024 = n4023 ^ n2086 ^ 1'b0 ;
  assign n4025 = n3765 | n3824 ;
  assign n4026 = n826 | n2276 ;
  assign n4027 = n4025 & ~n4026 ;
  assign n4028 = n2368 ^ n1945 ^ 1'b0 ;
  assign n4029 = ~n833 & n1230 ;
  assign n4030 = n2402 & n4029 ;
  assign n4031 = n1638 | n4030 ;
  assign n4032 = n4028 & ~n4031 ;
  assign n4033 = n589 & n644 ;
  assign n4034 = ~n1891 & n4033 ;
  assign n4035 = n984 & ~n3600 ;
  assign n4036 = n4034 & n4035 ;
  assign n4038 = n1770 & n2184 ;
  assign n4037 = n865 | n1951 ;
  assign n4039 = n4038 ^ n4037 ^ 1'b0 ;
  assign n4040 = n1904 ^ n1173 ^ 1'b0 ;
  assign n4041 = n22 & ~n4040 ;
  assign n4042 = n4041 ^ n3030 ^ 1'b0 ;
  assign n4043 = n3121 | n4042 ;
  assign n4044 = ~n2034 & n2192 ;
  assign n4045 = n1585 | n4044 ;
  assign n4046 = n725 & n2980 ;
  assign n4047 = n4046 ^ n2588 ^ 1'b0 ;
  assign n4048 = n3869 ^ n1858 ^ n272 ;
  assign n4049 = n4048 ^ n3235 ^ 1'b0 ;
  assign n4050 = n80 & ~n4049 ;
  assign n4051 = n1480 ^ n692 ^ 1'b0 ;
  assign n4052 = n3271 | n4051 ;
  assign n4053 = n4052 ^ n1198 ^ n496 ;
  assign n4054 = n744 ^ n469 ^ 1'b0 ;
  assign n4055 = n4054 ^ n1029 ^ n1004 ;
  assign n4056 = n4055 ^ n2436 ^ 1'b0 ;
  assign n4057 = n3097 ^ n2768 ^ 1'b0 ;
  assign n4062 = n3654 ^ n735 ^ 1'b0 ;
  assign n4063 = n4062 ^ n2752 ^ 1'b0 ;
  assign n4064 = ~n3313 & n4063 ;
  assign n4058 = n1779 ^ n525 ^ 1'b0 ;
  assign n4059 = n4058 ^ n1180 ^ 1'b0 ;
  assign n4060 = ( n757 & ~n3009 ) | ( n757 & n4059 ) | ( ~n3009 & n4059 ) ;
  assign n4061 = n2347 & n4060 ;
  assign n4065 = n4064 ^ n4061 ^ 1'b0 ;
  assign n4066 = n2225 ^ n2036 ^ 1'b0 ;
  assign n4067 = n1652 & ~n4066 ;
  assign n4068 = n766 & ~n4067 ;
  assign n4069 = n1959 & ~n4068 ;
  assign n4070 = ~n2618 & n4069 ;
  assign n4071 = n3133 ^ n2758 ^ 1'b0 ;
  assign n4072 = n1972 ^ n747 ^ 1'b0 ;
  assign n4073 = ~n1751 & n4072 ;
  assign n4074 = n1571 & n4073 ;
  assign n4076 = n702 & n712 ;
  assign n4077 = n4076 ^ n2030 ^ 1'b0 ;
  assign n4075 = n563 | n1619 ;
  assign n4078 = n4077 ^ n4075 ^ 1'b0 ;
  assign n4079 = n2653 ^ n764 ^ 1'b0 ;
  assign n4081 = ~n217 & n2964 ;
  assign n4082 = ~n1475 & n4081 ;
  assign n4080 = ~n260 & n889 ;
  assign n4083 = n4082 ^ n4080 ^ 1'b0 ;
  assign n4084 = n238 & ~n2732 ;
  assign n4091 = ~n1073 & n3394 ;
  assign n4086 = n719 ^ n35 ^ 1'b0 ;
  assign n4085 = n1248 ^ n481 ^ 1'b0 ;
  assign n4087 = n4086 ^ n4085 ^ 1'b0 ;
  assign n4088 = n1359 | n4087 ;
  assign n4089 = n238 | n4088 ;
  assign n4090 = n4089 ^ n1952 ^ 1'b0 ;
  assign n4092 = n4091 ^ n4090 ^ 1'b0 ;
  assign n4093 = n238 | n1563 ;
  assign n4094 = n3964 & n4093 ;
  assign n4095 = n4094 ^ n178 ^ 1'b0 ;
  assign n4096 = n3479 ^ n1386 ^ 1'b0 ;
  assign n4097 = ~n1771 & n4096 ;
  assign n4098 = ~n645 & n2660 ;
  assign n4099 = ~n803 & n4098 ;
  assign n4101 = n1717 & n2320 ;
  assign n4102 = ~n1260 & n4101 ;
  assign n4100 = ~n65 & n523 ;
  assign n4103 = n4102 ^ n4100 ^ 1'b0 ;
  assign n4104 = ~n1716 & n4103 ;
  assign n4106 = n633 ^ n197 ^ 1'b0 ;
  assign n4107 = ~n228 & n4106 ;
  assign n4108 = x10 & ~n691 ;
  assign n4109 = n1045 & n4108 ;
  assign n4110 = n1582 | n4109 ;
  assign n4111 = ( n1231 & ~n4107 ) | ( n1231 & n4110 ) | ( ~n4107 & n4110 ) ;
  assign n4105 = ( x10 & ~n1516 ) | ( x10 & n2387 ) | ( ~n1516 & n2387 ) ;
  assign n4112 = n4111 ^ n4105 ^ 1'b0 ;
  assign n4113 = n1980 & n4112 ;
  assign n4114 = n1149 & ~n2286 ;
  assign n4115 = n3566 ^ n510 ^ 1'b0 ;
  assign n4116 = n1641 ^ n1202 ^ 1'b0 ;
  assign n4117 = ~n2475 & n4116 ;
  assign n4118 = n2080 & n4117 ;
  assign n4119 = n4118 ^ n1363 ^ 1'b0 ;
  assign n4120 = n2505 & n4119 ;
  assign n4121 = n82 | n4120 ;
  assign n4122 = n1517 & n2425 ;
  assign n4123 = n2986 | n4122 ;
  assign n4124 = n2484 & n2761 ;
  assign n4127 = ~n788 & n1234 ;
  assign n4125 = n2687 ^ n2566 ^ 1'b0 ;
  assign n4126 = n3223 & ~n4125 ;
  assign n4128 = n4127 ^ n4126 ^ n2560 ;
  assign n4132 = n1959 ^ n744 ^ 1'b0 ;
  assign n4129 = n957 ^ n317 ^ n51 ;
  assign n4130 = n4129 ^ n57 ^ 1'b0 ;
  assign n4131 = n911 & ~n4130 ;
  assign n4133 = n4132 ^ n4131 ^ 1'b0 ;
  assign n4134 = n1902 & ~n4133 ;
  assign n4135 = n4134 ^ n1444 ^ n1175 ;
  assign n4138 = n1029 ^ n1022 ^ n852 ;
  assign n4139 = n4138 ^ n3043 ^ 1'b0 ;
  assign n4140 = n2539 & ~n4139 ;
  assign n4136 = n1779 ^ n135 ^ 1'b0 ;
  assign n4137 = n115 & n4136 ;
  assign n4141 = n4140 ^ n4137 ^ 1'b0 ;
  assign n4142 = ~n1521 & n2032 ;
  assign n4149 = n2610 | n2673 ;
  assign n4143 = n2694 ^ n1521 ^ 1'b0 ;
  assign n4144 = ( n462 & n3137 ) | ( n462 & n4143 ) | ( n3137 & n4143 ) ;
  assign n4145 = n364 | n480 ;
  assign n4146 = n4145 ^ n1839 ^ 1'b0 ;
  assign n4147 = n4146 ^ n2378 ^ 1'b0 ;
  assign n4148 = n4144 & n4147 ;
  assign n4150 = n4149 ^ n4148 ^ 1'b0 ;
  assign n4151 = n588 | n3790 ;
  assign n4152 = n137 & n2176 ;
  assign n4153 = n4152 ^ n1762 ^ 1'b0 ;
  assign n4154 = n611 | n4153 ;
  assign n4157 = n1303 & n2217 ;
  assign n4158 = ~n44 & n4157 ;
  assign n4159 = n1041 & ~n4158 ;
  assign n4155 = n481 | n2580 ;
  assign n4156 = n418 | n4155 ;
  assign n4160 = n4159 ^ n4156 ^ 1'b0 ;
  assign n4163 = ~n806 & n1470 ;
  assign n4164 = n4163 ^ n3633 ^ n846 ;
  assign n4161 = n3429 ^ n2963 ^ 1'b0 ;
  assign n4162 = n2282 & n4161 ;
  assign n4165 = n4164 ^ n4162 ^ 1'b0 ;
  assign n4166 = n142 | n3998 ;
  assign n4167 = n4166 ^ n2014 ^ 1'b0 ;
  assign n4168 = n2071 & n4167 ;
  assign n4169 = n3837 ^ n1387 ^ 1'b0 ;
  assign n4170 = n4168 | n4169 ;
  assign n4171 = n823 | n4170 ;
  assign n4172 = n976 ^ n735 ^ 1'b0 ;
  assign n4173 = n411 | n4172 ;
  assign n4174 = n4173 ^ n2384 ^ 1'b0 ;
  assign n4175 = n3554 | n4174 ;
  assign n4176 = n536 ^ n435 ^ 1'b0 ;
  assign n4177 = ~n511 & n4176 ;
  assign n4178 = ~n228 & n1526 ;
  assign n4179 = n4178 ^ n3569 ^ 1'b0 ;
  assign n4180 = n2727 ^ n2556 ^ n401 ;
  assign n4181 = ~n3229 & n4180 ;
  assign n4182 = n1260 ^ n750 ^ 1'b0 ;
  assign n4183 = ~n1386 & n4182 ;
  assign n4184 = n4183 ^ n1234 ^ 1'b0 ;
  assign n4185 = ~n4062 & n4184 ;
  assign n4186 = n2918 & ~n3100 ;
  assign n4187 = ( n400 & n848 ) | ( n400 & ~n3353 ) | ( n848 & ~n3353 ) ;
  assign n4188 = n881 & ~n2979 ;
  assign n4189 = n4188 ^ n916 ^ 1'b0 ;
  assign n4190 = n3517 ^ n2582 ^ 1'b0 ;
  assign n4191 = n4189 | n4190 ;
  assign n4192 = n3277 ^ n1025 ^ n246 ;
  assign n4193 = ~n3959 & n4192 ;
  assign n4194 = n4193 ^ n983 ^ 1'b0 ;
  assign n4195 = n2976 & ~n4194 ;
  assign n4196 = n740 ^ n682 ^ n220 ;
  assign n4197 = n1287 & n2828 ;
  assign n4199 = n887 | n1326 ;
  assign n4198 = n263 | n3435 ;
  assign n4200 = n4199 ^ n4198 ^ 1'b0 ;
  assign n4201 = ~n448 & n2190 ;
  assign n4202 = n1566 ^ x9 ^ 1'b0 ;
  assign n4203 = n2050 ^ n1402 ^ 1'b0 ;
  assign n4204 = n4203 ^ n1943 ^ n351 ;
  assign n4205 = ( n1243 & ~n4202 ) | ( n1243 & n4204 ) | ( ~n4202 & n4204 ) ;
  assign n4206 = n3410 & n4205 ;
  assign n4207 = n4201 & n4206 ;
  assign n4208 = ~n102 & n2207 ;
  assign n4209 = n4208 ^ n2733 ^ 1'b0 ;
  assign n4210 = n4123 | n4209 ;
  assign n4211 = n2413 ^ n884 ^ n265 ;
  assign n4212 = ~n1441 & n3720 ;
  assign n4213 = n309 & n4212 ;
  assign n4214 = ~n463 & n4213 ;
  assign n4215 = n4214 ^ n1942 ^ 1'b0 ;
  assign n4216 = n1585 | n2187 ;
  assign n4217 = n4216 ^ n1374 ^ 1'b0 ;
  assign n4218 = n1092 ^ n304 ^ 1'b0 ;
  assign n4219 = n3296 ^ n711 ^ 1'b0 ;
  assign n4220 = n2757 ^ n102 ^ 1'b0 ;
  assign n4221 = n532 ^ n202 ^ n44 ;
  assign n4222 = n525 & n4221 ;
  assign n4223 = n4220 | n4222 ;
  assign n4224 = n3484 ^ n2129 ^ 1'b0 ;
  assign n4225 = n3645 & ~n4224 ;
  assign n4226 = n1835 & ~n2755 ;
  assign n4227 = n4226 ^ n2034 ^ n1310 ;
  assign n4228 = n4227 ^ n582 ^ 1'b0 ;
  assign n4229 = n1699 & ~n2283 ;
  assign n4230 = ~n3413 & n4229 ;
  assign n4231 = n247 | n556 ;
  assign n4232 = n1781 & n3363 ;
  assign n4233 = ( n2911 & n4231 ) | ( n2911 & n4232 ) | ( n4231 & n4232 ) ;
  assign n4234 = x6 & n2344 ;
  assign n4235 = ( n1262 & n2750 ) | ( n1262 & ~n3241 ) | ( n2750 & ~n3241 ) ;
  assign n4236 = n4235 ^ n2565 ^ 1'b0 ;
  assign n4237 = n3636 | n4236 ;
  assign n4238 = ~n787 & n2173 ;
  assign n4239 = ~n2977 & n4238 ;
  assign n4240 = n1467 | n1800 ;
  assign n4241 = n4240 ^ n2345 ^ 1'b0 ;
  assign n4242 = n893 | n2571 ;
  assign n4244 = ~n639 & n771 ;
  assign n4245 = n3779 & n4244 ;
  assign n4246 = n4245 ^ n3202 ^ n1913 ;
  assign n4247 = n4246 ^ n349 ^ 1'b0 ;
  assign n4243 = n3120 ^ n897 ^ n790 ;
  assign n4248 = n4247 ^ n4243 ^ 1'b0 ;
  assign n4249 = n3615 & n4248 ;
  assign n4250 = ~n2385 & n2433 ;
  assign n4251 = n4250 ^ n3482 ^ n846 ;
  assign n4252 = n1948 | n2594 ;
  assign n4253 = n1285 ^ x10 ^ 1'b0 ;
  assign n4254 = n252 | n818 ;
  assign n4255 = n1720 | n4254 ;
  assign n4256 = n1171 & ~n4255 ;
  assign n4257 = ( n1134 & ~n1641 ) | ( n1134 & n2719 ) | ( ~n1641 & n2719 ) ;
  assign n4258 = n84 | n129 ;
  assign n4259 = n4258 ^ n1079 ^ 1'b0 ;
  assign n4260 = n80 | n1871 ;
  assign n4261 = n4260 ^ n1274 ^ 1'b0 ;
  assign n4262 = ~n637 & n4261 ;
  assign n4263 = n4262 ^ n1666 ^ 1'b0 ;
  assign n4264 = ~n603 & n1298 ;
  assign n4265 = ( ~n1355 & n2056 ) | ( ~n1355 & n2765 ) | ( n2056 & n2765 ) ;
  assign n4269 = n153 & n1842 ;
  assign n4270 = n1602 & n4269 ;
  assign n4266 = n3897 ^ n1040 ^ 1'b0 ;
  assign n4267 = n1133 | n4266 ;
  assign n4268 = n1952 | n4267 ;
  assign n4271 = n4270 ^ n4268 ^ 1'b0 ;
  assign n4272 = n4014 ^ n1451 ^ 1'b0 ;
  assign n4273 = n4272 ^ n1460 ^ n67 ;
  assign n4274 = n3750 & ~n4273 ;
  assign n4275 = ( ~n1121 & n1300 ) | ( ~n1121 & n2123 ) | ( n1300 & n2123 ) ;
  assign n4276 = n4275 ^ n4262 ^ n1828 ;
  assign n4277 = n4276 ^ n4273 ^ 1'b0 ;
  assign n4278 = n4277 ^ n1614 ^ n108 ;
  assign n4279 = ~n1516 & n3040 ;
  assign n4280 = ~n732 & n4279 ;
  assign n4282 = n2381 | n3310 ;
  assign n4283 = n1400 | n4282 ;
  assign n4281 = n1587 & ~n1820 ;
  assign n4284 = n4283 ^ n4281 ^ 1'b0 ;
  assign n4285 = n169 & n4284 ;
  assign n4286 = n153 & n2811 ;
  assign n4287 = n496 | n2113 ;
  assign n4288 = ~n37 & n1332 ;
  assign n4289 = ( n40 & n372 ) | ( n40 & n4288 ) | ( n372 & n4288 ) ;
  assign n4290 = n976 ^ n424 ^ n245 ;
  assign n4291 = n4290 ^ n926 ^ 1'b0 ;
  assign n4292 = ~n4289 & n4291 ;
  assign n4293 = n4292 ^ n1348 ^ 1'b0 ;
  assign n4294 = ~n3919 & n4293 ;
  assign n4296 = n1290 & ~n1533 ;
  assign n4295 = ~n3102 & n4257 ;
  assign n4297 = n4296 ^ n4295 ^ 1'b0 ;
  assign n4298 = ( n1568 & n1681 ) | ( n1568 & n3049 ) | ( n1681 & n3049 ) ;
  assign n4299 = n3973 & ~n4298 ;
  assign n4300 = ~n578 & n4299 ;
  assign n4301 = ~n1376 & n4300 ;
  assign n4302 = n4301 ^ n3456 ^ 1'b0 ;
  assign n4303 = n16 & n4302 ;
  assign n4304 = ( n1357 & n1957 ) | ( n1357 & n3819 ) | ( n1957 & n3819 ) ;
  assign n4305 = ~n1011 & n1731 ;
  assign n4306 = n107 & n168 ;
  assign n4307 = ~n1212 & n4306 ;
  assign n4308 = ~n159 & n4307 ;
  assign n4309 = ( n32 & n1274 ) | ( n32 & n2159 ) | ( n1274 & n2159 ) ;
  assign n4310 = n1402 | n4309 ;
  assign n4311 = n2021 & n4310 ;
  assign n4312 = n2666 & n4218 ;
  assign n4313 = n4312 ^ n1348 ^ 1'b0 ;
  assign n4314 = n1078 ^ n41 ^ 1'b0 ;
  assign n4315 = n637 | n4314 ;
  assign n4316 = n2221 ^ n1569 ^ 1'b0 ;
  assign n4317 = n4316 ^ n2808 ^ 1'b0 ;
  assign n4318 = n4317 ^ n1240 ^ n188 ;
  assign n4319 = n3016 ^ n532 ^ 1'b0 ;
  assign n4320 = ~n2313 & n4319 ;
  assign n4321 = n3127 ^ n627 ^ 1'b0 ;
  assign n4322 = ~n1525 & n4321 ;
  assign n4323 = ~n1168 & n4322 ;
  assign n4324 = n4323 ^ n2556 ^ 1'b0 ;
  assign n4325 = n89 & ~n4252 ;
  assign n4326 = n2403 | n3530 ;
  assign n4327 = ~n611 & n1188 ;
  assign n4328 = n4327 ^ n1403 ^ n1061 ;
  assign n4330 = n2281 ^ n1718 ^ n829 ;
  assign n4329 = n2915 | n3988 ;
  assign n4331 = n4330 ^ n4329 ^ 1'b0 ;
  assign n4332 = n1320 & n3755 ;
  assign n4333 = ~n835 & n4332 ;
  assign n4334 = n2241 | n4333 ;
  assign n4335 = n876 | n1950 ;
  assign n4336 = ( n2230 & n4319 ) | ( n2230 & n4335 ) | ( n4319 & n4335 ) ;
  assign n4337 = n1326 & ~n2832 ;
  assign n4338 = ( ~n98 & n652 ) | ( ~n98 & n722 ) | ( n652 & n722 ) ;
  assign n4339 = n1566 ^ n596 ^ n390 ;
  assign n4340 = n4339 ^ n1789 ^ n32 ;
  assign n4341 = n4340 ^ n1690 ^ 1'b0 ;
  assign n4342 = n596 & n1827 ;
  assign n4343 = ( n859 & n1400 ) | ( n859 & ~n3791 ) | ( n1400 & ~n3791 ) ;
  assign n4344 = n4343 ^ n1446 ^ 1'b0 ;
  assign n4345 = n4344 ^ n177 ^ 1'b0 ;
  assign n4346 = n1241 & n4345 ;
  assign n4347 = ~n3177 & n4346 ;
  assign n4348 = n728 & ~n2705 ;
  assign n4349 = n209 & ~n316 ;
  assign n4350 = n4349 ^ n999 ^ 1'b0 ;
  assign n4351 = n2758 ^ n1348 ^ 1'b0 ;
  assign n4352 = n4351 ^ n1262 ^ 1'b0 ;
  assign n4353 = n2779 | n4352 ;
  assign n4354 = n1357 | n4353 ;
  assign n4355 = n4114 ^ n2516 ^ 1'b0 ;
  assign n4356 = n2960 ^ n1232 ^ 1'b0 ;
  assign n4357 = n725 ^ n174 ^ 1'b0 ;
  assign n4358 = n4357 ^ n1875 ^ 1'b0 ;
  assign n4359 = n755 | n4358 ;
  assign n4360 = ~n1638 & n2282 ;
  assign n4361 = n4360 ^ n164 ^ 1'b0 ;
  assign n4362 = n4361 ^ n353 ^ 1'b0 ;
  assign n4363 = n1527 | n4362 ;
  assign n4364 = ( n1140 & n1852 ) | ( n1140 & n1962 ) | ( n1852 & n1962 ) ;
  assign n4365 = ~n635 & n3292 ;
  assign n4366 = n1112 & n1940 ;
  assign n4367 = n2476 & ~n4366 ;
  assign n4368 = ( ~n214 & n466 ) | ( ~n214 & n1666 ) | ( n466 & n1666 ) ;
  assign n4369 = n966 & n4368 ;
  assign n4370 = n3526 ^ n1744 ^ 1'b0 ;
  assign n4371 = n3939 | n4370 ;
  assign n4372 = n3863 | n4111 ;
  assign n4373 = n4235 ^ n3951 ^ 1'b0 ;
  assign n4376 = n261 | n406 ;
  assign n4377 = n2873 & n4376 ;
  assign n4378 = ( n706 & n2699 ) | ( n706 & n4377 ) | ( n2699 & n4377 ) ;
  assign n4374 = n1164 ^ n111 ^ 1'b0 ;
  assign n4375 = ~n480 & n4374 ;
  assign n4379 = n4378 ^ n4375 ^ 1'b0 ;
  assign n4380 = n13 & n4379 ;
  assign n4381 = n969 | n2951 ;
  assign n4382 = n848 | n3879 ;
  assign n4383 = n1405 & n2140 ;
  assign n4386 = n4082 ^ n1296 ^ 1'b0 ;
  assign n4387 = n711 & ~n4386 ;
  assign n4384 = n1550 & ~n2337 ;
  assign n4385 = ~n1902 & n4384 ;
  assign n4388 = n4387 ^ n4385 ^ n1355 ;
  assign n4389 = n1767 & n2122 ;
  assign n4390 = n349 & n4389 ;
  assign n4391 = ( ~x7 & n136 ) | ( ~x7 & n506 ) | ( n136 & n506 ) ;
  assign n4392 = n4391 ^ n2542 ^ 1'b0 ;
  assign n4393 = n334 | n4392 ;
  assign n4394 = n4393 ^ n3767 ^ 1'b0 ;
  assign n4395 = n168 & n3846 ;
  assign n4396 = n4395 ^ n1700 ^ 1'b0 ;
  assign n4397 = ( ~n1068 & n2885 ) | ( ~n1068 & n4396 ) | ( n2885 & n4396 ) ;
  assign n4402 = n2918 ^ n1783 ^ n1036 ;
  assign n4398 = n2034 ^ n965 ^ 1'b0 ;
  assign n4399 = n40 & ~n4398 ;
  assign n4400 = n2256 | n4399 ;
  assign n4401 = n2694 & n4400 ;
  assign n4403 = n4402 ^ n4401 ^ 1'b0 ;
  assign n4404 = n401 ^ x10 ^ 1'b0 ;
  assign n4405 = ( n308 & n1880 ) | ( n308 & n4404 ) | ( n1880 & n4404 ) ;
  assign n4406 = n1324 | n4405 ;
  assign n4407 = n1629 & ~n2789 ;
  assign n4408 = n202 & n4407 ;
  assign n4409 = n115 & n2662 ;
  assign n4410 = n4409 ^ n4006 ^ 1'b0 ;
  assign n4411 = n3555 | n4410 ;
  assign n4412 = n1909 & ~n3020 ;
  assign n4413 = n3359 ^ n1771 ^ 1'b0 ;
  assign n4414 = n4413 ^ n57 ^ 1'b0 ;
  assign n4415 = n1050 | n4414 ;
  assign n4416 = n545 | n4415 ;
  assign n4417 = n2570 & ~n4416 ;
  assign n4418 = ~n953 & n4417 ;
  assign n4419 = n1823 & n4418 ;
  assign n4420 = n2849 ^ n1535 ^ 1'b0 ;
  assign n4421 = n3655 & ~n4420 ;
  assign n4422 = n3088 ^ n2726 ^ 1'b0 ;
  assign n4423 = n1502 ^ n1272 ^ 1'b0 ;
  assign n4424 = n3500 | n4423 ;
  assign n4425 = n4424 ^ n2182 ^ 1'b0 ;
  assign n4426 = n2428 ^ n1407 ^ 1'b0 ;
  assign n4427 = n2917 ^ n2104 ^ 1'b0 ;
  assign n4428 = ( n769 & n2228 ) | ( n769 & ~n4427 ) | ( n2228 & ~n4427 ) ;
  assign n4429 = n4428 ^ n1223 ^ n1149 ;
  assign n4430 = n3720 ^ n2337 ^ 1'b0 ;
  assign n4431 = ~n102 & n4430 ;
  assign n4432 = n4431 ^ n3750 ^ 1'b0 ;
  assign n4433 = n77 & ~n1548 ;
  assign n4434 = n4433 ^ n1206 ^ 1'b0 ;
  assign n4435 = ( n1233 & n1930 ) | ( n1233 & n4434 ) | ( n1930 & n4434 ) ;
  assign n4436 = n4435 ^ n3165 ^ n3149 ;
  assign n4437 = n3687 ^ n202 ^ 1'b0 ;
  assign n4438 = n4436 | n4437 ;
  assign n4439 = n4432 | n4438 ;
  assign n4440 = n1614 & ~n2041 ;
  assign n4441 = n928 & n4440 ;
  assign n4442 = n4441 ^ n326 ^ 1'b0 ;
  assign n4443 = n1904 | n2225 ;
  assign n4444 = n125 | n4443 ;
  assign n4445 = n4444 ^ n2759 ^ 1'b0 ;
  assign n4446 = n813 & n2241 ;
  assign n4447 = n4445 & ~n4446 ;
  assign n4452 = ( n1046 & n1564 ) | ( n1046 & ~n2060 ) | ( n1564 & ~n2060 ) ;
  assign n4450 = ( n63 & n270 ) | ( n63 & ~n1662 ) | ( n270 & ~n1662 ) ;
  assign n4451 = n1351 | n4450 ;
  assign n4453 = n4452 ^ n4451 ^ 1'b0 ;
  assign n4449 = n3495 & n3557 ;
  assign n4454 = n4453 ^ n4449 ^ 1'b0 ;
  assign n4448 = n854 & n2877 ;
  assign n4455 = n4454 ^ n4448 ^ 1'b0 ;
  assign n4456 = n2370 & ~n3737 ;
  assign n4457 = n4456 ^ n3059 ^ 1'b0 ;
  assign n4458 = ( x8 & n145 ) | ( x8 & ~n4457 ) | ( n145 & ~n4457 ) ;
  assign n4459 = n4458 ^ n532 ^ 1'b0 ;
  assign n4460 = n4459 ^ n953 ^ 1'b0 ;
  assign n4462 = n1418 ^ n621 ^ 1'b0 ;
  assign n4463 = ( n1149 & ~n2505 ) | ( n1149 & n4343 ) | ( ~n2505 & n4343 ) ;
  assign n4464 = ( n3602 & n4462 ) | ( n3602 & ~n4463 ) | ( n4462 & ~n4463 ) ;
  assign n4461 = ~n1522 & n2525 ;
  assign n4465 = n4464 ^ n4461 ^ n2830 ;
  assign n4466 = n3782 ^ n368 ^ 1'b0 ;
  assign n4467 = n3446 | n4466 ;
  assign n4468 = n3608 | n4467 ;
  assign n4469 = n135 & n1664 ;
  assign n4470 = n4469 ^ n1439 ^ 1'b0 ;
  assign n4471 = n4468 | n4470 ;
  assign n4472 = n1800 | n4471 ;
  assign n4473 = n2980 | n4472 ;
  assign n4474 = n672 ^ n648 ^ 1'b0 ;
  assign n4475 = n1741 & ~n4474 ;
  assign n4476 = n4475 ^ n238 ^ 1'b0 ;
  assign n4477 = n2365 | n4476 ;
  assign n4478 = n2575 & ~n4477 ;
  assign n4479 = ~n3410 & n4478 ;
  assign n4480 = n1407 & n2225 ;
  assign n4481 = n903 & n4273 ;
  assign n4482 = ~n2625 & n4481 ;
  assign n4483 = n4482 ^ n3465 ^ 1'b0 ;
  assign n4484 = n927 | n3027 ;
  assign n4485 = n4484 ^ n3133 ^ 1'b0 ;
  assign n4486 = n4485 ^ n2147 ^ n276 ;
  assign n4487 = ~n3469 & n4486 ;
  assign n4488 = n3218 ^ n1336 ^ 1'b0 ;
  assign n4489 = n303 | n4488 ;
  assign n4490 = n2009 ^ n776 ^ 1'b0 ;
  assign n4491 = n4489 & ~n4490 ;
  assign n4492 = n32 | n603 ;
  assign n4493 = n4492 ^ n619 ^ 1'b0 ;
  assign n4494 = n4493 ^ n3351 ^ 1'b0 ;
  assign n4495 = ~n4491 & n4494 ;
  assign n4496 = ~n3399 & n4495 ;
  assign n4497 = n4496 ^ n3866 ^ 1'b0 ;
  assign n4498 = n601 & n2676 ;
  assign n4499 = n2154 & ~n4498 ;
  assign n4500 = n4499 ^ n1270 ^ 1'b0 ;
  assign n4502 = n1516 ^ n1255 ^ 1'b0 ;
  assign n4501 = n3105 | n3699 ;
  assign n4503 = n4502 ^ n4501 ^ 1'b0 ;
  assign n4504 = n4503 ^ n1302 ^ 1'b0 ;
  assign n4505 = n4500 | n4504 ;
  assign n4506 = n1054 & n2421 ;
  assign n4507 = n2354 & ~n2612 ;
  assign n4508 = n1991 ^ n1937 ^ n1875 ;
  assign n4509 = n4508 ^ n3750 ^ 1'b0 ;
  assign n4510 = ~n2429 & n4509 ;
  assign n4511 = n2241 & n2951 ;
  assign n4512 = n4511 ^ n1443 ^ n1412 ;
  assign n4513 = n809 | n4404 ;
  assign n4514 = n4513 ^ n1007 ^ 1'b0 ;
  assign n4515 = n4514 ^ n2062 ^ n1926 ;
  assign n4516 = n4515 ^ n1435 ^ 1'b0 ;
  assign n4519 = n35 & n426 ;
  assign n4520 = n4519 ^ n1676 ^ 1'b0 ;
  assign n4517 = n99 & ~n374 ;
  assign n4518 = n1031 & n4517 ;
  assign n4521 = n4520 ^ n4518 ^ n998 ;
  assign n4522 = ~n4095 & n4521 ;
  assign n4523 = n4522 ^ n788 ^ 1'b0 ;
  assign n4524 = n3225 | n3793 ;
  assign n4525 = n4524 ^ n647 ^ 1'b0 ;
  assign n4526 = ~n2887 & n4525 ;
  assign n4527 = n641 ^ n209 ^ 1'b0 ;
  assign n4528 = ~n4526 & n4527 ;
  assign n4529 = n2051 ^ n1056 ^ 1'b0 ;
  assign n4530 = n2202 ^ n1105 ^ 1'b0 ;
  assign n4531 = n1105 & n1220 ;
  assign n4532 = n1640 ^ n289 ^ 1'b0 ;
  assign n4533 = n3720 & ~n4532 ;
  assign n4534 = ( n667 & n1400 ) | ( n667 & n4533 ) | ( n1400 & n4533 ) ;
  assign n4535 = n3406 ^ n2537 ^ 1'b0 ;
  assign n4536 = n1600 & n4535 ;
  assign n4537 = ( n545 & ~n3544 ) | ( n545 & n4290 ) | ( ~n3544 & n4290 ) ;
  assign n4538 = n1303 | n1716 ;
  assign n4539 = n2134 & ~n2532 ;
  assign n4540 = n4539 ^ n2261 ^ n1261 ;
  assign n4541 = n4540 ^ n3584 ^ 1'b0 ;
  assign n4542 = ( n1247 & n4538 ) | ( n1247 & n4541 ) | ( n4538 & n4541 ) ;
  assign n4543 = n870 ^ n434 ^ 1'b0 ;
  assign n4544 = n1496 | n4543 ;
  assign n4545 = n126 | n4544 ;
  assign n4546 = n430 & ~n2837 ;
  assign n4547 = n1176 & n4546 ;
  assign n4548 = n4547 ^ n32 ^ 1'b0 ;
  assign n4551 = n1311 ^ n491 ^ 1'b0 ;
  assign n4549 = n1013 ^ n204 ^ 1'b0 ;
  assign n4550 = n220 & ~n4549 ;
  assign n4552 = n4551 ^ n4550 ^ 1'b0 ;
  assign n4553 = ~n4430 & n4552 ;
  assign n4554 = ~n2986 & n4292 ;
  assign n4555 = ~n1507 & n4554 ;
  assign n4556 = ~n2726 & n4258 ;
  assign n4557 = ~n2327 & n4556 ;
  assign n4558 = n3491 ^ n464 ^ 1'b0 ;
  assign n4559 = n2389 | n4072 ;
  assign n4560 = n4559 ^ n2661 ^ n525 ;
  assign n4561 = n622 & ~n1298 ;
  assign n4562 = n4561 ^ n1639 ^ 1'b0 ;
  assign n4563 = n620 | n957 ;
  assign n4564 = n98 | n4563 ;
  assign n4565 = n2270 | n4564 ;
  assign n4566 = n1105 & n4565 ;
  assign n4567 = ~n2148 & n4566 ;
  assign n4568 = ( n137 & n654 ) | ( n137 & ~n4567 ) | ( n654 & ~n4567 ) ;
  assign n4569 = n2684 & n4568 ;
  assign n4570 = n1820 ^ n795 ^ 1'b0 ;
  assign n4571 = n4570 ^ n3997 ^ 1'b0 ;
  assign n4572 = n1922 & ~n3812 ;
  assign n4577 = n2597 ^ n2094 ^ 1'b0 ;
  assign n4573 = n22 & ~n1290 ;
  assign n4574 = n1865 & n4573 ;
  assign n4575 = ( n1888 & ~n2828 ) | ( n1888 & n4574 ) | ( ~n2828 & n4574 ) ;
  assign n4576 = n4575 ^ n4072 ^ n3353 ;
  assign n4578 = n4577 ^ n4576 ^ 1'b0 ;
  assign n4579 = ( n3014 & ~n3173 ) | ( n3014 & n3700 ) | ( ~n3173 & n3700 ) ;
  assign n4580 = n4422 ^ n3409 ^ n2483 ;
  assign n4581 = n853 & n928 ;
  assign n4582 = n4581 ^ n2104 ^ 1'b0 ;
  assign n4583 = n4582 ^ n607 ^ 1'b0 ;
  assign n4584 = n1216 & ~n4583 ;
  assign n4585 = n3867 & n4584 ;
  assign n4586 = ~n4580 & n4585 ;
  assign n4587 = n1997 | n4586 ;
  assign n4588 = n878 ^ n566 ^ 1'b0 ;
  assign n4589 = n3064 & ~n4588 ;
  assign n4590 = n4589 ^ n1120 ^ 1'b0 ;
  assign n4593 = ( n451 & n913 ) | ( n451 & ~n2670 ) | ( n913 & ~n2670 ) ;
  assign n4594 = n3686 | n4593 ;
  assign n4595 = n2409 & ~n4594 ;
  assign n4591 = ( n430 & ~n1069 ) | ( n430 & n1168 ) | ( ~n1069 & n1168 ) ;
  assign n4592 = n1293 & ~n4591 ;
  assign n4596 = n4595 ^ n4592 ^ 1'b0 ;
  assign n4597 = n4078 ^ n1764 ^ 1'b0 ;
  assign n4598 = n4562 | n4597 ;
  assign n4599 = n1339 & n4598 ;
  assign n4601 = ~n481 & n777 ;
  assign n4602 = n1866 & n4601 ;
  assign n4603 = n1578 & ~n4602 ;
  assign n4604 = n4603 ^ n3127 ^ 1'b0 ;
  assign n4600 = n863 & n3560 ;
  assign n4605 = n4604 ^ n4600 ^ 1'b0 ;
  assign n4606 = n1686 ^ n369 ^ 1'b0 ;
  assign n4607 = n2913 | n4606 ;
  assign n4608 = n63 & n461 ;
  assign n4609 = ~n2851 & n4608 ;
  assign n4610 = n4607 & n4609 ;
  assign n4611 = n1207 | n1643 ;
  assign n4612 = n3614 | n4611 ;
  assign n4613 = n2328 & ~n2672 ;
  assign n4614 = n4613 ^ n183 ^ 1'b0 ;
  assign n4615 = n4614 ^ n3881 ^ 1'b0 ;
  assign n4616 = ~n2503 & n4278 ;
  assign n4617 = n3384 & n4616 ;
  assign n4618 = n4617 ^ n3882 ^ 1'b0 ;
  assign n4619 = n1893 | n3149 ;
  assign n4620 = n168 | n4619 ;
  assign n4625 = n1896 ^ n839 ^ 1'b0 ;
  assign n4626 = ~n921 & n4625 ;
  assign n4621 = n3195 ^ n1472 ^ 1'b0 ;
  assign n4622 = ~n2451 & n4621 ;
  assign n4623 = ~n162 & n4622 ;
  assign n4624 = ~n1017 & n4623 ;
  assign n4627 = n4626 ^ n4624 ^ 1'b0 ;
  assign n4628 = n4627 ^ n4252 ^ 1'b0 ;
  assign n4629 = ( ~n3882 & n4195 ) | ( ~n3882 & n4628 ) | ( n4195 & n4628 ) ;
  assign n4630 = n1881 & ~n3663 ;
  assign n4631 = ~n3555 & n4630 ;
  assign n4632 = n2539 & n2827 ;
  assign n4633 = n4632 ^ n117 ^ 1'b0 ;
  assign n4634 = n709 & n4633 ;
  assign n4635 = ~n1629 & n4634 ;
  assign n4636 = n614 & n887 ;
  assign n4637 = n4636 ^ n500 ^ 1'b0 ;
  assign n4638 = ( n1315 & n2757 ) | ( n1315 & ~n4637 ) | ( n2757 & ~n4637 ) ;
  assign n4639 = n3523 | n4638 ;
  assign n4640 = ( n108 & ~n2101 ) | ( n108 & n3229 ) | ( ~n2101 & n3229 ) ;
  assign n4641 = n3184 ^ n2012 ^ 1'b0 ;
  assign n4642 = n4641 ^ n328 ^ n100 ;
  assign n4643 = n1642 ^ n315 ^ 1'b0 ;
  assign n4644 = n547 | n4643 ;
  assign n4645 = ( ~n403 & n926 ) | ( ~n403 & n1741 ) | ( n926 & n1741 ) ;
  assign n4646 = n4645 ^ n2531 ^ 1'b0 ;
  assign n4647 = n4646 ^ n719 ^ 1'b0 ;
  assign n4648 = n2216 ^ n98 ^ 1'b0 ;
  assign n4649 = n1336 & n1578 ;
  assign n4650 = n4649 ^ n276 ^ 1'b0 ;
  assign n4651 = ~n570 & n1253 ;
  assign n4652 = n2857 & n4651 ;
  assign n4653 = ~n1378 & n4652 ;
  assign n4654 = n1137 | n4653 ;
  assign n4655 = n1167 & n1674 ;
  assign n4656 = n4655 ^ n3802 ^ 1'b0 ;
  assign n4657 = ~n2072 & n4656 ;
  assign n4658 = n1746 ^ n966 ^ 1'b0 ;
  assign n4661 = n1768 ^ n78 ^ 1'b0 ;
  assign n4660 = ( n237 & n2170 ) | ( n237 & ~n2528 ) | ( n2170 & ~n2528 ) ;
  assign n4659 = ~n889 & n1234 ;
  assign n4662 = n4661 ^ n4660 ^ n4659 ;
  assign n4663 = ~n255 & n1764 ;
  assign n4664 = n766 ^ n126 ^ 1'b0 ;
  assign n4665 = n3057 & ~n4664 ;
  assign n4666 = ~n955 & n4665 ;
  assign n4667 = ~n3465 & n4666 ;
  assign n4668 = n1175 | n2137 ;
  assign n4669 = n316 | n863 ;
  assign n4670 = n777 | n4669 ;
  assign n4672 = n352 & ~n3988 ;
  assign n4673 = n4672 ^ n1320 ^ 1'b0 ;
  assign n4671 = n3531 ^ n951 ^ 1'b0 ;
  assign n4674 = n4673 ^ n4671 ^ n1361 ;
  assign n4675 = n2749 ^ n523 ^ n174 ;
  assign n4676 = n1748 ^ n1250 ^ 1'b0 ;
  assign n4677 = n4675 & n4676 ;
  assign n4684 = ( n326 & n1751 ) | ( n326 & ~n3261 ) | ( n1751 & ~n3261 ) ;
  assign n4678 = ( ~n817 & n1038 ) | ( ~n817 & n2054 ) | ( n1038 & n2054 ) ;
  assign n4679 = n352 ^ n158 ^ 1'b0 ;
  assign n4680 = n4679 ^ n2752 ^ 1'b0 ;
  assign n4681 = n4678 & ~n4680 ;
  assign n4682 = ~n1351 & n4681 ;
  assign n4683 = n4682 ^ n4008 ^ 1'b0 ;
  assign n4685 = n4684 ^ n4683 ^ n411 ;
  assign n4687 = n506 & n556 ;
  assign n4688 = n2784 & n4687 ;
  assign n4686 = n1052 & n2831 ;
  assign n4689 = n4688 ^ n4686 ^ n1360 ;
  assign n4690 = ( ~n790 & n2203 ) | ( ~n790 & n3922 ) | ( n2203 & n3922 ) ;
  assign n4691 = n3158 & n4690 ;
  assign n4694 = n2135 & ~n3709 ;
  assign n4695 = ~n840 & n4694 ;
  assign n4692 = n1206 ^ n20 ^ 1'b0 ;
  assign n4693 = ~n3812 & n4692 ;
  assign n4696 = n4695 ^ n4693 ^ n582 ;
  assign n4697 = n4696 ^ n1382 ^ 1'b0 ;
  assign n4698 = n4697 ^ n889 ^ 1'b0 ;
  assign n4699 = n1480 ^ n177 ^ 1'b0 ;
  assign n4700 = n4699 ^ n729 ^ 1'b0 ;
  assign n4701 = n4700 ^ n3109 ^ 1'b0 ;
  assign n4702 = n3508 ^ n2901 ^ 1'b0 ;
  assign n4703 = n757 ^ n521 ^ 1'b0 ;
  assign n4704 = n4703 ^ n240 ^ 1'b0 ;
  assign n4705 = ~n1122 & n4704 ;
  assign n4706 = n4705 ^ n1051 ^ 1'b0 ;
  assign n4707 = n4706 ^ n4240 ^ 1'b0 ;
  assign n4708 = n241 & n4707 ;
  assign n4709 = n2059 & n3726 ;
  assign n4710 = ~n757 & n4709 ;
  assign n4711 = ( n3544 & n4708 ) | ( n3544 & n4710 ) | ( n4708 & n4710 ) ;
  assign n4712 = n4344 ^ n3973 ^ n336 ;
  assign n4713 = n2505 ^ n1827 ^ 1'b0 ;
  assign n4714 = n3211 ^ n1225 ^ 1'b0 ;
  assign n4715 = n4260 & n4714 ;
  assign n4716 = n3398 ^ n2180 ^ 1'b0 ;
  assign n4717 = n3040 & n4716 ;
  assign n4718 = x6 & ~n2088 ;
  assign n4719 = n4718 ^ n2006 ^ 1'b0 ;
  assign n4720 = n2105 | n4719 ;
  assign n4721 = n4720 ^ n4528 ^ n2786 ;
  assign n4737 = n2910 ^ n2281 ^ 1'b0 ;
  assign n4735 = n361 & ~n2148 ;
  assign n4736 = ( ~n428 & n1341 ) | ( ~n428 & n4735 ) | ( n1341 & n4735 ) ;
  assign n4738 = n4737 ^ n4736 ^ 1'b0 ;
  assign n4739 = n4738 ^ n2587 ^ 1'b0 ;
  assign n4740 = n628 | n4739 ;
  assign n4741 = n4740 ^ n1849 ^ n159 ;
  assign n4722 = ~n1487 & n2343 ;
  assign n4723 = n2769 & n4722 ;
  assign n4727 = n998 | n1256 ;
  assign n4724 = n792 ^ n41 ^ 1'b0 ;
  assign n4725 = n2423 & n4724 ;
  assign n4726 = n1426 & ~n4725 ;
  assign n4728 = n4727 ^ n4726 ^ 1'b0 ;
  assign n4729 = n4434 & n4728 ;
  assign n4730 = n4729 ^ n664 ^ n37 ;
  assign n4731 = n3648 & ~n4730 ;
  assign n4732 = n4723 & n4731 ;
  assign n4733 = n2145 & n2177 ;
  assign n4734 = ~n4732 & n4733 ;
  assign n4742 = n4741 ^ n4734 ^ 1'b0 ;
  assign n4743 = n467 ^ n96 ^ 1'b0 ;
  assign n4744 = n3231 ^ n1093 ^ 1'b0 ;
  assign n4745 = n4743 & ~n4744 ;
  assign n4746 = n125 | n1267 ;
  assign n4747 = n2370 | n4746 ;
  assign n4748 = n2390 ^ n70 ^ 1'b0 ;
  assign n4749 = n656 | n4748 ;
  assign n4750 = n2104 ^ n285 ^ x0 ;
  assign n4751 = n4750 ^ n2094 ^ 1'b0 ;
  assign n4752 = ( n2286 & n2702 ) | ( n2286 & ~n4751 ) | ( n2702 & ~n4751 ) ;
  assign n4754 = n2040 ^ n1071 ^ n437 ;
  assign n4755 = n448 & ~n4754 ;
  assign n4756 = n1046 & n4755 ;
  assign n4757 = n4226 & ~n4756 ;
  assign n4753 = ~n2808 & n4545 ;
  assign n4758 = n4757 ^ n4753 ^ 1'b0 ;
  assign n4759 = n171 | n730 ;
  assign n4760 = n1218 | n4759 ;
  assign n4761 = ( n171 & n1276 ) | ( n171 & n1617 ) | ( n1276 & n1617 ) ;
  assign n4762 = n3201 | n4761 ;
  assign n4763 = n4760 | n4762 ;
  assign n4764 = ~n3702 & n4763 ;
  assign n4765 = n4764 ^ n3253 ^ 1'b0 ;
  assign n4766 = n4352 | n4765 ;
  assign n4767 = n2006 & ~n4766 ;
  assign n4768 = n729 | n3868 ;
  assign n4769 = ( n1095 & ~n4767 ) | ( n1095 & n4768 ) | ( ~n4767 & n4768 ) ;
  assign n4770 = n2720 ^ n184 ^ n151 ;
  assign n4771 = n631 | n2966 ;
  assign n4772 = n4272 | n4771 ;
  assign n4774 = n2373 ^ n172 ^ 1'b0 ;
  assign n4775 = n464 & n4774 ;
  assign n4776 = n3144 & n4775 ;
  assign n4777 = ~n2907 & n4776 ;
  assign n4778 = n4777 ^ n594 ^ 1'b0 ;
  assign n4773 = ( n1071 & ~n1286 ) | ( n1071 & n3207 ) | ( ~n1286 & n3207 ) ;
  assign n4779 = n4778 ^ n4773 ^ 1'b0 ;
  assign n4780 = n3971 | n4756 ;
  assign n4781 = n596 | n2840 ;
  assign n4785 = ( ~n309 & n383 ) | ( ~n309 & n469 ) | ( n383 & n469 ) ;
  assign n4782 = n55 & n1312 ;
  assign n4783 = n2464 & n4782 ;
  assign n4784 = n4783 ^ n1522 ^ 1'b0 ;
  assign n4786 = n4785 ^ n4784 ^ 1'b0 ;
  assign n4787 = n3176 ^ n1805 ^ 1'b0 ;
  assign n4788 = n3483 ^ n1079 ^ 1'b0 ;
  assign n4789 = ( n2568 & ~n3232 ) | ( n2568 & n4788 ) | ( ~n3232 & n4788 ) ;
  assign n4790 = n3140 ^ n461 ^ 1'b0 ;
  assign n4791 = n4789 | n4790 ;
  assign n4792 = n4787 & ~n4791 ;
  assign n4793 = ( n763 & n800 ) | ( n763 & ~n2089 ) | ( n800 & ~n2089 ) ;
  assign n4794 = n1786 & n4458 ;
  assign n4795 = n3395 | n4794 ;
  assign n4796 = n1084 ^ n600 ^ n383 ;
  assign n4797 = n4796 ^ n1666 ^ n1384 ;
  assign n4798 = n4797 ^ n2128 ^ 1'b0 ;
  assign n4799 = n1658 | n4798 ;
  assign n4801 = n4377 ^ n503 ^ 1'b0 ;
  assign n4800 = ~n1515 & n3148 ;
  assign n4802 = n4801 ^ n4800 ^ 1'b0 ;
  assign n4803 = ( n3089 & n4799 ) | ( n3089 & ~n4802 ) | ( n4799 & ~n4802 ) ;
  assign n4804 = ( n4793 & ~n4795 ) | ( n4793 & n4803 ) | ( ~n4795 & n4803 ) ;
  assign n4805 = n583 & ~n694 ;
  assign n4806 = ~n74 & n4805 ;
  assign n4807 = n4806 ^ n1611 ^ 1'b0 ;
  assign n4809 = n180 | n411 ;
  assign n4808 = n1190 | n3387 ;
  assign n4810 = n4809 ^ n4808 ^ 1'b0 ;
  assign n4811 = n23 & ~n686 ;
  assign n4812 = n4811 ^ n2084 ^ 1'b0 ;
  assign n4813 = n4812 ^ n51 ^ 1'b0 ;
  assign n4814 = n725 ^ n615 ^ 1'b0 ;
  assign n4815 = n4813 | n4814 ;
  assign n4816 = n293 | n961 ;
  assign n4817 = n4815 & ~n4816 ;
  assign n4818 = n1365 | n4743 ;
  assign n4819 = ( n1006 & n1436 ) | ( n1006 & n4818 ) | ( n1436 & n4818 ) ;
  assign n4821 = n4188 ^ n2716 ^ n437 ;
  assign n4822 = n4821 ^ n1961 ^ 1'b0 ;
  assign n4823 = ~n202 & n4822 ;
  assign n4824 = n4405 & n4823 ;
  assign n4825 = n4824 ^ n394 ^ 1'b0 ;
  assign n4820 = n77 & ~n3014 ;
  assign n4826 = n4825 ^ n4820 ^ 1'b0 ;
  assign n4827 = n132 | n2192 ;
  assign n4828 = n109 & n1791 ;
  assign n4829 = n4828 ^ n2123 ^ 1'b0 ;
  assign n4830 = ~n241 & n712 ;
  assign n4831 = n2551 & ~n4830 ;
  assign n4832 = ~n4829 & n4831 ;
  assign n4833 = n4053 & n4301 ;
  assign n4834 = n1905 & n4833 ;
  assign n4835 = n1103 | n1232 ;
  assign n4836 = n3714 ^ n374 ^ 1'b0 ;
  assign n4837 = ~n231 & n4836 ;
  assign n4838 = n4835 | n4837 ;
  assign n4839 = n818 | n1223 ;
  assign n4840 = n1178 | n4839 ;
  assign n4841 = n4840 ^ n1488 ^ n892 ;
  assign n4842 = ( n2419 & n4425 ) | ( n2419 & n4841 ) | ( n4425 & n4841 ) ;
  assign n4843 = n654 & ~n954 ;
  assign n4844 = n4843 ^ n269 ^ 1'b0 ;
  assign n4845 = n4844 ^ n4758 ^ 1'b0 ;
  assign n4846 = n2198 ^ n1047 ^ n585 ;
  assign n4847 = ~n2835 & n4846 ;
  assign n4848 = n237 & n738 ;
  assign n4849 = n4848 ^ n1279 ^ 1'b0 ;
  assign n4850 = n426 | n4849 ;
  assign n4851 = n4847 & ~n4850 ;
  assign n4852 = n3149 & ~n4801 ;
  assign n4853 = n4852 ^ n1282 ^ 1'b0 ;
  assign n4854 = n2062 & n4853 ;
  assign n4855 = n3512 ^ n2312 ^ 1'b0 ;
  assign n4856 = n4719 & n4855 ;
  assign n4857 = n1885 & n4050 ;
  assign n4858 = n1300 & n2319 ;
  assign n4859 = n4858 ^ n2231 ^ 1'b0 ;
  assign n4860 = n4859 ^ n506 ^ 1'b0 ;
  assign n4861 = n2604 ^ n1405 ^ n886 ;
  assign n4862 = ( n250 & n2019 ) | ( n250 & ~n4861 ) | ( n2019 & ~n4861 ) ;
  assign n4863 = n2602 & ~n4862 ;
  assign n4864 = ~n2764 & n3395 ;
  assign n4865 = ~n471 & n1400 ;
  assign n4866 = n4865 ^ n2466 ^ 1'b0 ;
  assign n4872 = n1231 & n2482 ;
  assign n4869 = ~n1263 & n3681 ;
  assign n4867 = n2250 ^ n1249 ^ n49 ;
  assign n4868 = n1878 & ~n4867 ;
  assign n4870 = n4869 ^ n4868 ^ 1'b0 ;
  assign n4871 = n1348 & ~n4870 ;
  assign n4873 = n4872 ^ n4871 ^ 1'b0 ;
  assign n4874 = n4866 & ~n4873 ;
  assign n4875 = n4874 ^ n744 ^ 1'b0 ;
  assign n4876 = n788 & n4573 ;
  assign n4877 = ~n1450 & n4876 ;
  assign n4878 = n1515 & ~n4877 ;
  assign n4879 = n1957 | n2044 ;
  assign n4880 = n4879 ^ n3541 ^ 1'b0 ;
  assign n4881 = n2806 ^ n1697 ^ 1'b0 ;
  assign n4882 = n336 & ~n4881 ;
  assign n4883 = ~n4880 & n4882 ;
  assign n4884 = n4883 ^ n995 ^ 1'b0 ;
  assign n4885 = n4368 ^ n1457 ^ 1'b0 ;
  assign n4886 = n4884 | n4885 ;
  assign n4889 = ~n255 & n2236 ;
  assign n4887 = n4502 ^ n813 ^ n648 ;
  assign n4888 = n4887 ^ n3221 ^ 1'b0 ;
  assign n4890 = n4889 ^ n4888 ^ 1'b0 ;
  assign n4891 = x1 & ~n563 ;
  assign n4892 = n4891 ^ n1773 ^ 1'b0 ;
  assign n4893 = n4890 | n4892 ;
  assign n4894 = n4893 ^ n263 ^ 1'b0 ;
  assign n4896 = n493 & n647 ;
  assign n4895 = n1357 & n1793 ;
  assign n4897 = n4896 ^ n4895 ^ 1'b0 ;
  assign n4898 = n4897 ^ n2815 ^ 1'b0 ;
  assign n4899 = n4743 & ~n4898 ;
  assign n4900 = n3981 ^ n113 ^ 1'b0 ;
  assign n4901 = n1302 ^ n42 ^ 1'b0 ;
  assign n4902 = n3475 ^ n3190 ^ 1'b0 ;
  assign n4903 = n4901 & n4902 ;
  assign n4904 = ~n1569 & n3868 ;
  assign n4905 = ~n627 & n1861 ;
  assign n4906 = n4905 ^ n3445 ^ 1'b0 ;
  assign n4907 = ~n902 & n2461 ;
  assign n4908 = ~n2243 & n4907 ;
  assign n4909 = n4402 ^ n2873 ^ 1'b0 ;
  assign n4910 = n1082 & n4909 ;
  assign n4911 = n4910 ^ n1681 ^ 1'b0 ;
  assign n4914 = n1140 ^ n33 ^ 1'b0 ;
  assign n4915 = n4914 ^ n3033 ^ n2636 ;
  assign n4912 = n242 | n1823 ;
  assign n4913 = n1726 | n4912 ;
  assign n4916 = n4915 ^ n4913 ^ 1'b0 ;
  assign n4917 = n1816 & ~n2070 ;
  assign n4918 = n4917 ^ n1100 ^ n794 ;
  assign n4920 = n1522 & ~n1754 ;
  assign n4921 = n4920 ^ n773 ^ 1'b0 ;
  assign n4922 = ~n2375 & n4921 ;
  assign n4919 = ~n1442 & n4810 ;
  assign n4923 = n4922 ^ n4919 ^ 1'b0 ;
  assign n4924 = ~n2695 & n4894 ;
  assign n4925 = n4924 ^ n2676 ^ 1'b0 ;
  assign n4926 = n1476 & ~n3973 ;
  assign n4927 = n4926 ^ n1294 ^ 1'b0 ;
  assign n4928 = ( n20 & ~n2986 ) | ( n20 & n4927 ) | ( ~n2986 & n4927 ) ;
  assign n4929 = ~n852 & n1145 ;
  assign n4930 = n3581 & n4929 ;
  assign n4931 = n4114 | n4930 ;
  assign n4932 = n394 & n2438 ;
  assign n4933 = ~n1171 & n4932 ;
  assign n4935 = n4563 ^ n3115 ^ 1'b0 ;
  assign n4936 = n1721 & ~n4935 ;
  assign n4934 = ~n373 & n2652 ;
  assign n4937 = n4936 ^ n4934 ^ 1'b0 ;
  assign n4938 = n4674 ^ n1376 ^ 1'b0 ;
  assign n4939 = n3326 & n4938 ;
  assign n4940 = n4736 ^ n2246 ^ 1'b0 ;
  assign n4941 = n28 | n4940 ;
  assign n4942 = n356 & n2939 ;
  assign n4943 = n3939 & n4942 ;
  assign n4944 = n4283 & n4943 ;
  assign n4945 = n2119 ^ n1235 ^ n332 ;
  assign n4946 = n3029 ^ n1453 ^ 1'b0 ;
  assign n4947 = n927 | n4946 ;
  assign n4948 = n4200 ^ n1641 ^ 1'b0 ;
  assign n4949 = ( n4488 & n4947 ) | ( n4488 & n4948 ) | ( n4947 & n4948 ) ;
  assign n4950 = n318 & ~n978 ;
  assign n4951 = n1066 & n4950 ;
  assign n4952 = n4951 ^ n3109 ^ 1'b0 ;
  assign n4953 = n577 & n4952 ;
  assign n4954 = ~n91 & n1288 ;
  assign n4955 = n4954 ^ n156 ^ 1'b0 ;
  assign n4956 = n2640 | n4955 ;
  assign n4957 = n4723 & ~n4956 ;
  assign n4958 = n4957 ^ n720 ^ 1'b0 ;
  assign n4959 = n2020 & n4958 ;
  assign n4960 = n4959 ^ n2123 ^ 1'b0 ;
  assign n4961 = n1185 | n4960 ;
  assign n4962 = n2705 ^ n2165 ^ 1'b0 ;
  assign n4963 = ~n1845 & n4962 ;
  assign n4964 = ~n3260 & n4963 ;
  assign n4965 = n1723 & n2488 ;
  assign n4966 = n620 & ~n628 ;
  assign n4967 = n575 & ~n4966 ;
  assign n4968 = n4673 ^ n1307 ^ n803 ;
  assign n4969 = x10 | n3093 ;
  assign n4970 = n4055 ^ n3486 ^ 1'b0 ;
  assign n4975 = n139 | n1931 ;
  assign n4973 = n538 | n1505 ;
  assign n4974 = n1216 | n4973 ;
  assign n4971 = n838 ^ n82 ^ 1'b0 ;
  assign n4972 = n37 & ~n4971 ;
  assign n4976 = n4975 ^ n4974 ^ n4972 ;
  assign n4977 = n4801 ^ n2714 ^ n1812 ;
  assign n4978 = ~n342 & n4325 ;
  assign n4979 = n136 & n340 ;
  assign n4980 = ~n4962 & n4979 ;
  assign n4981 = n2372 & n4913 ;
  assign n4982 = n4882 ^ n1175 ^ 1'b0 ;
  assign n4983 = n1075 & ~n4982 ;
  assign n4985 = n375 & n1280 ;
  assign n4984 = n2951 | n3005 ;
  assign n4986 = n4985 ^ n4984 ^ 1'b0 ;
  assign n4987 = n1368 | n3041 ;
  assign n4988 = n3033 & ~n3805 ;
  assign n4989 = ~n4987 & n4988 ;
  assign n4990 = n4986 & n4989 ;
  assign n4991 = n223 & n2214 ;
  assign n4992 = n4991 ^ n2209 ^ 1'b0 ;
  assign n4993 = n1746 ^ n1281 ^ 1'b0 ;
  assign n4994 = ( n63 & n448 ) | ( n63 & ~n848 ) | ( n448 & ~n848 ) ;
  assign n4995 = n4994 ^ n1424 ^ 1'b0 ;
  assign n4996 = n1459 & ~n4995 ;
  assign n4997 = ( ~n1133 & n4547 ) | ( ~n1133 & n4996 ) | ( n4547 & n4996 ) ;
  assign n4998 = n1253 & n4997 ;
  assign n4999 = n3076 ^ n108 ^ 1'b0 ;
  assign n5000 = n1777 ^ n534 ^ 1'b0 ;
  assign n5001 = n784 & ~n5000 ;
  assign n5002 = n3744 | n4240 ;
  assign n5003 = n5001 | n5002 ;
  assign n5004 = n5003 ^ n3541 ^ 1'b0 ;
  assign n5006 = n2460 ^ n1124 ^ 1'b0 ;
  assign n5005 = ~n499 & n4743 ;
  assign n5007 = n5006 ^ n5005 ^ 1'b0 ;
  assign n5008 = n1684 ^ n421 ^ 1'b0 ;
  assign n5009 = n5008 ^ n3188 ^ 1'b0 ;
  assign n5010 = n578 | n4390 ;
  assign n5011 = n5010 ^ n1311 ^ 1'b0 ;
  assign n5012 = ~n778 & n3123 ;
  assign n5013 = n5012 ^ n3505 ^ 1'b0 ;
  assign n5014 = n1934 ^ n1918 ^ 1'b0 ;
  assign n5015 = n4913 ^ n498 ^ 1'b0 ;
  assign n5016 = ~n966 & n5015 ;
  assign n5017 = n447 & ~n3897 ;
  assign n5018 = n5017 ^ n3709 ^ 1'b0 ;
  assign n5019 = n4226 ^ n1540 ^ 1'b0 ;
  assign n5020 = ~n261 & n5019 ;
  assign n5021 = n962 & n1167 ;
  assign n5022 = ~n5020 & n5021 ;
  assign n5023 = n23 | n5022 ;
  assign n5024 = n5023 ^ n2288 ^ 1'b0 ;
  assign n5025 = n453 ^ n420 ^ 1'b0 ;
  assign n5026 = n553 | n5025 ;
  assign n5027 = n1095 & ~n5026 ;
  assign n5028 = n5024 & n5027 ;
  assign n5029 = n5028 ^ n1317 ^ 1'b0 ;
  assign n5036 = n655 ^ n342 ^ n80 ;
  assign n5035 = n1272 & n3682 ;
  assign n5037 = n5036 ^ n5035 ^ 1'b0 ;
  assign n5031 = n532 & n1348 ;
  assign n5032 = n2604 & n5031 ;
  assign n5033 = n5032 ^ n2328 ^ n1876 ;
  assign n5034 = ~n3305 & n5033 ;
  assign n5038 = n5037 ^ n5034 ^ 1'b0 ;
  assign n5039 = n1332 & ~n5038 ;
  assign n5030 = n1116 | n1345 ;
  assign n5040 = n5039 ^ n5030 ^ 1'b0 ;
  assign n5041 = n4887 ^ n1179 ^ 1'b0 ;
  assign n5042 = ~n5024 & n5041 ;
  assign n5043 = n829 | n1010 ;
  assign n5044 = ~n2207 & n3314 ;
  assign n5045 = n3879 & ~n5044 ;
  assign n5046 = ~n500 & n696 ;
  assign n5047 = n5046 ^ n1775 ^ 1'b0 ;
  assign n5048 = n5047 ^ n4058 ^ 1'b0 ;
  assign n5049 = n4001 ^ n1960 ^ 1'b0 ;
  assign n5050 = n1000 | n5049 ;
  assign n5051 = n5050 ^ n3392 ^ n2172 ;
  assign n5052 = n490 ^ n362 ^ 1'b0 ;
  assign n5053 = n203 & ~n2776 ;
  assign n5054 = n5052 | n5053 ;
  assign n5055 = n5054 ^ n3984 ^ n1424 ;
  assign n5056 = ~n4794 & n5055 ;
  assign n5057 = n4239 & n5056 ;
  assign n5058 = ( n267 & n1907 ) | ( n267 & ~n4972 ) | ( n1907 & ~n4972 ) ;
  assign n5059 = ( n341 & n866 ) | ( n341 & n2431 ) | ( n866 & n2431 ) ;
  assign n5060 = n5059 ^ n1213 ^ 1'b0 ;
  assign n5061 = n2412 & n5060 ;
  assign n5062 = n5061 ^ n850 ^ 1'b0 ;
  assign n5063 = n4699 & ~n5062 ;
  assign n5064 = ~n281 & n5063 ;
  assign n5065 = n5064 ^ n5053 ^ 1'b0 ;
  assign n5066 = ~n3700 & n5065 ;
  assign n5070 = ( n102 & n344 ) | ( n102 & ~n790 ) | ( n344 & ~n790 ) ;
  assign n5068 = ( n2072 & n2423 ) | ( n2072 & n3306 ) | ( n2423 & n3306 ) ;
  assign n5067 = n782 & ~n4118 ;
  assign n5069 = n5068 ^ n5067 ^ 1'b0 ;
  assign n5071 = n5070 ^ n5069 ^ 1'b0 ;
  assign n5072 = n5066 & n5071 ;
  assign n5073 = n5072 ^ n3308 ^ 1'b0 ;
  assign n5078 = n4584 ^ n3785 ^ n944 ;
  assign n5079 = n900 ^ n448 ^ 1'b0 ;
  assign n5080 = ~n5078 & n5079 ;
  assign n5074 = n3142 ^ n993 ^ 1'b0 ;
  assign n5075 = n5074 ^ n3354 ^ 1'b0 ;
  assign n5076 = n2885 & ~n5075 ;
  assign n5077 = ~n2445 & n5076 ;
  assign n5081 = n5080 ^ n5077 ^ 1'b0 ;
  assign n5082 = n953 & n5081 ;
  assign n5083 = n1071 ^ n98 ^ 1'b0 ;
  assign n5084 = n5083 ^ n994 ^ 1'b0 ;
  assign n5085 = n2944 ^ n790 ^ n571 ;
  assign n5086 = n5085 ^ n2209 ^ n1808 ;
  assign n5087 = n1320 ^ n35 ^ 1'b0 ;
  assign n5088 = n1484 & n5087 ;
  assign n5089 = ( n291 & n5086 ) | ( n291 & n5088 ) | ( n5086 & n5088 ) ;
  assign n5090 = n2169 ^ n1114 ^ 1'b0 ;
  assign n5091 = ( n33 & ~n137 ) | ( n33 & n5090 ) | ( ~n137 & n5090 ) ;
  assign n5094 = n1453 ^ n1370 ^ 1'b0 ;
  assign n5095 = n5094 ^ n3098 ^ n43 ;
  assign n5092 = n63 & n1037 ;
  assign n5093 = ~n4180 & n5092 ;
  assign n5096 = n5095 ^ n5093 ^ 1'b0 ;
  assign n5097 = n3394 | n5096 ;
  assign n5098 = n609 | n4333 ;
  assign n5099 = ~n3156 & n4399 ;
  assign n5100 = n2060 & n5099 ;
  assign n5101 = ~n5098 & n5100 ;
  assign n5102 = n3581 ^ n1518 ^ 1'b0 ;
  assign n5103 = n727 ^ n707 ^ 1'b0 ;
  assign n5104 = n2896 | n5103 ;
  assign n5105 = n5104 ^ n2178 ^ 1'b0 ;
  assign n5106 = n5102 & n5105 ;
  assign n5107 = n3858 ^ n145 ^ 1'b0 ;
  assign n5108 = n5106 & ~n5107 ;
  assign n5109 = n2423 ^ n1824 ^ n1167 ;
  assign n5110 = n723 ^ n448 ^ 1'b0 ;
  assign n5111 = ~n521 & n2588 ;
  assign n5112 = n1943 | n5111 ;
  assign n5113 = ( n631 & ~n1122 ) | ( n631 & n2949 ) | ( ~n1122 & n2949 ) ;
  assign n5114 = n305 | n2245 ;
  assign n5115 = n3193 & n5114 ;
  assign n5116 = ~n804 & n1632 ;
  assign n5117 = n5116 ^ n1943 ^ 1'b0 ;
  assign n5118 = ~n4488 & n5117 ;
  assign n5119 = ( n2736 & n5115 ) | ( n2736 & ~n5118 ) | ( n5115 & ~n5118 ) ;
  assign n5120 = ~n1848 & n4071 ;
  assign n5121 = n2849 & n3205 ;
  assign n5122 = n5121 ^ n4834 ^ 1'b0 ;
  assign n5123 = n2529 ^ n1748 ^ n756 ;
  assign n5124 = n5123 ^ n4324 ^ 1'b0 ;
  assign n5125 = n1095 ^ n108 ^ 1'b0 ;
  assign n5126 = n1684 & ~n5125 ;
  assign n5127 = n3759 & n5126 ;
  assign n5130 = n2679 ^ n1176 ^ 1'b0 ;
  assign n5128 = n902 ^ n736 ^ 1'b0 ;
  assign n5129 = n5128 ^ n929 ^ 1'b0 ;
  assign n5131 = n5130 ^ n5129 ^ 1'b0 ;
  assign n5132 = ( ~n145 & n1762 ) | ( ~n145 & n2494 ) | ( n1762 & n2494 ) ;
  assign n5133 = n5132 ^ n4019 ^ 1'b0 ;
  assign n5134 = n4859 | n5133 ;
  assign n5135 = n5134 ^ n1838 ^ 1'b0 ;
  assign n5136 = n1181 & ~n2735 ;
  assign n5137 = ( ~x10 & n1273 ) | ( ~x10 & n3108 ) | ( n1273 & n3108 ) ;
  assign n5138 = n3157 ^ n1665 ^ 1'b0 ;
  assign n5139 = n5137 | n5138 ;
  assign n5140 = n3151 | n5139 ;
  assign n5141 = n99 & ~n2422 ;
  assign n5142 = n2165 & n5141 ;
  assign n5143 = ( n612 & ~n826 ) | ( n612 & n5142 ) | ( ~n826 & n5142 ) ;
  assign n5144 = ( n805 & n1614 ) | ( n805 & ~n5143 ) | ( n1614 & ~n5143 ) ;
  assign n5146 = n5107 ^ n1225 ^ 1'b0 ;
  assign n5145 = n3370 ^ n3038 ^ n3030 ;
  assign n5147 = n5146 ^ n5145 ^ 1'b0 ;
  assign n5148 = n2684 ^ n263 ^ 1'b0 ;
  assign n5149 = n797 & ~n5148 ;
  assign n5150 = ( n2432 & n2511 ) | ( n2432 & ~n5149 ) | ( n2511 & ~n5149 ) ;
  assign n5151 = n4523 ^ n3057 ^ 1'b0 ;
  assign n5152 = n5151 ^ n226 ^ 1'b0 ;
  assign n5153 = n5150 | n5152 ;
  assign n5154 = n645 & ~n908 ;
  assign n5155 = n5154 ^ n1918 ^ 1'b0 ;
  assign n5156 = n5155 ^ n2382 ^ 1'b0 ;
  assign n5157 = n5156 ^ n1826 ^ n734 ;
  assign n5159 = n1613 & ~n1630 ;
  assign n5158 = n2423 | n3116 ;
  assign n5160 = n5159 ^ n5158 ^ 1'b0 ;
  assign n5161 = n1522 & n5160 ;
  assign n5162 = n1915 ^ n298 ^ 1'b0 ;
  assign n5163 = n772 | n933 ;
  assign n5164 = n5162 & ~n5163 ;
  assign n5165 = n3579 | n5164 ;
  assign n5166 = ( n3106 & n4303 ) | ( n3106 & ~n4533 ) | ( n4303 & ~n4533 ) ;
  assign n5167 = n2327 ^ n795 ^ 1'b0 ;
  assign n5168 = n1285 & n5167 ;
  assign n5172 = n1538 ^ n1526 ^ n706 ;
  assign n5173 = n5172 ^ n37 ^ 1'b0 ;
  assign n5169 = n3125 ^ n2339 ^ n147 ;
  assign n5170 = n4300 | n5169 ;
  assign n5171 = n105 | n5170 ;
  assign n5174 = n5173 ^ n5171 ^ n2181 ;
  assign n5175 = n5168 & n5174 ;
  assign n5176 = n1623 ^ n181 ^ 1'b0 ;
  assign n5177 = n32 | n3037 ;
  assign n5178 = n299 & ~n5177 ;
  assign n5179 = n2844 ^ n2489 ^ n2408 ;
  assign n5180 = n5179 ^ n4675 ^ 1'b0 ;
  assign n5181 = n780 & n1554 ;
  assign n5182 = n5181 ^ n265 ^ 1'b0 ;
  assign n5183 = n2913 ^ n1812 ^ n126 ;
  assign n5184 = ~n2928 & n5183 ;
  assign n5185 = ~n4405 & n5184 ;
  assign n5186 = ( ~n947 & n3429 ) | ( ~n947 & n5185 ) | ( n3429 & n5185 ) ;
  assign n5187 = n3874 & n4897 ;
  assign n5188 = n5187 ^ n1079 ^ 1'b0 ;
  assign n5189 = n2571 ^ x3 ^ 1'b0 ;
  assign n5190 = n84 | n1104 ;
  assign n5191 = n1931 | n5190 ;
  assign n5192 = n1623 & n5191 ;
  assign n5193 = ~n100 & n5192 ;
  assign n5194 = n5193 ^ n2897 ^ 1'b0 ;
  assign n5195 = n3175 & n5194 ;
  assign n5196 = ~n601 & n5195 ;
  assign n5197 = ~n2570 & n5196 ;
  assign n5198 = n1793 | n5197 ;
  assign n5199 = n5198 ^ n1840 ^ 1'b0 ;
  assign n5200 = n3636 ^ n2650 ^ 1'b0 ;
  assign n5202 = ( n2198 & ~n3359 ) | ( n2198 & n4552 ) | ( ~n3359 & n4552 ) ;
  assign n5201 = n141 & ~n2869 ;
  assign n5203 = n5202 ^ n5201 ^ 1'b0 ;
  assign n5204 = n2277 & ~n5203 ;
  assign n5205 = n1496 & ~n1533 ;
  assign n5206 = ( n695 & ~n2405 ) | ( n695 & n5205 ) | ( ~n2405 & n5205 ) ;
  assign n5207 = n4406 ^ n105 ^ 1'b0 ;
  assign n5208 = n1122 ^ n236 ^ 1'b0 ;
  assign n5209 = n3127 | n5208 ;
  assign n5210 = n5209 ^ n1155 ^ 1'b0 ;
  assign n5211 = n2073 ^ n1393 ^ 1'b0 ;
  assign n5212 = n1450 & ~n5211 ;
  assign n5213 = n3024 & n5212 ;
  assign n5214 = ~n5210 & n5213 ;
  assign n5219 = n35 & n279 ;
  assign n5216 = n3652 ^ n1843 ^ 1'b0 ;
  assign n5217 = n4848 & n5216 ;
  assign n5215 = n28 | n2034 ;
  assign n5218 = n5217 ^ n5215 ^ 1'b0 ;
  assign n5220 = n5219 ^ n5218 ^ 1'b0 ;
  assign n5221 = n154 & ~n1255 ;
  assign n5222 = n5221 ^ n5163 ^ 1'b0 ;
  assign n5223 = n5222 ^ n197 ^ 1'b0 ;
  assign n5224 = ~n3048 & n5223 ;
  assign n5225 = ~n105 & n794 ;
  assign n5226 = n4012 | n5044 ;
  assign n5227 = n214 & ~n5226 ;
  assign n5228 = ~n1848 & n5227 ;
  assign n5229 = ( n1038 & ~n2604 ) | ( n1038 & n4956 ) | ( ~n2604 & n4956 ) ;
  assign n5230 = n5229 ^ n1940 ^ 1'b0 ;
  assign n5231 = ~n1024 & n5230 ;
  assign n5232 = ~n620 & n5231 ;
  assign n5233 = n5232 ^ n534 ^ 1'b0 ;
  assign n5234 = n5233 ^ n626 ^ 1'b0 ;
  assign n5235 = ~n44 & n1457 ;
  assign n5236 = ~n5234 & n5235 ;
  assign n5237 = n5236 ^ n3120 ^ 1'b0 ;
  assign n5239 = n500 & ~n839 ;
  assign n5238 = ~n2664 & n2993 ;
  assign n5240 = n5239 ^ n5238 ^ 1'b0 ;
  assign n5241 = n1238 & n1262 ;
  assign n5242 = ( n2194 & n2217 ) | ( n2194 & ~n5241 ) | ( n2217 & ~n5241 ) ;
  assign n5243 = n490 & ~n2631 ;
  assign n5244 = n5243 ^ n2696 ^ 1'b0 ;
  assign n5245 = n1244 ^ n886 ^ 1'b0 ;
  assign n5246 = n2977 & ~n5245 ;
  assign n5247 = n5246 ^ n3833 ^ n2557 ;
  assign n5248 = n191 | n3676 ;
  assign n5249 = n5248 ^ n72 ^ 1'b0 ;
  assign n5250 = n4779 & n5249 ;
  assign n5251 = n2325 ^ n984 ^ 1'b0 ;
  assign n5252 = n4706 & n5251 ;
  assign n5253 = ( ~n953 & n1089 ) | ( ~n953 & n2025 ) | ( n1089 & n2025 ) ;
  assign n5254 = n2360 ^ n572 ^ 1'b0 ;
  assign n5255 = n3362 ^ n1202 ^ n176 ;
  assign n5256 = n4110 ^ n3030 ^ 1'b0 ;
  assign n5257 = n1612 & ~n5256 ;
  assign n5258 = n5257 ^ n3961 ^ 1'b0 ;
  assign n5259 = n5083 ^ n141 ^ 1'b0 ;
  assign n5260 = n2793 | n5259 ;
  assign n5261 = n5260 ^ n221 ^ 1'b0 ;
  assign n5262 = ( ~n2262 & n4614 ) | ( ~n2262 & n5261 ) | ( n4614 & n5261 ) ;
  assign n5267 = n1264 & n4399 ;
  assign n5268 = n2309 & n5267 ;
  assign n5269 = n2552 | n5268 ;
  assign n5263 = n3737 ^ n3375 ^ n2944 ;
  assign n5264 = n5263 ^ n3969 ^ 1'b0 ;
  assign n5265 = ( ~n105 & n2326 ) | ( ~n105 & n3009 ) | ( n2326 & n3009 ) ;
  assign n5266 = ~n5264 & n5265 ;
  assign n5270 = n5269 ^ n5266 ^ 1'b0 ;
  assign n5271 = n3154 ^ n150 ^ 1'b0 ;
  assign n5272 = n4330 & n5271 ;
  assign n5273 = n3304 & n5047 ;
  assign n5274 = ( n2422 & ~n4795 ) | ( n2422 & n5273 ) | ( ~n4795 & n5273 ) ;
  assign n5275 = n1848 ^ n933 ^ 1'b0 ;
  assign n5276 = n2176 & ~n5275 ;
  assign n5277 = ~n223 & n5276 ;
  assign n5278 = n3382 ^ n3193 ^ 1'b0 ;
  assign n5279 = ~n1787 & n5278 ;
  assign n5280 = n4382 ^ n3284 ^ n2294 ;
  assign n5283 = ~n177 & n2618 ;
  assign n5284 = n5283 ^ n40 ^ 1'b0 ;
  assign n5285 = ~n2918 & n5284 ;
  assign n5281 = n2708 & n3260 ;
  assign n5282 = n5281 ^ n2845 ^ 1'b0 ;
  assign n5286 = n5285 ^ n5282 ^ 1'b0 ;
  assign n5287 = n5061 ^ n619 ^ 1'b0 ;
  assign n5288 = n498 & n3486 ;
  assign n5289 = n5288 ^ n100 ^ 1'b0 ;
  assign n5290 = n5289 ^ n2886 ^ 1'b0 ;
  assign n5291 = n409 & ~n5290 ;
  assign n5292 = n5291 ^ n4120 ^ 1'b0 ;
  assign n5293 = n3343 | n5292 ;
  assign n5294 = n4088 & ~n5293 ;
  assign n5295 = n1940 & ~n5294 ;
  assign n5296 = n5295 ^ n4016 ^ 1'b0 ;
  assign n5297 = n3128 & n5296 ;
  assign n5298 = n637 & n5297 ;
  assign n5300 = ( ~n124 & n1856 ) | ( ~n124 & n2778 ) | ( n1856 & n2778 ) ;
  assign n5299 = n1124 & n2378 ;
  assign n5301 = n5300 ^ n5299 ^ 1'b0 ;
  assign n5302 = n5301 ^ n2951 ^ 1'b0 ;
  assign n5303 = n5302 ^ n848 ^ 1'b0 ;
  assign n5304 = n1746 | n5303 ;
  assign n5305 = ( n1959 & n3069 ) | ( n1959 & n3904 ) | ( n3069 & n3904 ) ;
  assign n5306 = n5305 ^ n3123 ^ 1'b0 ;
  assign n5307 = ~n3737 & n5306 ;
  assign n5308 = n102 | n1081 ;
  assign n5309 = n637 & ~n5308 ;
  assign n5310 = n3059 & n3410 ;
  assign n5311 = ~n141 & n4694 ;
  assign n5312 = n1815 & ~n3408 ;
  assign n5317 = n1468 & ~n3698 ;
  assign n5318 = ~n2030 & n5317 ;
  assign n5314 = n3181 ^ n1723 ^ n1462 ;
  assign n5313 = ( n644 & n1630 ) | ( n644 & n3676 ) | ( n1630 & n3676 ) ;
  assign n5315 = n5314 ^ n5313 ^ 1'b0 ;
  assign n5316 = n5315 ^ n319 ^ 1'b0 ;
  assign n5319 = n5318 ^ n5316 ^ 1'b0 ;
  assign n5320 = n1967 & n5319 ;
  assign n5321 = n3506 & ~n5320 ;
  assign n5322 = n5066 ^ n2545 ^ n395 ;
  assign n5323 = n3019 ^ n824 ^ 1'b0 ;
  assign n5324 = n5323 ^ n2459 ^ 1'b0 ;
  assign n5325 = n1247 ^ n524 ^ 1'b0 ;
  assign n5326 = n3361 ^ n1521 ^ 1'b0 ;
  assign n5327 = n3375 | n5326 ;
  assign n5328 = n1880 & ~n5327 ;
  assign n5329 = ~n5325 & n5328 ;
  assign n5330 = n2065 ^ n1448 ^ 1'b0 ;
  assign n5331 = ~n3597 & n5330 ;
  assign n5332 = n4643 ^ n1959 ^ 1'b0 ;
  assign n5333 = ~n1980 & n5332 ;
  assign n5334 = n1360 | n1403 ;
  assign n5335 = n4733 | n5334 ;
  assign n5336 = n150 & n5335 ;
  assign n5337 = n4338 & n5336 ;
  assign n5338 = n2045 ^ n1789 ^ 1'b0 ;
  assign n5339 = ~n243 & n714 ;
  assign n5340 = n5338 & ~n5339 ;
  assign n5341 = n2769 & n5340 ;
  assign n5342 = n2335 ^ n2110 ^ 1'b0 ;
  assign n5343 = n4827 ^ n1378 ^ 1'b0 ;
  assign n5344 = n5333 & n5343 ;
  assign n5345 = n3786 ^ n527 ^ 1'b0 ;
  assign n5346 = ~n1779 & n5345 ;
  assign n5347 = n3687 ^ n226 ^ 1'b0 ;
  assign n5348 = n1781 & ~n5347 ;
  assign n5349 = n1298 ^ n63 ^ 1'b0 ;
  assign n5350 = n23 & n5349 ;
  assign n5351 = x3 & ~n484 ;
  assign n5352 = n518 | n5351 ;
  assign n5353 = n5350 & n5352 ;
  assign n5354 = n5348 & n5353 ;
  assign n5355 = n5354 ^ n1318 ^ 1'b0 ;
  assign n5356 = n201 & ~n4383 ;
  assign n5357 = n1679 & n2808 ;
  assign n5358 = n202 | n372 ;
  assign n5359 = n5358 ^ n2623 ^ 1'b0 ;
  assign n5360 = n5359 ^ n1329 ^ 1'b0 ;
  assign n5361 = n4042 & n5360 ;
  assign n5362 = n2113 ^ n249 ^ 1'b0 ;
  assign n5363 = ~n3343 & n5362 ;
  assign n5364 = n4847 | n5363 ;
  assign n5365 = n4462 ^ n1746 ^ n190 ;
  assign n5366 = n2791 ^ n515 ^ 1'b0 ;
  assign n5367 = n4071 ^ n876 ^ 1'b0 ;
  assign n5368 = n2686 & ~n5367 ;
  assign n5369 = n4357 & ~n5290 ;
  assign n5370 = n1425 & n5369 ;
  assign n5371 = n1890 & ~n5370 ;
  assign n5372 = n5371 ^ n2848 ^ 1'b0 ;
  assign n5373 = n4725 ^ n3006 ^ n2495 ;
  assign n5374 = n3651 | n5373 ;
  assign n5375 = n208 ^ n98 ^ 1'b0 ;
  assign n5376 = n4804 & n5375 ;
  assign n5377 = n3663 ^ n3526 ^ n3368 ;
  assign n5378 = n1184 & ~n5377 ;
  assign n5379 = n771 & n2524 ;
  assign n5380 = n5379 ^ n491 ^ 1'b0 ;
  assign n5381 = n4674 & ~n5380 ;
  assign n5382 = n2469 ^ n1232 ^ 1'b0 ;
  assign n5383 = n3699 ^ n3467 ^ 1'b0 ;
  assign n5384 = n5382 | n5383 ;
  assign n5385 = n1156 & n1822 ;
  assign n5386 = n5385 ^ n719 ^ 1'b0 ;
  assign n5387 = n1525 & ~n2107 ;
  assign n5388 = n3983 ^ n2055 ^ 1'b0 ;
  assign n5389 = n1365 | n1706 ;
  assign n5390 = n5388 & n5389 ;
  assign n5391 = n5387 & n5390 ;
  assign n5392 = n41 & ~n1896 ;
  assign n5393 = ~n1290 & n2412 ;
  assign n5394 = n2048 & n5393 ;
  assign n5395 = n1926 ^ n231 ^ x6 ;
  assign n5396 = n2303 | n5395 ;
  assign n5397 = ( n100 & n1527 ) | ( n100 & ~n2032 ) | ( n1527 & ~n2032 ) ;
  assign n5398 = n5397 ^ n2017 ^ 1'b0 ;
  assign n5399 = n4945 & n5398 ;
  assign n5400 = n505 & n3633 ;
  assign n5401 = n5400 ^ n4941 ^ 1'b0 ;
  assign n5402 = n2672 | n5401 ;
  assign n5413 = n97 | n1095 ;
  assign n5414 = n603 & ~n5413 ;
  assign n5408 = n1560 | n2857 ;
  assign n5409 = n2229 & n5212 ;
  assign n5410 = n2128 & n5409 ;
  assign n5411 = n5408 & ~n5410 ;
  assign n5412 = n5411 ^ n2296 ^ 1'b0 ;
  assign n5415 = n5414 ^ n5412 ^ n1336 ;
  assign n5416 = n2797 | n5415 ;
  assign n5403 = n2917 & n3187 ;
  assign n5404 = n5403 ^ n2807 ^ 1'b0 ;
  assign n5405 = n2794 ^ n2583 ^ 1'b0 ;
  assign n5406 = n5404 & ~n5405 ;
  assign n5407 = ~n2609 & n5406 ;
  assign n5417 = n5416 ^ n5407 ^ 1'b0 ;
  assign n5418 = n1468 ^ n118 ^ 1'b0 ;
  assign n5419 = n341 & n2374 ;
  assign n5420 = ( n5338 & n5418 ) | ( n5338 & n5419 ) | ( n5418 & n5419 ) ;
  assign n5421 = n5420 ^ n1015 ^ 1'b0 ;
  assign n5426 = n2117 | n3059 ;
  assign n5427 = n875 & ~n5426 ;
  assign n5424 = n450 & ~n1645 ;
  assign n5422 = n1324 | n2854 ;
  assign n5423 = n3541 & ~n5422 ;
  assign n5425 = n5424 ^ n5423 ^ 1'b0 ;
  assign n5428 = n5427 ^ n5425 ^ 1'b0 ;
  assign n5429 = n5428 ^ n4308 ^ 1'b0 ;
  assign n5430 = n4773 | n5429 ;
  assign n5431 = n91 | n1691 ;
  assign n5432 = n1490 | n5431 ;
  assign n5433 = n2541 & ~n5432 ;
  assign n5434 = ~n2268 & n3466 ;
  assign n5435 = n5434 ^ n149 ^ 1'b0 ;
  assign n5436 = n276 & n455 ;
  assign n5437 = n3295 ^ n448 ^ 1'b0 ;
  assign n5438 = n998 & ~n2858 ;
  assign n5439 = ~n2213 & n5438 ;
  assign n5440 = n5439 ^ n2646 ^ 1'b0 ;
  assign n5441 = ( n1490 & n3168 ) | ( n1490 & ~n3704 ) | ( n3168 & ~n3704 ) ;
  assign n5442 = ( ~n3330 & n4516 ) | ( ~n3330 & n5441 ) | ( n4516 & n5441 ) ;
  assign n5443 = n2810 ^ n2484 ^ 1'b0 ;
  assign n5444 = n3406 ^ n1240 ^ 1'b0 ;
  assign n5445 = n5444 ^ n780 ^ 1'b0 ;
  assign n5446 = ~n5443 & n5445 ;
  assign n5447 = n154 & ~n2090 ;
  assign n5448 = n995 & ~n5447 ;
  assign n5449 = n5448 ^ n4626 ^ 1'b0 ;
  assign n5450 = ( n354 & ~n1942 ) | ( n354 & n5449 ) | ( ~n1942 & n5449 ) ;
  assign n5451 = n5450 ^ n1064 ^ 1'b0 ;
  assign n5452 = ~n1403 & n2507 ;
  assign n5453 = n91 & n5452 ;
  assign n5454 = n5453 ^ n1562 ^ 1'b0 ;
  assign n5455 = n5451 & ~n5454 ;
  assign n5456 = n5455 ^ n4862 ^ n3843 ;
  assign n5457 = ~n4359 & n5456 ;
  assign n5459 = n5408 ^ n1024 ^ 1'b0 ;
  assign n5458 = n2486 ^ n2160 ^ 1'b0 ;
  assign n5460 = n5459 ^ n5458 ^ 1'b0 ;
  assign n5461 = ~n5457 & n5460 ;
  assign n5462 = n291 & ~n3184 ;
  assign n5463 = n5462 ^ n1472 ^ 1'b0 ;
  assign n5464 = n3115 & ~n5463 ;
  assign n5466 = n1115 ^ n954 ^ 1'b0 ;
  assign n5465 = n1311 ^ n1029 ^ 1'b0 ;
  assign n5467 = n5466 ^ n5465 ^ 1'b0 ;
  assign n5468 = n5464 & n5467 ;
  assign n5469 = ~n2616 & n5397 ;
  assign n5470 = n2561 ^ n951 ^ 1'b0 ;
  assign n5477 = n1153 ^ n105 ^ 1'b0 ;
  assign n5471 = n417 & n1140 ;
  assign n5472 = ~n214 & n5471 ;
  assign n5473 = n5472 ^ n1910 ^ 1'b0 ;
  assign n5474 = ~n3540 & n5473 ;
  assign n5475 = ~n656 & n5474 ;
  assign n5476 = n3774 | n5475 ;
  assign n5478 = n5477 ^ n5476 ^ 1'b0 ;
  assign n5479 = n5470 | n5478 ;
  assign n5480 = n1332 | n2583 ;
  assign n5481 = n4181 | n5480 ;
  assign n5483 = n443 & n962 ;
  assign n5484 = n5483 ^ n186 ^ 1'b0 ;
  assign n5485 = n5484 ^ n1506 ^ 1'b0 ;
  assign n5482 = n1605 ^ n1572 ^ 1'b0 ;
  assign n5486 = n5485 ^ n5482 ^ n3608 ;
  assign n5487 = n334 & ~n376 ;
  assign n5488 = n5487 ^ n3098 ^ 1'b0 ;
  assign n5489 = n5488 ^ n2427 ^ 1'b0 ;
  assign n5490 = ~n3603 & n5489 ;
  assign n5491 = ~n1295 & n5490 ;
  assign n5492 = n897 ^ n854 ^ 1'b0 ;
  assign n5493 = ~n2634 & n5492 ;
  assign n5494 = n4214 ^ n3496 ^ 1'b0 ;
  assign n5495 = n5494 ^ n3926 ^ 1'b0 ;
  assign n5496 = ~n1362 & n2810 ;
  assign n5497 = ~n250 & n4678 ;
  assign n5498 = n5496 & n5497 ;
  assign n5499 = n2322 ^ n2246 ^ 1'b0 ;
  assign n5500 = n3372 & n5499 ;
  assign n5501 = n5500 ^ n709 ^ 1'b0 ;
  assign n5502 = n1728 | n3240 ;
  assign n5503 = n1348 & n5502 ;
  assign n5504 = n5503 ^ n3948 ^ 1'b0 ;
  assign n5505 = n4432 & n5504 ;
  assign n5506 = n5501 & n5505 ;
  assign n5507 = n4196 ^ n1695 ^ n1694 ;
  assign n5508 = ( n1665 & n2139 ) | ( n1665 & n5507 ) | ( n2139 & n5507 ) ;
  assign n5509 = n63 & ~n2828 ;
  assign n5510 = n2067 ^ n541 ^ 1'b0 ;
  assign n5511 = n63 | n5510 ;
  assign n5512 = ( n2896 & ~n5509 ) | ( n2896 & n5511 ) | ( ~n5509 & n5511 ) ;
  assign n5513 = n1766 | n2312 ;
  assign n5514 = n186 ^ n73 ^ 1'b0 ;
  assign n5515 = n1503 | n5514 ;
  assign n5516 = n1693 | n5515 ;
  assign n5517 = n5516 ^ n547 ^ 1'b0 ;
  assign n5518 = n1079 & ~n4149 ;
  assign n5519 = n5517 & n5518 ;
  assign n5520 = n1805 | n2783 ;
  assign n5521 = n1213 & ~n5520 ;
  assign n5522 = n2811 ^ n1869 ^ n1500 ;
  assign n5523 = n358 & n5522 ;
  assign n5524 = ~n1149 & n5523 ;
  assign n5525 = n4799 | n5524 ;
  assign n5526 = n5525 ^ n3964 ^ 1'b0 ;
  assign n5527 = ( n109 & ~n152 ) | ( n109 & n5526 ) | ( ~n152 & n5526 ) ;
  assign n5528 = n5521 & n5527 ;
  assign n5529 = n5519 & n5528 ;
  assign n5530 = n804 | n5529 ;
  assign n5531 = n3495 | n5530 ;
  assign n5532 = ~n802 & n5531 ;
  assign n5533 = n5532 ^ n1647 ^ 1'b0 ;
  assign n5534 = n5222 ^ n4272 ^ 1'b0 ;
  assign n5535 = n2296 & ~n2954 ;
  assign n5536 = n902 | n5535 ;
  assign n5537 = ~n1427 & n3651 ;
  assign n5538 = ~n2090 & n2844 ;
  assign n5539 = n5537 & ~n5538 ;
  assign n5540 = ~n1560 & n5539 ;
  assign n5548 = n2698 ^ n965 ^ 1'b0 ;
  assign n5549 = n609 & n5548 ;
  assign n5545 = ( n2542 & n3084 ) | ( n2542 & n3940 ) | ( n3084 & n3940 ) ;
  assign n5541 = n583 | n849 ;
  assign n5542 = n2909 ^ n2657 ^ n733 ;
  assign n5543 = n5542 ^ n455 ^ 1'b0 ;
  assign n5544 = ~n5541 & n5543 ;
  assign n5546 = n5545 ^ n5544 ^ 1'b0 ;
  assign n5547 = ~n2451 & n5546 ;
  assign n5550 = n5549 ^ n5547 ^ 1'b0 ;
  assign n5551 = n48 & n5388 ;
  assign n5552 = n5551 ^ n713 ^ n709 ;
  assign n5553 = ~n32 & n1800 ;
  assign n5554 = n5553 ^ n824 ^ 1'b0 ;
  assign n5555 = ~n4280 & n5554 ;
  assign n5556 = ~n2826 & n5555 ;
  assign n5557 = n296 & n1629 ;
  assign n5558 = n5557 ^ n1634 ^ 1'b0 ;
  assign n5559 = n1011 & n5558 ;
  assign n5560 = n5559 ^ n1812 ^ 1'b0 ;
  assign n5561 = ~n1080 & n5560 ;
  assign n5562 = ~n4223 & n5561 ;
  assign n5563 = n98 & ~n2055 ;
  assign n5564 = ( n949 & n2597 ) | ( n949 & n5561 ) | ( n2597 & n5561 ) ;
  assign n5565 = ( n1387 & ~n2630 ) | ( n1387 & n3614 ) | ( ~n2630 & n3614 ) ;
  assign n5566 = ~n829 & n1400 ;
  assign n5567 = n5566 ^ n2785 ^ 1'b0 ;
  assign n5568 = n5565 & n5567 ;
  assign n5569 = n2989 ^ n984 ^ 1'b0 ;
  assign n5570 = n5569 ^ n3922 ^ n358 ;
  assign n5571 = n557 & n1350 ;
  assign n5572 = n2413 & ~n5502 ;
  assign n5573 = n5572 ^ n3162 ^ n2954 ;
  assign n5574 = ( n1320 & ~n3373 ) | ( n1320 & n3824 ) | ( ~n3373 & n3824 ) ;
  assign n5575 = n929 & ~n5574 ;
  assign n5576 = n4411 & n5575 ;
  assign n5584 = n802 ^ n680 ^ 1'b0 ;
  assign n5582 = n4058 ^ n1462 ^ 1'b0 ;
  assign n5577 = n983 & ~n1435 ;
  assign n5578 = n139 & n5577 ;
  assign n5579 = n963 & ~n5578 ;
  assign n5580 = n5197 & n5579 ;
  assign n5581 = ~n2966 & n5580 ;
  assign n5583 = n5582 ^ n5581 ^ 1'b0 ;
  assign n5585 = n5584 ^ n5583 ^ 1'b0 ;
  assign n5586 = n774 & ~n4204 ;
  assign n5587 = n5586 ^ n176 ^ 1'b0 ;
  assign n5588 = n5587 ^ n4008 ^ 1'b0 ;
  assign n5589 = n1405 & n5588 ;
  assign n5590 = n709 & ~n3429 ;
  assign n5591 = n5538 | n5590 ;
  assign n5592 = ( n3040 & ~n3179 ) | ( n3040 & n4056 ) | ( ~n3179 & n4056 ) ;
  assign n5593 = ~n1386 & n5592 ;
  assign n5594 = n5591 & n5593 ;
  assign n5595 = n5594 ^ n5264 ^ n4347 ;
  assign n5596 = n2610 ^ n2576 ^ 1'b0 ;
  assign n5597 = n2078 | n2804 ;
  assign n5598 = n3628 & n5597 ;
  assign n5599 = n5598 ^ n2729 ^ 1'b0 ;
  assign n5600 = n5596 & n5599 ;
  assign n5601 = ~n1455 & n5600 ;
  assign n5602 = n998 ^ n379 ^ 1'b0 ;
  assign n5603 = n5602 ^ n762 ^ 1'b0 ;
  assign n5604 = n5603 ^ n1926 ^ 1'b0 ;
  assign n5605 = n918 & n2595 ;
  assign n5606 = n826 & n5605 ;
  assign n5607 = ~n902 & n2307 ;
  assign n5608 = ( n82 & n5606 ) | ( n82 & n5607 ) | ( n5606 & n5607 ) ;
  assign n5609 = n5608 ^ n5240 ^ 1'b0 ;
  assign n5610 = n2090 & ~n5609 ;
  assign n5611 = n1686 & n3544 ;
  assign n5612 = n39 & n5611 ;
  assign n5613 = n1195 | n5612 ;
  assign n5614 = n5522 | n5613 ;
  assign n5615 = n5614 ^ n641 ^ 1'b0 ;
  assign n5619 = n4357 ^ n3027 ^ 1'b0 ;
  assign n5620 = n4654 & ~n5619 ;
  assign n5617 = ~n604 & n1314 ;
  assign n5616 = n400 & n3192 ;
  assign n5618 = n5617 ^ n5616 ^ n1455 ;
  assign n5621 = n5620 ^ n5618 ^ 1'b0 ;
  assign n5622 = n5217 & n5621 ;
  assign n5623 = n3742 ^ n3255 ^ n1467 ;
  assign n5624 = n270 | n4889 ;
  assign n5625 = n5624 ^ n527 ^ 1'b0 ;
  assign n5626 = ~n41 & n177 ;
  assign n5627 = n5626 ^ n2636 ^ n918 ;
  assign n5628 = ~n1641 & n2815 ;
  assign n5629 = n827 ^ n439 ^ 1'b0 ;
  assign n5630 = n1895 | n5629 ;
  assign n5631 = n960 & n5630 ;
  assign n5632 = n1488 & n2242 ;
  assign n5634 = n231 & n2618 ;
  assign n5633 = n892 & n4741 ;
  assign n5635 = n5634 ^ n5633 ^ 1'b0 ;
  assign n5640 = ~n1538 & n2179 ;
  assign n5636 = n1348 & n1614 ;
  assign n5637 = n5636 ^ n1717 ^ 1'b0 ;
  assign n5638 = n2303 & ~n5637 ;
  assign n5639 = n5638 ^ n836 ^ 1'b0 ;
  assign n5641 = n5640 ^ n5639 ^ 1'b0 ;
  assign n5647 = n51 | n5064 ;
  assign n5648 = n5647 ^ n1282 ^ 1'b0 ;
  assign n5649 = ( n4083 & ~n4435 ) | ( n4083 & n5648 ) | ( ~n4435 & n5648 ) ;
  assign n5642 = n245 & n424 ;
  assign n5643 = n1282 & n5642 ;
  assign n5644 = n2953 ^ n2943 ^ 1'b0 ;
  assign n5645 = n960 & ~n5644 ;
  assign n5646 = ~n5643 & n5645 ;
  assign n5650 = n5649 ^ n5646 ^ 1'b0 ;
  assign n5651 = n1071 | n4514 ;
  assign n5652 = n493 & n5651 ;
  assign n5653 = n5652 ^ n3183 ^ n3180 ;
  assign n5654 = n4560 ^ n3167 ^ 1'b0 ;
  assign n5655 = n5654 ^ n3435 ^ 1'b0 ;
  assign n5657 = n1793 ^ n1427 ^ 1'b0 ;
  assign n5656 = n3603 ^ n2203 ^ n366 ;
  assign n5658 = n5657 ^ n5656 ^ n4342 ;
  assign n5659 = n611 ^ n79 ^ 1'b0 ;
  assign n5660 = n5059 & ~n5659 ;
  assign n5661 = n5660 ^ n1493 ^ 1'b0 ;
  assign n5662 = n3575 & n5661 ;
  assign n5663 = n4688 ^ n4120 ^ 1'b0 ;
  assign n5665 = n172 | n3625 ;
  assign n5664 = n91 | n3630 ;
  assign n5666 = n5665 ^ n5664 ^ 1'b0 ;
  assign n5667 = ~n734 & n1225 ;
  assign n5668 = ( ~n2350 & n5666 ) | ( ~n2350 & n5667 ) | ( n5666 & n5667 ) ;
  assign n5671 = n3445 ^ n341 ^ 1'b0 ;
  assign n5672 = n3856 | n5671 ;
  assign n5669 = n1531 & ~n2915 ;
  assign n5670 = ~n2818 & n5669 ;
  assign n5673 = n5672 ^ n5670 ^ 1'b0 ;
  assign n5674 = n3602 ^ n1124 ^ 1'b0 ;
  assign n5675 = n1741 & ~n5674 ;
  assign n5676 = ( ~n916 & n1167 ) | ( ~n916 & n5675 ) | ( n1167 & n5675 ) ;
  assign n5677 = n5335 & n5676 ;
  assign n5678 = n5673 & n5677 ;
  assign n5679 = n747 & ~n5678 ;
  assign n5682 = n1745 & ~n2146 ;
  assign n5683 = ~n1303 & n5682 ;
  assign n5684 = n3597 ^ n1045 ^ 1'b0 ;
  assign n5685 = n5684 ^ n2036 ^ 1'b0 ;
  assign n5686 = n5683 & n5685 ;
  assign n5681 = n3686 | n4526 ;
  assign n5687 = n5686 ^ n5681 ^ 1'b0 ;
  assign n5680 = n3196 & n4974 ;
  assign n5688 = n5687 ^ n5680 ^ 1'b0 ;
  assign n5689 = n5557 ^ n1332 ^ 1'b0 ;
  assign n5690 = x5 & ~n5689 ;
  assign n5691 = ( n156 & n179 ) | ( n156 & ~n882 ) | ( n179 & ~n882 ) ;
  assign n5692 = n5691 ^ n4107 ^ 1'b0 ;
  assign n5693 = ~n172 & n5692 ;
  assign n5694 = n319 | n340 ;
  assign n5695 = n5694 ^ n4493 ^ 1'b0 ;
  assign n5696 = n1517 | n5695 ;
  assign n5697 = n3837 & n5696 ;
  assign n5698 = n263 & ~n529 ;
  assign n5699 = n5698 ^ n647 ^ 1'b0 ;
  assign n5700 = ( ~n1167 & n1348 ) | ( ~n1167 & n3082 ) | ( n1348 & n3082 ) ;
  assign n5701 = ~n2471 & n5700 ;
  assign n5702 = n5699 & n5701 ;
  assign n5703 = n401 | n5702 ;
  assign n5704 = n5703 ^ n674 ^ 1'b0 ;
  assign n5705 = n442 & n2925 ;
  assign n5706 = n5705 ^ n954 ^ 1'b0 ;
  assign n5707 = ( ~n587 & n3229 ) | ( ~n587 & n5706 ) | ( n3229 & n5706 ) ;
  assign n5708 = n1332 | n5707 ;
  assign n5709 = n451 & n4258 ;
  assign n5710 = ~n169 & n2916 ;
  assign n5711 = n3973 ^ n3898 ^ n2674 ;
  assign n5712 = ( n4310 & n5710 ) | ( n4310 & ~n5711 ) | ( n5710 & ~n5711 ) ;
  assign n5713 = n790 ^ n63 ^ 1'b0 ;
  assign n5714 = n5713 ^ n4004 ^ n2795 ;
  assign n5715 = ( ~n2616 & n3824 ) | ( ~n2616 & n5714 ) | ( n3824 & n5714 ) ;
  assign n5716 = n5715 ^ n1175 ^ 1'b0 ;
  assign n5717 = n3673 ^ n2203 ^ n1233 ;
  assign n5718 = ~n4491 & n5717 ;
  assign n5719 = ( n2892 & n5716 ) | ( n2892 & n5718 ) | ( n5716 & n5718 ) ;
  assign n5720 = n1381 | n2165 ;
  assign n5721 = n608 | n5720 ;
  assign n5722 = n3774 & ~n5721 ;
  assign n5723 = n448 | n4673 ;
  assign n5724 = n2993 | n5723 ;
  assign n5725 = ~n5722 & n5724 ;
  assign n5728 = n5143 ^ n753 ^ 1'b0 ;
  assign n5729 = n3193 & ~n5728 ;
  assign n5726 = n2885 & ~n3307 ;
  assign n5727 = ~n2282 & n5726 ;
  assign n5730 = n5729 ^ n5727 ^ 1'b0 ;
  assign n5731 = n3465 & ~n3892 ;
  assign n5732 = n523 & n5731 ;
  assign n5733 = n203 & ~n2047 ;
  assign n5734 = n5732 & n5733 ;
  assign n5735 = n5388 ^ n2775 ^ 1'b0 ;
  assign n5736 = n5735 ^ n5001 ^ 1'b0 ;
  assign n5737 = n4231 ^ n2807 ^ n1335 ;
  assign n5738 = ( n84 & n2595 ) | ( n84 & ~n5737 ) | ( n2595 & ~n5737 ) ;
  assign n5739 = n2131 | n4723 ;
  assign n5740 = n4985 & ~n5739 ;
  assign n5741 = ( n3773 & n4793 ) | ( n3773 & n5740 ) | ( n4793 & n5740 ) ;
  assign n5742 = n2161 ^ n876 ^ 1'b0 ;
  assign n5743 = n5742 ^ n2987 ^ 1'b0 ;
  assign n5744 = n2944 | n3271 ;
  assign n5745 = ~n1842 & n2925 ;
  assign n5746 = n3867 | n3884 ;
  assign n5747 = n3684 | n5746 ;
  assign n5748 = ~n2117 & n2449 ;
  assign n5749 = n5748 ^ n2811 ^ n2500 ;
  assign n5750 = n524 | n5749 ;
  assign n5751 = n1260 ^ n514 ^ 1'b0 ;
  assign n5752 = n5751 ^ n4490 ^ 1'b0 ;
  assign n5753 = n3203 & n5752 ;
  assign n5754 = n2401 ^ n899 ^ n626 ;
  assign n5755 = ~n566 & n1028 ;
  assign n5756 = n3759 & n5755 ;
  assign n5757 = ( n829 & ~n5754 ) | ( n829 & n5756 ) | ( ~n5754 & n5756 ) ;
  assign n5758 = n4706 & n5143 ;
  assign n5759 = ~n222 & n1472 ;
  assign n5760 = n1175 ^ n1167 ^ n906 ;
  assign n5761 = ~n2047 & n5760 ;
  assign n5762 = n3203 & n5761 ;
  assign n5763 = n5759 & n5762 ;
  assign n5764 = ~n4542 & n5763 ;
  assign n5768 = n2650 & ~n2805 ;
  assign n5766 = n3552 ^ n1876 ^ n141 ;
  assign n5767 = n1587 & ~n5766 ;
  assign n5769 = n5768 ^ n5767 ^ 1'b0 ;
  assign n5770 = n5769 ^ n955 ^ 1'b0 ;
  assign n5765 = ~n1403 & n1734 ;
  assign n5771 = n5770 ^ n5765 ^ 1'b0 ;
  assign n5772 = n3658 ^ n1419 ^ 1'b0 ;
  assign n5773 = n1122 | n5772 ;
  assign n5774 = n3085 | n5773 ;
  assign n5775 = n3925 ^ n1679 ^ 1'b0 ;
  assign n5776 = n5774 & ~n5775 ;
  assign n5777 = n3418 & n5776 ;
  assign n5778 = n5777 ^ n3009 ^ 1'b0 ;
  assign n5779 = ~n987 & n3726 ;
  assign n5780 = n93 & n5779 ;
  assign n5781 = n2142 & ~n5780 ;
  assign n5782 = n2784 ^ n2032 ^ 1'b0 ;
  assign n5783 = n5782 ^ n2387 ^ 1'b0 ;
  assign n5784 = n5783 ^ n5776 ^ 1'b0 ;
  assign n5785 = n3227 | n5784 ;
  assign n5786 = ( n4221 & n4270 ) | ( n4221 & n5241 ) | ( n4270 & n5241 ) ;
  assign n5787 = ~n1746 & n3020 ;
  assign n5788 = n102 & n5787 ;
  assign n5789 = n2653 ^ n1789 ^ 1'b0 ;
  assign n5790 = n5688 | n5789 ;
  assign n5791 = n644 & ~n1276 ;
  assign n5793 = n3521 ^ n136 ^ n26 ;
  assign n5792 = ~n1820 & n2481 ;
  assign n5794 = n5793 ^ n5792 ^ 1'b0 ;
  assign n5795 = ( n2086 & n3295 ) | ( n2086 & ~n5794 ) | ( n3295 & ~n5794 ) ;
  assign n5796 = ( n73 & n1249 ) | ( n73 & ~n5795 ) | ( n1249 & ~n5795 ) ;
  assign n5797 = ~n1133 & n1328 ;
  assign n5798 = n5797 ^ n1592 ^ 1'b0 ;
  assign n5799 = ~n1875 & n5798 ;
  assign n5801 = n439 | n2635 ;
  assign n5802 = n5801 ^ n2173 ^ 1'b0 ;
  assign n5800 = n134 | n1493 ;
  assign n5803 = n5802 ^ n5800 ^ n2509 ;
  assign n5804 = n171 | n5440 ;
  assign n5805 = n435 & ~n4515 ;
  assign n5806 = n5805 ^ n3761 ^ 1'b0 ;
  assign n5807 = ~n1666 & n1839 ;
  assign n5808 = ~n4548 & n5807 ;
  assign n5809 = n5691 ^ n2971 ^ 1'b0 ;
  assign n5810 = n1022 & n5809 ;
  assign n5811 = n863 & n5810 ;
  assign n5812 = n2727 & ~n5811 ;
  assign n5813 = n5812 ^ n3192 ^ 1'b0 ;
  assign n5814 = ( n252 & n963 ) | ( n252 & ~n5455 ) | ( n963 & ~n5455 ) ;
  assign n5815 = n5814 ^ n3351 ^ n3271 ;
  assign n5821 = ~n949 & n2098 ;
  assign n5822 = ~n201 & n5821 ;
  assign n5817 = n2986 ^ n1647 ^ n443 ;
  assign n5818 = n5817 ^ n2513 ^ 1'b0 ;
  assign n5816 = n3168 | n4233 ;
  assign n5819 = n5818 ^ n5816 ^ 1'b0 ;
  assign n5820 = n2105 | n5819 ;
  assign n5823 = n5822 ^ n5820 ^ n3158 ;
  assign n5824 = n3271 ^ n3053 ^ n2073 ;
  assign n5825 = n3967 ^ n2640 ^ n188 ;
  assign n5826 = ~n3365 & n5825 ;
  assign n5827 = ~n800 & n5826 ;
  assign n5828 = n1441 ^ n255 ^ 1'b0 ;
  assign n5829 = ~n769 & n5828 ;
  assign n5830 = n5827 & n5829 ;
  assign n5831 = n4154 ^ n989 ^ 1'b0 ;
  assign n5832 = n30 & ~n563 ;
  assign n5833 = n1791 & n2447 ;
  assign n5834 = ~n5832 & n5833 ;
  assign n5835 = n5831 | n5834 ;
  assign n5836 = n5835 ^ n3149 ^ 1'b0 ;
  assign n5837 = ( n4116 & ~n4807 ) | ( n4116 & n5200 ) | ( ~n4807 & n5200 ) ;
  assign n5838 = n596 & n2946 ;
  assign n5839 = n1419 ^ n221 ^ 1'b0 ;
  assign n5840 = n5838 | n5839 ;
  assign n5841 = ( n1660 & ~n3149 ) | ( n1660 & n3810 ) | ( ~n3149 & n3810 ) ;
  assign n5842 = ~n5840 & n5841 ;
  assign n5843 = n5842 ^ n1383 ^ 1'b0 ;
  assign n5844 = n5843 ^ n1746 ^ 1'b0 ;
  assign n5845 = n2237 ^ n1207 ^ 1'b0 ;
  assign n5846 = n5845 ^ n3004 ^ 1'b0 ;
  assign n5847 = n4357 | n5846 ;
  assign n5848 = n2326 ^ n999 ^ n308 ;
  assign n5849 = n3634 & n5848 ;
  assign n5850 = n5849 ^ n1826 ^ 1'b0 ;
  assign n5851 = ( n2854 & n4602 ) | ( n2854 & n4983 ) | ( n4602 & n4983 ) ;
  assign n5852 = n991 ^ n455 ^ 1'b0 ;
  assign n5853 = n5852 ^ n1043 ^ 1'b0 ;
  assign n5854 = ( ~n1898 & n2589 ) | ( ~n1898 & n5853 ) | ( n2589 & n5853 ) ;
  assign n5855 = n3105 | n3604 ;
  assign n5856 = n67 | n5855 ;
  assign n5857 = n3469 | n5856 ;
  assign n5858 = n5857 ^ n4199 ^ 1'b0 ;
  assign n5859 = n837 ^ n581 ^ 1'b0 ;
  assign n5860 = n5859 ^ n5251 ^ 1'b0 ;
  assign n5861 = n4904 ^ n3770 ^ 1'b0 ;
  assign n5862 = n3567 ^ n3137 ^ 1'b0 ;
  assign n5863 = n3088 & ~n3421 ;
  assign n5864 = ~n18 & n5863 ;
  assign n5865 = ~n1917 & n2596 ;
  assign n5866 = ~x6 & n5865 ;
  assign n5867 = n5866 ^ n3985 ^ n949 ;
  assign n5868 = n150 & ~n2712 ;
  assign n5869 = n560 & ~n1249 ;
  assign n5870 = n3699 & ~n5869 ;
  assign n5871 = n3295 | n5870 ;
  assign n5872 = n3848 & ~n5871 ;
  assign n5873 = n63 & ~n1807 ;
  assign n5874 = ( n358 & ~n863 ) | ( n358 & n1591 ) | ( ~n863 & n1591 ) ;
  assign n5875 = n4988 & ~n5874 ;
  assign n5876 = n5875 ^ n4366 ^ 1'b0 ;
  assign n5877 = ( n4006 & n5873 ) | ( n4006 & n5876 ) | ( n5873 & n5876 ) ;
  assign n5878 = n4048 ^ n54 ^ 1'b0 ;
  assign n5879 = n5878 ^ n4294 ^ 1'b0 ;
  assign n5881 = n2070 ^ n864 ^ 1'b0 ;
  assign n5880 = n2259 & ~n3364 ;
  assign n5882 = n5881 ^ n5880 ^ 1'b0 ;
  assign n5884 = n1443 & ~n3029 ;
  assign n5885 = ~n3379 & n5884 ;
  assign n5883 = n2870 ^ n62 ^ 1'b0 ;
  assign n5886 = n5885 ^ n5883 ^ 1'b0 ;
  assign n5887 = n5886 ^ n5822 ^ 1'b0 ;
  assign n5888 = n2541 & ~n5887 ;
  assign n5895 = n238 & ~n786 ;
  assign n5889 = n1439 ^ n1019 ^ 1'b0 ;
  assign n5890 = n928 & ~n5889 ;
  assign n5891 = n2313 ^ n991 ^ n100 ;
  assign n5892 = n5891 ^ n3348 ^ 1'b0 ;
  assign n5893 = n5890 & n5892 ;
  assign n5894 = ~n3744 & n5893 ;
  assign n5896 = n5895 ^ n5894 ^ 1'b0 ;
  assign n5898 = ( ~n151 & n605 ) | ( ~n151 & n2447 ) | ( n605 & n2447 ) ;
  assign n5897 = n4809 ^ n759 ^ 1'b0 ;
  assign n5899 = n5898 ^ n5897 ^ 1'b0 ;
  assign n5900 = n2701 | n5899 ;
  assign n5901 = n5900 ^ n172 ^ 1'b0 ;
  assign n5902 = n4262 & ~n5901 ;
  assign n5903 = n3671 & ~n5322 ;
  assign n5904 = n5797 ^ n4629 ^ 1'b0 ;
  assign n5905 = ~n1330 & n2492 ;
  assign n5906 = n5905 ^ n1832 ^ 1'b0 ;
  assign n5907 = n5906 ^ n5696 ^ n1489 ;
  assign n5908 = n2568 | n3195 ;
  assign n5909 = n2041 & ~n5908 ;
  assign n5910 = n5909 ^ n4242 ^ n1606 ;
  assign n5911 = n5910 ^ n259 ^ 1'b0 ;
  assign n5912 = n137 | n2138 ;
  assign n5913 = n2640 ^ n63 ^ n15 ;
  assign n5914 = ~n3122 & n5913 ;
  assign n5915 = n1848 | n4366 ;
  assign n5916 = n4147 & ~n5384 ;
  assign n5917 = n2124 ^ n2034 ^ 1'b0 ;
  assign n5918 = n2021 & ~n5917 ;
  assign n5919 = n1942 & n5918 ;
  assign n5920 = n4099 | n5919 ;
  assign n5921 = n4276 & ~n4847 ;
  assign n5922 = ~n5678 & n5921 ;
  assign n5923 = ~n2799 & n5922 ;
  assign n5924 = ~n732 & n1713 ;
  assign n5925 = n3209 & ~n5924 ;
  assign n5926 = n946 | n2841 ;
  assign n5927 = n4674 & ~n5926 ;
  assign n5928 = n5890 ^ n3372 ^ n2677 ;
  assign n5930 = n4167 ^ n259 ^ 1'b0 ;
  assign n5929 = n1897 & ~n5053 ;
  assign n5931 = n5930 ^ n5929 ^ 1'b0 ;
  assign n5932 = n5761 ^ n2213 ^ 1'b0 ;
  assign n5933 = n1198 & ~n5028 ;
  assign n5934 = n1878 & n2693 ;
  assign n5935 = ~n4254 & n5934 ;
  assign n5936 = n5935 ^ n641 ^ 1'b0 ;
  assign n5937 = n974 ^ n417 ^ n312 ;
  assign n5938 = n4719 & n5937 ;
  assign n5939 = ( n2986 & ~n5936 ) | ( n2986 & n5938 ) | ( ~n5936 & n5938 ) ;
  assign n5940 = n5939 ^ n3067 ^ 1'b0 ;
  assign n5941 = ~n723 & n5940 ;
  assign n5942 = n3508 ^ n656 ^ x11 ;
  assign n5943 = n698 | n5942 ;
  assign n5944 = n5943 ^ n2746 ^ 1'b0 ;
  assign n5945 = ~n4216 & n5944 ;
  assign n5946 = n5684 & n5945 ;
  assign n5947 = n3111 & ~n3582 ;
  assign n5948 = n5946 & n5947 ;
  assign n5949 = ~n332 & n4523 ;
  assign n5950 = n2524 ^ n1108 ^ 1'b0 ;
  assign n5951 = n105 & n5950 ;
  assign n5952 = n3201 & n5759 ;
  assign n5953 = ( n4310 & n5951 ) | ( n4310 & n5952 ) | ( n5951 & n5952 ) ;
  assign n5954 = n2378 ^ n1942 ^ 1'b0 ;
  assign n5955 = n5954 ^ n1818 ^ 1'b0 ;
  assign n5956 = n208 | n2471 ;
  assign n5957 = n556 | n5956 ;
  assign n5958 = ( n720 & ~n4904 ) | ( n720 & n5957 ) | ( ~n4904 & n5957 ) ;
  assign n5959 = n5234 | n5845 ;
  assign n5960 = n2682 & n5222 ;
  assign n5961 = n1800 & n5960 ;
  assign n5962 = n346 ^ n91 ^ 1'b0 ;
  assign n5963 = n5961 | n5962 ;
  assign n5967 = n5078 ^ n2535 ^ 1'b0 ;
  assign n5968 = ~n921 & n5967 ;
  assign n5964 = n2935 & ~n4159 ;
  assign n5965 = n400 & n5964 ;
  assign n5966 = n5965 ^ n3663 ^ 1'b0 ;
  assign n5969 = n5968 ^ n5966 ^ 1'b0 ;
  assign n5970 = n3383 ^ n998 ^ 1'b0 ;
  assign n5971 = n4458 & ~n5970 ;
  assign n5972 = ~n4273 & n5971 ;
  assign n5973 = n5070 ^ n4539 ^ n4289 ;
  assign n5974 = ~n3170 & n4319 ;
  assign n5975 = ( n5509 & ~n5973 ) | ( n5509 & n5974 ) | ( ~n5973 & n5974 ) ;
  assign n5976 = n1722 & n2463 ;
  assign n5977 = ~n1457 & n5976 ;
  assign n5978 = n5977 ^ n2876 ^ 1'b0 ;
  assign n5979 = n1169 & n3151 ;
  assign n5980 = ~n2537 & n2935 ;
  assign n5981 = ~n597 & n5980 ;
  assign n5982 = n5981 ^ n1845 ^ 1'b0 ;
  assign n5984 = ~n177 & n1586 ;
  assign n5985 = n1346 & n5984 ;
  assign n5986 = n1290 ^ n597 ^ 1'b0 ;
  assign n5987 = ( n1786 & n5985 ) | ( n1786 & n5986 ) | ( n5985 & n5986 ) ;
  assign n5983 = n1216 & ~n3170 ;
  assign n5988 = n5987 ^ n5983 ^ 1'b0 ;
  assign n5989 = n260 & ~n2044 ;
  assign n5990 = n5989 ^ n1996 ^ 1'b0 ;
  assign n5991 = ~n59 & n5782 ;
  assign n5992 = n5991 ^ n989 ^ 1'b0 ;
  assign n5993 = n5992 ^ n2758 ^ 1'b0 ;
  assign n5994 = n5990 & ~n5993 ;
  assign n5995 = n5994 ^ n1766 ^ n272 ;
  assign n5996 = n3824 ^ n1666 ^ 1'b0 ;
  assign n5997 = n5758 ^ n3979 ^ n3662 ;
  assign n5998 = n1602 | n4127 ;
  assign n5999 = n556 ^ n523 ^ 1'b0 ;
  assign n6000 = n5088 & n5999 ;
  assign n6001 = n6000 ^ n4322 ^ n1640 ;
  assign n6002 = n2830 & n6001 ;
  assign n6003 = ~n2083 & n6002 ;
  assign n6004 = n1408 ^ n1051 ^ 1'b0 ;
  assign n6005 = n633 & ~n654 ;
  assign n6008 = n1882 ^ n989 ^ n698 ;
  assign n6009 = n6008 ^ n2511 ^ n42 ;
  assign n6006 = n2836 & ~n5458 ;
  assign n6007 = n6006 ^ n4267 ^ 1'b0 ;
  assign n6010 = n6009 ^ n6007 ^ n624 ;
  assign n6011 = ~n459 & n1315 ;
  assign n6012 = n6011 ^ n411 ^ 1'b0 ;
  assign n6013 = n1432 & n6012 ;
  assign n6014 = n6013 ^ n2514 ^ n601 ;
  assign n6015 = n2270 & ~n2986 ;
  assign n6016 = n1424 & n6015 ;
  assign n6017 = n2170 ^ n129 ^ 1'b0 ;
  assign n6018 = n692 | n6017 ;
  assign n6019 = n6018 ^ n3919 ^ 1'b0 ;
  assign n6020 = n2402 ^ n1600 ^ 1'b0 ;
  assign n6021 = n3437 ^ n865 ^ n318 ;
  assign n6022 = n5088 | n6021 ;
  assign n6023 = n1167 ^ n1076 ^ 1'b0 ;
  assign n6024 = ~n378 & n6023 ;
  assign n6025 = ( n1896 & ~n3479 ) | ( n1896 & n6024 ) | ( ~n3479 & n6024 ) ;
  assign n6026 = n6025 ^ n4703 ^ n169 ;
  assign n6027 = n888 & n1586 ;
  assign n6028 = n57 & n1784 ;
  assign n6029 = n6028 ^ n1605 ^ 1'b0 ;
  assign n6030 = n1052 & ~n6029 ;
  assign n6031 = n260 | n3083 ;
  assign n6032 = n1135 & ~n6031 ;
  assign n6033 = n2483 & ~n6032 ;
  assign n6034 = ~n4845 & n6033 ;
  assign n6035 = n2833 ^ n713 ^ 1'b0 ;
  assign n6036 = n3443 | n6035 ;
  assign n6037 = n6036 ^ n5602 ^ 1'b0 ;
  assign n6038 = ~n513 & n3967 ;
  assign n6039 = ~n6037 & n6038 ;
  assign n6040 = n6039 ^ n694 ^ 1'b0 ;
  assign n6041 = n97 | n4138 ;
  assign n6042 = ( ~n1944 & n3953 ) | ( ~n1944 & n6041 ) | ( n3953 & n6041 ) ;
  assign n6043 = n5738 ^ n2262 ^ 1'b0 ;
  assign n6044 = n1660 | n4549 ;
  assign n6045 = n6044 ^ n910 ^ 1'b0 ;
  assign n6046 = ~n5820 & n6045 ;
  assign n6047 = n6046 ^ n3725 ^ 1'b0 ;
  assign n6048 = n4612 ^ n3275 ^ 1'b0 ;
  assign n6049 = ~n6047 & n6048 ;
  assign n6050 = n5132 ^ n5114 ^ 1'b0 ;
  assign n6057 = ~n585 & n4760 ;
  assign n6058 = ~n209 & n6057 ;
  assign n6051 = n991 | n4030 ;
  assign n6052 = ( n168 & n1143 ) | ( n168 & n6051 ) | ( n1143 & n6051 ) ;
  assign n6053 = n1373 & ~n1918 ;
  assign n6054 = n6053 ^ n145 ^ 1'b0 ;
  assign n6055 = ~n6052 & n6054 ;
  assign n6056 = n2324 & n6055 ;
  assign n6059 = n6058 ^ n6056 ^ 1'b0 ;
  assign n6060 = ( n1869 & n3336 ) | ( n1869 & ~n6059 ) | ( n3336 & ~n6059 ) ;
  assign n6061 = n5773 ^ n1022 ^ 1'b0 ;
  assign n6062 = n4815 | n6061 ;
  assign n6063 = n3691 ^ n2344 ^ 1'b0 ;
  assign n6064 = ~n6062 & n6063 ;
  assign n6067 = n4457 ^ n3506 ^ n2218 ;
  assign n6065 = n2563 | n4327 ;
  assign n6066 = n6065 ^ n1081 ^ 1'b0 ;
  assign n6068 = n6067 ^ n6066 ^ 1'b0 ;
  assign n6069 = n1220 | n6068 ;
  assign n6070 = n2023 | n2123 ;
  assign n6071 = n6070 ^ n2631 ^ 1'b0 ;
  assign n6072 = n1649 & ~n6071 ;
  assign n6073 = ~n3414 & n6072 ;
  assign n6074 = n2902 | n6073 ;
  assign n6075 = n3339 ^ n152 ^ 1'b0 ;
  assign n6077 = n1051 & ~n5557 ;
  assign n6078 = n6077 ^ n1635 ^ 1'b0 ;
  assign n6076 = n5415 ^ n4163 ^ 1'b0 ;
  assign n6079 = n6078 ^ n6076 ^ 1'b0 ;
  assign n6080 = n6079 ^ n252 ^ 1'b0 ;
  assign n6081 = n2080 ^ n1533 ^ x3 ;
  assign n6082 = ~n2649 & n6081 ;
  assign n6083 = n991 ^ n334 ^ 1'b0 ;
  assign n6084 = ~n3671 & n6083 ;
  assign n6085 = ~n381 & n6084 ;
  assign n6086 = n6085 ^ n4801 ^ 1'b0 ;
  assign n6087 = ~n1279 & n6086 ;
  assign n6088 = n6087 ^ n1764 ^ 1'b0 ;
  assign n6089 = n6088 ^ n2186 ^ 1'b0 ;
  assign n6090 = ~n1956 & n2433 ;
  assign n6091 = n101 & n6090 ;
  assign n6092 = n5582 ^ n3027 ^ 1'b0 ;
  assign n6093 = n4240 | n6092 ;
  assign n6094 = n4048 ^ n1439 ^ 1'b0 ;
  assign n6095 = n4399 ^ n2778 ^ 1'b0 ;
  assign n6096 = n1037 & ~n6095 ;
  assign n6097 = n1459 | n2720 ;
  assign n6098 = ~n873 & n1256 ;
  assign n6099 = n1010 ^ n360 ^ 1'b0 ;
  assign n6100 = n1339 & ~n6099 ;
  assign n6101 = n945 & n5742 ;
  assign n6102 = n135 | n2025 ;
  assign n6103 = n91 & n6102 ;
  assign n6104 = ~n2053 & n6103 ;
  assign n6105 = n89 | n6104 ;
  assign n6106 = n6105 ^ n5244 ^ 1'b0 ;
  assign n6107 = ~n3922 & n6106 ;
  assign n6113 = n551 | n2107 ;
  assign n6114 = n6113 ^ n1800 ^ 1'b0 ;
  assign n6112 = n1760 & ~n4192 ;
  assign n6115 = n6114 ^ n6112 ^ 1'b0 ;
  assign n6108 = ~n2138 & n3301 ;
  assign n6109 = n6108 ^ n3389 ^ 1'b0 ;
  assign n6110 = n1948 & ~n6109 ;
  assign n6111 = n1079 | n6110 ;
  assign n6116 = n6115 ^ n6111 ^ n1360 ;
  assign n6120 = n2806 | n3294 ;
  assign n6117 = n654 | n772 ;
  assign n6118 = n2170 & ~n6117 ;
  assign n6119 = n4216 & ~n6118 ;
  assign n6121 = n6120 ^ n6119 ^ 1'b0 ;
  assign n6122 = n719 & n3207 ;
  assign n6123 = n469 & n1436 ;
  assign n6124 = n1628 ^ n1421 ^ 1'b0 ;
  assign n6125 = n6123 & ~n6124 ;
  assign n6126 = ~n603 & n6125 ;
  assign n6127 = ~n2005 & n6126 ;
  assign n6128 = n6127 ^ n6008 ^ 1'b0 ;
  assign n6129 = n6128 ^ n601 ^ 1'b0 ;
  assign n6130 = n878 ^ n443 ^ 1'b0 ;
  assign n6131 = n79 & ~n6130 ;
  assign n6132 = n63 | n581 ;
  assign n6133 = n5318 & ~n6132 ;
  assign n6134 = n2859 | n6133 ;
  assign n6135 = n379 & ~n3580 ;
  assign n6136 = n3599 ^ n1168 ^ 1'b0 ;
  assign n6137 = n2958 & n6136 ;
  assign n6138 = n6137 ^ n2751 ^ 1'b0 ;
  assign n6142 = ~n57 & n1334 ;
  assign n6143 = n6142 ^ n345 ^ 1'b0 ;
  assign n6139 = n1896 ^ n1845 ^ 1'b0 ;
  assign n6140 = n6139 ^ n3336 ^ 1'b0 ;
  assign n6141 = n1766 | n6140 ;
  assign n6144 = n6143 ^ n6141 ^ 1'b0 ;
  assign n6145 = n6144 ^ n2142 ^ 1'b0 ;
  assign n6146 = n1762 & ~n6145 ;
  assign n6147 = n2885 | n6146 ;
  assign n6148 = n2763 ^ n1809 ^ 1'b0 ;
  assign n6149 = ~n1118 & n6148 ;
  assign n6154 = n1522 ^ n1324 ^ n202 ;
  assign n6150 = n1164 & ~n3959 ;
  assign n6151 = n6150 ^ n503 ^ 1'b0 ;
  assign n6152 = n1138 & n6151 ;
  assign n6153 = n6152 ^ n5535 ^ n1563 ;
  assign n6155 = n6154 ^ n6153 ^ 1'b0 ;
  assign n6156 = n305 & n1560 ;
  assign n6157 = n178 | n6156 ;
  assign n6158 = ~n1412 & n6157 ;
  assign n6159 = ~n1647 & n6158 ;
  assign n6160 = n6049 ^ n4614 ^ n3371 ;
  assign n6161 = n4633 & n5088 ;
  assign n6162 = n3413 ^ n3156 ^ 1'b0 ;
  assign n6163 = n6161 & n6162 ;
  assign n6164 = n636 ^ n459 ^ 1'b0 ;
  assign n6165 = n3180 | n6164 ;
  assign n6166 = n2328 | n6165 ;
  assign n6167 = ( n5527 & n5540 ) | ( n5527 & n6166 ) | ( n5540 & n6166 ) ;
  assign n6168 = ( ~n867 & n1287 ) | ( ~n867 & n4567 ) | ( n1287 & n4567 ) ;
  assign n6169 = n2005 ^ n1282 ^ n865 ;
  assign n6170 = n2867 & n6169 ;
  assign n6171 = n5658 & n6170 ;
  assign n6172 = n5012 ^ n3053 ^ 1'b0 ;
  assign n6173 = n1810 & ~n6172 ;
  assign n6174 = n3242 & ~n4567 ;
  assign n6175 = n1904 & ~n2461 ;
  assign n6176 = n5057 | n6175 ;
  assign n6177 = ~n1276 & n2493 ;
  assign n6178 = n6177 ^ n1373 ^ 1'b0 ;
  assign n6179 = n976 | n1403 ;
  assign n6180 = n6179 ^ n2225 ^ 1'b0 ;
  assign n6181 = ( n195 & n2622 ) | ( n195 & n6180 ) | ( n2622 & n6180 ) ;
  assign n6182 = n1162 | n6181 ;
  assign n6183 = n5236 & ~n5656 ;
  assign n6184 = n5222 ^ n2005 ^ 1'b0 ;
  assign n6185 = n973 & ~n6184 ;
  assign n6186 = ( n261 & n4399 ) | ( n261 & n6185 ) | ( n4399 & n6185 ) ;
  assign n6187 = ( n172 & ~n2723 ) | ( n172 & n2886 ) | ( ~n2723 & n2886 ) ;
  assign n6188 = n6187 ^ n1885 ^ 1'b0 ;
  assign n6189 = ( n1253 & ~n2546 ) | ( n1253 & n4503 ) | ( ~n2546 & n4503 ) ;
  assign n6190 = n2082 | n6189 ;
  assign n6191 = n6190 ^ n1225 ^ 1'b0 ;
  assign n6192 = n3853 ^ n261 ^ 1'b0 ;
  assign n6193 = ~n3519 & n6192 ;
  assign n6197 = n216 & n784 ;
  assign n6196 = ( n65 & n1474 ) | ( n65 & ~n4560 ) | ( n1474 & ~n4560 ) ;
  assign n6194 = n2752 | n4193 ;
  assign n6195 = n6194 ^ n742 ^ 1'b0 ;
  assign n6198 = n6197 ^ n6196 ^ n6195 ;
  assign n6199 = n228 & ~n5596 ;
  assign n6200 = ~n5203 & n5590 ;
  assign n6201 = ~n5070 & n6200 ;
  assign n6202 = n5457 ^ n4465 ^ n4434 ;
  assign n6203 = ~n6201 & n6202 ;
  assign n6204 = n247 & n6203 ;
  assign n6205 = n2843 & n3256 ;
  assign n6206 = ~n157 & n6205 ;
  assign n6207 = n4801 ^ n524 ^ 1'b0 ;
  assign n6208 = n4425 & ~n6207 ;
  assign n6209 = ~n159 & n6208 ;
  assign n6210 = ~n1744 & n6209 ;
  assign n6211 = n3477 | n3660 ;
  assign n6212 = ~n1071 & n5430 ;
  assign n6213 = n2871 & n4763 ;
  assign n6214 = n122 & ~n6213 ;
  assign n6216 = ~n61 & n1108 ;
  assign n6217 = ~n835 & n6216 ;
  assign n6215 = n686 & ~n2432 ;
  assign n6218 = n6217 ^ n6215 ^ 1'b0 ;
  assign n6219 = n5197 ^ n411 ^ 1'b0 ;
  assign n6220 = n5483 ^ n2755 ^ n654 ;
  assign n6221 = n6220 ^ n2650 ^ 1'b0 ;
  assign n6222 = ( n3486 & ~n5451 ) | ( n3486 & n6221 ) | ( ~n5451 & n6221 ) ;
  assign n6223 = ~n2354 & n3708 ;
  assign n6224 = n881 & n2157 ;
  assign n6225 = n4904 ^ n145 ^ 1'b0 ;
  assign n6226 = n342 & ~n4761 ;
  assign n6227 = n6226 ^ n32 ^ 1'b0 ;
  assign n6228 = ~n261 & n3148 ;
  assign n6229 = n6228 ^ n3466 ^ 1'b0 ;
  assign n6230 = n1487 ^ n344 ^ n36 ;
  assign n6231 = n6230 ^ n5281 ^ 1'b0 ;
  assign n6233 = n3962 ^ n1934 ^ 1'b0 ;
  assign n6234 = n2049 & ~n6233 ;
  assign n6232 = n174 & n2443 ;
  assign n6235 = n6234 ^ n6232 ^ 1'b0 ;
  assign n6236 = n1373 & n6235 ;
  assign n6237 = n3090 ^ n1103 ^ 1'b0 ;
  assign n6238 = n1984 & n6237 ;
  assign n6239 = n6238 ^ n4792 ^ n1131 ;
  assign n6241 = n817 & ~n3861 ;
  assign n6240 = n1353 ^ n1248 ^ 1'b0 ;
  assign n6242 = n6241 ^ n6240 ^ n893 ;
  assign n6243 = n1122 ^ n1100 ^ 1'b0 ;
  assign n6244 = n1526 ^ n156 ^ 1'b0 ;
  assign n6245 = n6243 & ~n6244 ;
  assign n6246 = ~n338 & n6245 ;
  assign n6247 = n6246 ^ n2006 ^ 1'b0 ;
  assign n6248 = n6247 ^ n1142 ^ 1'b0 ;
  assign n6249 = n1876 & ~n6248 ;
  assign n6250 = n1432 & n6249 ;
  assign n6251 = n6250 ^ n3985 ^ 1'b0 ;
  assign n6252 = n434 & ~n4359 ;
  assign n6253 = ~n1874 & n6252 ;
  assign n6254 = n1520 & ~n3179 ;
  assign n6255 = ( ~n134 & n293 ) | ( ~n134 & n1447 ) | ( n293 & n1447 ) ;
  assign n6256 = n36 | n2344 ;
  assign n6257 = n6255 & ~n6256 ;
  assign n6258 = n6257 ^ n1197 ^ 1'b0 ;
  assign n6259 = n1929 & n6258 ;
  assign n6260 = n498 | n2104 ;
  assign n6261 = n1931 | n6260 ;
  assign n6262 = n6261 ^ n5155 ^ n4495 ;
  assign n6263 = ( n37 & n1104 ) | ( n37 & n2327 ) | ( n1104 & n2327 ) ;
  assign n6264 = n3290 | n6263 ;
  assign n6265 = n6264 ^ n2567 ^ 1'b0 ;
  assign n6266 = ( n4725 & n6262 ) | ( n4725 & n6265 ) | ( n6262 & n6265 ) ;
  assign n6267 = n2733 & ~n6266 ;
  assign n6268 = ~n797 & n1596 ;
  assign n6269 = ~n2757 & n6268 ;
  assign n6270 = n4502 ^ n1201 ^ 1'b0 ;
  assign n6271 = ~n6269 & n6270 ;
  assign n6272 = ~n5712 & n6271 ;
  assign n6273 = ~n2067 & n2176 ;
  assign n6274 = n3510 ^ n2236 ^ 1'b0 ;
  assign n6275 = ~n2436 & n6150 ;
  assign n6276 = n1818 ^ n1332 ^ 1'b0 ;
  assign n6277 = n209 & n6276 ;
  assign n6278 = n4156 ^ n3084 ^ n1169 ;
  assign n6279 = n6278 ^ n1318 ^ 1'b0 ;
  assign n6280 = n822 | n6279 ;
  assign n6281 = n2119 | n6280 ;
  assign n6282 = n6277 | n6281 ;
  assign n6283 = n1186 & ~n2044 ;
  assign n6284 = n723 & n6283 ;
  assign n6285 = n6284 ^ n6205 ^ 1'b0 ;
  assign n6286 = n386 & n3612 ;
  assign n6287 = n676 ^ n519 ^ 1'b0 ;
  assign n6288 = n6286 & n6287 ;
  assign n6289 = ( n279 & n1623 ) | ( n279 & ~n2271 ) | ( n1623 & ~n2271 ) ;
  assign n6290 = n6289 ^ n4869 ^ 1'b0 ;
  assign n6291 = n6288 & n6290 ;
  assign n6292 = x6 & ~n2904 ;
  assign n6293 = n2916 & ~n6292 ;
  assign n6294 = n1459 & ~n5143 ;
  assign n6295 = n1234 & ~n4904 ;
  assign n6296 = ~n2904 & n6295 ;
  assign n6297 = n2858 ^ n220 ^ 1'b0 ;
  assign n6298 = n4678 & n6297 ;
  assign n6299 = n6298 ^ n4617 ^ 1'b0 ;
  assign n6300 = n1539 & n5353 ;
  assign n6301 = n6300 ^ n633 ^ 1'b0 ;
  assign n6302 = n1944 ^ n1630 ^ 1'b0 ;
  assign n6303 = ~n1045 & n6302 ;
  assign n6304 = n1856 & n6303 ;
  assign n6305 = n6304 ^ n4812 ^ 1'b0 ;
  assign n6306 = n2034 & n6305 ;
  assign n6307 = n6306 ^ n51 ^ 1'b0 ;
  assign n6308 = ( n3906 & n5099 ) | ( n3906 & n5837 ) | ( n5099 & n5837 ) ;
  assign n6309 = n1695 | n3575 ;
  assign n6310 = n6309 ^ n3237 ^ 1'b0 ;
  assign n6311 = n622 & n2115 ;
  assign n6312 = ~n2332 & n6311 ;
  assign n6313 = n6312 ^ n680 ^ 1'b0 ;
  assign n6315 = n260 | n1976 ;
  assign n6316 = n1786 | n6315 ;
  assign n6314 = n3888 & ~n6071 ;
  assign n6317 = n6316 ^ n6314 ^ 1'b0 ;
  assign n6318 = n2999 & n5099 ;
  assign n6319 = n6318 ^ n1962 ^ 1'b0 ;
  assign n6320 = n1868 | n4146 ;
  assign n6321 = n6320 ^ n1300 ^ 1'b0 ;
  assign n6322 = n2262 & n6321 ;
  assign n6323 = n4568 & n6322 ;
  assign n6324 = n6323 ^ n3698 ^ 1'b0 ;
  assign n6325 = n350 & n1228 ;
  assign n6326 = n6325 ^ n2213 ^ 1'b0 ;
  assign n6327 = ~n2101 & n6326 ;
  assign n6328 = n6327 ^ n1849 ^ 1'b0 ;
  assign n6329 = ~n2668 & n4163 ;
  assign n6330 = n6329 ^ n1382 ^ 1'b0 ;
  assign n6331 = n3500 ^ n2939 ^ 1'b0 ;
  assign n6332 = n221 | n6331 ;
  assign n6333 = ( ~n260 & n1883 ) | ( ~n260 & n2428 ) | ( n1883 & n2428 ) ;
  assign n6334 = n1972 & n6333 ;
  assign n6335 = n3348 & n6334 ;
  assign n6336 = n627 & n4763 ;
  assign n6337 = n130 & ~n2362 ;
  assign n6338 = n6337 ^ n2612 ^ 1'b0 ;
  assign n6339 = n3886 | n6338 ;
  assign n6340 = ( n4126 & ~n5239 ) | ( n4126 & n6339 ) | ( ~n5239 & n6339 ) ;
  assign n6341 = n1761 ^ n1210 ^ 1'b0 ;
  assign n6342 = ( ~n2720 & n3585 ) | ( ~n2720 & n6341 ) | ( n3585 & n6341 ) ;
  assign n6343 = n6342 ^ n3609 ^ 1'b0 ;
  assign n6344 = n360 | n5882 ;
  assign n6345 = n6344 ^ n35 ^ 1'b0 ;
  assign n6346 = ~n889 & n2124 ;
  assign n6347 = n471 | n3144 ;
  assign n6348 = n4573 | n6347 ;
  assign n6349 = n6348 ^ n3404 ^ 1'b0 ;
  assign n6350 = n5312 | n6349 ;
  assign n6351 = ~n3252 & n6350 ;
  assign n6352 = n3302 & n3312 ;
  assign n6353 = n35 | n700 ;
  assign n6355 = n957 | n3642 ;
  assign n6354 = n2781 & n5526 ;
  assign n6356 = n6355 ^ n6354 ^ 1'b0 ;
  assign n6357 = n1315 & n3432 ;
  assign n6358 = ( n4252 & n6356 ) | ( n4252 & ~n6357 ) | ( n6356 & ~n6357 ) ;
  assign n6359 = n6353 | n6358 ;
  assign n6360 = n6359 ^ n3395 ^ 1'b0 ;
  assign n6363 = ( ~n137 & n776 ) | ( ~n137 & n5107 ) | ( n776 & n5107 ) ;
  assign n6364 = n6363 ^ n3569 ^ 1'b0 ;
  assign n6365 = n5954 & n6364 ;
  assign n6361 = n2971 ^ n1953 ^ 1'b0 ;
  assign n6362 = ( n780 & n1048 ) | ( n780 & ~n6361 ) | ( n1048 & ~n6361 ) ;
  assign n6366 = n6365 ^ n6362 ^ n1522 ;
  assign n6367 = n884 | n3554 ;
  assign n6368 = n2427 & ~n6367 ;
  assign n6369 = n3489 | n6368 ;
  assign n6370 = n6369 ^ n3149 ^ n517 ;
  assign n6372 = n1246 & ~n4781 ;
  assign n6373 = n1040 | n6372 ;
  assign n6374 = n6373 ^ n2319 ^ 1'b0 ;
  assign n6371 = ~n102 & n2076 ;
  assign n6375 = n6374 ^ n6371 ^ 1'b0 ;
  assign n6376 = n4752 ^ n2745 ^ 1'b0 ;
  assign n6377 = n104 ^ n65 ^ 1'b0 ;
  assign n6378 = ~n1619 & n3749 ;
  assign n6379 = n6378 ^ n2289 ^ 1'b0 ;
  assign n6380 = ( n506 & n765 ) | ( n506 & ~n3244 ) | ( n765 & ~n3244 ) ;
  assign n6381 = n710 & n6380 ;
  assign n6382 = n4937 ^ n4653 ^ 1'b0 ;
  assign n6383 = n5796 ^ n1429 ^ n698 ;
  assign n6384 = n966 & ~n4887 ;
  assign n6385 = n4429 & ~n6384 ;
  assign n6386 = n2923 | n4467 ;
  assign n6387 = n1767 ^ n1262 ^ 1'b0 ;
  assign n6388 = n2170 & ~n5318 ;
  assign n6389 = ~n1507 & n4475 ;
  assign n6390 = n5037 & ~n6389 ;
  assign n6395 = n3059 ^ n2447 ^ 1'b0 ;
  assign n6396 = n408 & n6395 ;
  assign n6391 = n1232 | n3179 ;
  assign n6392 = n6391 ^ n3742 ^ 1'b0 ;
  assign n6393 = n1249 & n6392 ;
  assign n6394 = n5175 & n6393 ;
  assign n6397 = n6396 ^ n6394 ^ 1'b0 ;
  assign n6398 = n6105 & ~n6397 ;
  assign n6401 = ~n1723 & n6265 ;
  assign n6402 = ~n4002 & n6401 ;
  assign n6399 = ~n5142 & n5515 ;
  assign n6400 = n1464 | n6399 ;
  assign n6403 = n6402 ^ n6400 ^ 1'b0 ;
  assign n6404 = n1459 & n2821 ;
  assign n6405 = n2630 | n6404 ;
  assign n6406 = n3276 | n6405 ;
  assign n6407 = n5421 ^ n2674 ^ 1'b0 ;
  assign n6408 = n4445 ^ n2558 ^ 1'b0 ;
  assign n6409 = n1195 & n2421 ;
  assign n6410 = n2904 & ~n6409 ;
  assign n6411 = n6410 ^ n1764 ^ 1'b0 ;
  assign n6412 = n3479 ^ n3149 ^ n2591 ;
  assign n6413 = ( n1706 & n1736 ) | ( n1706 & ~n3260 ) | ( n1736 & ~n3260 ) ;
  assign n6414 = ~n871 & n6413 ;
  assign n6415 = n6412 | n6414 ;
  assign n6416 = n1751 | n3946 ;
  assign n6417 = n6416 ^ n2633 ^ 1'b0 ;
  assign n6418 = n4633 & n5139 ;
  assign n6419 = n4650 & n4711 ;
  assign n6420 = n6419 ^ n2535 ^ 1'b0 ;
  assign n6421 = n1024 & ~n2776 ;
  assign n6422 = n1335 ^ n1177 ^ 1'b0 ;
  assign n6423 = n3107 ^ n2190 ^ 1'b0 ;
  assign n6429 = n1124 & n3119 ;
  assign n6430 = n1746 & n6429 ;
  assign n6424 = ( x8 & x10 ) | ( x8 & n1339 ) | ( x10 & n1339 ) ;
  assign n6425 = n276 | n6424 ;
  assign n6426 = n6425 ^ n1875 ^ 1'b0 ;
  assign n6427 = ~n1768 & n6426 ;
  assign n6428 = n6427 ^ n4896 ^ 1'b0 ;
  assign n6431 = n6430 ^ n6428 ^ n3185 ;
  assign n6432 = n4880 ^ n2570 ^ 1'b0 ;
  assign n6433 = n1383 & ~n6432 ;
  assign n6440 = n4132 ^ n873 ^ n696 ;
  assign n6434 = n742 & n808 ;
  assign n6435 = ~n37 & n6434 ;
  assign n6436 = n848 & ~n6435 ;
  assign n6437 = n6436 ^ n6088 ^ 1'b0 ;
  assign n6438 = n3575 ^ n141 ^ 1'b0 ;
  assign n6439 = n6437 & ~n6438 ;
  assign n6441 = n6440 ^ n6439 ^ 1'b0 ;
  assign n6442 = n4002 ^ n2729 ^ 1'b0 ;
  assign n6443 = n3119 & ~n6442 ;
  assign n6444 = n5377 | n6443 ;
  assign n6445 = n1290 & ~n6368 ;
  assign n6446 = n6445 ^ n1371 ^ 1'b0 ;
  assign n6447 = n1616 & n4452 ;
  assign n6448 = n6447 ^ n1348 ^ 1'b0 ;
  assign n6449 = n696 & n6448 ;
  assign n6450 = n5631 & n6398 ;
  assign n6451 = n3248 & ~n3777 ;
  assign n6452 = n6451 ^ n438 ^ 1'b0 ;
  assign n6453 = n3934 ^ n3005 ^ 1'b0 ;
  assign n6454 = n1787 | n6453 ;
  assign n6455 = n151 & ~n3045 ;
  assign n6456 = n2541 ^ n1326 ^ 1'b0 ;
  assign n6457 = n6456 ^ n6013 ^ 1'b0 ;
  assign n6458 = n1825 & n4681 ;
  assign n6459 = n1104 | n3341 ;
  assign n6460 = n143 & ~n6459 ;
  assign n6461 = n6460 ^ n5128 ^ 1'b0 ;
  assign n6462 = n1823 | n6461 ;
  assign n6463 = n6458 & ~n6462 ;
  assign n6464 = n6463 ^ n3680 ^ 1'b0 ;
  assign n6465 = n736 ^ n126 ^ 1'b0 ;
  assign n6466 = n1737 & ~n6465 ;
  assign n6467 = ~n63 & n1959 ;
  assign n6468 = ~n947 & n6467 ;
  assign n6469 = ~n1327 & n3531 ;
  assign n6470 = ~n2294 & n6469 ;
  assign n6471 = n6470 ^ n2750 ^ 1'b0 ;
  assign n6472 = ~n6468 & n6471 ;
  assign n6473 = ~n6466 & n6472 ;
  assign n6476 = n2833 ^ n1346 ^ 1'b0 ;
  assign n6477 = n3333 & ~n6476 ;
  assign n6474 = n2561 ^ n1360 ^ n188 ;
  assign n6475 = n2790 | n6474 ;
  assign n6478 = n6477 ^ n6475 ^ 1'b0 ;
  assign n6479 = n2878 ^ n1841 ^ 1'b0 ;
  assign n6480 = n3693 & ~n6479 ;
  assign n6481 = n1155 & n1310 ;
  assign n6482 = n6481 ^ n3119 ^ n778 ;
  assign n6484 = ~n249 & n2699 ;
  assign n6485 = n6484 ^ n332 ^ 1'b0 ;
  assign n6486 = n811 & n2413 ;
  assign n6487 = ~n6485 & n6486 ;
  assign n6483 = ~n4698 & n4812 ;
  assign n6488 = n6487 ^ n6483 ^ 1'b0 ;
  assign n6489 = n278 & n4679 ;
  assign n6490 = n6489 ^ n3045 ^ 1'b0 ;
  assign n6491 = n6490 ^ n2827 ^ 1'b0 ;
  assign n6492 = ~n6424 & n6491 ;
  assign n6493 = n6492 ^ n1616 ^ 1'b0 ;
  assign n6494 = n5416 ^ n1824 ^ 1'b0 ;
  assign n6495 = n6493 | n6494 ;
  assign n6496 = n4988 ^ n3984 ^ n368 ;
  assign n6497 = n3825 ^ n3778 ^ 1'b0 ;
  assign n6498 = n5690 ^ n587 ^ 1'b0 ;
  assign n6499 = n4454 ^ n2810 ^ 1'b0 ;
  assign n6500 = n5036 & n6499 ;
  assign n6501 = n3805 ^ n1628 ^ 1'b0 ;
  assign n6502 = n2776 ^ n2474 ^ 1'b0 ;
  assign n6503 = n3909 & ~n6502 ;
  assign n6504 = ~n2123 & n6503 ;
  assign n6505 = n1839 & ~n6504 ;
  assign n6506 = n5224 | n6505 ;
  assign n6507 = n4381 ^ n3020 ^ 1'b0 ;
  assign n6508 = n166 & ~n6507 ;
  assign n6509 = n5559 ^ n2472 ^ 1'b0 ;
  assign n6510 = n5915 ^ n750 ^ 1'b0 ;
  assign n6511 = ~n6182 & n6510 ;
  assign n6512 = n6128 ^ n2231 ^ 1'b0 ;
  assign n6513 = n3719 & ~n6512 ;
  assign n6518 = n2199 | n6008 ;
  assign n6514 = n4204 ^ n2874 ^ n1974 ;
  assign n6515 = n5602 | n6514 ;
  assign n6516 = n1339 & ~n6515 ;
  assign n6517 = n6516 ^ n5781 ^ n5311 ;
  assign n6519 = n6518 ^ n6517 ^ 1'b0 ;
  assign n6520 = n5419 & n6519 ;
  assign n6521 = n6513 & n6520 ;
  assign n6522 = n2999 ^ n966 ^ 1'b0 ;
  assign n6523 = n2945 & ~n6522 ;
  assign n6524 = ~x10 & n368 ;
  assign n6525 = n5583 ^ n63 ^ 1'b0 ;
  assign n6526 = n803 & ~n6525 ;
  assign n6527 = n3835 & n6454 ;
  assign n6528 = n1402 ^ n37 ^ 1'b0 ;
  assign n6529 = n4084 & n6528 ;
  assign n6530 = n6529 ^ n3663 ^ 1'b0 ;
  assign n6531 = n6530 ^ n6336 ^ n143 ;
  assign n6532 = n4363 ^ n3591 ^ n2567 ;
  assign n6545 = ~n2360 & n2886 ;
  assign n6540 = n1179 ^ n999 ^ 1'b0 ;
  assign n6541 = n4608 & ~n6540 ;
  assign n6542 = n2653 | n6541 ;
  assign n6533 = ( n533 & n1210 ) | ( n533 & n4158 ) | ( n1210 & n4158 ) ;
  assign n6534 = n2596 & n5676 ;
  assign n6535 = ~n6533 & n6534 ;
  assign n6536 = n1112 ^ n294 ^ 1'b0 ;
  assign n6537 = n2413 | n6536 ;
  assign n6538 = n825 & n6537 ;
  assign n6539 = n6535 & n6538 ;
  assign n6543 = n6542 ^ n6539 ^ 1'b0 ;
  assign n6544 = n738 & ~n6543 ;
  assign n6546 = n6545 ^ n6544 ^ 1'b0 ;
  assign n6547 = n3478 | n6546 ;
  assign n6548 = ( ~n411 & n4812 ) | ( ~n411 & n5696 ) | ( n4812 & n5696 ) ;
  assign n6549 = ~n195 & n6548 ;
  assign n6550 = n6415 ^ n1367 ^ n1041 ;
  assign n6551 = n1861 | n3461 ;
  assign n6552 = n6551 ^ n6180 ^ 1'b0 ;
  assign n6553 = n744 ^ n341 ^ 1'b0 ;
  assign n6554 = n4976 & n6553 ;
  assign n6555 = n5561 ^ n4445 ^ n366 ;
  assign n6556 = n801 | n6555 ;
  assign n6557 = n1898 ^ n676 ^ 1'b0 ;
  assign n6558 = n38 & ~n2935 ;
  assign n6559 = n1709 | n6558 ;
  assign n6560 = n6559 ^ n5169 ^ 1'b0 ;
  assign n6561 = ( n2374 & ~n2855 ) | ( n2374 & n6560 ) | ( ~n2855 & n6560 ) ;
  assign n6563 = n2289 ^ n486 ^ 1'b0 ;
  assign n6564 = n884 | n6563 ;
  assign n6565 = ~n572 & n776 ;
  assign n6566 = n366 & n6565 ;
  assign n6567 = n6566 ^ n2104 ^ 1'b0 ;
  assign n6568 = n6564 & ~n6567 ;
  assign n6562 = ( n1357 & n1553 ) | ( n1357 & ~n4368 ) | ( n1553 & ~n4368 ) ;
  assign n6569 = n6568 ^ n6562 ^ n5461 ;
  assign n6571 = ( n886 & n1276 ) | ( n886 & n2692 ) | ( n1276 & n2692 ) ;
  assign n6570 = n4252 ^ n4149 ^ n3843 ;
  assign n6572 = n6571 ^ n6570 ^ n260 ;
  assign n6573 = ~n3661 & n6572 ;
  assign n6574 = n2836 & n6573 ;
  assign n6575 = n1079 | n6574 ;
  assign n6579 = n3236 | n4376 ;
  assign n6576 = ~n1503 & n2870 ;
  assign n6577 = n5331 ^ n375 ^ 1'b0 ;
  assign n6578 = n6576 & ~n6577 ;
  assign n6580 = n6579 ^ n6578 ^ 1'b0 ;
  assign n6581 = ~n3007 & n6580 ;
  assign n6582 = n6575 ^ n4846 ^ 1'b0 ;
  assign n6583 = n3548 ^ n951 ^ 1'b0 ;
  assign n6584 = ( n611 & ~n1340 ) | ( n611 & n2804 ) | ( ~n1340 & n2804 ) ;
  assign n6585 = ( n1279 & n6583 ) | ( n1279 & n6584 ) | ( n6583 & n6584 ) ;
  assign n6586 = n255 | n6585 ;
  assign n6587 = n6586 ^ n5985 ^ 1'b0 ;
  assign n6588 = n3217 ^ n2705 ^ 1'b0 ;
  assign n6589 = n1166 | n6588 ;
  assign n6590 = ( n2355 & n4097 ) | ( n2355 & n6589 ) | ( n4097 & n6589 ) ;
  assign n6591 = ( n186 & n3307 ) | ( n186 & n6590 ) | ( n3307 & n6590 ) ;
  assign n6592 = n6591 ^ n6503 ^ 1'b0 ;
  assign n6593 = n1262 & n6592 ;
  assign n6594 = n1456 ^ n263 ^ 1'b0 ;
  assign n6595 = n100 & ~n6594 ;
  assign n6596 = n6229 & n6595 ;
  assign n6597 = ( n744 & ~n759 ) | ( n744 & n1079 ) | ( ~n759 & n1079 ) ;
  assign n6598 = n3361 | n6597 ;
  assign n6599 = n6598 ^ n6126 ^ n637 ;
  assign n6600 = n3890 & ~n6599 ;
  assign n6601 = ~n957 & n4025 ;
  assign n6602 = ~n2903 & n5714 ;
  assign n6603 = n6602 ^ n4737 ^ n3762 ;
  assign n6604 = ~n209 & n6603 ;
  assign n6605 = n6604 ^ n780 ^ 1'b0 ;
  assign n6606 = n6167 ^ n3201 ^ 1'b0 ;
  assign n6607 = n554 & n3281 ;
  assign n6608 = n136 & ~n2242 ;
  assign n6609 = n4880 ^ n3749 ^ 1'b0 ;
  assign n6610 = ~n6608 & n6609 ;
  assign n6611 = n6610 ^ n1893 ^ 1'b0 ;
  assign n6612 = ( n4543 & ~n6607 ) | ( n4543 & n6611 ) | ( ~n6607 & n6611 ) ;
  assign n6613 = ( n184 & n5483 ) | ( n184 & ~n6612 ) | ( n5483 & ~n6612 ) ;
  assign n6614 = n4545 ^ n2854 ^ 1'b0 ;
  assign n6615 = ( n2729 & n2844 ) | ( n2729 & ~n6614 ) | ( n2844 & ~n6614 ) ;
  assign n6616 = n5934 ^ n1951 ^ n908 ;
  assign n6617 = ~n4956 & n6616 ;
  assign n6618 = n6018 & n6617 ;
  assign n6619 = n510 & n4056 ;
  assign n6620 = n6619 ^ n2868 ^ 1'b0 ;
  assign n6621 = n5941 ^ n2934 ^ 1'b0 ;
  assign n6622 = n6620 | n6621 ;
  assign n6623 = ( n710 & n1081 ) | ( n710 & ~n4443 ) | ( n1081 & ~n4443 ) ;
  assign n6624 = n5109 & n6623 ;
  assign n6625 = n6624 ^ n2307 ^ 1'b0 ;
  assign n6626 = ~n3698 & n6625 ;
  assign n6627 = n6626 ^ n4877 ^ 1'b0 ;
  assign n6628 = n6562 ^ n6236 ^ 1'b0 ;
  assign n6629 = ~n1302 & n5016 ;
  assign n6630 = n381 & n2261 ;
  assign n6631 = n6527 ^ n2729 ^ 1'b0 ;
  assign n6632 = ~n104 & n6631 ;
  assign n6633 = n89 & n1579 ;
  assign n6634 = n6633 ^ n1315 ^ 1'b0 ;
  assign n6635 = n13 & ~n6634 ;
  assign n6636 = ~n131 & n6635 ;
  assign n6637 = n1124 ^ n1017 ^ 1'b0 ;
  assign n6638 = n875 & n6637 ;
  assign n6639 = n2631 | n6638 ;
  assign n6640 = ~n2232 & n3121 ;
  assign n6641 = n1234 & n1525 ;
  assign n6642 = n3740 & n5603 ;
  assign n6643 = n6642 ^ n2428 ^ 1'b0 ;
  assign n6644 = n2676 ^ n220 ^ 1'b0 ;
  assign n6645 = n6275 | n6644 ;
  assign n6646 = n6643 & ~n6645 ;
  assign n6647 = n2577 & ~n6646 ;
  assign n6648 = ( n2798 & ~n4099 ) | ( n2798 & n6647 ) | ( ~n4099 & n6647 ) ;
  assign n6649 = n6648 ^ n2951 ^ 1'b0 ;
  assign n6650 = n6632 & n6649 ;
  assign n6651 = n2986 & ~n3891 ;
  assign n6652 = n6651 ^ n4568 ^ 1'b0 ;
  assign n6653 = ( ~n1026 & n2022 ) | ( ~n1026 & n4563 ) | ( n2022 & n4563 ) ;
  assign n6654 = n6653 ^ n5447 ^ 1'b0 ;
  assign n6655 = n204 | n991 ;
  assign n6656 = n2544 | n6655 ;
  assign n6657 = n6654 & n6656 ;
  assign n6658 = ( n3800 & n5861 ) | ( n3800 & n6657 ) | ( n5861 & n6657 ) ;
  assign n6659 = n2868 & ~n5255 ;
  assign n6660 = n3528 ^ n957 ^ 1'b0 ;
  assign n6661 = n1365 | n1628 ;
  assign n6662 = n604 | n2229 ;
  assign n6663 = n1704 & n2826 ;
  assign n6664 = n6663 ^ n1461 ^ 1'b0 ;
  assign n6665 = n4747 & ~n6664 ;
  assign n6666 = n6665 ^ n5259 ^ 1'b0 ;
  assign n6667 = n421 & n5848 ;
  assign n6668 = n3824 ^ n763 ^ 1'b0 ;
  assign n6669 = n6668 ^ n6599 ^ 1'b0 ;
  assign n6670 = n5205 & ~n6669 ;
  assign n6671 = n1836 ^ n394 ^ 1'b0 ;
  assign n6672 = ~n4397 & n5599 ;
  assign n6673 = n6672 ^ n5769 ^ 1'b0 ;
  assign n6674 = n940 & n3710 ;
  assign n6675 = n6674 ^ n2257 ^ 1'b0 ;
  assign n6676 = n6675 ^ n5628 ^ 1'b0 ;
  assign n6677 = n656 ^ n411 ^ 1'b0 ;
  assign n6678 = ~n4540 & n6677 ;
  assign n6679 = ( n698 & n1213 ) | ( n698 & n1439 ) | ( n1213 & n1439 ) ;
  assign n6680 = ~n32 & n6679 ;
  assign n6681 = ~n6678 & n6680 ;
  assign n6682 = ~n2233 & n5603 ;
  assign n6683 = n1520 & ~n6682 ;
  assign n6684 = n1854 ^ n249 ^ 1'b0 ;
  assign n6685 = n1523 & ~n6684 ;
  assign n6686 = n2889 & n6685 ;
  assign n6687 = n886 & ~n5501 ;
  assign n6688 = n1861 & ~n3170 ;
  assign n6689 = n6688 ^ n3033 ^ 1'b0 ;
  assign n6690 = n6689 ^ n2006 ^ 1'b0 ;
  assign n6691 = n1621 ^ n498 ^ n315 ;
  assign n6692 = n1463 | n6691 ;
  assign n6693 = n2064 & ~n6692 ;
  assign n6694 = ~n3730 & n6693 ;
  assign n6695 = ~n452 & n6694 ;
  assign n6696 = ~n906 & n957 ;
  assign n6697 = n57 & ~n3235 ;
  assign n6698 = n6697 ^ n2432 ^ 1'b0 ;
  assign n6699 = n6696 & ~n6698 ;
  assign n6700 = n2971 ^ n1241 ^ 1'b0 ;
  assign n6701 = n6700 ^ n612 ^ 1'b0 ;
  assign n6702 = n6699 | n6701 ;
  assign n6703 = ~n4153 & n4251 ;
  assign n6704 = n122 | n3592 ;
  assign n6705 = n1813 & ~n6704 ;
  assign n6706 = ~n3781 & n6705 ;
  assign n6707 = n3292 & n6706 ;
  assign n6708 = n4250 ^ n2034 ^ 1'b0 ;
  assign n6709 = n4700 & ~n6708 ;
  assign n6710 = x9 & n1454 ;
  assign n6711 = n521 | n4551 ;
  assign n6712 = n1895 & ~n6711 ;
  assign n6713 = n6712 ^ n194 ^ 1'b0 ;
  assign n6714 = n4889 ^ n1241 ^ 1'b0 ;
  assign n6715 = n6713 & ~n6714 ;
  assign n6716 = n6715 ^ n4925 ^ 1'b0 ;
  assign n6717 = n3004 & ~n3375 ;
  assign n6718 = n6717 ^ n5164 ^ n328 ;
  assign n6719 = n3850 ^ n2864 ^ 1'b0 ;
  assign n6720 = n3734 & n6719 ;
  assign n6721 = n6718 & n6720 ;
  assign n6722 = n6721 ^ n6392 ^ 1'b0 ;
  assign n6723 = n1177 ^ n261 ^ 1'b0 ;
  assign n6724 = n2192 | n5024 ;
  assign n6725 = n5645 | n6724 ;
  assign n6726 = ~n2339 & n5103 ;
  assign n6727 = n6726 ^ n1489 ^ 1'b0 ;
  assign n6728 = n3634 & n5898 ;
  assign n6729 = n6727 & n6728 ;
  assign n6730 = n5631 ^ n1527 ^ 1'b0 ;
  assign n6731 = n1093 | n6730 ;
  assign n6732 = n6716 ^ n3046 ^ n2156 ;
  assign n6735 = n2482 ^ n1131 ^ 1'b0 ;
  assign n6736 = n2582 & n6735 ;
  assign n6737 = n6736 ^ n4741 ^ n589 ;
  assign n6738 = n5930 & ~n6737 ;
  assign n6733 = n3861 | n5997 ;
  assign n6734 = n1226 & n6733 ;
  assign n6739 = n6738 ^ n6734 ^ 1'b0 ;
  assign n6740 = n4067 ^ n3357 ^ 1'b0 ;
  assign n6741 = n6740 ^ n2186 ^ 1'b0 ;
  assign n6742 = ~n886 & n3385 ;
  assign n6743 = n6742 ^ n3684 ^ 1'b0 ;
  assign n6744 = n6743 ^ n3393 ^ 1'b0 ;
  assign n6745 = ~n6741 & n6744 ;
  assign n6746 = n5022 | n6745 ;
  assign n6747 = n4663 ^ n20 ^ 1'b0 ;
  assign n6748 = n1453 & n5209 ;
  assign n6749 = n4018 ^ n2731 ^ 1'b0 ;
  assign n6750 = n2065 | n6749 ;
  assign n6751 = n6750 ^ n803 ^ 1'b0 ;
  assign n6752 = n3811 | n6751 ;
  assign n6753 = ( n3792 & ~n4446 ) | ( n3792 & n6752 ) | ( ~n4446 & n6752 ) ;
  assign n6754 = n3307 & n6753 ;
  assign n6755 = n4966 ^ n1805 ^ 1'b0 ;
  assign n6756 = n3332 & ~n6755 ;
  assign n6760 = n3372 & ~n3469 ;
  assign n6761 = ~n2799 & n6760 ;
  assign n6762 = n6761 ^ n1889 ^ 1'b0 ;
  assign n6757 = ~n2732 & n4559 ;
  assign n6758 = n249 & n6757 ;
  assign n6759 = n6758 ^ n3523 ^ 1'b0 ;
  assign n6763 = n6762 ^ n6759 ^ 1'b0 ;
  assign n6764 = n6756 & n6763 ;
  assign n6765 = n6764 ^ n2652 ^ 1'b0 ;
  assign n6766 = n101 & n6765 ;
  assign n6767 = ~n529 & n1200 ;
  assign n6768 = n3062 ^ n1326 ^ 1'b0 ;
  assign n6769 = ~n1891 & n5729 ;
  assign n6770 = n176 & n6769 ;
  assign n6771 = n4140 | n6770 ;
  assign n6773 = n4735 & n6638 ;
  assign n6774 = ~n6187 & n6773 ;
  assign n6772 = n4072 & n4637 ;
  assign n6775 = n6774 ^ n6772 ^ 1'b0 ;
  assign n6776 = n6775 ^ n2775 ^ n1412 ;
  assign n6777 = n3902 | n5870 ;
  assign n6778 = n6777 ^ n3769 ^ 1'b0 ;
  assign n6779 = ( n5139 & n6531 ) | ( n5139 & n6778 ) | ( n6531 & n6778 ) ;
  assign n6780 = n4727 ^ n996 ^ 1'b0 ;
  assign n6781 = ( n2666 & ~n5131 ) | ( n2666 & n6780 ) | ( ~n5131 & n6780 ) ;
  assign n6782 = n1503 | n3737 ;
  assign n6783 = n3365 & ~n6782 ;
  assign n6784 = n2906 & n6783 ;
  assign n6785 = n3295 ^ n1175 ^ 1'b0 ;
  assign n6786 = ~n1148 & n6785 ;
  assign n6787 = n6786 ^ n5419 ^ 1'b0 ;
  assign n6788 = n263 | n1682 ;
  assign n6789 = n6788 ^ n2405 ^ n1462 ;
  assign n6790 = n6789 ^ n2387 ^ n601 ;
  assign n6791 = n6790 ^ n1535 ^ 1'b0 ;
  assign n6792 = n2561 & n6791 ;
  assign n6793 = n2346 ^ n987 ^ n617 ;
  assign n6794 = n2492 & n6426 ;
  assign n6795 = ~n6793 & n6794 ;
  assign n6796 = n6795 ^ n5280 ^ 1'b0 ;
  assign n6797 = n1153 & n1355 ;
  assign n6798 = n6797 ^ n5285 ^ 1'b0 ;
  assign n6799 = n51 | n6798 ;
  assign n6800 = n661 & ~n6799 ;
  assign n6801 = n5896 & n6800 ;
  assign n6802 = n1461 ^ x11 ^ 1'b0 ;
  assign n6803 = ~n2451 & n6802 ;
  assign n6804 = ~n605 & n6803 ;
  assign n6805 = n2457 | n5678 ;
  assign n6806 = ~n6804 & n6805 ;
  assign n6807 = n493 & n1803 ;
  assign n6808 = n4120 ^ n2076 ^ 1'b0 ;
  assign n6809 = ( n4138 & n4781 ) | ( n4138 & ~n6808 ) | ( n4781 & ~n6808 ) ;
  assign n6815 = n369 ^ n151 ^ 1'b0 ;
  assign n6814 = n557 & n1056 ;
  assign n6816 = n6815 ^ n6814 ^ n5169 ;
  assign n6810 = ~n2732 & n5582 ;
  assign n6811 = n1148 & n6810 ;
  assign n6812 = n6811 ^ n829 ^ 1'b0 ;
  assign n6813 = n5289 | n6812 ;
  assign n6817 = n6816 ^ n6813 ^ 1'b0 ;
  assign n6818 = ~n6809 & n6817 ;
  assign n6819 = ~n6807 & n6818 ;
  assign n6820 = ~n1983 & n2701 ;
  assign n6821 = n2531 ^ n46 ^ 1'b0 ;
  assign n6822 = n2787 & ~n4841 ;
  assign n6823 = n6822 ^ n5140 ^ 1'b0 ;
  assign n6824 = n165 & n1706 ;
  assign n6825 = ~n530 & n6824 ;
  assign n6826 = n255 & n609 ;
  assign n6827 = n6825 & n6826 ;
  assign n6828 = n1818 | n6827 ;
  assign n6829 = n6828 ^ n5877 ^ 1'b0 ;
  assign n6830 = n6094 & n6249 ;
  assign n6831 = n1135 & n6830 ;
  assign n6834 = n664 & n1932 ;
  assign n6835 = ~n475 & n6834 ;
  assign n6832 = n491 & n1647 ;
  assign n6833 = n206 & n6832 ;
  assign n6836 = n6835 ^ n6833 ^ 1'b0 ;
  assign n6837 = ~n4044 & n6836 ;
  assign n6838 = n42 | n710 ;
  assign n6839 = n6837 | n6838 ;
  assign n6840 = n5103 ^ n1169 ^ 1'b0 ;
  assign n6841 = n5760 & n6840 ;
  assign n6842 = n6215 ^ n2816 ^ 1'b0 ;
  assign n6843 = n694 | n6842 ;
  assign n6844 = n3946 & ~n6843 ;
  assign n6845 = n4954 ^ n2446 ^ n1095 ;
  assign n6846 = n1288 & ~n6845 ;
  assign n6847 = n2084 | n2277 ;
  assign n6848 = n6847 ^ n2286 ^ 1'b0 ;
  assign n6849 = n1900 & ~n4215 ;
  assign n6850 = n2469 ^ n1048 ^ 1'b0 ;
  assign n6851 = n5106 | n6850 ;
  assign n6852 = n6575 ^ n2779 ^ 1'b0 ;
  assign n6853 = n3214 ^ n2181 ^ 1'b0 ;
  assign n6854 = n5724 ^ n1140 ^ 1'b0 ;
  assign n6855 = n919 | n6854 ;
  assign n6856 = n471 & ~n6855 ;
  assign n6857 = n5638 & ~n6856 ;
  assign n6858 = ~x10 & n6857 ;
  assign n6864 = n2885 ^ n2806 ^ n631 ;
  assign n6859 = x9 & n958 ;
  assign n6860 = ~n3566 & n6859 ;
  assign n6861 = n4447 | n6860 ;
  assign n6862 = n6861 ^ n1597 ^ 1'b0 ;
  assign n6863 = n2886 & n6862 ;
  assign n6865 = n6864 ^ n6863 ^ 1'b0 ;
  assign n6871 = n1185 & ~n4796 ;
  assign n6868 = n5020 ^ n435 ^ 1'b0 ;
  assign n6869 = n5918 & ~n6868 ;
  assign n6866 = n3365 ^ n2058 ^ n235 ;
  assign n6867 = n6866 ^ n788 ^ 1'b0 ;
  assign n6870 = n6869 ^ n6867 ^ n1157 ;
  assign n6872 = n6871 ^ n6870 ^ n3064 ;
  assign n6873 = n3812 | n6206 ;
  assign n6874 = n4053 | n6215 ;
  assign n6877 = n3696 ^ n1189 ^ 1'b0 ;
  assign n6875 = n4632 ^ n2980 ^ 1'b0 ;
  assign n6876 = n6776 & ~n6875 ;
  assign n6878 = n6877 ^ n6876 ^ 1'b0 ;
  assign n6879 = n1100 | n3872 ;
  assign n6880 = ~n235 & n6879 ;
  assign n6881 = n5850 | n6880 ;
  assign n6882 = n6871 & ~n6881 ;
  assign n6883 = n971 ^ n43 ^ 1'b0 ;
  assign n6884 = n824 | n4915 ;
  assign n6885 = n6884 ^ n3158 ^ 1'b0 ;
  assign n6886 = n4286 | n6700 ;
  assign n6887 = n113 | n4202 ;
  assign n6888 = n6887 ^ n4331 ^ 1'b0 ;
  assign n6889 = n5919 ^ n5795 ^ n296 ;
  assign n6890 = n2021 | n6866 ;
  assign n6891 = ~n242 & n997 ;
  assign n6892 = n1276 & n6891 ;
  assign n6893 = n6890 & n6892 ;
  assign n6897 = n3876 & n6558 ;
  assign n6894 = ~n157 & n5325 ;
  assign n6895 = ~n6603 & n6894 ;
  assign n6896 = n6895 ^ n459 ^ 1'b0 ;
  assign n6898 = n6897 ^ n6896 ^ 1'b0 ;
  assign n6899 = n3698 ^ n3680 ^ 1'b0 ;
  assign n6900 = n5424 ^ n935 ^ 1'b0 ;
  assign n6901 = n6899 & n6900 ;
  assign n6902 = n4769 ^ n3034 ^ 1'b0 ;
  assign n6903 = n3284 ^ n2971 ^ 1'b0 ;
  assign n6904 = n98 | n303 ;
  assign n6905 = n3696 | n6904 ;
  assign n6906 = n6905 ^ n1436 ^ 1'b0 ;
  assign n6907 = ~n1081 & n3407 ;
  assign n6908 = ~n1762 & n6907 ;
  assign n6909 = ( n1028 & n5382 ) | ( n1028 & ~n6908 ) | ( n5382 & ~n6908 ) ;
  assign n6910 = n6909 ^ n4542 ^ 1'b0 ;
  assign n6913 = n592 & n1450 ;
  assign n6914 = n6913 ^ n1568 ^ 1'b0 ;
  assign n6911 = ~n576 & n1906 ;
  assign n6912 = n2059 & n6911 ;
  assign n6915 = n6914 ^ n6912 ^ 1'b0 ;
  assign n6916 = n3285 ^ n2650 ^ 1'b0 ;
  assign n6917 = ~n672 & n5447 ;
  assign n6918 = n491 & n911 ;
  assign n6919 = n6918 ^ n188 ^ 1'b0 ;
  assign n6920 = n6917 & ~n6919 ;
  assign n6921 = n844 & n6920 ;
  assign n6922 = ( n5119 & n5490 ) | ( n5119 & n6921 ) | ( n5490 & n6921 ) ;
  assign n6923 = n3180 ^ n100 ^ 1'b0 ;
  assign n6924 = n2828 ^ n1654 ^ 1'b0 ;
  assign n6925 = n3013 ^ n2722 ^ 1'b0 ;
  assign n6926 = n2696 ^ n485 ^ 1'b0 ;
  assign n6927 = ~n2986 & n6926 ;
  assign n6931 = n6553 ^ n1312 ^ 1'b0 ;
  assign n6932 = n1773 & ~n6931 ;
  assign n6933 = n6932 ^ n6802 ^ 1'b0 ;
  assign n6934 = n6933 ^ n3101 ^ 1'b0 ;
  assign n6929 = n3113 ^ n1751 ^ n364 ;
  assign n6928 = n464 & ~n4086 ;
  assign n6930 = n6929 ^ n6928 ^ 1'b0 ;
  assign n6935 = n6934 ^ n6930 ^ 1'b0 ;
  assign n6936 = n6935 ^ n5958 ^ 1'b0 ;
  assign n6937 = n6927 & n6936 ;
  assign n6938 = n6937 ^ n2813 ^ 1'b0 ;
  assign n6939 = n2811 ^ n1407 ^ n866 ;
  assign n6940 = ( n3658 & n3928 ) | ( n3658 & n6939 ) | ( n3928 & n6939 ) ;
  assign n6941 = n6940 ^ n5978 ^ n2429 ;
  assign n6942 = n3690 ^ n3636 ^ 1'b0 ;
  assign n6943 = n4769 & n4880 ;
  assign n6944 = n951 | n6943 ;
  assign n6945 = n6944 ^ n1740 ^ 1'b0 ;
  assign n6946 = n4425 ^ n2002 ^ 1'b0 ;
  assign n6947 = n6856 | n6946 ;
  assign n6948 = n2813 | n6947 ;
  assign n6949 = n3738 ^ n3592 ^ 1'b0 ;
  assign n6950 = n1423 | n3772 ;
  assign n6951 = n6949 & ~n6950 ;
  assign n6952 = n6951 ^ n1928 ^ 1'b0 ;
  assign n6953 = n82 & n6952 ;
  assign n6954 = n2697 & n6953 ;
  assign n6955 = n2177 | n2808 ;
  assign n6956 = n6142 ^ n3293 ^ 1'b0 ;
  assign n6957 = n6956 ^ n3637 ^ n2794 ;
  assign n6958 = n6957 ^ n2201 ^ n510 ;
  assign n6959 = n1178 & n2431 ;
  assign n6960 = n6959 ^ n2906 ^ 1'b0 ;
  assign n6961 = n6438 | n6960 ;
  assign n6962 = n3237 | n6961 ;
  assign n6963 = n2821 ^ n2048 ^ 1'b0 ;
  assign n6964 = n1668 | n6963 ;
  assign n6965 = n6964 ^ n2807 ^ 1'b0 ;
  assign n6966 = n3051 & ~n4340 ;
  assign n6967 = n5106 & ~n6966 ;
  assign n6968 = n6967 ^ n6676 ^ 1'b0 ;
  assign n6969 = n6247 ^ n4403 ^ n2145 ;
  assign n6970 = n2635 ^ n2446 ^ 1'b0 ;
  assign n6971 = n2049 & n6970 ;
  assign n6972 = ~n230 & n6971 ;
  assign n6973 = n6972 ^ n1245 ^ 1'b0 ;
  assign n6976 = n3305 ^ n205 ^ 1'b0 ;
  assign n6974 = n1921 | n6643 ;
  assign n6975 = n2836 | n6974 ;
  assign n6977 = n6976 ^ n6975 ^ 1'b0 ;
  assign n6978 = n4267 ^ n4191 ^ 1'b0 ;
  assign n6979 = ~n3567 & n6520 ;
  assign n6980 = n3255 | n6251 ;
  assign n6981 = n3898 | n6980 ;
  assign n6982 = n612 & ~n1662 ;
  assign n6983 = n6982 ^ n837 ^ 1'b0 ;
  assign n6984 = ~n4276 & n4574 ;
  assign n6985 = ~n6983 & n6984 ;
  assign n6986 = n513 | n5722 ;
  assign n6987 = n6985 & ~n6986 ;
  assign n6988 = n6987 ^ n1871 ^ 1'b0 ;
  assign n6991 = ~n841 & n3837 ;
  assign n6989 = n1817 & ~n3445 ;
  assign n6990 = n6989 ^ n2399 ^ 1'b0 ;
  assign n6992 = n6991 ^ n6990 ^ 1'b0 ;
  assign n6993 = n2783 ^ n473 ^ 1'b0 ;
  assign n6994 = ( n1581 & n1728 ) | ( n1581 & ~n6931 ) | ( n1728 & ~n6931 ) ;
  assign n6995 = n2944 & n3390 ;
  assign n6996 = n364 & ~n6995 ;
  assign n6997 = n3749 & ~n6996 ;
  assign n6998 = ~n6994 & n6997 ;
  assign n6999 = n6993 | n6998 ;
  assign n7000 = n6999 ^ n6931 ^ 1'b0 ;
  assign n7002 = n2405 ^ n1209 ^ 1'b0 ;
  assign n7003 = n7002 ^ n2651 ^ 1'b0 ;
  assign n7004 = n7003 ^ n3727 ^ 1'b0 ;
  assign n7001 = n1094 & ~n1240 ;
  assign n7005 = n7004 ^ n7001 ^ n838 ;
  assign n7006 = n1279 | n5526 ;
  assign n7007 = n3221 & ~n7006 ;
  assign n7008 = ~n4856 & n7007 ;
  assign n7009 = n2147 & n4345 ;
  assign n7010 = n299 | n7009 ;
  assign n7011 = n5471 ^ n4150 ^ n1848 ;
  assign n7012 = n7011 ^ n1630 ^ 1'b0 ;
  assign n7013 = ~n2445 & n7012 ;
  assign n7014 = n272 | n7013 ;
  assign n7015 = n1965 ^ n752 ^ 1'b0 ;
  assign n7016 = ~n2023 & n7015 ;
  assign n7017 = n586 & ~n761 ;
  assign n7018 = n7017 ^ n3290 ^ 1'b0 ;
  assign n7019 = n7016 & n7018 ;
  assign n7020 = n7019 ^ n165 ^ n57 ;
  assign n7021 = n601 & n7020 ;
  assign n7022 = n1622 ^ n744 ^ 1'b0 ;
  assign n7023 = n6435 & n7022 ;
  assign n7031 = n41 | n2538 ;
  assign n7024 = n2032 & n6674 ;
  assign n7025 = n7024 ^ n2036 ^ 1'b0 ;
  assign n7026 = n5191 ^ n1459 ^ 1'b0 ;
  assign n7027 = n7025 & ~n7026 ;
  assign n7028 = n7027 ^ n5107 ^ 1'b0 ;
  assign n7029 = n7028 ^ n5557 ^ 1'b0 ;
  assign n7030 = ~n4373 & n7029 ;
  assign n7032 = n7031 ^ n7030 ^ 1'b0 ;
  assign n7033 = n723 & ~n7032 ;
  assign n7034 = n317 & n1181 ;
  assign n7035 = n7034 ^ n5443 ^ n2858 ;
  assign n7036 = n3521 | n4713 ;
  assign n7037 = n7036 ^ n3633 ^ 1'b0 ;
  assign n7038 = n7037 ^ n3096 ^ 1'b0 ;
  assign n7039 = n4373 | n7038 ;
  assign n7040 = n4435 ^ n714 ^ 1'b0 ;
  assign n7041 = n2915 & ~n4785 ;
  assign n7042 = n5447 ^ n1171 ^ 1'b0 ;
  assign n7043 = ~n1487 & n7042 ;
  assign n7044 = n3245 ^ n2223 ^ 1'b0 ;
  assign n7045 = n656 | n7044 ;
  assign n7046 = n7045 ^ n1818 ^ 1'b0 ;
  assign n7047 = n4754 & ~n5282 ;
  assign n7050 = ~n1093 & n3398 ;
  assign n7051 = ~n1382 & n7050 ;
  assign n7052 = ( n1100 & ~n4118 ) | ( n1100 & n7051 ) | ( ~n4118 & n7051 ) ;
  assign n7048 = ~n3512 & n4127 ;
  assign n7049 = n7048 ^ n6098 ^ 1'b0 ;
  assign n7053 = n7052 ^ n7049 ^ 1'b0 ;
  assign n7054 = n381 & ~n7053 ;
  assign n7055 = n408 | n1213 ;
  assign n7056 = n7055 ^ n3326 ^ 1'b0 ;
  assign n7057 = n4056 ^ n3429 ^ 1'b0 ;
  assign n7058 = n4303 & n7057 ;
  assign n7059 = n7058 ^ n2239 ^ 1'b0 ;
  assign n7060 = n2081 & n7059 ;
  assign n7061 = n4099 ^ n1709 ^ 1'b0 ;
  assign n7062 = n2671 | n5855 ;
  assign n7063 = ~n7061 & n7062 ;
  assign n7064 = n5233 & n7063 ;
  assign n7065 = ( ~n1885 & n2445 ) | ( ~n1885 & n4207 ) | ( n2445 & n4207 ) ;
  assign n7066 = n6449 ^ n3087 ^ 1'b0 ;
  assign n7067 = n7065 | n7066 ;
  assign n7068 = n6535 ^ n1539 ^ 1'b0 ;
  assign n7069 = n46 & ~n7068 ;
  assign n7070 = n4199 & n7069 ;
  assign n7071 = n2337 | n7070 ;
  assign n7072 = n3911 & ~n7071 ;
  assign n7073 = n1596 & n3203 ;
  assign n7074 = n6510 & n7073 ;
  assign n7075 = n5402 ^ n3231 ^ 1'b0 ;
  assign n7076 = n491 & ~n7075 ;
  assign n7077 = ~n25 & n2291 ;
  assign n7078 = n5282 ^ n1249 ^ 1'b0 ;
  assign n7079 = n6075 ^ n4171 ^ 1'b0 ;
  assign n7080 = n2770 & ~n7079 ;
  assign n7081 = n2503 ^ n2027 ^ n1734 ;
  assign n7082 = ( n135 & ~n2461 ) | ( n135 & n3415 ) | ( ~n2461 & n3415 ) ;
  assign n7083 = n7081 | n7082 ;
  assign n7084 = n2966 & ~n7083 ;
  assign n7085 = ~n1000 & n4770 ;
  assign n7086 = n7084 & n7085 ;
  assign n7087 = n656 | n2826 ;
  assign n7088 = n2176 & ~n7087 ;
  assign n7089 = n7088 ^ n5033 ^ 1'b0 ;
  assign n7090 = n355 | n7089 ;
  assign n7091 = n937 | n7090 ;
  assign n7092 = n4890 ^ n4426 ^ 1'b0 ;
  assign n7093 = n2529 & ~n4646 ;
  assign n7094 = n2107 & n7093 ;
  assign n7095 = n3671 | n6707 ;
  assign n7096 = n7095 ^ n4497 ^ 1'b0 ;
  assign n7097 = ( n4545 & n7094 ) | ( n4545 & n7096 ) | ( n7094 & n7096 ) ;
  assign n7098 = ( n4397 & n7092 ) | ( n4397 & ~n7097 ) | ( n7092 & ~n7097 ) ;
  assign n7099 = ( n530 & n3310 ) | ( n530 & n3749 ) | ( n3310 & n3749 ) ;
  assign n7100 = n5661 & n7099 ;
  assign n7101 = n756 & n7100 ;
  assign n7102 = ~n6516 & n7101 ;
  assign n7103 = n7069 ^ n1751 ^ n1612 ;
  assign n7113 = n6125 ^ n3179 ^ 1'b0 ;
  assign n7112 = n3610 ^ n1724 ^ n652 ;
  assign n7105 = n1293 ^ n1286 ^ 1'b0 ;
  assign n7106 = n2237 | n7105 ;
  assign n7107 = n1993 | n7106 ;
  assign n7108 = n7107 ^ n3704 ^ 1'b0 ;
  assign n7109 = n3382 & ~n7108 ;
  assign n7110 = n375 & n7109 ;
  assign n7104 = n1068 ^ n334 ^ 1'b0 ;
  assign n7111 = n7110 ^ n7104 ^ 1'b0 ;
  assign n7114 = n7113 ^ n7112 ^ n7111 ;
  assign n7115 = n2347 ^ n2067 ^ 1'b0 ;
  assign n7116 = n5354 ^ n3010 ^ 1'b0 ;
  assign n7117 = ~n7115 & n7116 ;
  assign n7118 = n5760 & n7117 ;
  assign n7119 = ( n777 & n2414 ) | ( n777 & ~n2546 ) | ( n2414 & ~n2546 ) ;
  assign n7120 = n510 & n4047 ;
  assign n7121 = ( n631 & n1467 ) | ( n631 & ~n2080 ) | ( n1467 & ~n2080 ) ;
  assign n7122 = n7121 ^ n48 ^ 1'b0 ;
  assign n7123 = n7122 ^ n1698 ^ 1'b0 ;
  assign n7124 = n7123 ^ n1877 ^ 1'b0 ;
  assign n7125 = n2495 | n7124 ;
  assign n7132 = n1940 & n5599 ;
  assign n7133 = n749 & n7132 ;
  assign n7126 = n165 & ~n742 ;
  assign n7127 = n1664 & ~n7126 ;
  assign n7128 = n7127 ^ n1262 ^ 1'b0 ;
  assign n7129 = n7128 ^ n3634 ^ 1'b0 ;
  assign n7130 = n6243 | n7129 ;
  assign n7131 = ~n4690 & n7130 ;
  assign n7134 = n7133 ^ n7131 ^ 1'b0 ;
  assign n7135 = ~n1317 & n4232 ;
  assign n7136 = n3125 & ~n7025 ;
  assign n7137 = n7136 ^ n2836 ^ n2556 ;
  assign n7138 = n1419 | n7137 ;
  assign n7139 = n2241 & ~n5641 ;
  assign n7140 = ~n780 & n7139 ;
  assign n7141 = n1035 ^ n734 ^ 1'b0 ;
  assign n7142 = n5814 | n7141 ;
  assign n7143 = n256 ^ x8 ^ 1'b0 ;
  assign n7144 = n1843 & n7143 ;
  assign n7145 = n6899 & n7144 ;
  assign n7146 = ~n2747 & n7145 ;
  assign n7147 = n1499 & ~n1505 ;
  assign n7148 = n249 & ~n7098 ;
  assign n7149 = ~n7147 & n7148 ;
  assign n7150 = n1807 & ~n2556 ;
  assign n7151 = n3397 ^ n1506 ^ 1'b0 ;
  assign n7152 = n3313 & ~n7151 ;
  assign n7153 = n7152 ^ n1859 ^ 1'b0 ;
  assign n7154 = n7153 ^ n5088 ^ 1'b0 ;
  assign n7155 = n4435 ^ n644 ^ 1'b0 ;
  assign n7156 = n1367 | n7155 ;
  assign n7157 = n4647 & ~n7156 ;
  assign n7158 = n7154 & n7157 ;
  assign n7159 = n2334 & ~n2974 ;
  assign n7160 = n500 | n4072 ;
  assign n7161 = n7159 & ~n7160 ;
  assign n7162 = n3773 & n5389 ;
  assign n7163 = ~n2828 & n7162 ;
  assign n7164 = n1237 & n2541 ;
  assign n7165 = n7163 | n7164 ;
  assign n7166 = ( n2561 & ~n3775 ) | ( n2561 & n5436 ) | ( ~n3775 & n5436 ) ;
  assign n7167 = n7166 ^ n1718 ^ n409 ;
  assign n7168 = ( n276 & n1175 ) | ( n276 & ~n3296 ) | ( n1175 & ~n3296 ) ;
  assign n7169 = n2384 & n7168 ;
  assign n7170 = n4654 & ~n4877 ;
  assign n7171 = n7170 ^ n2806 ^ 1'b0 ;
  assign n7172 = ~n787 & n7171 ;
  assign n7173 = n3912 & n7172 ;
  assign n7174 = n7169 & n7173 ;
  assign n7175 = n204 | n513 ;
  assign n7176 = n7175 ^ x0 ^ 1'b0 ;
  assign n7177 = n4173 ^ n2297 ^ 1'b0 ;
  assign n7178 = n7176 & n7177 ;
  assign n7179 = n7178 ^ n3318 ^ 1'b0 ;
  assign n7180 = n2510 & ~n7179 ;
  assign n7181 = ( n2859 & n5348 ) | ( n2859 & n6722 ) | ( n5348 & n6722 ) ;
  assign n7182 = ( n4523 & ~n5229 ) | ( n4523 & n7181 ) | ( ~n5229 & n7181 ) ;
  assign n7183 = n777 & n2972 ;
  assign n7184 = ~n1944 & n7183 ;
  assign n7185 = ~n5526 & n7184 ;
  assign n7186 = n6337 ^ n833 ^ 1'b0 ;
  assign n7187 = n7186 ^ n1167 ^ 1'b0 ;
  assign n7188 = n2736 & ~n7187 ;
  assign n7189 = ~n4980 & n6765 ;
  assign n7191 = ~n745 & n2636 ;
  assign n7192 = n1360 & n7191 ;
  assign n7190 = n4728 ^ n1031 ^ 1'b0 ;
  assign n7193 = n7192 ^ n7190 ^ 1'b0 ;
  assign n7194 = n1419 & n3521 ;
  assign n7195 = n1754 | n4529 ;
  assign n7196 = n2181 ^ n1241 ^ 1'b0 ;
  assign n7197 = n588 & n1506 ;
  assign n7198 = ~n306 & n1934 ;
  assign n7199 = n7198 ^ n1433 ^ 1'b0 ;
  assign n7200 = n6412 | n7199 ;
  assign n7201 = n4745 | n7200 ;
  assign n7202 = n7201 ^ n818 ^ 1'b0 ;
  assign n7203 = n7197 & ~n7202 ;
  assign n7204 = n7203 ^ n2492 ^ 1'b0 ;
  assign n7205 = n6289 & n7204 ;
  assign n7206 = n1959 & n3874 ;
  assign n7207 = ~n7205 & n7206 ;
  assign n7208 = ( n3784 & ~n5239 ) | ( n3784 & n7207 ) | ( ~n5239 & n7207 ) ;
  assign n7209 = n2496 & n6157 ;
  assign n7210 = n2195 & n7209 ;
  assign n7211 = n7210 ^ n1412 ^ 1'b0 ;
  assign n7212 = n3607 & n7211 ;
  assign n7213 = n7212 ^ n5785 ^ 1'b0 ;
  assign n7214 = n4237 & ~n4939 ;
  assign n7215 = n1958 ^ n1278 ^ n1063 ;
  assign n7216 = ~n6146 & n7215 ;
  assign n7217 = n4343 ^ n1527 ^ 1'b0 ;
  assign n7218 = n3561 | n7217 ;
  assign n7219 = n6243 ^ n3842 ^ 1'b0 ;
  assign n7220 = n464 & n1348 ;
  assign n7221 = n2452 & n7220 ;
  assign n7222 = n4786 ^ n1216 ^ x10 ;
  assign n7223 = n7222 ^ n3799 ^ 1'b0 ;
  assign n7224 = n4214 ^ n221 ^ 1'b0 ;
  assign n7225 = n5107 & ~n7224 ;
  assign n7226 = n2906 & n4799 ;
  assign n7227 = n157 | n1531 ;
  assign n7228 = ~n142 & n6503 ;
  assign n7229 = n7227 & n7228 ;
  assign n7230 = ~n866 & n7229 ;
  assign n7231 = n150 | n2246 ;
  assign n7232 = n4275 ^ n3119 ^ 1'b0 ;
  assign n7233 = n283 & n7232 ;
  assign n7234 = n6205 & n7233 ;
  assign n7235 = n7234 ^ n4390 ^ 1'b0 ;
  assign n7236 = n4552 ^ n2055 ^ n1627 ;
  assign n7237 = n2731 ^ n1181 ^ 1'b0 ;
  assign n7238 = n7236 & n7237 ;
  assign n7239 = n7238 ^ n171 ^ 1'b0 ;
  assign n7240 = ( n698 & n809 ) | ( n698 & ~n2532 ) | ( n809 & ~n2532 ) ;
  assign n7241 = n3073 ^ n1022 ^ 1'b0 ;
  assign n7242 = ~n7240 & n7241 ;
  assign n7243 = n7242 ^ n5004 ^ n517 ;
  assign n7247 = n2902 ^ n2378 ^ 1'b0 ;
  assign n7248 = n6985 | n7247 ;
  assign n7244 = n1771 | n4018 ;
  assign n7245 = ( n356 & n383 ) | ( n356 & ~n706 ) | ( n383 & ~n706 ) ;
  assign n7246 = ~n7244 & n7245 ;
  assign n7249 = n7248 ^ n7246 ^ 1'b0 ;
  assign n7250 = n1917 & n7249 ;
  assign n7251 = n1734 & ~n1804 ;
  assign n7252 = n3851 ^ n572 ^ 1'b0 ;
  assign n7253 = n1051 & ~n4345 ;
  assign n7254 = n1710 & ~n1907 ;
  assign n7255 = n7254 ^ n5996 ^ 1'b0 ;
  assign n7256 = ~n705 & n3753 ;
  assign n7257 = n3663 & ~n6029 ;
  assign n7258 = ~n7256 & n7257 ;
  assign n7259 = ~n3294 & n7258 ;
  assign n7260 = n1826 & ~n2325 ;
  assign n7261 = ~n2786 & n4487 ;
  assign n7262 = n5748 ^ n3483 ^ 1'b0 ;
  assign n7263 = n7262 ^ n2162 ^ 1'b0 ;
  assign n7264 = n7261 & n7263 ;
  assign n7265 = n2055 ^ n870 ^ 1'b0 ;
  assign n7266 = n4285 ^ n1794 ^ 1'b0 ;
  assign n7267 = n7265 & n7266 ;
  assign n7268 = n5781 ^ n2592 ^ 1'b0 ;
  assign n7269 = n6864 ^ n1092 ^ 1'b0 ;
  assign n7270 = n1036 & ~n1410 ;
  assign n7271 = n882 | n7270 ;
  assign n7272 = ~n1677 & n2330 ;
  assign n7273 = ~n61 & n7272 ;
  assign n7274 = n7273 ^ n4402 ^ 1'b0 ;
  assign n7275 = n2922 & ~n7274 ;
  assign n7276 = n7275 ^ n2047 ^ n1518 ;
  assign n7277 = n6748 ^ n2483 ^ 1'b0 ;
  assign n7278 = n7276 | n7277 ;
  assign n7279 = n1484 ^ n590 ^ 1'b0 ;
  assign n7280 = n1348 & ~n7279 ;
  assign n7281 = n191 | n2971 ;
  assign n7282 = n7281 ^ n2495 ^ 1'b0 ;
  assign n7283 = n7282 ^ n4067 ^ 1'b0 ;
  assign n7284 = n2595 ^ n840 ^ 1'b0 ;
  assign n7285 = n7284 ^ n4405 ^ n104 ;
  assign n7286 = n839 & n3409 ;
  assign n7287 = ( n4512 & n5276 ) | ( n4512 & n7286 ) | ( n5276 & n7286 ) ;
  assign n7288 = ( ~n7283 & n7285 ) | ( ~n7283 & n7287 ) | ( n7285 & n7287 ) ;
  assign n7291 = ~n2405 & n2411 ;
  assign n7289 = ( ~n477 & n548 ) | ( ~n477 & n3413 ) | ( n548 & n3413 ) ;
  assign n7290 = n2169 & n7289 ;
  assign n7292 = n7291 ^ n7290 ^ 1'b0 ;
  assign n7293 = ~n112 & n5713 ;
  assign n7294 = ~n968 & n3298 ;
  assign n7295 = n716 & n7294 ;
  assign n7296 = n6348 ^ n6319 ^ n4549 ;
  assign n7297 = n5969 & ~n6178 ;
  assign n7298 = n4777 | n6030 ;
  assign n7299 = n3909 ^ n63 ^ 1'b0 ;
  assign n7300 = n1169 & n7299 ;
  assign n7301 = n7300 ^ n1166 ^ 1'b0 ;
  assign n7302 = n6272 | n7301 ;
  assign n7303 = n4617 ^ n2489 ^ 1'b0 ;
  assign n7304 = n1115 | n2699 ;
  assign n7305 = n7304 ^ n816 ^ 1'b0 ;
  assign n7306 = n6914 & ~n7305 ;
  assign n7307 = n7306 ^ n1200 ^ 1'b0 ;
  assign n7308 = ~n1772 & n2827 ;
  assign n7309 = n1237 & n4793 ;
  assign n7310 = n7309 ^ n5580 ^ 1'b0 ;
  assign n7311 = ~n7308 & n7310 ;
  assign n7312 = n7311 ^ n4147 ^ 1'b0 ;
  assign n7313 = n7312 ^ n2471 ^ 1'b0 ;
  assign n7314 = n4140 & n7313 ;
  assign n7317 = n6384 ^ n2207 ^ n865 ;
  assign n7315 = n318 & ~n5692 ;
  assign n7316 = n750 | n7315 ;
  assign n7318 = n7317 ^ n7316 ^ 1'b0 ;
  assign n7319 = n2092 & n6871 ;
  assign n7320 = n5174 ^ n4138 ^ n2680 ;
  assign n7321 = n4432 & n7320 ;
  assign n7322 = n7321 ^ n7106 ^ 1'b0 ;
  assign n7323 = ~n738 & n7322 ;
  assign n7324 = ~n7319 & n7323 ;
  assign n7325 = n1035 ^ n771 ^ n718 ;
  assign n7326 = n5475 & ~n7325 ;
  assign n7327 = n4844 & ~n7326 ;
  assign n7328 = n7327 ^ n2583 ^ n624 ;
  assign n7329 = n1553 | n4315 ;
  assign n7330 = n7329 ^ n4469 ^ 1'b0 ;
  assign n7331 = n275 ^ n122 ^ 1'b0 ;
  assign n7332 = ~n888 & n7331 ;
  assign n7333 = n5037 | n7332 ;
  assign n7334 = n3505 | n7333 ;
  assign n7335 = n2808 ^ n1728 ^ 1'b0 ;
  assign n7336 = n1710 & ~n2027 ;
  assign n7337 = ~n2463 & n7336 ;
  assign n7338 = n506 | n2655 ;
  assign n7339 = ~n946 & n7338 ;
  assign n7340 = n1374 & n7339 ;
  assign n7341 = n2731 & ~n7340 ;
  assign n7342 = n7337 & n7341 ;
  assign n7343 = n3579 ^ n596 ^ 1'b0 ;
  assign n7344 = n7342 | n7343 ;
  assign n7345 = n7335 | n7344 ;
  assign n7346 = ~n63 & n1167 ;
  assign n7347 = n7346 ^ n1809 ^ 1'b0 ;
  assign n7348 = n7347 ^ n2435 ^ n53 ;
  assign n7349 = n7348 ^ n3193 ^ n496 ;
  assign n7350 = ( ~n169 & n2257 ) | ( ~n169 & n4475 ) | ( n2257 & n4475 ) ;
  assign n7351 = n99 & ~n411 ;
  assign n7352 = n7351 ^ n525 ^ 1'b0 ;
  assign n7353 = n7352 ^ n1832 ^ 1'b0 ;
  assign n7354 = n1415 & ~n7353 ;
  assign n7355 = n2799 & ~n6993 ;
  assign n7356 = ~n7354 & n7355 ;
  assign n7357 = n473 & ~n7356 ;
  assign n7359 = n4233 ^ n2152 ^ 1'b0 ;
  assign n7360 = n4538 & ~n7359 ;
  assign n7358 = ~n4434 & n6471 ;
  assign n7361 = n7360 ^ n7358 ^ n4285 ;
  assign n7362 = ~n1702 & n3732 ;
  assign n7363 = n7362 ^ n271 ^ 1'b0 ;
  assign n7364 = n7363 ^ n5418 ^ n4144 ;
  assign n7365 = ( n7357 & n7361 ) | ( n7357 & ~n7364 ) | ( n7361 & ~n7364 ) ;
  assign n7366 = n2176 ^ n2048 ^ n1716 ;
  assign n7367 = ~n7256 & n7366 ;
  assign n7368 = n3632 | n7367 ;
  assign n7369 = n6135 | n7368 ;
  assign n7370 = n7365 | n7369 ;
  assign n7371 = n436 & n6666 ;
  assign n7372 = n2853 ^ n1179 ^ 1'b0 ;
  assign n7373 = n3006 & ~n7372 ;
  assign n7374 = n7373 ^ n983 ^ 1'b0 ;
  assign n7375 = n3457 & ~n5637 ;
  assign n7376 = ~n7374 & n7375 ;
  assign n7377 = n2880 & ~n3567 ;
  assign n7378 = n3842 ^ n134 ^ 1'b0 ;
  assign n7379 = n6222 ^ n4204 ^ 1'b0 ;
  assign n7380 = n7378 & ~n7379 ;
  assign n7382 = ~n561 & n5913 ;
  assign n7383 = n7382 ^ n4493 ^ 1'b0 ;
  assign n7384 = n7383 ^ n2618 ^ n1397 ;
  assign n7381 = ~n376 & n582 ;
  assign n7385 = n7384 ^ n7381 ^ 1'b0 ;
  assign n7386 = n7385 ^ n4617 ^ 1'b0 ;
  assign n7387 = ~n80 & n256 ;
  assign n7388 = ( n666 & ~n3774 ) | ( n666 & n7387 ) | ( ~n3774 & n7387 ) ;
  assign n7389 = n1134 & ~n5163 ;
  assign n7390 = n7389 ^ n5037 ^ 1'b0 ;
  assign n7391 = n3365 | n7390 ;
  assign n7392 = ~n1712 & n2142 ;
  assign n7393 = ( ~n4202 & n4987 ) | ( ~n4202 & n7392 ) | ( n4987 & n7392 ) ;
  assign n7394 = n2657 | n6951 ;
  assign n7395 = n7393 & ~n7394 ;
  assign n7396 = n2012 & ~n7395 ;
  assign n7397 = n7396 ^ n2044 ^ 1'b0 ;
  assign n7398 = n2695 | n3432 ;
  assign n7399 = n7398 ^ n6555 ^ n2140 ;
  assign n7400 = ( n76 & ~n145 ) | ( n76 & n7399 ) | ( ~n145 & n7399 ) ;
  assign n7401 = n2164 & ~n7400 ;
  assign n7402 = n3642 ^ n2368 ^ 1'b0 ;
  assign n7403 = n2184 & n7402 ;
  assign n7404 = n7403 ^ n3680 ^ 1'b0 ;
  assign n7412 = n1324 | n1786 ;
  assign n7413 = n7412 ^ n2135 ^ 1'b0 ;
  assign n7408 = n3051 ^ n742 ^ 1'b0 ;
  assign n7409 = n922 & n1387 ;
  assign n7410 = ~n1851 & n7409 ;
  assign n7411 = n7408 & n7410 ;
  assign n7405 = n2892 ^ n536 ^ 1'b0 ;
  assign n7406 = n2995 & n3088 ;
  assign n7407 = n7405 & ~n7406 ;
  assign n7414 = n7413 ^ n7411 ^ n7407 ;
  assign n7415 = n999 | n4220 ;
  assign n7416 = n7415 ^ n4104 ^ 1'b0 ;
  assign n7417 = ~n3722 & n7416 ;
  assign n7418 = n63 | n394 ;
  assign n7419 = ( n1575 & ~n2758 ) | ( n1575 & n7418 ) | ( ~n2758 & n7418 ) ;
  assign n7420 = n1681 ^ n1231 ^ 1'b0 ;
  assign n7421 = n1073 | n7420 ;
  assign n7422 = n3790 | n7421 ;
  assign n7423 = n2264 & ~n7422 ;
  assign n7425 = n4555 & ~n5740 ;
  assign n7424 = n526 & n3932 ;
  assign n7426 = n7425 ^ n7424 ^ 1'b0 ;
  assign n7427 = n1959 & n3739 ;
  assign n7428 = n1426 & n2825 ;
  assign n7429 = n5391 | n6783 ;
  assign n7430 = n4195 | n7429 ;
  assign n7431 = n4641 ^ n965 ^ 1'b0 ;
  assign n7432 = n3797 | n7431 ;
  assign n7433 = n2418 & ~n6987 ;
  assign n7434 = ( n416 & n5806 ) | ( n416 & n5990 ) | ( n5806 & n5990 ) ;
  assign n7435 = n7434 ^ n3523 ^ n639 ;
  assign n7436 = x4 & ~n7435 ;
  assign n7437 = n3034 ^ n702 ^ 1'b0 ;
  assign n7438 = ~n6230 & n7437 ;
  assign n7441 = x10 | n1273 ;
  assign n7442 = n2460 & n2940 ;
  assign n7443 = n7442 ^ n611 ^ 1'b0 ;
  assign n7444 = ~n7441 & n7443 ;
  assign n7445 = n4563 & n7444 ;
  assign n7439 = n2584 ^ n702 ^ 1'b0 ;
  assign n7440 = n3567 | n7439 ;
  assign n7446 = n7445 ^ n7440 ^ n4143 ;
  assign n7447 = n6743 ^ n4757 ^ 1'b0 ;
  assign n7449 = n4204 ^ n947 ^ n639 ;
  assign n7450 = n2330 & n7449 ;
  assign n7448 = n3577 | n4270 ;
  assign n7451 = n7450 ^ n7448 ^ 1'b0 ;
  assign n7454 = n6246 ^ n4264 ^ n1223 ;
  assign n7452 = n1856 ^ n1744 ^ 1'b0 ;
  assign n7453 = n3584 & ~n7452 ;
  assign n7455 = n7454 ^ n7453 ^ 1'b0 ;
  assign n7456 = n5239 | n7455 ;
  assign n7457 = n7456 ^ n1562 ^ 1'b0 ;
  assign n7458 = n3191 & n7457 ;
  assign n7459 = ~n4120 & n7458 ;
  assign n7461 = ~n1311 & n4643 ;
  assign n7462 = n7461 ^ n3652 ^ 1'b0 ;
  assign n7463 = ~n3469 & n7462 ;
  assign n7460 = n5515 ^ n4537 ^ n4252 ;
  assign n7464 = n7463 ^ n7460 ^ n652 ;
  assign n7465 = ~n272 & n4914 ;
  assign n7466 = n1245 & ~n2403 ;
  assign n7467 = n1830 & n7466 ;
  assign n7468 = n7467 ^ n3784 ^ 1'b0 ;
  assign n7469 = n7062 & ~n7468 ;
  assign n7470 = ( n656 & n4232 ) | ( n656 & ~n5980 ) | ( n4232 & ~n5980 ) ;
  assign n7471 = n329 & ~n2304 ;
  assign n7472 = n728 ^ n154 ^ 1'b0 ;
  assign n7473 = n1280 & ~n7472 ;
  assign n7474 = n1621 & ~n7473 ;
  assign n7475 = ~n7471 & n7474 ;
  assign n7476 = n841 | n3541 ;
  assign n7477 = n7476 ^ n637 ^ 1'b0 ;
  assign n7478 = ~n4947 & n7477 ;
  assign n7479 = n772 | n1775 ;
  assign n7480 = n711 | n2672 ;
  assign n7481 = n5935 | n7480 ;
  assign n7482 = n7481 ^ n1387 ^ n650 ;
  assign n7483 = ( n6819 & n7479 ) | ( n6819 & ~n7482 ) | ( n7479 & ~n7482 ) ;
  assign n7484 = n1441 & n5314 ;
  assign n7485 = n4436 & ~n4730 ;
  assign n7486 = n6255 | n7485 ;
  assign n7487 = n7486 ^ n3539 ^ 1'b0 ;
  assign n7488 = n590 & ~n3573 ;
  assign n7489 = ( n368 & ~n556 ) | ( n368 & n2397 ) | ( ~n556 & n2397 ) ;
  assign n7490 = n6078 ^ n461 ^ 1'b0 ;
  assign n7491 = n7489 & ~n7490 ;
  assign n7492 = ~n5270 & n7491 ;
  assign n7493 = n294 | n7492 ;
  assign n7494 = n355 ^ n209 ^ 1'b0 ;
  assign n7495 = n7494 ^ n5515 ^ 1'b0 ;
  assign n7496 = ~x8 & n4288 ;
  assign n7497 = ~n1368 & n3505 ;
  assign n7498 = n7496 & n7497 ;
  assign n7499 = n5068 | n5255 ;
  assign n7500 = n1327 & n2073 ;
  assign n7501 = n7500 ^ n736 ^ 1'b0 ;
  assign n7502 = n177 & n7501 ;
  assign n7503 = ( n2037 & n4060 ) | ( n2037 & ~n7502 ) | ( n4060 & ~n7502 ) ;
  assign n7504 = n2504 | n5018 ;
  assign n7505 = n7503 | n7504 ;
  assign n7506 = n4715 ^ n753 ^ 1'b0 ;
  assign n7507 = n2080 | n6384 ;
  assign n7508 = n7507 ^ n6122 ^ 1'b0 ;
  assign n7511 = ( n260 & n4889 ) | ( n260 & ~n5618 ) | ( n4889 & ~n5618 ) ;
  assign n7509 = n6264 ^ n1878 ^ 1'b0 ;
  assign n7510 = n5478 | n7509 ;
  assign n7512 = n7511 ^ n7510 ^ 1'b0 ;
  assign n7513 = n4347 ^ n2944 ^ n814 ;
  assign n7514 = n7513 ^ n987 ^ 1'b0 ;
  assign n7515 = n887 ^ n777 ^ 1'b0 ;
  assign n7516 = n5059 & n7515 ;
  assign n7517 = n1490 & n7516 ;
  assign n7518 = ~n4322 & n7517 ;
  assign n7519 = n7518 ^ n7010 ^ 1'b0 ;
  assign n7520 = n3461 | n7519 ;
  assign n7521 = ~n43 & n368 ;
  assign n7522 = n7521 ^ n4608 ^ 1'b0 ;
  assign n7523 = ( ~n48 & n2602 ) | ( ~n48 & n7522 ) | ( n2602 & n7522 ) ;
  assign n7524 = n7523 ^ n4226 ^ 1'b0 ;
  assign n7525 = ~n2321 & n7524 ;
  assign n7526 = n7383 ^ n978 ^ n756 ;
  assign n7527 = n2657 & n3274 ;
  assign n7528 = n1824 & ~n5699 ;
  assign n7529 = n7528 ^ n2447 ^ 1'b0 ;
  assign n7530 = n7529 ^ n6660 ^ 1'b0 ;
  assign n7531 = n890 | n7290 ;
  assign n7532 = ( n526 & n1653 ) | ( n526 & ~n1798 ) | ( n1653 & ~n1798 ) ;
  assign n7533 = n4042 & n7532 ;
  assign n7534 = n4656 & n7533 ;
  assign n7538 = n4343 & n5750 ;
  assign n7539 = n7538 ^ n596 ^ 1'b0 ;
  assign n7535 = n1401 & ~n2348 ;
  assign n7536 = n7535 ^ n177 ^ 1'b0 ;
  assign n7537 = n813 | n7536 ;
  assign n7540 = n7539 ^ n7537 ^ 1'b0 ;
  assign n7541 = n1604 | n5578 ;
  assign n7542 = n4085 | n7541 ;
  assign n7543 = ( n1988 & ~n3217 ) | ( n1988 & n7542 ) | ( ~n3217 & n7542 ) ;
  assign n7544 = n4602 & ~n7118 ;
  assign n7545 = n3570 ^ n2156 ^ n1699 ;
  assign n7546 = ~n2768 & n7545 ;
  assign n7547 = n7546 ^ n5840 ^ 1'b0 ;
  assign n7548 = ~n153 & n7547 ;
  assign n7549 = n6135 & n7548 ;
  assign n7550 = n7549 ^ n7122 ^ 1'b0 ;
  assign n7551 = n3558 & ~n3630 ;
  assign n7552 = n448 ^ n23 ^ 1'b0 ;
  assign n7553 = ~n4210 & n7552 ;
  assign n7554 = ( n2747 & n4627 ) | ( n2747 & n7553 ) | ( n4627 & n7553 ) ;
  assign n7555 = ~n1505 & n3263 ;
  assign n7556 = n7555 ^ n1506 ^ 1'b0 ;
  assign n7557 = n334 | n999 ;
  assign n7558 = ( ~n3305 & n3923 ) | ( ~n3305 & n6380 ) | ( n3923 & n6380 ) ;
  assign n7559 = n7558 ^ n3998 ^ 1'b0 ;
  assign n7560 = n7557 | n7559 ;
  assign n7561 = n2710 | n7560 ;
  assign n7562 = n2552 ^ n1967 ^ 1'b0 ;
  assign n7563 = n1296 & n7562 ;
  assign n7564 = ~n570 & n1069 ;
  assign n7565 = n7564 ^ n702 ^ 1'b0 ;
  assign n7566 = n7565 ^ n2925 ^ 1'b0 ;
  assign n7567 = n4794 | n7566 ;
  assign n7568 = n581 & ~n7567 ;
  assign n7569 = n2374 & ~n2435 ;
  assign n7570 = n374 | n2712 ;
  assign n7571 = n7317 | n7570 ;
  assign n7572 = n7571 ^ n7081 ^ 1'b0 ;
  assign n7573 = n57 & n3120 ;
  assign n7574 = n670 & n7573 ;
  assign n7575 = ~n392 & n3925 ;
  assign n7576 = n3966 & n7575 ;
  assign n7577 = n7576 ^ n107 ^ 1'b0 ;
  assign n7578 = n484 | n1279 ;
  assign n7579 = n611 & ~n7578 ;
  assign n7580 = n7579 ^ n4024 ^ 1'b0 ;
  assign n7581 = n7580 ^ n2846 ^ 1'b0 ;
  assign n7582 = n38 & ~n3651 ;
  assign n7583 = ~x1 & n7582 ;
  assign n7584 = n7583 ^ n604 ^ 1'b0 ;
  assign n7585 = n2874 & ~n7584 ;
  assign n7586 = ( n7577 & n7581 ) | ( n7577 & ~n7585 ) | ( n7581 & ~n7585 ) ;
  assign n7587 = ~n874 & n7340 ;
  assign n7588 = ( n299 & ~n2177 ) | ( n299 & n7587 ) | ( ~n2177 & n7587 ) ;
  assign n7589 = ~n2569 & n3863 ;
  assign n7590 = n7589 ^ n1628 ^ 1'b0 ;
  assign n7591 = n1149 & ~n2815 ;
  assign n7592 = ~n4830 & n7591 ;
  assign n7593 = n7592 ^ n7013 ^ 1'b0 ;
  assign n7594 = n4770 & ~n7593 ;
  assign n7600 = n760 ^ n260 ^ 1'b0 ;
  assign n7601 = n7600 ^ n3146 ^ n73 ;
  assign n7595 = n2030 & ~n2039 ;
  assign n7596 = n1684 & n7595 ;
  assign n7597 = n4650 & ~n7596 ;
  assign n7598 = n7597 ^ n4690 ^ 1'b0 ;
  assign n7599 = n285 & n7598 ;
  assign n7602 = n7601 ^ n7599 ^ 1'b0 ;
  assign n7603 = ~n5941 & n7602 ;
  assign n7604 = n7603 ^ n5774 ^ 1'b0 ;
  assign n7605 = ~n3131 & n7604 ;
  assign n7606 = n3749 & ~n7285 ;
  assign n7607 = ~n1614 & n7606 ;
  assign n7608 = n82 & n4852 ;
  assign n7609 = ~n1193 & n7608 ;
  assign n7610 = n7607 & n7609 ;
  assign n7611 = n604 | n2857 ;
  assign n7612 = n7611 ^ n2446 ^ 1'b0 ;
  assign n7613 = n4115 & ~n4361 ;
  assign n7614 = n4250 ^ n1288 ^ 1'b0 ;
  assign n7615 = ~n471 & n2357 ;
  assign n7616 = n7615 ^ n4614 ^ 1'b0 ;
  assign n7617 = n7017 & n7616 ;
  assign n7618 = n1013 & ~n1903 ;
  assign n7619 = n7618 ^ n4010 ^ 1'b0 ;
  assign n7620 = n5182 & n7619 ;
  assign n7621 = n3812 ^ n2694 ^ 1'b0 ;
  assign n7622 = n7621 ^ n2474 ^ 1'b0 ;
  assign n7623 = n2241 & n6551 ;
  assign n7624 = n7623 ^ n2114 ^ 1'b0 ;
  assign n7625 = n7624 ^ n1548 ^ 1'b0 ;
  assign n7626 = ~n7622 & n7625 ;
  assign n7627 = n6355 ^ n5164 ^ n428 ;
  assign n7628 = n6488 ^ n1704 ^ 1'b0 ;
  assign n7629 = ~n3567 & n7628 ;
  assign n7630 = n5572 & n6205 ;
  assign n7631 = n213 & n890 ;
  assign n7632 = n360 | n5092 ;
  assign n7633 = n7632 ^ n959 ^ 1'b0 ;
  assign n7634 = ( n1292 & n2294 ) | ( n1292 & n4849 ) | ( n2294 & n4849 ) ;
  assign n7635 = n7634 ^ n1861 ^ 1'b0 ;
  assign n7637 = ~n523 & n1810 ;
  assign n7638 = n7637 ^ n1959 ^ 1'b0 ;
  assign n7636 = ~n448 & n7087 ;
  assign n7639 = n7638 ^ n7636 ^ 1'b0 ;
  assign n7640 = n1471 & n2758 ;
  assign n7641 = n7640 ^ n1538 ^ 1'b0 ;
  assign n7642 = n1327 & ~n4880 ;
  assign n7643 = ( n7622 & ~n7641 ) | ( n7622 & n7642 ) | ( ~n7641 & n7642 ) ;
  assign n7644 = n7643 ^ n4001 ^ 1'b0 ;
  assign n7645 = n4016 ^ n533 ^ 1'b0 ;
  assign n7646 = ( n3397 & n5554 ) | ( n3397 & n7645 ) | ( n5554 & n7645 ) ;
  assign n7647 = ~n1695 & n7646 ;
  assign n7648 = n7647 ^ n2949 ^ 1'b0 ;
  assign n7649 = x4 & n951 ;
  assign n7650 = n648 & n7649 ;
  assign n7651 = n7648 & n7650 ;
  assign n7652 = n7651 ^ n761 ^ 1'b0 ;
  assign n7653 = n4171 & n5756 ;
  assign n7654 = n2081 ^ n1240 ^ 1'b0 ;
  assign n7655 = n1919 ^ n799 ^ 1'b0 ;
  assign n7656 = n780 & ~n7655 ;
  assign n7657 = n108 & ~n3075 ;
  assign n7658 = n1245 | n1766 ;
  assign n7659 = ( n254 & n7657 ) | ( n254 & n7658 ) | ( n7657 & n7658 ) ;
  assign n7660 = n1666 & ~n4153 ;
  assign n7661 = n7660 ^ n6759 ^ 1'b0 ;
  assign n7662 = n893 & ~n6205 ;
  assign n7663 = n7662 ^ n2214 ^ 1'b0 ;
  assign n7664 = n1781 & ~n3565 ;
  assign n7665 = n7664 ^ n276 ^ 1'b0 ;
  assign n7666 = ( n2101 & ~n7122 ) | ( n2101 & n7665 ) | ( ~n7122 & n7665 ) ;
  assign n7667 = n2092 & ~n7666 ;
  assign n7668 = n7667 ^ n358 ^ 1'b0 ;
  assign n7669 = n7557 | n7668 ;
  assign n7670 = n3902 & ~n7669 ;
  assign n7671 = n890 | n7670 ;
  assign n7672 = n7663 & ~n7671 ;
  assign n7673 = n7672 ^ n1412 ^ 1'b0 ;
  assign n7674 = n4425 & n7673 ;
  assign n7675 = n826 ^ n362 ^ 1'b0 ;
  assign n7676 = n180 & ~n7675 ;
  assign n7677 = n925 & n1380 ;
  assign n7678 = ~n2419 & n7677 ;
  assign n7679 = n3770 | n7678 ;
  assign n7680 = n3035 | n7679 ;
  assign n7681 = n7680 ^ n3763 ^ n1940 ;
  assign n7682 = ( n2391 & ~n5679 ) | ( n2391 & n7681 ) | ( ~n5679 & n7681 ) ;
  assign n7683 = n1777 | n5736 ;
  assign n7684 = n4397 & ~n7683 ;
  assign n7685 = n5569 & ~n7684 ;
  assign n7686 = n7685 ^ n2876 ^ 1'b0 ;
  assign n7687 = ( n318 & ~n6298 ) | ( n318 & n6509 ) | ( ~n6298 & n6509 ) ;
  assign n7688 = n1801 & ~n3304 ;
  assign n7689 = n7688 ^ n1461 ^ 1'b0 ;
  assign n7690 = n7689 ^ n6447 ^ 1'b0 ;
  assign n7696 = n5424 ^ n3140 ^ n2602 ;
  assign n7691 = n98 | n1796 ;
  assign n7692 = n1489 | n7691 ;
  assign n7693 = n4860 ^ n1026 ^ 1'b0 ;
  assign n7694 = n7692 & n7693 ;
  assign n7695 = n2335 & n7694 ;
  assign n7697 = n7696 ^ n7695 ^ 1'b0 ;
  assign n7698 = n5183 ^ n2595 ^ n2327 ;
  assign n7699 = n1426 & ~n7698 ;
  assign n7700 = ~x10 & n7516 ;
  assign n7701 = n7700 ^ n2810 ^ 1'b0 ;
  assign n7702 = ( n1511 & n3557 ) | ( n1511 & ~n7701 ) | ( n3557 & ~n7701 ) ;
  assign n7703 = n7702 ^ n7661 ^ 1'b0 ;
  assign n7704 = n7699 & n7703 ;
  assign n7705 = ~n542 & n6717 ;
  assign n7710 = ~n139 & n2152 ;
  assign n7706 = ( n2213 & n3561 ) | ( n2213 & n4343 ) | ( n3561 & n4343 ) ;
  assign n7707 = n2296 & n7706 ;
  assign n7708 = n7707 ^ n3180 ^ n115 ;
  assign n7709 = ~n4786 & n7708 ;
  assign n7711 = n7710 ^ n7709 ^ 1'b0 ;
  assign n7712 = n2855 ^ n891 ^ 1'b0 ;
  assign n7713 = n2176 & ~n7712 ;
  assign n7714 = n7054 & n7713 ;
  assign n7715 = ~n7711 & n7714 ;
  assign n7716 = n5191 ^ n596 ^ 1'b0 ;
  assign n7717 = n2241 | n7716 ;
  assign n7718 = ( n4322 & ~n5039 ) | ( n4322 & n6257 ) | ( ~n5039 & n6257 ) ;
  assign n7719 = n263 | n871 ;
  assign n7720 = ~n1110 & n7719 ;
  assign n7721 = n4756 & n7720 ;
  assign n7722 = n1345 | n7721 ;
  assign n7723 = n278 & n6187 ;
  assign n7724 = n7723 ^ n3608 ^ 1'b0 ;
  assign n7725 = n6808 & n7724 ;
  assign n7726 = n7725 ^ n7724 ^ 1'b0 ;
  assign n7727 = n63 & ~n852 ;
  assign n7728 = ~n611 & n7727 ;
  assign n7729 = n1428 & ~n3807 ;
  assign n7730 = n7729 ^ n1562 ^ 1'b0 ;
  assign n7731 = n5549 ^ n2216 ^ 1'b0 ;
  assign n7732 = n4508 & n7731 ;
  assign n7733 = n2281 & n3130 ;
  assign n7734 = ~n7732 & n7733 ;
  assign n7735 = n6111 ^ n803 ^ 1'b0 ;
  assign n7736 = n1802 ^ n887 ^ 1'b0 ;
  assign n7737 = n2203 & ~n7736 ;
  assign n7738 = n154 & n3385 ;
  assign n7739 = ~n1906 & n2140 ;
  assign n7740 = n7739 ^ n1619 ^ 1'b0 ;
  assign n7741 = ( n2521 & n7738 ) | ( n2521 & ~n7740 ) | ( n7738 & ~n7740 ) ;
  assign n7742 = n983 & n2482 ;
  assign n7743 = ~n4662 & n7742 ;
  assign n7744 = n5289 & n7743 ;
  assign n7745 = n6044 | n7744 ;
  assign n7746 = n7745 ^ n1262 ^ 1'b0 ;
  assign n7750 = n1462 ^ n396 ^ 1'b0 ;
  assign n7751 = n7750 ^ n2278 ^ 1'b0 ;
  assign n7752 = n7751 ^ n1945 ^ 1'b0 ;
  assign n7753 = ( ~n428 & n7198 ) | ( ~n428 & n7752 ) | ( n7198 & n7752 ) ;
  assign n7748 = n4813 ^ n287 ^ 1'b0 ;
  assign n7749 = ~n3138 & n7748 ;
  assign n7747 = ( n1019 & ~n4054 ) | ( n1019 & n7069 ) | ( ~n4054 & n7069 ) ;
  assign n7754 = n7753 ^ n7749 ^ n7747 ;
  assign n7755 = n3758 & ~n4536 ;
  assign n7756 = n614 & n3362 ;
  assign n7757 = n7756 ^ n1346 ^ 1'b0 ;
  assign n7758 = n5378 ^ n4889 ^ 1'b0 ;
  assign n7759 = ~n221 & n7758 ;
  assign n7760 = ( n2179 & ~n4727 ) | ( n2179 & n7071 ) | ( ~n4727 & n7071 ) ;
  assign n7761 = n505 & ~n4058 ;
  assign n7762 = ( ~n2567 & n3696 ) | ( ~n2567 & n7761 ) | ( n3696 & n7761 ) ;
  assign n7763 = n4107 ^ n918 ^ 1'b0 ;
  assign n7764 = n4281 & n7763 ;
  assign n7765 = ~n7762 & n7764 ;
  assign n7766 = n7765 ^ n2379 ^ 1'b0 ;
  assign n7767 = n4543 | n7756 ;
  assign n7768 = n7641 ^ n1424 ^ 1'b0 ;
  assign n7769 = n7768 ^ n436 ^ 1'b0 ;
  assign n7770 = n580 & ~n7769 ;
  assign n7771 = n7770 ^ n3198 ^ n2586 ;
  assign n7772 = n3155 ^ n147 ^ 1'b0 ;
  assign n7773 = n7771 & n7772 ;
  assign n7774 = n5082 ^ n879 ^ 1'b0 ;
  assign n7775 = n7774 ^ n5451 ^ 1'b0 ;
  assign n7776 = ( ~n1880 & n4143 ) | ( ~n1880 & n5797 ) | ( n4143 & n5797 ) ;
  assign n7777 = n2966 ^ n999 ^ 1'b0 ;
  assign n7778 = n2746 & n7777 ;
  assign n7779 = ( n51 & n854 ) | ( n51 & ~n7778 ) | ( n854 & ~n7778 ) ;
  assign n7780 = n7779 ^ n7238 ^ n5323 ;
  assign n7781 = n5844 | n6842 ;
  assign n7782 = n7780 & ~n7781 ;
  assign n7784 = n1082 & ~n2547 ;
  assign n7783 = ~n1691 & n2122 ;
  assign n7785 = n7784 ^ n7783 ^ 1'b0 ;
  assign n7786 = n7337 ^ n1464 ^ 1'b0 ;
  assign n7787 = n7786 ^ n6743 ^ n4465 ;
  assign n7789 = n5047 ^ n3236 ^ 1'b0 ;
  assign n7790 = n7467 | n7789 ;
  assign n7788 = n4978 | n5353 ;
  assign n7791 = n7790 ^ n7788 ^ n424 ;
  assign n7792 = n5817 ^ n2830 ^ 1'b0 ;
  assign n7793 = n291 & ~n7792 ;
  assign n7794 = n7793 ^ n3709 ^ 1'b0 ;
  assign n7795 = ( n135 & n2649 ) | ( n135 & ~n7794 ) | ( n2649 & ~n7794 ) ;
  assign n7797 = n6246 ^ n2207 ^ 1'b0 ;
  assign n7798 = n577 & n7797 ;
  assign n7796 = n4086 ^ n1139 ^ 1'b0 ;
  assign n7799 = n7798 ^ n7796 ^ 1'b0 ;
  assign n7800 = n860 & n1969 ;
  assign n7801 = n7800 ^ n2499 ^ 1'b0 ;
  assign n7802 = n3832 ^ n3446 ^ 1'b0 ;
  assign n7803 = n129 & n1812 ;
  assign n7804 = n7803 ^ n372 ^ 1'b0 ;
  assign n7805 = n3833 | n7804 ;
  assign n7806 = n7805 ^ n5284 ^ 1'b0 ;
  assign n7807 = n5102 & n7806 ;
  assign n7808 = n940 & n2195 ;
  assign n7809 = n7807 & ~n7808 ;
  assign n7810 = n502 & n7809 ;
  assign n7811 = n1600 & n2345 ;
  assign n7812 = ~n1507 & n7811 ;
  assign n7813 = n1824 & ~n4772 ;
  assign n7814 = n7813 ^ n1500 ^ 1'b0 ;
  assign n7815 = ~n949 & n7814 ;
  assign n7818 = n423 ^ n101 ^ 1'b0 ;
  assign n7819 = n6583 ^ n965 ^ 1'b0 ;
  assign n7820 = ~n7818 & n7819 ;
  assign n7816 = n3125 ^ n2479 ^ 1'b0 ;
  assign n7817 = ~n2071 & n7816 ;
  assign n7821 = n7820 ^ n7817 ^ 1'b0 ;
  assign n7822 = ~n2326 & n7821 ;
  assign n7823 = ~n4754 & n5262 ;
  assign n7824 = n441 & ~n3848 ;
  assign n7825 = ~n4041 & n7824 ;
  assign n7826 = n445 & n2868 ;
  assign n7827 = ~n5036 & n7826 ;
  assign n7828 = n5400 & n7827 ;
  assign n7829 = ~n7290 & n7828 ;
  assign n7830 = n5329 & n7829 ;
  assign n7831 = n5453 ^ n2203 ^ 1'b0 ;
  assign n7832 = n7831 ^ n2504 ^ 1'b0 ;
  assign n7833 = ~n890 & n7322 ;
  assign n7834 = n7833 ^ n700 ^ 1'b0 ;
  assign n7842 = n77 ^ x9 ^ 1'b0 ;
  assign n7837 = ~n1437 & n5348 ;
  assign n7838 = n1632 & n7837 ;
  assign n7835 = ~n2330 & n2573 ;
  assign n7836 = n7835 ^ n397 ^ 1'b0 ;
  assign n7839 = n7838 ^ n7836 ^ n383 ;
  assign n7840 = n771 & n2816 ;
  assign n7841 = ~n7839 & n7840 ;
  assign n7843 = n7842 ^ n7841 ^ 1'b0 ;
  assign n7844 = n2923 | n7843 ;
  assign n7845 = n5594 | n7844 ;
  assign n7846 = n7845 ^ n749 ^ 1'b0 ;
  assign n7847 = n3401 ^ n1463 ^ 1'b0 ;
  assign n7848 = ( n3101 & ~n7642 ) | ( n3101 & n7847 ) | ( ~n7642 & n7847 ) ;
  assign n7850 = n1073 | n2971 ;
  assign n7849 = n44 & ~n6368 ;
  assign n7851 = n7850 ^ n7849 ^ 1'b0 ;
  assign n7854 = n1686 & n4959 ;
  assign n7852 = n2833 | n4149 ;
  assign n7853 = n1032 & n7852 ;
  assign n7855 = n7854 ^ n7853 ^ 1'b0 ;
  assign n7856 = ~n1751 & n7855 ;
  assign n7857 = ~n3082 & n3119 ;
  assign n7858 = ~n2904 & n7857 ;
  assign n7859 = ( n3370 & ~n4584 ) | ( n3370 & n7858 ) | ( ~n4584 & n7858 ) ;
  assign n7860 = n7327 ^ n2266 ^ 1'b0 ;
  assign n7861 = ~n33 & n6978 ;
  assign n7862 = n7861 ^ n1988 ^ 1'b0 ;
  assign n7863 = n7860 | n7862 ;
  assign n7864 = ( n65 & n1262 ) | ( n65 & n2054 ) | ( n1262 & n2054 ) ;
  assign n7865 = n5038 & n7864 ;
  assign n7866 = n7865 ^ n1838 ^ 1'b0 ;
  assign n7867 = n3710 & ~n5526 ;
  assign n7868 = n5241 ^ n1353 ^ 1'b0 ;
  assign n7869 = n7868 ^ n7802 ^ 1'b0 ;
  assign n7870 = n3998 ^ n3456 ^ n1489 ;
  assign n7871 = n1367 & ~n4515 ;
  assign n7872 = n7871 ^ n2650 ^ 1'b0 ;
  assign n7873 = n7870 & ~n7872 ;
  assign n7874 = n7873 ^ n1507 ^ 1'b0 ;
  assign n7875 = n607 & n4514 ;
  assign n7876 = n2605 ^ n1628 ^ n183 ;
  assign n7877 = ~n676 & n7876 ;
  assign n7878 = n7135 & n7877 ;
  assign n7880 = n260 | n2755 ;
  assign n7879 = n6195 ^ n5850 ^ 1'b0 ;
  assign n7881 = n7880 ^ n7879 ^ n4772 ;
  assign n7882 = n2106 & ~n2911 ;
  assign n7883 = ~n627 & n2961 ;
  assign n7884 = ~x1 & n7883 ;
  assign n7885 = n7884 ^ n6126 ^ 1'b0 ;
  assign n7886 = n3038 ^ n1824 ^ 1'b0 ;
  assign n7887 = n6596 & ~n7886 ;
  assign n7888 = n5052 & n7887 ;
  assign n7889 = n534 & n4988 ;
  assign n7890 = ~n3872 & n7889 ;
  assign n7891 = n7890 ^ n686 ^ 1'b0 ;
  assign n7892 = ( n1858 & ~n6778 ) | ( n1858 & n7465 ) | ( ~n6778 & n7465 ) ;
  assign n7893 = n139 & n767 ;
  assign n7894 = n336 & ~n7893 ;
  assign n7895 = n7894 ^ n1628 ^ 1'b0 ;
  assign n7896 = n7895 ^ n3755 ^ 1'b0 ;
  assign n7901 = n1196 | n1225 ;
  assign n7902 = n7901 ^ n1265 ^ 1'b0 ;
  assign n7897 = n5809 ^ n255 ^ 1'b0 ;
  assign n7898 = n251 | n7897 ;
  assign n7899 = n645 | n5249 ;
  assign n7900 = n7898 & ~n7899 ;
  assign n7903 = n7902 ^ n7900 ^ n1491 ;
  assign n7904 = n2076 & ~n7903 ;
  assign n7905 = n2348 & ~n4396 ;
  assign n7906 = ~n3506 & n7905 ;
  assign n7907 = n1023 & n3271 ;
  assign n7910 = n3382 & ~n3945 ;
  assign n7911 = n7910 ^ n916 ^ 1'b0 ;
  assign n7908 = n5754 ^ n3671 ^ 1'b0 ;
  assign n7909 = n728 & ~n7908 ;
  assign n7912 = n7911 ^ n7909 ^ 1'b0 ;
  assign n7913 = n6415 ^ n1716 ^ n870 ;
  assign n7914 = n1865 ^ n1827 ^ 1'b0 ;
  assign n7915 = n2216 & ~n7914 ;
  assign n7916 = ~n7913 & n7915 ;
  assign n7918 = n2367 ^ n883 ^ 1'b0 ;
  assign n7917 = ( n1209 & ~n3037 ) | ( n1209 & n5453 ) | ( ~n3037 & n5453 ) ;
  assign n7919 = n7918 ^ n7917 ^ 1'b0 ;
  assign n7920 = n4525 & ~n7919 ;
  assign n7921 = ( n498 & n4273 ) | ( n498 & n7920 ) | ( n4273 & n7920 ) ;
  assign n7922 = n7921 ^ n1457 ^ 1'b0 ;
  assign n7923 = n6991 & n7922 ;
  assign n7924 = n4457 ^ n727 ^ 1'b0 ;
  assign n7925 = ~n3632 & n7924 ;
  assign n7926 = n130 & n7925 ;
  assign n7927 = n7926 ^ n5977 ^ 1'b0 ;
  assign n7928 = n1083 & n1305 ;
  assign n7929 = n7928 ^ n607 ^ 1'b0 ;
  assign n7930 = n4070 | n7929 ;
  assign n7931 = n6576 ^ n214 ^ 1'b0 ;
  assign n7932 = n1647 ^ n1425 ^ n186 ;
  assign n7933 = ~n3389 & n3788 ;
  assign n7934 = ~n411 & n3840 ;
  assign n7935 = n7934 ^ n1581 ^ 1'b0 ;
  assign n7936 = ~n102 & n381 ;
  assign n7937 = ~n7935 & n7936 ;
  assign n7938 = n5797 & ~n7937 ;
  assign n7939 = n6384 ^ n884 ^ 1'b0 ;
  assign n7940 = n46 & ~n126 ;
  assign n7941 = ( n5504 & n6503 ) | ( n5504 & ~n7940 ) | ( n6503 & ~n7940 ) ;
  assign n7942 = n1758 & ~n7244 ;
  assign n7943 = n7942 ^ n5797 ^ 1'b0 ;
  assign n7944 = n3869 ^ n3802 ^ 1'b0 ;
  assign n7945 = n1720 | n7875 ;
  assign n7946 = n35 & n4901 ;
  assign n7947 = n6699 & n7946 ;
  assign n7948 = n7534 ^ n3530 ^ 1'b0 ;
  assign n7949 = n4096 | n7948 ;
  assign n7950 = n3383 ^ n2405 ^ 1'b0 ;
  assign n7951 = ~n2747 & n7950 ;
  assign n7952 = ( n119 & n3034 ) | ( n119 & ~n7951 ) | ( n3034 & ~n7951 ) ;
  assign n7953 = n7450 ^ n5310 ^ 1'b0 ;
  assign n7954 = n7903 & n7953 ;
  assign n7955 = ~n1660 & n2053 ;
  assign n7956 = n190 & n7955 ;
  assign n7957 = ~n1627 & n2354 ;
  assign n7958 = n7957 ^ n4686 ^ n2795 ;
  assign n7959 = n7958 ^ n4422 ^ 1'b0 ;
  assign n7960 = n7956 | n7959 ;
  assign n7961 = n2879 ^ n1516 ^ 1'b0 ;
  assign n7962 = n3908 & n7961 ;
  assign n7963 = n1223 & n7962 ;
  assign n7964 = ~n7960 & n7963 ;
  assign n7965 = n7964 ^ n1127 ^ 1'b0 ;
  assign n7967 = n879 | n2434 ;
  assign n7968 = n816 | n7967 ;
  assign n7966 = n105 & n2964 ;
  assign n7969 = n7968 ^ n7966 ^ 1'b0 ;
  assign n7970 = n7965 & n7969 ;
  assign n7973 = ( n684 & ~n3443 ) | ( n684 & n4656 ) | ( ~n3443 & n4656 ) ;
  assign n7971 = n6808 ^ n2546 ^ 1'b0 ;
  assign n7972 = ~n2892 & n7971 ;
  assign n7974 = n7973 ^ n7972 ^ 1'b0 ;
  assign n7975 = n7648 ^ n6299 ^ n442 ;
  assign n7976 = n1062 & n1169 ;
  assign n7977 = n2446 ^ n1737 ^ n204 ;
  assign n7978 = n7977 ^ n3421 ^ 1'b0 ;
  assign n7979 = n4251 ^ n1809 ^ n324 ;
  assign n7980 = ~n6014 & n7979 ;
  assign n7981 = n1666 & n7368 ;
  assign n7982 = n7981 ^ n628 ^ 1'b0 ;
  assign n7983 = n2666 & n3681 ;
  assign n7984 = n7983 ^ n1134 ^ 1'b0 ;
  assign n7985 = ~n1527 & n7984 ;
  assign n7986 = ~n834 & n7985 ;
  assign n7987 = ~n7654 & n7986 ;
  assign n7988 = n694 & ~n740 ;
  assign n7989 = n4525 ^ n3802 ^ 1'b0 ;
  assign n7990 = n1270 & n7989 ;
  assign n7991 = n7990 ^ n589 ^ 1'b0 ;
  assign n7992 = n4663 & ~n7304 ;
  assign n7993 = ~n7991 & n7992 ;
  assign n7994 = n7988 | n7993 ;
  assign n7995 = x6 & ~n1945 ;
  assign n7996 = n7995 ^ n3866 ^ 1'b0 ;
  assign n7997 = n7996 ^ n6699 ^ 1'b0 ;
  assign n7998 = n676 ^ n390 ^ 1'b0 ;
  assign n7999 = n265 | n7998 ;
  assign n8000 = n1267 & ~n7999 ;
  assign n8001 = n8000 ^ n4205 ^ 1'b0 ;
  assign n8007 = ( n844 & n2229 ) | ( n844 & n4608 ) | ( n2229 & n4608 ) ;
  assign n8008 = n3190 | n8007 ;
  assign n8002 = ~n63 & n7638 ;
  assign n8003 = n6603 & n8002 ;
  assign n8004 = n8003 ^ n5223 ^ 1'b0 ;
  assign n8005 = n4939 & ~n8004 ;
  assign n8006 = n839 & n8005 ;
  assign n8009 = n8008 ^ n8006 ^ 1'b0 ;
  assign n8010 = n8009 ^ n7879 ^ 1'b0 ;
  assign n8011 = n5226 ^ n2615 ^ 1'b0 ;
  assign n8012 = n4004 & ~n8011 ;
  assign n8013 = ~n6370 & n8012 ;
  assign n8014 = n8013 ^ n4969 ^ 1'b0 ;
  assign n8015 = ( ~n1169 & n4903 ) | ( ~n1169 & n8014 ) | ( n4903 & n8014 ) ;
  assign n8016 = n4961 ^ n1387 ^ n97 ;
  assign n8017 = n6581 ^ n944 ^ n125 ;
  assign n8018 = n8017 ^ n517 ^ 1'b0 ;
  assign n8019 = n3916 ^ n1182 ^ 1'b0 ;
  assign n8020 = ~n209 & n8019 ;
  assign n8021 = n8020 ^ n5649 ^ n2557 ;
  assign n8022 = n7658 ^ n3720 ^ 1'b0 ;
  assign n8023 = n1600 & ~n8022 ;
  assign n8024 = n26 & ~n2483 ;
  assign n8025 = n154 & n1695 ;
  assign n8026 = ( ~n2599 & n8024 ) | ( ~n2599 & n8025 ) | ( n8024 & n8025 ) ;
  assign n8027 = n8026 ^ n5762 ^ 1'b0 ;
  assign n8028 = n5799 ^ n4132 ^ n966 ;
  assign n8029 = n180 & n491 ;
  assign n8030 = n1426 & ~n7273 ;
  assign n8031 = n8030 ^ n5134 ^ 1'b0 ;
  assign n8032 = n2328 & ~n5197 ;
  assign n8033 = n1000 & ~n8032 ;
  assign n8034 = n6423 ^ n1426 ^ 1'b0 ;
  assign n8035 = n2402 ^ n607 ^ 1'b0 ;
  assign n8036 = ~n676 & n1918 ;
  assign n8037 = n8036 ^ n2806 ^ 1'b0 ;
  assign n8038 = ~n744 & n7761 ;
  assign n8039 = ~n8037 & n8038 ;
  assign n8040 = n6058 ^ n3067 ^ 1'b0 ;
  assign n8041 = ~n8039 & n8040 ;
  assign n8042 = n5458 ^ n3408 ^ 1'b0 ;
  assign n8043 = n8041 & ~n8042 ;
  assign n8044 = ~n8035 & n8043 ;
  assign n8045 = n8044 ^ n3985 ^ 1'b0 ;
  assign n8052 = n7920 ^ n3912 ^ n3456 ;
  assign n8046 = n772 ^ n734 ^ 1'b0 ;
  assign n8047 = n345 & n1202 ;
  assign n8048 = n1423 ^ n1232 ^ 1'b0 ;
  assign n8049 = ( ~n6087 & n8047 ) | ( ~n6087 & n8048 ) | ( n8047 & n8048 ) ;
  assign n8050 = ~n3459 & n8049 ;
  assign n8051 = n8046 & n8050 ;
  assign n8053 = n8052 ^ n8051 ^ 1'b0 ;
  assign n8054 = n5648 | n8053 ;
  assign n8055 = n947 ^ n523 ^ 1'b0 ;
  assign n8056 = n750 & ~n4933 ;
  assign n8057 = ( n134 & ~n1891 ) | ( n134 & n3195 ) | ( ~n1891 & n3195 ) ;
  assign n8058 = n8057 ^ n6024 ^ 1'b0 ;
  assign n8059 = n3027 ^ n2667 ^ 1'b0 ;
  assign n8060 = n1367 | n8059 ;
  assign n8061 = n8060 ^ n3615 ^ n3046 ;
  assign n8062 = n1461 ^ n1055 ^ 1'b0 ;
  assign n8063 = ~n2006 & n8062 ;
  assign n8064 = ~n4086 & n8063 ;
  assign n8065 = n8061 & n8064 ;
  assign n8066 = n4927 ^ n944 ^ 1'b0 ;
  assign n8067 = ( ~n577 & n2106 ) | ( ~n577 & n8066 ) | ( n2106 & n8066 ) ;
  assign n8068 = ( n773 & n2115 ) | ( n773 & ~n7701 ) | ( n2115 & ~n7701 ) ;
  assign n8069 = n6136 & ~n8068 ;
  assign n8070 = n8069 ^ n2165 ^ 1'b0 ;
  assign n8071 = n8070 ^ n3195 ^ 1'b0 ;
  assign n8072 = ( n2705 & n2925 ) | ( n2705 & ~n4719 ) | ( n2925 & ~n4719 ) ;
  assign n8073 = ( n1470 & n1746 ) | ( n1470 & ~n8072 ) | ( n1746 & ~n8072 ) ;
  assign n8074 = n101 | n2184 ;
  assign n8075 = n8074 ^ n2050 ^ 1'b0 ;
  assign n8076 = ~n8073 & n8075 ;
  assign n8077 = n1512 & n4376 ;
  assign n8078 = ~n5650 & n8077 ;
  assign n8079 = n8078 ^ n1081 ^ 1'b0 ;
  assign n8080 = n3313 ^ n141 ^ 1'b0 ;
  assign n8081 = ~n396 & n2922 ;
  assign n8082 = ~n2887 & n8081 ;
  assign n8083 = x3 | n5977 ;
  assign n8084 = n864 | n7726 ;
  assign n8085 = n281 & n597 ;
  assign n8086 = n2414 ^ n186 ^ 1'b0 ;
  assign n8087 = n6736 ^ n3923 ^ 1'b0 ;
  assign n8088 = n338 & n8087 ;
  assign n8089 = n7106 ^ n6564 ^ n453 ;
  assign n8090 = ( ~n752 & n947 ) | ( ~n752 & n1922 ) | ( n947 & n1922 ) ;
  assign n8091 = n2932 ^ n1258 ^ 1'b0 ;
  assign n8092 = n7530 ^ n5649 ^ 1'b0 ;
  assign n8093 = ~n8091 & n8092 ;
  assign n8094 = ~n115 & n1447 ;
  assign n8095 = ~n1880 & n7029 ;
  assign n8097 = n1890 | n2309 ;
  assign n8096 = n132 | n5469 ;
  assign n8098 = n8097 ^ n8096 ^ n1762 ;
  assign n8099 = n2291 ^ n759 ^ 1'b0 ;
  assign n8100 = n5388 & ~n6904 ;
  assign n8101 = ~n8099 & n8100 ;
  assign n8102 = n7927 | n8101 ;
  assign n8103 = n8102 ^ n2160 ^ 1'b0 ;
  assign n8104 = n4688 ^ n2216 ^ 1'b0 ;
  assign n8105 = n5694 | n8104 ;
  assign n8106 = n4273 & ~n5384 ;
  assign n8107 = n8106 ^ n3926 ^ n648 ;
  assign n8108 = n8105 & ~n8107 ;
  assign n8109 = ( ~n1088 & n1185 ) | ( ~n1088 & n5893 ) | ( n1185 & n5893 ) ;
  assign n8110 = n4303 ^ n1715 ^ 1'b0 ;
  assign n8111 = n8110 ^ n769 ^ 1'b0 ;
  assign n8112 = n44 & ~n8111 ;
  assign n8113 = n2399 ^ n1898 ^ 1'b0 ;
  assign n8114 = n4551 ^ n1182 ^ 1'b0 ;
  assign n8115 = n8114 ^ n6315 ^ n2307 ;
  assign n8116 = ~n882 & n8115 ;
  assign n8117 = n191 & n8116 ;
  assign n8118 = n3975 & ~n8117 ;
  assign n8119 = n8118 ^ n6698 ^ 1'b0 ;
  assign n8120 = n8119 ^ n3510 ^ 1'b0 ;
  assign n8121 = n2186 & ~n4390 ;
  assign n8122 = ~n6288 & n8121 ;
  assign n8123 = n1305 & n2101 ;
  assign n8124 = n2307 | n3189 ;
  assign n8125 = n8124 ^ n1309 ^ 1'b0 ;
  assign n8126 = n2615 & n7998 ;
  assign n8127 = n6443 ^ n434 ^ 1'b0 ;
  assign n8128 = n8127 ^ n2264 ^ 1'b0 ;
  assign n8130 = n1561 ^ n174 ^ n101 ;
  assign n8131 = n661 ^ n37 ^ 1'b0 ;
  assign n8132 = n5088 & ~n8131 ;
  assign n8133 = n8130 & n8132 ;
  assign n8129 = n6245 ^ n3416 ^ 1'b0 ;
  assign n8134 = n8133 ^ n8129 ^ 1'b0 ;
  assign n8135 = n3123 & n8076 ;
  assign n8136 = n8122 ^ n3128 ^ 1'b0 ;
  assign n8137 = n5716 | n8136 ;
  assign n8138 = n435 & ~n6612 ;
  assign n8139 = n4647 ^ n3100 ^ 1'b0 ;
  assign n8140 = n8139 ^ n2190 ^ 1'b0 ;
  assign n8141 = n4146 & n4754 ;
  assign n8142 = n2378 ^ n342 ^ 1'b0 ;
  assign n8143 = ( n998 & n1891 ) | ( n998 & ~n8142 ) | ( n1891 & ~n8142 ) ;
  assign n8144 = n8143 ^ n3367 ^ 1'b0 ;
  assign n8145 = ~n8141 & n8144 ;
  assign n8146 = n8145 ^ n3467 ^ 1'b0 ;
  assign n8147 = n8146 ^ n1038 ^ 1'b0 ;
  assign n8148 = ~n2015 & n5735 ;
  assign n8149 = ( n1003 & n2623 ) | ( n1003 & ~n8148 ) | ( n2623 & ~n8148 ) ;
  assign n8152 = x4 & ~n7233 ;
  assign n8150 = n4742 ^ n3763 ^ 1'b0 ;
  assign n8151 = n7710 | n8150 ;
  assign n8153 = n8152 ^ n8151 ^ 1'b0 ;
  assign n8154 = n4062 ^ n443 ^ 1'b0 ;
  assign n8155 = n3959 | n8154 ;
  assign n8156 = n4737 | n8155 ;
  assign n8157 = n8156 ^ n5219 ^ 1'b0 ;
  assign n8158 = n7171 & ~n8157 ;
  assign n8160 = n3198 ^ n3067 ^ 1'b0 ;
  assign n8159 = n4793 ^ n2397 ^ 1'b0 ;
  assign n8161 = n8160 ^ n8159 ^ 1'b0 ;
  assign n8162 = ~n6460 & n8161 ;
  assign n8163 = n750 | n2766 ;
  assign n8164 = n2813 ^ n1040 ^ 1'b0 ;
  assign n8165 = ( n1970 & n8163 ) | ( n1970 & n8164 ) | ( n8163 & n8164 ) ;
  assign n8166 = n8165 ^ n2898 ^ 1'b0 ;
  assign n8167 = n2843 ^ n780 ^ x9 ;
  assign n8170 = n4307 ^ n3061 ^ 1'b0 ;
  assign n8168 = ~n2649 & n7215 ;
  assign n8169 = n2431 & ~n8168 ;
  assign n8171 = n8170 ^ n8169 ^ 1'b0 ;
  assign n8172 = n8171 ^ n6504 ^ x8 ;
  assign n8173 = n2286 & n5599 ;
  assign n8174 = n6212 ^ n4653 ^ 1'b0 ;
  assign n8175 = ~n3460 & n8174 ;
  assign n8176 = ( n1475 & n5165 ) | ( n1475 & ~n5443 ) | ( n5165 & ~n5443 ) ;
  assign n8177 = n2976 ^ n1789 ^ 1'b0 ;
  assign n8178 = n2177 | n4019 ;
  assign n8179 = n8178 ^ n1694 ^ 1'b0 ;
  assign n8180 = n8177 | n8179 ;
  assign n8181 = n8180 ^ n8039 ^ 1'b0 ;
  assign n8182 = n5515 ^ n1856 ^ 1'b0 ;
  assign n8183 = n5720 ^ n5682 ^ n3128 ;
  assign n8184 = n8183 ^ n1891 ^ n816 ;
  assign n8185 = n4971 ^ n1125 ^ 1'b0 ;
  assign n8186 = n1279 ^ n249 ^ 1'b0 ;
  assign n8187 = n5051 & n8186 ;
  assign n8188 = n2569 | n4086 ;
  assign n8189 = n1443 ^ n1400 ^ 1'b0 ;
  assign n8190 = ~n8188 & n8189 ;
  assign n8191 = n8190 ^ n4168 ^ n2164 ;
  assign n8192 = ~n3053 & n3655 ;
  assign n8193 = n386 ^ n216 ^ 1'b0 ;
  assign n8194 = ~n1970 & n6143 ;
  assign n8195 = n8193 & n8194 ;
  assign n8196 = n4060 & n8195 ;
  assign n8197 = ~n8192 & n8196 ;
  assign n8198 = n5395 & ~n7347 ;
  assign n8199 = n583 | n8198 ;
  assign n8200 = n7427 & n8199 ;
  assign n8201 = ~n5376 & n8200 ;
  assign n8203 = n6073 ^ n1278 ^ 1'b0 ;
  assign n8202 = n2332 & ~n3713 ;
  assign n8204 = n8203 ^ n8202 ^ 1'b0 ;
  assign n8205 = n3558 | n5136 ;
  assign n8206 = n2906 ^ n773 ^ 1'b0 ;
  assign n8207 = n8206 ^ n240 ^ 1'b0 ;
  assign n8208 = ~n7362 & n8207 ;
  assign n8209 = n381 & ~n2177 ;
  assign n8210 = n4992 ^ n3246 ^ 1'b0 ;
  assign n8211 = n8209 | n8210 ;
  assign n8212 = n2819 & ~n6479 ;
  assign n8213 = n4553 | n6369 ;
  assign n8214 = n2913 & ~n8213 ;
  assign n8215 = ( n523 & ~n1314 ) | ( n523 & n2597 ) | ( ~n1314 & n2597 ) ;
  assign n8216 = n6490 & ~n8215 ;
  assign n8217 = n846 & ~n915 ;
  assign n8218 = ~n1784 & n8217 ;
  assign n8219 = ~n1201 & n2575 ;
  assign n8220 = n1491 & n8219 ;
  assign n8221 = n2282 & ~n8220 ;
  assign n8222 = n30 & n8221 ;
  assign n8223 = n8222 ^ n4100 ^ 1'b0 ;
  assign n8224 = n8218 | n8223 ;
  assign n8225 = n4787 | n8224 ;
  assign n8226 = n213 & ~n6386 ;
  assign n8227 = ( n524 & n1930 ) | ( n524 & n3457 ) | ( n1930 & n3457 ) ;
  assign n8228 = n5531 & ~n8227 ;
  assign n8229 = n5845 ^ n437 ^ 1'b0 ;
  assign n8230 = n7019 ^ n186 ^ 1'b0 ;
  assign n8231 = n8229 & n8230 ;
  assign n8232 = n1905 | n3035 ;
  assign n8233 = ~n3791 & n8232 ;
  assign n8234 = n8233 ^ n603 ^ 1'b0 ;
  assign n8235 = n8234 ^ n7977 ^ 1'b0 ;
  assign n8236 = n41 & ~n8235 ;
  assign n8237 = n803 & ~n5163 ;
  assign n8238 = n2316 ^ n334 ^ 1'b0 ;
  assign n8239 = n8237 & n8238 ;
  assign n8240 = n7329 ^ n1871 ^ 1'b0 ;
  assign n8241 = n8240 ^ n7706 ^ 1'b0 ;
  assign n8242 = ~n1090 & n1409 ;
  assign n8243 = n8159 ^ n2798 ^ 1'b0 ;
  assign n8244 = ( ~n2225 & n7864 ) | ( ~n2225 & n8243 ) | ( n7864 & n8243 ) ;
  assign n8245 = n4681 ^ n301 ^ 1'b0 ;
  assign n8246 = n1495 & n4319 ;
  assign n8247 = n8246 ^ n1424 ^ 1'b0 ;
  assign n8248 = ( ~n3470 & n5207 ) | ( ~n3470 & n5900 ) | ( n5207 & n5900 ) ;
  assign n8249 = ( n376 & ~n5234 ) | ( n376 & n5639 ) | ( ~n5234 & n5639 ) ;
  assign n8250 = ~n2802 & n3454 ;
  assign n8251 = n8250 ^ n5083 ^ 1'b0 ;
  assign n8252 = n8251 ^ n5742 ^ 1'b0 ;
  assign n8253 = ~n2274 & n8252 ;
  assign n8254 = n8249 & ~n8253 ;
  assign n8255 = n2100 | n6597 ;
  assign n8256 = n8255 ^ n5104 ^ 1'b0 ;
  assign n8257 = n845 & ~n8256 ;
  assign n8258 = ( n113 & n1078 ) | ( n113 & n8257 ) | ( n1078 & n8257 ) ;
  assign n8259 = n2198 & ~n6166 ;
  assign n8260 = ( n2041 & n5284 ) | ( n2041 & ~n6289 ) | ( n5284 & ~n6289 ) ;
  assign n8261 = ~n740 & n8260 ;
  assign n8262 = n8259 & n8261 ;
  assign n8263 = n969 | n7893 ;
  assign n8264 = n1107 | n8263 ;
  assign n8265 = ( n791 & n1155 ) | ( n791 & n2274 ) | ( n1155 & n2274 ) ;
  assign n8266 = ~n8264 & n8265 ;
  assign n8267 = n1173 | n4288 ;
  assign n8268 = ~n1783 & n8267 ;
  assign n8269 = n1642 ^ n87 ^ 1'b0 ;
  assign n8270 = n386 & ~n4558 ;
  assign n8271 = n4334 & n8270 ;
  assign n8272 = n179 & n2073 ;
  assign n8273 = n8272 ^ n5699 ^ 1'b0 ;
  assign n8274 = ~n5241 & n8273 ;
  assign n8275 = ~n2062 & n8274 ;
  assign n8276 = ~n5163 & n5217 ;
  assign n8277 = n8276 ^ n5974 ^ 1'b0 ;
  assign n8278 = n633 & n1210 ;
  assign n8279 = ( n1854 & n6445 ) | ( n1854 & n8278 ) | ( n6445 & n8278 ) ;
  assign n8280 = n2750 ^ n1103 ^ 1'b0 ;
  assign n8281 = n5296 & n8280 ;
  assign n8282 = n2139 | n5083 ;
  assign n8283 = n8282 ^ n814 ^ 1'b0 ;
  assign n8284 = n5563 & n8283 ;
  assign n8285 = n4039 ^ n230 ^ 1'b0 ;
  assign n8286 = n2094 & ~n5115 ;
  assign n8287 = n8285 & n8286 ;
  assign n8288 = n6144 | n8287 ;
  assign n8289 = ~n3140 & n7713 ;
  assign n8290 = n3029 | n8289 ;
  assign n8291 = n8288 & ~n8290 ;
  assign n8292 = n6653 ^ n2289 ^ n963 ;
  assign n8293 = n1513 ^ n499 ^ 1'b0 ;
  assign n8294 = ~n1103 & n8293 ;
  assign n8295 = n8294 ^ n5488 ^ 1'b0 ;
  assign n8296 = n5406 & ~n8295 ;
  assign n8297 = n8296 ^ n2696 ^ n1783 ;
  assign n8298 = n8292 & ~n8297 ;
  assign n8302 = n6150 ^ n4223 ^ n3795 ;
  assign n8301 = n5178 & ~n5650 ;
  assign n8303 = n8302 ^ n8301 ^ 1'b0 ;
  assign n8299 = n773 ^ x3 ^ 1'b0 ;
  assign n8300 = ( n2728 & n4914 ) | ( n2728 & n8299 ) | ( n4914 & n8299 ) ;
  assign n8304 = n8303 ^ n8300 ^ n2561 ;
  assign n8305 = ~n4852 & n8304 ;
  assign n8306 = ( ~n2989 & n7475 ) | ( ~n2989 & n8305 ) | ( n7475 & n8305 ) ;
  assign n8307 = n893 ^ n866 ^ 1'b0 ;
  assign n8308 = ~n216 & n8307 ;
  assign n8309 = n5348 ^ n256 ^ 1'b0 ;
  assign n8310 = ~n2452 & n8309 ;
  assign n8311 = n8226 ^ n5870 ^ n5716 ;
  assign n8312 = n4782 ^ n2365 ^ 1'b0 ;
  assign n8313 = n1166 & ~n3455 ;
  assign n8314 = ( ~n1039 & n3094 ) | ( ~n1039 & n8313 ) | ( n3094 & n8313 ) ;
  assign n8315 = n7344 ^ n4558 ^ 1'b0 ;
  assign n8316 = n6563 & n8315 ;
  assign n8317 = n5203 | n5796 ;
  assign n8318 = n8317 ^ n1841 ^ 1'b0 ;
  assign n8321 = n5848 ^ n1636 ^ n126 ;
  assign n8322 = n221 | n334 ;
  assign n8323 = n8322 ^ n2039 ^ 1'b0 ;
  assign n8324 = n8323 ^ n119 ^ 1'b0 ;
  assign n8325 = n107 & n8324 ;
  assign n8326 = n8321 & n8325 ;
  assign n8319 = n8207 ^ n6403 ^ 1'b0 ;
  assign n8320 = n7354 & n8319 ;
  assign n8327 = n8326 ^ n8320 ^ 1'b0 ;
  assign n8328 = n4275 & ~n5337 ;
  assign n8329 = n7908 & n8328 ;
  assign n8330 = n6770 | n8329 ;
  assign n8331 = ~n619 & n4072 ;
  assign n8332 = n2179 & n3973 ;
  assign n8333 = ~n4434 & n8332 ;
  assign n8334 = n5186 ^ n2605 ^ n2157 ;
  assign n8335 = n224 | n3891 ;
  assign n8336 = n5948 ^ n1110 ^ 1'b0 ;
  assign n8337 = n8335 & ~n8336 ;
  assign n8338 = n6333 ^ n79 ^ 1'b0 ;
  assign n8339 = n122 & ~n3704 ;
  assign n8340 = n8339 ^ n4337 ^ 1'b0 ;
  assign n8341 = n3686 ^ n263 ^ 1'b0 ;
  assign n8342 = ( n8338 & n8340 ) | ( n8338 & ~n8341 ) | ( n8340 & ~n8341 ) ;
  assign n8343 = n8342 ^ n5517 ^ 1'b0 ;
  assign n8344 = n4622 ^ n4507 ^ 1'b0 ;
  assign n8345 = n3709 ^ n543 ^ 1'b0 ;
  assign n8346 = n164 & n8345 ;
  assign n8347 = ( n3174 & n8344 ) | ( n3174 & ~n8346 ) | ( n8344 & ~n8346 ) ;
  assign n8348 = ( n5052 & ~n5771 ) | ( n5052 & n8347 ) | ( ~n5771 & n8347 ) ;
  assign n8349 = n3775 ^ n561 ^ 1'b0 ;
  assign n8350 = n8165 & n8349 ;
  assign n8351 = ( n6204 & n7383 ) | ( n6204 & n8350 ) | ( n7383 & n8350 ) ;
  assign n8352 = n3238 | n8351 ;
  assign n8353 = n8352 ^ n1028 ^ 1'b0 ;
  assign n8354 = n609 & ~n2088 ;
  assign n8355 = n585 & ~n597 ;
  assign n8356 = n8355 ^ n2011 ^ 1'b0 ;
  assign n8357 = n1525 & ~n4195 ;
  assign n8358 = n4071 | n5886 ;
  assign n8359 = n169 | n8358 ;
  assign n8360 = n8359 ^ n5373 ^ 1'b0 ;
  assign n8361 = n827 | n8360 ;
  assign n8362 = ( n408 & n3961 ) | ( n408 & n5214 ) | ( n3961 & n5214 ) ;
  assign n8363 = ~n2202 & n8362 ;
  assign n8364 = n8363 ^ n5284 ^ 1'b0 ;
  assign n8365 = ( n1822 & ~n2032 ) | ( n1822 & n2471 ) | ( ~n2032 & n2471 ) ;
  assign n8366 = n6796 | n8365 ;
  assign n8367 = n8366 ^ n6199 ^ 1'b0 ;
  assign n8368 = n6496 ^ n2209 ^ n53 ;
  assign n8369 = n8368 ^ n332 ^ 1'b0 ;
  assign n8373 = ( ~n98 & n411 ) | ( ~n98 & n1635 ) | ( n411 & n1635 ) ;
  assign n8370 = n791 & n5246 ;
  assign n8371 = n8370 ^ n1389 ^ 1'b0 ;
  assign n8372 = n8371 ^ n4359 ^ 1'b0 ;
  assign n8374 = n8373 ^ n8372 ^ 1'b0 ;
  assign n8375 = n3801 ^ n3238 ^ 1'b0 ;
  assign n8376 = n4062 & n5564 ;
  assign n8377 = n8375 | n8376 ;
  assign n8378 = n8377 ^ n2759 ^ 1'b0 ;
  assign n8379 = n316 & n1446 ;
  assign n8381 = n2286 | n3134 ;
  assign n8382 = n8381 ^ n2036 ^ 1'b0 ;
  assign n8383 = n8382 ^ n7413 ^ n925 ;
  assign n8380 = x7 & ~n6392 ;
  assign n8384 = n8383 ^ n8380 ^ 1'b0 ;
  assign n8385 = ~n8379 & n8384 ;
  assign n8386 = n6608 | n6842 ;
  assign n8387 = n8386 ^ n7227 ^ 1'b0 ;
  assign n8388 = n3326 & n5559 ;
  assign n8389 = n8388 ^ n1345 ^ 1'b0 ;
  assign n8390 = n8389 ^ n7389 ^ n5799 ;
  assign n8391 = ~n581 & n8325 ;
  assign n8392 = n8390 & n8391 ;
  assign n8393 = n484 & n5089 ;
  assign n8394 = n1072 & ~n8393 ;
  assign n8395 = n8394 ^ n1439 ^ 1'b0 ;
  assign n8396 = n134 & ~n2341 ;
  assign n8397 = n8396 ^ n1736 ^ 1'b0 ;
  assign n8398 = n8039 | n8397 ;
  assign n8399 = n1820 | n8398 ;
  assign n8400 = n3469 & ~n8399 ;
  assign n8401 = n8057 | n8400 ;
  assign n8402 = n3669 ^ n3452 ^ 1'b0 ;
  assign n8403 = n4948 & n8402 ;
  assign n8404 = n3554 ^ n1931 ^ n378 ;
  assign n8405 = n2012 & ~n8404 ;
  assign n8406 = ~n102 & n8405 ;
  assign n8408 = n1139 & ~n2071 ;
  assign n8409 = n8408 ^ n3454 ^ n2128 ;
  assign n8410 = n8409 ^ n49 ^ 1'b0 ;
  assign n8411 = n2313 & n8410 ;
  assign n8407 = n5036 & ~n7329 ;
  assign n8412 = n8411 ^ n8407 ^ 1'b0 ;
  assign n8413 = ~n8406 & n8412 ;
  assign n8414 = ( n900 & n1361 ) | ( n900 & n8142 ) | ( n1361 & n8142 ) ;
  assign n8415 = n766 & n8414 ;
  assign n8416 = n2389 & n8415 ;
  assign n8417 = n6666 ^ n727 ^ 1'b0 ;
  assign n8418 = n1712 | n8417 ;
  assign n8419 = n360 & n7776 ;
  assign n8420 = ~n8418 & n8419 ;
  assign n8421 = n8420 ^ n1400 ^ 1'b0 ;
  assign n8422 = n1316 & ~n1517 ;
  assign n8423 = n269 & n8422 ;
  assign n8424 = ( n2302 & n5543 ) | ( n2302 & n8423 ) | ( n5543 & n8423 ) ;
  assign n8425 = n8424 ^ x10 ^ 1'b0 ;
  assign n8426 = n3163 | n8425 ;
  assign n8427 = n8426 ^ n6014 ^ 1'b0 ;
  assign n8428 = n1147 ^ n1024 ^ x10 ;
  assign n8429 = n4044 & ~n8428 ;
  assign n8430 = n42 | n6929 ;
  assign n8431 = n893 & ~n8430 ;
  assign n8432 = ( n2296 & ~n2918 ) | ( n2296 & n4340 ) | ( ~n2918 & n4340 ) ;
  assign n8433 = n6102 & ~n8432 ;
  assign n8434 = n8433 ^ n2517 ^ 1'b0 ;
  assign n8435 = n5399 & ~n7169 ;
  assign n8436 = ~n3045 & n3713 ;
  assign n8437 = n8436 ^ n3882 ^ 1'b0 ;
  assign n8438 = n7434 & n8437 ;
  assign n8440 = n1928 & n5565 ;
  assign n8439 = ~n147 & n3257 ;
  assign n8441 = n8440 ^ n8439 ^ 1'b0 ;
  assign n8442 = n8441 ^ n4971 ^ 1'b0 ;
  assign n8443 = n2885 & ~n5670 ;
  assign n8444 = ~n1974 & n8443 ;
  assign n8445 = ~n4743 & n8444 ;
  assign n8446 = n8445 ^ n2413 ^ 1'b0 ;
  assign n8447 = n2546 ^ n906 ^ 1'b0 ;
  assign n8448 = n8447 ^ n7197 ^ n1311 ;
  assign n8449 = ( n1877 & n7796 ) | ( n1877 & n8448 ) | ( n7796 & n8448 ) ;
  assign n8450 = n8446 & ~n8449 ;
  assign n8451 = n5220 ^ n259 ^ n188 ;
  assign n8452 = n4235 | n4252 ;
  assign n8453 = n8452 ^ n5570 ^ 1'b0 ;
  assign n8454 = n3040 | n8453 ;
  assign n8455 = n190 & ~n8454 ;
  assign n8456 = n4849 ^ n4608 ^ n1566 ;
  assign n8457 = n4767 & ~n8456 ;
  assign n8458 = ~n2596 & n6581 ;
  assign n8459 = n2076 ^ n1483 ^ 1'b0 ;
  assign n8460 = ~n8458 & n8459 ;
  assign n8461 = ~n2080 & n6320 ;
  assign n8462 = n2971 & n8461 ;
  assign n8463 = x3 & ~n6689 ;
  assign n8464 = ~n1184 & n8463 ;
  assign n8465 = n8462 & n8464 ;
  assign n8471 = n2869 & n3006 ;
  assign n8466 = n1357 ^ n318 ^ x0 ;
  assign n8467 = n5735 ^ n5559 ^ 1'b0 ;
  assign n8468 = ~n5241 & n8467 ;
  assign n8469 = ~n3321 & n8468 ;
  assign n8470 = n8466 & ~n8469 ;
  assign n8472 = n8471 ^ n8470 ^ n1607 ;
  assign n8477 = n4971 ^ n745 ^ 1'b0 ;
  assign n8478 = n97 | n8477 ;
  assign n8479 = n4134 | n8478 ;
  assign n8480 = n808 & ~n8479 ;
  assign n8473 = n1419 & ~n4044 ;
  assign n8474 = n8473 ^ n5450 ^ 1'b0 ;
  assign n8475 = n1272 & n8474 ;
  assign n8476 = n8475 ^ n5111 ^ 1'b0 ;
  assign n8481 = n8480 ^ n8476 ^ 1'b0 ;
  assign n8482 = ~n7559 & n8481 ;
  assign n8483 = n8482 ^ n5012 ^ 1'b0 ;
  assign n8484 = ~n883 & n1888 ;
  assign n8485 = n8484 ^ n93 ^ 1'b0 ;
  assign n8486 = n8485 ^ n6914 ^ 1'b0 ;
  assign n8488 = ~n72 & n1109 ;
  assign n8489 = n4154 & n8488 ;
  assign n8487 = n654 & n3840 ;
  assign n8490 = n8489 ^ n8487 ^ 1'b0 ;
  assign n8491 = n8490 ^ n881 ^ 1'b0 ;
  assign n8492 = ~n2432 & n8143 ;
  assign n8493 = n1535 & n8492 ;
  assign n8494 = n8491 | n8493 ;
  assign n8495 = n8486 & n8494 ;
  assign n8496 = n8495 ^ n4280 ^ 1'b0 ;
  assign n8497 = n4010 ^ n3307 ^ n1290 ;
  assign n8498 = ( n1296 & ~n2408 ) | ( n1296 & n3911 ) | ( ~n2408 & n3911 ) ;
  assign n8499 = n8498 ^ n1533 ^ 1'b0 ;
  assign n8500 = n8497 & n8499 ;
  assign n8501 = n8500 ^ n6119 ^ 1'b0 ;
  assign n8502 = n4383 & n8501 ;
  assign n8503 = ~n5563 & n8502 ;
  assign n8504 = ~n3660 & n8503 ;
  assign n8505 = n8504 ^ n170 ^ 1'b0 ;
  assign n8506 = n1061 & n8505 ;
  assign n8507 = n619 & n8506 ;
  assign n8508 = n8507 ^ n139 ^ 1'b0 ;
  assign n8509 = n629 & n4195 ;
  assign n8510 = ~n617 & n7338 ;
  assign n8511 = n8510 ^ n411 ^ 1'b0 ;
  assign n8512 = n8511 ^ n1766 ^ 1'b0 ;
  assign n8513 = n2738 & n8512 ;
  assign n8514 = n8513 ^ n676 ^ 1'b0 ;
  assign n8517 = ~n2259 & n4939 ;
  assign n8518 = n8517 ^ n4797 ^ n2387 ;
  assign n8516 = n959 & ~n2055 ;
  assign n8515 = n7785 ^ n1984 ^ 1'b0 ;
  assign n8519 = n8518 ^ n8516 ^ n8515 ;
  assign n8520 = n1516 ^ n1069 ^ 1'b0 ;
  assign n8521 = n2367 & n8520 ;
  assign n8522 = n8187 & ~n8521 ;
  assign n8523 = n6795 ^ n3971 ^ 1'b0 ;
  assign n8524 = n310 & ~n6139 ;
  assign n8525 = n151 | n6230 ;
  assign n8526 = n411 | n8525 ;
  assign n8527 = n6428 ^ n2882 ^ 1'b0 ;
  assign n8528 = ( n657 & ~n7348 ) | ( n657 & n8527 ) | ( ~n7348 & n8527 ) ;
  assign n8529 = n35 & ~n276 ;
  assign n8530 = n3302 ^ n242 ^ 1'b0 ;
  assign n8531 = ~n3229 & n8530 ;
  assign n8532 = ~n8529 & n8531 ;
  assign n8533 = ( ~n5568 & n5796 ) | ( ~n5568 & n6736 ) | ( n5796 & n6736 ) ;
  assign n8534 = n8532 | n8533 ;
  assign n8535 = n8534 ^ n269 ^ 1'b0 ;
  assign n8536 = ~n2860 & n8535 ;
  assign n8537 = n5599 & n7218 ;
  assign n8539 = n826 | n4298 ;
  assign n8540 = n23 & n8539 ;
  assign n8538 = n619 & n6506 ;
  assign n8541 = n8540 ^ n8538 ^ 1'b0 ;
  assign n8542 = n505 & ~n590 ;
  assign n8543 = n7006 & ~n8542 ;
  assign n8544 = n361 | n8543 ;
  assign n8545 = ~n1393 & n3064 ;
  assign n8546 = n8545 ^ n5823 ^ 1'b0 ;
  assign n8547 = ~n7968 & n8546 ;
  assign n8548 = n1796 ^ n1296 ^ 1'b0 ;
  assign n8549 = n2584 & ~n8548 ;
  assign n8550 = n4380 ^ n435 ^ 1'b0 ;
  assign n8551 = n4906 | n8550 ;
  assign n8552 = n5068 ^ n2758 ^ 1'b0 ;
  assign n8553 = n3192 & ~n8552 ;
  assign n8554 = ~n7891 & n8553 ;
  assign n8555 = ~n110 & n2591 ;
  assign n8556 = n8555 ^ n1380 ^ 1'b0 ;
  assign n8557 = n3483 & n4703 ;
  assign n8558 = ( n791 & ~n1865 ) | ( n791 & n3500 ) | ( ~n1865 & n3500 ) ;
  assign n8559 = ~n1045 & n8558 ;
  assign n8560 = n2145 & n8559 ;
  assign n8561 = n7888 | n8560 ;
  assign n8562 = n7624 & ~n8561 ;
  assign n8563 = n2956 & n3626 ;
  assign n8564 = n2918 & ~n6121 ;
  assign n8565 = n8563 & n8564 ;
  assign n8568 = n1531 & n2233 ;
  assign n8569 = n8568 ^ n77 ^ 1'b0 ;
  assign n8566 = n6801 ^ n4647 ^ 1'b0 ;
  assign n8567 = n6660 & ~n8566 ;
  assign n8570 = n8569 ^ n8567 ^ 1'b0 ;
  assign n8571 = n2990 & ~n8570 ;
  assign n8572 = n1419 | n5938 ;
  assign n8573 = ~n4703 & n8572 ;
  assign n8574 = n8573 ^ n5237 ^ 1'b0 ;
  assign n8575 = n1064 & ~n7425 ;
  assign n8576 = n6428 ^ n5607 ^ 1'b0 ;
  assign n8577 = n8576 ^ n5815 ^ 1'b0 ;
  assign n8579 = ~n1690 & n6756 ;
  assign n8580 = n7347 & n8579 ;
  assign n8578 = n1138 | n5378 ;
  assign n8581 = n8580 ^ n8578 ^ 1'b0 ;
  assign n8584 = n279 & ~n1402 ;
  assign n8585 = n8584 ^ n3019 ^ 1'b0 ;
  assign n8582 = n5570 ^ n1781 ^ 1'b0 ;
  assign n8583 = n2472 | n8582 ;
  assign n8586 = n8585 ^ n8583 ^ 1'b0 ;
  assign n8587 = n7707 ^ n3877 ^ 1'b0 ;
  assign n8588 = n3916 & ~n8587 ;
  assign n8589 = n8588 ^ n5162 ^ 1'b0 ;
  assign n8590 = n4643 & ~n8589 ;
  assign n8591 = ( ~n126 & n1033 ) | ( ~n126 & n2039 ) | ( n1033 & n2039 ) ;
  assign n8592 = n4257 | n8591 ;
  assign n8593 = n570 & ~n1999 ;
  assign n8594 = n4214 ^ n1079 ^ 1'b0 ;
  assign n8595 = n4617 & ~n8594 ;
  assign n8596 = ~n1351 & n8595 ;
  assign n8597 = n8596 ^ n5149 ^ 1'b0 ;
  assign n8598 = n8593 & n8597 ;
  assign n8599 = n8598 ^ n2110 ^ 1'b0 ;
  assign n8600 = n1953 | n8599 ;
  assign n8601 = n6607 & n8173 ;
  assign n8602 = n2551 & n6638 ;
  assign n8603 = ~n2845 & n8602 ;
  assign n8604 = ~n888 & n8603 ;
  assign n8605 = n8604 ^ n7921 ^ n2345 ;
  assign n8606 = n7938 ^ n1170 ^ 1'b0 ;
  assign n8607 = ( n1153 & ~n2135 ) | ( n1153 & n5155 ) | ( ~n2135 & n5155 ) ;
  assign n8608 = ( n524 & ~n908 ) | ( n524 & n7121 ) | ( ~n908 & n7121 ) ;
  assign n8609 = n1957 | n3043 ;
  assign n8610 = n8608 | n8609 ;
  assign n8611 = ~n1412 & n8610 ;
  assign n8612 = n8607 & n8611 ;
  assign n8613 = n6778 | n7033 ;
  assign n8614 = n8613 ^ n3244 ^ 1'b0 ;
  assign n8615 = n7283 | n8614 ;
  assign n8616 = n6215 ^ n2644 ^ 1'b0 ;
  assign n8617 = n2640 ^ n636 ^ 1'b0 ;
  assign n8618 = ~n125 & n8617 ;
  assign n8619 = n1453 & n8618 ;
  assign n8620 = n6638 ^ x4 ^ 1'b0 ;
  assign n8621 = n8619 & n8620 ;
  assign n8622 = n8621 ^ n5603 ^ n1196 ;
  assign n8623 = n8622 ^ n183 ^ 1'b0 ;
  assign n8624 = n6142 & ~n8623 ;
  assign n8625 = n8624 ^ n1734 ^ 1'b0 ;
  assign n8626 = n3190 | n8625 ;
  assign n8627 = n8626 ^ n5561 ^ 1'b0 ;
  assign n8628 = n4951 | n8627 ;
  assign n8629 = n7610 ^ n3650 ^ 1'b0 ;
  assign n8630 = n3392 ^ n1600 ^ n280 ;
  assign n8631 = n6149 & n8630 ;
  assign n8632 = ~n1368 & n1650 ;
  assign n8633 = n8632 ^ n162 ^ 1'b0 ;
  assign n8634 = n1650 & n8633 ;
  assign n8635 = ~n8631 & n8634 ;
  assign n8636 = n4201 ^ n1279 ^ 1'b0 ;
  assign n8637 = ~n1525 & n6471 ;
  assign n8638 = n3093 & n8637 ;
  assign n8639 = n8638 ^ n922 ^ 1'b0 ;
  assign n8640 = n3353 ^ n461 ^ 1'b0 ;
  assign n8643 = n532 & ~n2075 ;
  assign n8644 = n8643 ^ n3020 ^ 1'b0 ;
  assign n8645 = ~n2584 & n8644 ;
  assign n8646 = ~n3440 & n8645 ;
  assign n8647 = n8646 ^ n3898 ^ 1'b0 ;
  assign n8648 = n1898 & n2280 ;
  assign n8649 = ( n5061 & n5244 ) | ( n5061 & ~n8648 ) | ( n5244 & ~n8648 ) ;
  assign n8650 = n8647 & n8649 ;
  assign n8651 = n7265 & n8650 ;
  assign n8641 = n221 & n1698 ;
  assign n8642 = ~n6454 & n8641 ;
  assign n8652 = n8651 ^ n8642 ^ 1'b0 ;
  assign n8653 = n8640 & n8652 ;
  assign n8654 = ~n2339 & n8653 ;
  assign n8655 = n5122 ^ n4930 ^ 1'b0 ;
  assign n8656 = ( n2997 & ~n4280 ) | ( n2997 & n8655 ) | ( ~n4280 & n8655 ) ;
  assign n8657 = n3824 ^ n2182 ^ 1'b0 ;
  assign n8658 = n4539 & ~n8657 ;
  assign n8659 = n392 & n8658 ;
  assign n8660 = ( n1209 & n8346 ) | ( n1209 & ~n8659 ) | ( n8346 & ~n8659 ) ;
  assign n8661 = n5292 ^ n4745 ^ 1'b0 ;
  assign n8662 = n4385 | n6970 ;
  assign n8663 = n1367 & ~n6595 ;
  assign n8665 = n4307 ^ n1726 ^ 1'b0 ;
  assign n8666 = ~n360 & n8665 ;
  assign n8667 = n6855 & n8666 ;
  assign n8668 = n3437 | n8667 ;
  assign n8669 = n2765 | n8668 ;
  assign n8664 = n3261 & n3510 ;
  assign n8670 = n8669 ^ n8664 ^ 1'b0 ;
  assign n8671 = n5200 & ~n8670 ;
  assign n8672 = n6526 ^ n2058 ^ 1'b0 ;
  assign n8673 = n587 & ~n3828 ;
  assign n8674 = ~n8285 & n8572 ;
  assign n8675 = n4459 ^ n378 ^ 1'b0 ;
  assign n8676 = n1125 & n8675 ;
  assign n8677 = ~n4917 & n8676 ;
  assign n8678 = n8677 ^ n2094 ^ 1'b0 ;
  assign n8679 = n108 & n3261 ;
  assign n8680 = n8679 ^ n1150 ^ 1'b0 ;
  assign n8681 = n7271 & n8680 ;
  assign n8682 = n5953 ^ n395 ^ 1'b0 ;
  assign n8683 = ~n572 & n1156 ;
  assign n8684 = n355 | n8683 ;
  assign n8685 = x0 & ~n1917 ;
  assign n8686 = n8685 ^ n1022 ^ 1'b0 ;
  assign n8687 = ~n44 & n2952 ;
  assign n8688 = n8687 ^ n6737 ^ 1'b0 ;
  assign n8689 = n8688 ^ n6098 ^ 1'b0 ;
  assign n8690 = n8686 | n8689 ;
  assign n8691 = ~n8379 & n8690 ;
  assign n8692 = ( ~n2811 & n3082 ) | ( ~n2811 & n7034 ) | ( n3082 & n7034 ) ;
  assign n8693 = n4180 ^ n1207 ^ 1'b0 ;
  assign n8694 = n451 & n8693 ;
  assign n8695 = ~n7215 & n8694 ;
  assign n8696 = ~n8692 & n8695 ;
  assign n8697 = ( n1448 & ~n1525 ) | ( n1448 & n2635 ) | ( ~n1525 & n2635 ) ;
  assign n8698 = n7111 | n8697 ;
  assign n8699 = n1088 & n8698 ;
  assign n8700 = ~n6612 & n8699 ;
  assign n8701 = n8700 ^ n5463 ^ 1'b0 ;
  assign n8702 = n2990 ^ n1425 ^ 1'b0 ;
  assign n8703 = n4230 | n8702 ;
  assign n8704 = n8703 ^ n6262 ^ 1'b0 ;
  assign n8705 = n1824 & ~n4110 ;
  assign n8706 = ~n2986 & n8705 ;
  assign n8707 = n4431 ^ n2201 ^ n1463 ;
  assign n8708 = ~n8706 & n8707 ;
  assign n8709 = n8708 ^ n2609 ^ 1'b0 ;
  assign n8710 = n2689 & ~n5084 ;
  assign n8711 = ~n8709 & n8710 ;
  assign n8712 = n8711 ^ n8635 ^ 1'b0 ;
  assign n8713 = ( ~n712 & n3461 ) | ( ~n712 & n3577 ) | ( n3461 & n3577 ) ;
  assign n8714 = ( n2482 & n3914 ) | ( n2482 & ~n3967 ) | ( n3914 & ~n3967 ) ;
  assign n8715 = ( ~n5053 & n8713 ) | ( ~n5053 & n8714 ) | ( n8713 & n8714 ) ;
  assign n8716 = n7831 & ~n8715 ;
  assign n8717 = n989 & n8716 ;
  assign n8718 = n3450 | n7916 ;
  assign n8719 = n8718 ^ n4778 ^ 1'b0 ;
  assign n8720 = n3780 ^ n1766 ^ 1'b0 ;
  assign n8721 = n3088 ^ n1539 ^ 1'b0 ;
  assign n8722 = n5392 ^ n1760 ^ 1'b0 ;
  assign n8723 = n8721 & ~n8722 ;
  assign n8724 = n8720 & n8723 ;
  assign n8725 = n5145 & ~n5251 ;
  assign n8726 = ( n1245 & ~n3382 ) | ( n1245 & n4688 ) | ( ~n3382 & n4688 ) ;
  assign n8727 = n8726 ^ n6716 ^ 1'b0 ;
  assign n8728 = n5759 ^ n2769 ^ 1'b0 ;
  assign n8729 = n1804 & ~n2128 ;
  assign n8730 = n7692 ^ n1996 ^ n928 ;
  assign n8731 = ( n466 & n8729 ) | ( n466 & n8730 ) | ( n8729 & n8730 ) ;
  assign n8737 = n1876 & ~n3307 ;
  assign n8738 = n8737 ^ n2502 ^ 1'b0 ;
  assign n8739 = n4593 ^ n145 ^ 1'b0 ;
  assign n8740 = n8738 & ~n8739 ;
  assign n8741 = ( ~n982 & n2817 ) | ( ~n982 & n8740 ) | ( n2817 & n8740 ) ;
  assign n8732 = n1564 & n5817 ;
  assign n8733 = n8732 ^ n1421 ^ 1'b0 ;
  assign n8734 = n341 & ~n2274 ;
  assign n8735 = n8734 ^ n1166 ^ 1'b0 ;
  assign n8736 = ( n6288 & ~n8733 ) | ( n6288 & n8735 ) | ( ~n8733 & n8735 ) ;
  assign n8742 = n8741 ^ n8736 ^ 1'b0 ;
  assign n8743 = n8731 & ~n8742 ;
  assign n8744 = n4596 & ~n4920 ;
  assign n8745 = ~n8268 & n8744 ;
  assign n8746 = ~n3127 & n4507 ;
  assign n8747 = n8310 & ~n8746 ;
  assign n8751 = n4645 ^ n3890 ^ 1'b0 ;
  assign n8752 = ~n3138 & n6564 ;
  assign n8753 = n8751 & n8752 ;
  assign n8754 = n864 & ~n8753 ;
  assign n8748 = ~n1197 & n1532 ;
  assign n8749 = ~n7818 & n8748 ;
  assign n8750 = ~n5320 & n8749 ;
  assign n8755 = n8754 ^ n8750 ^ 1'b0 ;
  assign n8756 = n3923 ^ n3133 ^ 1'b0 ;
  assign n8757 = n8755 | n8756 ;
  assign n8758 = n8757 ^ n5073 ^ 1'b0 ;
  assign n8759 = n5675 ^ n3006 ^ 1'b0 ;
  assign n8760 = n8759 ^ n4567 ^ 1'b0 ;
  assign n8761 = ~n1818 & n8760 ;
  assign n8762 = n6291 & n8761 ;
  assign n8763 = n7506 & n8762 ;
  assign n8764 = ~n842 & n5479 ;
  assign n8765 = n1075 | n7207 ;
  assign n8766 = n6736 ^ n2110 ^ n251 ;
  assign n8767 = n8766 ^ n4558 ^ 1'b0 ;
  assign n8768 = n5114 & ~n8767 ;
  assign n8769 = ( ~n925 & n7503 ) | ( ~n925 & n8768 ) | ( n7503 & n8768 ) ;
  assign n8770 = ~n4336 & n7242 ;
  assign n8771 = n2798 | n8770 ;
  assign n8772 = n6240 & ~n8771 ;
  assign n8773 = n1104 | n3394 ;
  assign n8774 = n523 & ~n8773 ;
  assign n8775 = n6188 ^ n646 ^ n450 ;
  assign n8776 = ~n859 & n3464 ;
  assign n8777 = ~n4580 & n8776 ;
  assign n8779 = n1582 & n2514 ;
  assign n8780 = n8779 ^ n2009 ^ 1'b0 ;
  assign n8778 = n7752 ^ n7600 ^ n3284 ;
  assign n8781 = n8780 ^ n8778 ^ 1'b0 ;
  assign n8782 = ~n6025 & n8781 ;
  assign n8783 = ~n5595 & n8782 ;
  assign n8784 = ~n668 & n6692 ;
  assign n8785 = ~n2075 & n2661 ;
  assign n8786 = n8785 ^ n48 ^ 1'b0 ;
  assign n8787 = n8784 & ~n8786 ;
  assign n8792 = ( n2858 & n3552 ) | ( n2858 & ~n6081 ) | ( n3552 & ~n6081 ) ;
  assign n8793 = n8792 ^ n2176 ^ 1'b0 ;
  assign n8788 = n403 & ~n1292 ;
  assign n8789 = n8788 ^ n4574 ^ 1'b0 ;
  assign n8790 = n230 & ~n8789 ;
  assign n8791 = ~n5538 & n8790 ;
  assign n8794 = n8793 ^ n8791 ^ 1'b0 ;
  assign n8795 = n8794 ^ n3135 ^ 1'b0 ;
  assign n8796 = n3236 ^ n1512 ^ 1'b0 ;
  assign n8797 = ~n1414 & n8796 ;
  assign n8798 = n3706 ^ n2262 ^ 1'b0 ;
  assign n8799 = n6608 ^ n157 ^ 1'b0 ;
  assign n8800 = n459 | n8799 ;
  assign n8805 = n383 | n1110 ;
  assign n8806 = n4189 & ~n8805 ;
  assign n8801 = n2247 ^ n2195 ^ 1'b0 ;
  assign n8802 = n8801 ^ n3578 ^ n65 ;
  assign n8803 = n4367 ^ n265 ^ 1'b0 ;
  assign n8804 = n8802 & n8803 ;
  assign n8807 = n8806 ^ n8804 ^ 1'b0 ;
  assign n8808 = n1142 | n3985 ;
  assign n8809 = n8808 ^ n4957 ^ 1'b0 ;
  assign n8810 = n5504 | n8809 ;
  assign n8811 = n3398 | n5414 ;
  assign n8812 = n3823 & ~n8811 ;
  assign n8813 = n2435 & ~n5225 ;
  assign n8814 = n7880 ^ n1076 ^ 1'b0 ;
  assign n8815 = n2839 & n8814 ;
  assign n8816 = n1851 & n2731 ;
  assign n8817 = n1962 & n8816 ;
  assign n8818 = n8817 ^ n118 ^ 1'b0 ;
  assign n8819 = n8815 & ~n8818 ;
  assign n8820 = n5545 & n8819 ;
  assign n8821 = n7513 ^ n5972 ^ n3604 ;
  assign n8822 = n2704 & n6243 ;
  assign n8823 = n3408 ^ n313 ^ 1'b0 ;
  assign n8824 = n494 & n8823 ;
  assign n8825 = n2081 & n8271 ;
  assign n8826 = ~n4869 & n8825 ;
  assign n8827 = n443 & ~n5006 ;
  assign n8828 = ~n6485 & n8827 ;
  assign n8830 = n6181 ^ n2736 ^ 1'b0 ;
  assign n8831 = n5393 & n8335 ;
  assign n8832 = n8831 ^ n2108 ^ 1'b0 ;
  assign n8833 = ( n5143 & n8830 ) | ( n5143 & ~n8832 ) | ( n8830 & ~n8832 ) ;
  assign n8829 = n1407 ^ n395 ^ 1'b0 ;
  assign n8834 = n8833 ^ n8829 ^ 1'b0 ;
  assign n8835 = n2615 & n8834 ;
  assign n8837 = n5637 | n6743 ;
  assign n8838 = n8837 ^ n4488 ^ 1'b0 ;
  assign n8839 = n1262 & n8497 ;
  assign n8840 = n6585 & n8839 ;
  assign n8841 = n8840 ^ n5758 ^ 1'b0 ;
  assign n8842 = ( n2262 & n8838 ) | ( n2262 & n8841 ) | ( n8838 & n8841 ) ;
  assign n8843 = n8842 ^ n1231 ^ 1'b0 ;
  assign n8836 = n1054 | n1511 ;
  assign n8844 = n8843 ^ n8836 ^ 1'b0 ;
  assign n8845 = n8844 ^ n4298 ^ n3505 ;
  assign n8846 = n4058 ^ n63 ^ 1'b0 ;
  assign n8848 = n6212 ^ n5163 ^ 1'b0 ;
  assign n8847 = ~n3824 & n8555 ;
  assign n8849 = n8848 ^ n8847 ^ n6246 ;
  assign n8850 = n8846 & ~n8849 ;
  assign n8851 = ~n4052 & n8131 ;
  assign n8852 = ~n607 & n8851 ;
  assign n8853 = n999 & ~n1337 ;
  assign n8854 = n8853 ^ n5665 ^ 1'b0 ;
  assign n8855 = ~n521 & n6126 ;
  assign n8856 = n8855 ^ n5072 ^ 1'b0 ;
  assign n8857 = n8854 & ~n8856 ;
  assign n8858 = ( n2745 & n4177 ) | ( n2745 & n8857 ) | ( n4177 & n8857 ) ;
  assign n8859 = n8858 ^ n2001 ^ n1888 ;
  assign n8860 = n5852 ^ n1523 ^ 1'b0 ;
  assign n8861 = n2969 & n3195 ;
  assign n8862 = ~n1693 & n5102 ;
  assign n8863 = n1500 & n8862 ;
  assign n8864 = n4574 ^ n4394 ^ n3181 ;
  assign n8865 = n8864 ^ n2485 ^ 1'b0 ;
  assign n8866 = ~n8863 & n8865 ;
  assign n8867 = n3428 ^ n3073 ^ 1'b0 ;
  assign n8868 = n3477 | n8867 ;
  assign n8869 = n7391 ^ n3817 ^ 1'b0 ;
  assign n8870 = n8869 ^ n5469 ^ 1'b0 ;
  assign n8871 = n6208 & n8870 ;
  assign n8872 = n8871 ^ n799 ^ 1'b0 ;
  assign n8873 = ~n844 & n3202 ;
  assign n8874 = ~n7449 & n8873 ;
  assign n8875 = ~n7467 & n8874 ;
  assign n8876 = n8875 ^ n4175 ^ 1'b0 ;
  assign n8877 = n8012 ^ n6238 ^ 1'b0 ;
  assign n8878 = n249 & n7434 ;
  assign n8879 = n3714 ^ n695 ^ n527 ;
  assign n8880 = n8879 ^ n7864 ^ n4683 ;
  assign n8881 = n8880 ^ n7767 ^ n1830 ;
  assign n8882 = n8344 ^ n5036 ^ n234 ;
  assign n8883 = n8882 ^ n2718 ^ 1'b0 ;
  assign n8884 = n2729 & n8883 ;
  assign n8885 = n2692 ^ n1213 ^ 1'b0 ;
  assign n8886 = n7867 ^ n6297 ^ n206 ;
  assign n8887 = n8886 ^ n6379 ^ 1'b0 ;
  assign n8888 = n36 & n8887 ;
  assign n8889 = n481 | n1315 ;
  assign n8890 = n8889 ^ n7283 ^ 1'b0 ;
  assign n8891 = n4965 ^ n63 ^ 1'b0 ;
  assign n8892 = n4508 & ~n8891 ;
  assign n8893 = n2108 & n8892 ;
  assign n8894 = n1105 ^ n176 ^ x3 ;
  assign n8895 = n8894 ^ n5881 ^ n5310 ;
  assign n8896 = n5545 ^ n506 ^ 1'b0 ;
  assign n8897 = x7 & n3165 ;
  assign n8898 = n287 ^ n195 ^ 1'b0 ;
  assign n8899 = n8897 & ~n8898 ;
  assign n8900 = n8899 ^ n6547 ^ 1'b0 ;
  assign n8901 = n5526 & ~n8900 ;
  assign n8902 = n8896 & n8901 ;
  assign n8903 = ( n458 & n5691 ) | ( n458 & n6389 ) | ( n5691 & n6389 ) ;
  assign n8904 = ~n91 & n2122 ;
  assign n8905 = n3515 & n8904 ;
  assign n8906 = n8903 & n8905 ;
  assign n8907 = n2134 | n2387 ;
  assign n8908 = n8907 ^ n8143 ^ 1'b0 ;
  assign n8909 = ~n8906 & n8908 ;
  assign n8910 = n3962 & ~n4760 ;
  assign n8911 = n963 | n1294 ;
  assign n8912 = n1405 & ~n8911 ;
  assign n8913 = n8912 ^ n3894 ^ n3397 ;
  assign n8914 = n4149 ^ n895 ^ 1'b0 ;
  assign n8915 = n4167 & n8914 ;
  assign n8916 = n1412 | n3443 ;
  assign n8917 = n5039 | n8916 ;
  assign n8918 = ( n5685 & ~n8915 ) | ( n5685 & n8917 ) | ( ~n8915 & n8917 ) ;
  assign n8919 = ~n4595 & n5859 ;
  assign n8920 = n8919 ^ n4607 ^ 1'b0 ;
  assign n8921 = n8918 & n8920 ;
  assign n8922 = n3708 & n7426 ;
  assign n8923 = n6060 & n8922 ;
  assign n8924 = n101 | n7391 ;
  assign n8925 = n5803 | n8924 ;
  assign n8926 = n5329 ^ n3241 ^ 1'b0 ;
  assign n8927 = n8770 ^ n3868 ^ n2088 ;
  assign n8928 = ~n442 & n3351 ;
  assign n8929 = ~n5276 & n8928 ;
  assign n8930 = n4918 | n8929 ;
  assign n8931 = n8930 ^ n2254 ^ 1'b0 ;
  assign n8932 = n395 & n2736 ;
  assign n8933 = n1084 & n8932 ;
  assign n8934 = n4607 ^ n4429 ^ 1'b0 ;
  assign n8935 = n3005 ^ n392 ^ 1'b0 ;
  assign n8936 = n8934 & n8935 ;
  assign n8937 = n7852 | n8587 ;
  assign n8938 = n938 & ~n1823 ;
  assign n8939 = ~n2567 & n8938 ;
  assign n8941 = ( n187 & ~n471 ) | ( n187 & n661 ) | ( ~n471 & n661 ) ;
  assign n8940 = n2082 | n6493 ;
  assign n8942 = n8941 ^ n8940 ^ 1'b0 ;
  assign n8943 = n6101 ^ n1513 ^ 1'b0 ;
  assign n8944 = n8942 & n8943 ;
  assign n8945 = ~n5033 & n8944 ;
  assign n8946 = n381 & ~n411 ;
  assign n8947 = ~n695 & n8946 ;
  assign n8948 = n2587 & ~n8947 ;
  assign n8949 = n5828 & n6983 ;
  assign n8950 = n7188 & n8949 ;
  assign n8953 = ~n1233 & n2218 ;
  assign n8951 = n814 & ~n1693 ;
  assign n8952 = ~n4150 & n8951 ;
  assign n8954 = n8953 ^ n8952 ^ 1'b0 ;
  assign n8955 = n8954 ^ n1828 ^ 1'b0 ;
  assign n8956 = n5941 ^ n4880 ^ 1'b0 ;
  assign n8957 = ~n8955 & n8956 ;
  assign n8958 = ( n803 & n3628 ) | ( n803 & ~n8957 ) | ( n3628 & ~n8957 ) ;
  assign n8959 = n4146 & ~n4971 ;
  assign n8960 = n5339 | n8959 ;
  assign n8961 = n6039 ^ n1824 ^ n561 ;
  assign n8962 = ~n8960 & n8961 ;
  assign n8963 = n5832 & n8962 ;
  assign n8964 = ~n4778 & n8963 ;
  assign n8965 = ( n1478 & n5253 ) | ( n1478 & ~n8964 ) | ( n5253 & ~n8964 ) ;
  assign n8967 = n4325 ^ n1270 ^ 1'b0 ;
  assign n8968 = n8967 ^ n350 ^ 1'b0 ;
  assign n8969 = n508 | n933 ;
  assign n8970 = n8969 ^ n448 ^ 1'b0 ;
  assign n8971 = n5183 & ~n8970 ;
  assign n8972 = n8968 & n8971 ;
  assign n8966 = ~n1628 & n5444 ;
  assign n8973 = n8972 ^ n8966 ^ 1'b0 ;
  assign n8975 = n184 | n2505 ;
  assign n8974 = n1606 & ~n2208 ;
  assign n8976 = n8975 ^ n8974 ^ n2076 ;
  assign n8977 = n8976 ^ n5782 ^ n611 ;
  assign n8978 = ~n3212 & n5806 ;
  assign n8979 = n8978 ^ n7605 ^ n7543 ;
  assign n8984 = n3692 & ~n4320 ;
  assign n8985 = n8984 ^ n329 ^ 1'b0 ;
  assign n8980 = ~n1407 & n2333 ;
  assign n8981 = n2338 ^ n991 ^ 1'b0 ;
  assign n8982 = n8980 | n8981 ;
  assign n8983 = n931 & ~n8982 ;
  assign n8986 = n8985 ^ n8983 ^ 1'b0 ;
  assign n8987 = n2280 | n4754 ;
  assign n8988 = n8987 ^ n4750 ^ 1'b0 ;
  assign n8989 = n1326 | n8068 ;
  assign n8990 = n159 | n8989 ;
  assign n8991 = n8923 & ~n8990 ;
  assign n8992 = n5311 ^ n1996 ^ 1'b0 ;
  assign n8993 = n727 & n8992 ;
  assign n8994 = n8071 | n8993 ;
  assign n8995 = n7237 ^ n6360 ^ 1'b0 ;
  assign n8996 = n8995 ^ n8945 ^ 1'b0 ;
  assign n8997 = ~n2770 & n8555 ;
  assign n8998 = n8997 ^ n7836 ^ 1'b0 ;
  assign n8999 = n8998 ^ n6452 ^ 1'b0 ;
  assign n9000 = n8996 & n8999 ;
  assign n9002 = n36 & n6413 ;
  assign n9001 = n2288 | n4575 ;
  assign n9003 = n9002 ^ n9001 ^ 1'b0 ;
  assign n9004 = ( n574 & n1647 ) | ( n574 & n2202 ) | ( n1647 & n2202 ) ;
  assign n9005 = n9004 ^ n5858 ^ 1'b0 ;
  assign n9006 = n9005 ^ n1468 ^ 1'b0 ;
  assign n9007 = n70 & n846 ;
  assign n9008 = n9007 ^ n2784 ^ 1'b0 ;
  assign n9009 = n9008 ^ n6899 ^ 1'b0 ;
  assign n9024 = n5156 | n7784 ;
  assign n9021 = x10 & ~n3162 ;
  assign n9010 = ~n1532 & n2242 ;
  assign n9011 = n3690 & n9010 ;
  assign n9018 = n640 & n7354 ;
  assign n9012 = n817 | n2208 ;
  assign n9013 = ~n2854 & n9012 ;
  assign n9014 = n8145 ^ n6468 ^ n1845 ;
  assign n9015 = ~n3363 & n9014 ;
  assign n9016 = n882 | n9015 ;
  assign n9017 = n9013 & ~n9016 ;
  assign n9019 = n9018 ^ n9017 ^ 1'b0 ;
  assign n9020 = ( n7181 & n9011 ) | ( n7181 & ~n9019 ) | ( n9011 & ~n9019 ) ;
  assign n9022 = n9021 ^ n9020 ^ 1'b0 ;
  assign n9023 = n9022 ^ n6292 ^ 1'b0 ;
  assign n9025 = n9024 ^ n9023 ^ 1'b0 ;
  assign n9026 = n7449 & n9025 ;
  assign n9027 = n2327 ^ n723 ^ 1'b0 ;
  assign n9028 = ~n112 & n845 ;
  assign n9029 = n9028 ^ n909 ^ 1'b0 ;
  assign n9030 = n734 ^ n466 ^ 1'b0 ;
  assign n9031 = ~n9029 & n9030 ;
  assign n9032 = ~n838 & n9031 ;
  assign n9033 = n9032 ^ n5146 ^ n3387 ;
  assign n9034 = n9033 ^ n6536 ^ 1'b0 ;
  assign n9035 = n2846 ^ n142 ^ 1'b0 ;
  assign n9036 = n2496 & ~n9035 ;
  assign n9038 = n3708 & n4317 ;
  assign n9039 = n9038 ^ n2944 ^ 1'b0 ;
  assign n9037 = n2876 & ~n3573 ;
  assign n9040 = n9039 ^ n9037 ^ 1'b0 ;
  assign n9041 = n9036 & ~n9040 ;
  assign n9042 = n3998 | n4147 ;
  assign n9043 = n102 & ~n2095 ;
  assign n9044 = n5986 ^ n1105 ^ 1'b0 ;
  assign n9045 = n4413 | n9044 ;
  assign n9046 = n9045 ^ n8527 ^ 1'b0 ;
  assign n9047 = n6404 | n9046 ;
  assign n9048 = n9047 ^ n2332 ^ 1'b0 ;
  assign n9049 = n5006 & ~n9048 ;
  assign n9050 = n5700 ^ n2387 ^ 1'b0 ;
  assign n9051 = n9050 ^ n8802 ^ 1'b0 ;
  assign n9052 = n5252 ^ n211 ^ 1'b0 ;
  assign n9053 = n9052 ^ n2990 ^ 1'b0 ;
  assign n9054 = n5387 | n9053 ;
  assign n9055 = ~n825 & n2964 ;
  assign n9056 = n9055 ^ n6878 ^ 1'b0 ;
  assign n9057 = ~n2776 & n9056 ;
  assign n9058 = n1803 ^ n1079 ^ 1'b0 ;
  assign n9059 = n2412 & n9058 ;
  assign n9060 = n6658 ^ n2431 ^ 1'b0 ;
  assign n9061 = n2081 | n2706 ;
  assign n9062 = n8813 | n9061 ;
  assign n9063 = n9062 ^ n6352 ^ 1'b0 ;
  assign n9064 = n1751 & ~n5127 ;
  assign n9065 = ~n678 & n9064 ;
  assign n9066 = n9065 ^ n5233 ^ 1'b0 ;
  assign n9067 = n3330 ^ n2202 ^ 1'b0 ;
  assign n9068 = ~n5975 & n9067 ;
  assign n9069 = n543 & n5471 ;
  assign n9070 = ~n9068 & n9069 ;
  assign n9071 = n557 | n1363 ;
  assign n9072 = n1166 & ~n9071 ;
  assign n9073 = n4977 ^ n165 ^ 1'b0 ;
  assign n9074 = ( ~n849 & n9072 ) | ( ~n849 & n9073 ) | ( n9072 & n9073 ) ;
  assign n9075 = ( n177 & n2650 ) | ( n177 & ~n6389 ) | ( n2650 & ~n6389 ) ;
  assign n9076 = n1437 & ~n3466 ;
  assign n9077 = n445 & ~n2195 ;
  assign n9078 = ~n3124 & n9077 ;
  assign n9079 = ( n5651 & ~n9076 ) | ( n5651 & n9078 ) | ( ~n9076 & n9078 ) ;
  assign n9080 = n9079 ^ n1784 ^ 1'b0 ;
  assign n9081 = n4542 & ~n9080 ;
  assign n9082 = n9081 ^ n3412 ^ 1'b0 ;
  assign n9083 = n9075 | n9082 ;
  assign n9084 = n9083 ^ n6954 ^ 1'b0 ;
  assign n9085 = ( n2687 & ~n3263 ) | ( n2687 & n3896 ) | ( ~n3263 & n3896 ) ;
  assign n9086 = n4735 & n9085 ;
  assign n9087 = ~n7303 & n9086 ;
  assign n9092 = n8008 & n8380 ;
  assign n9093 = n9092 ^ n3335 ^ 1'b0 ;
  assign n9094 = ( n1934 & n6336 ) | ( n1934 & ~n9093 ) | ( n6336 & ~n9093 ) ;
  assign n9088 = n3304 | n4471 ;
  assign n9089 = n9088 ^ n3844 ^ 1'b0 ;
  assign n9090 = n2350 | n6783 ;
  assign n9091 = n9089 & ~n9090 ;
  assign n9095 = n9094 ^ n9091 ^ n962 ;
  assign n9096 = n2471 | n7228 ;
  assign n9097 = ~n2953 & n6705 ;
  assign n9098 = n9097 ^ n1523 ^ 1'b0 ;
  assign n9099 = ~n3532 & n9098 ;
  assign n9105 = n8335 ^ n5878 ^ 1'b0 ;
  assign n9106 = ~n6750 & n9105 ;
  assign n9107 = n9106 ^ n2779 ^ 1'b0 ;
  assign n9100 = n4533 | n5538 ;
  assign n9101 = ( n563 & n1880 ) | ( n563 & ~n1881 ) | ( n1880 & ~n1881 ) ;
  assign n9102 = n6021 | n7112 ;
  assign n9103 = n9101 | n9102 ;
  assign n9104 = n9100 & n9103 ;
  assign n9108 = n9107 ^ n9104 ^ 1'b0 ;
  assign n9109 = n3181 ^ x10 ^ 1'b0 ;
  assign n9110 = n6867 | n9109 ;
  assign n9111 = ( n3761 & ~n6972 ) | ( n3761 & n9110 ) | ( ~n6972 & n9110 ) ;
  assign n9112 = n990 & n2541 ;
  assign n9113 = n9112 ^ n2729 ^ 1'b0 ;
  assign n9114 = n5324 ^ n3901 ^ 1'b0 ;
  assign n9115 = ~n6205 & n9114 ;
  assign n9116 = ~n6353 & n9115 ;
  assign n9117 = n2528 | n5620 ;
  assign n9118 = n9116 & ~n9117 ;
  assign n9119 = n5979 ^ n792 ^ n694 ;
  assign n9120 = n2510 ^ n948 ^ 1'b0 ;
  assign n9121 = ~n2469 & n9120 ;
  assign n9122 = n965 & n9121 ;
  assign n9123 = n931 & ~n9122 ;
  assign n9124 = n8130 & n9123 ;
  assign n9125 = n1647 | n2553 ;
  assign n9126 = ~n51 & n585 ;
  assign n9127 = n9126 ^ n1237 ^ 1'b0 ;
  assign n9128 = n9127 ^ n4985 ^ 1'b0 ;
  assign n9129 = ~n7352 & n9128 ;
  assign n9130 = n9129 ^ n7615 ^ 1'b0 ;
  assign n9131 = n5541 ^ n3489 ^ n1612 ;
  assign n9132 = ( n4057 & n5806 ) | ( n4057 & n9131 ) | ( n5806 & n9131 ) ;
  assign n9133 = n4962 & ~n6774 ;
  assign n9134 = n9133 ^ n1322 ^ 1'b0 ;
  assign n9135 = n1295 & n9134 ;
  assign n9136 = n9132 & n9135 ;
  assign n9137 = ~n4530 & n9136 ;
  assign n9138 = ( ~n5195 & n5820 ) | ( ~n5195 & n5957 ) | ( n5820 & n5957 ) ;
  assign n9139 = n890 & n9138 ;
  assign n9140 = n3645 ^ n2209 ^ 1'b0 ;
  assign n9141 = n9140 ^ n9126 ^ 1'b0 ;
  assign n9142 = n9141 ^ n2422 ^ 1'b0 ;
  assign n9143 = ( n1602 & ~n3133 ) | ( n1602 & n3195 ) | ( ~n3133 & n3195 ) ;
  assign n9144 = n1693 ^ n20 ^ 1'b0 ;
  assign n9145 = n9144 ^ n6528 ^ n5356 ;
  assign n9146 = n3931 & ~n6788 ;
  assign n9147 = ~n3686 & n9146 ;
  assign n9148 = n9147 ^ n1241 ^ n811 ;
  assign n9149 = n667 & n8871 ;
  assign n9150 = n9149 ^ n1256 ^ n164 ;
  assign n9151 = ( n401 & ~n661 ) | ( n401 & n3563 ) | ( ~n661 & n3563 ) ;
  assign n9152 = n9151 ^ n134 ^ 1'b0 ;
  assign n9155 = n2216 & n3027 ;
  assign n9153 = n4819 & ~n8141 ;
  assign n9154 = n946 & n9153 ;
  assign n9156 = n9155 ^ n9154 ^ 1'b0 ;
  assign n9157 = n3470 | n4099 ;
  assign n9158 = n9157 ^ n2288 ^ 1'b0 ;
  assign n9159 = ~n6611 & n8128 ;
  assign n9160 = n5443 ^ n3626 ^ 1'b0 ;
  assign n9161 = n4454 & n9160 ;
  assign n9162 = ~n3543 & n3581 ;
  assign n9163 = n1560 & ~n9162 ;
  assign n9164 = n4641 & n9163 ;
  assign n9165 = n4986 ^ n3610 ^ 1'b0 ;
  assign n9166 = n122 | n7223 ;
  assign n9167 = n3891 & ~n9166 ;
  assign n9168 = ~n9165 & n9167 ;
  assign n9169 = n694 & n3402 ;
  assign n9170 = ~n98 & n9169 ;
  assign n9171 = n2646 & n9170 ;
  assign n9172 = n252 & n5107 ;
  assign n9173 = n9172 ^ n795 ^ 1'b0 ;
  assign n9174 = n176 | n7631 ;
  assign n9175 = n7778 | n9174 ;
  assign n9176 = n2614 | n7641 ;
  assign n9177 = ~n2108 & n2370 ;
  assign n9178 = n9177 ^ n7581 ^ 1'b0 ;
  assign n9179 = ( n7213 & n8057 ) | ( n7213 & ~n9178 ) | ( n8057 & ~n9178 ) ;
  assign n9180 = n2425 & n2625 ;
  assign n9181 = n9180 ^ n7796 ^ 1'b0 ;
  assign n9182 = n1595 & ~n3988 ;
  assign n9183 = n772 & n9182 ;
  assign n9184 = n287 | n915 ;
  assign n9185 = n9184 ^ n3466 ^ 1'b0 ;
  assign n9186 = n2723 & ~n9185 ;
  assign n9187 = n2728 ^ n122 ^ 1'b0 ;
  assign n9188 = n9186 & ~n9187 ;
  assign n9189 = ( n2253 & n9183 ) | ( n2253 & n9188 ) | ( n9183 & n9188 ) ;
  assign n9190 = n5242 ^ n2370 ^ 1'b0 ;
  assign n9191 = n5932 & n9190 ;
  assign n9192 = n9191 ^ n310 ^ 1'b0 ;
  assign n9193 = n4937 ^ n1286 ^ 1'b0 ;
  assign n9196 = n3102 | n7197 ;
  assign n9195 = n2648 ^ n1614 ^ 1'b0 ;
  assign n9194 = ( n68 & n5870 ) | ( n68 & ~n6752 ) | ( n5870 & ~n6752 ) ;
  assign n9197 = n9196 ^ n9195 ^ n9194 ;
  assign n9198 = ~n3122 & n3508 ;
  assign n9199 = n6700 & n9198 ;
  assign n9200 = n3962 ^ n3031 ^ 1'b0 ;
  assign n9201 = ( ~n5483 & n9199 ) | ( ~n5483 & n9200 ) | ( n9199 & n9200 ) ;
  assign n9202 = n7023 ^ n5485 ^ 1'b0 ;
  assign n9203 = n7350 & ~n9202 ;
  assign n9204 = n9201 & n9203 ;
  assign n9205 = n70 & ~n3299 ;
  assign n9206 = n7455 & n9205 ;
  assign n9209 = n178 & n5648 ;
  assign n9207 = ~n817 & n2214 ;
  assign n9208 = ~n1474 & n9207 ;
  assign n9210 = n9209 ^ n9208 ^ 1'b0 ;
  assign n9211 = n6366 | n9210 ;
  assign n9212 = n3345 | n8301 ;
  assign n9213 = n1568 & ~n9212 ;
  assign n9214 = n9211 | n9213 ;
  assign n9215 = n9206 & ~n9214 ;
  assign n9216 = ~n4391 & n7600 ;
  assign n9217 = n59 | n3686 ;
  assign n9218 = ( n2280 & n6868 ) | ( n2280 & n9217 ) | ( n6868 & n9217 ) ;
  assign n9219 = ~n2718 & n9218 ;
  assign n9220 = n645 & n9219 ;
  assign n9221 = n9220 ^ n3885 ^ n3241 ;
  assign n9222 = ~n1997 & n2925 ;
  assign n9223 = n1282 & n9222 ;
  assign n9224 = n3615 ^ n1290 ^ 1'b0 ;
  assign n9225 = n9224 ^ n7356 ^ 1'b0 ;
  assign n9226 = ~n8017 & n9225 ;
  assign n9227 = ( n999 & n1153 ) | ( n999 & n2320 ) | ( n1153 & n2320 ) ;
  assign n9228 = n3906 | n9227 ;
  assign n9229 = ~n6182 & n9228 ;
  assign n9230 = n9229 ^ n4862 ^ 1'b0 ;
  assign n9231 = n6011 & n6887 ;
  assign n9232 = n9231 ^ n8072 ^ n1170 ;
  assign n9233 = n493 & ~n1116 ;
  assign n9234 = n9233 ^ n8195 ^ 1'b0 ;
  assign n9235 = n1487 | n9234 ;
  assign n9236 = ~n3703 & n9235 ;
  assign n9237 = ~n722 & n5925 ;
  assign n9238 = n5678 & n9237 ;
  assign n9239 = n3967 & n8976 ;
  assign n9240 = n9239 ^ n3157 ^ 1'b0 ;
  assign n9241 = n649 ^ n532 ^ 1'b0 ;
  assign n9242 = n9241 ^ n3254 ^ n1056 ;
  assign n9243 = n9242 ^ n5502 ^ 1'b0 ;
  assign n9244 = ~n7452 & n9243 ;
  assign n9245 = n7490 ^ n732 ^ n256 ;
  assign n9246 = ~n9244 & n9245 ;
  assign n9247 = n9246 ^ n6934 ^ 1'b0 ;
  assign n9248 = ~n2181 & n9247 ;
  assign n9249 = n5289 ^ n1246 ^ 1'b0 ;
  assign n9250 = ~n3565 & n9249 ;
  assign n9251 = n2471 ^ n1518 ^ 1'b0 ;
  assign n9252 = n9251 ^ n4857 ^ 1'b0 ;
  assign n9253 = n9250 & n9252 ;
  assign n9254 = n3040 & n9253 ;
  assign n9255 = n9254 ^ n356 ^ 1'b0 ;
  assign n9256 = n5570 ^ n2586 ^ 1'b0 ;
  assign n9257 = n70 & n9256 ;
  assign n9258 = n3269 ^ n2848 ^ 1'b0 ;
  assign n9259 = n5766 ^ n3989 ^ 1'b0 ;
  assign n9260 = n3995 & ~n9259 ;
  assign n9261 = ( n3435 & n5420 ) | ( n3435 & n9260 ) | ( n5420 & n9260 ) ;
  assign n9262 = ~n9258 & n9261 ;
  assign n9263 = ( ~n6886 & n7154 ) | ( ~n6886 & n9262 ) | ( n7154 & n9262 ) ;
  assign n9264 = n1124 & ~n3755 ;
  assign n9265 = n9264 ^ n8543 ^ n4181 ;
  assign n9266 = ~n3270 & n9265 ;
  assign n9267 = ~n9263 & n9266 ;
  assign n9268 = n4686 & n5535 ;
  assign n9269 = n9268 ^ n2375 ^ 1'b0 ;
  assign n9270 = n89 & n2164 ;
  assign n9271 = ~n6583 & n9270 ;
  assign n9272 = n9271 ^ n57 ^ 1'b0 ;
  assign n9273 = n9272 ^ n3478 ^ 1'b0 ;
  assign n9274 = ( ~n214 & n890 ) | ( ~n214 & n4799 ) | ( n890 & n4799 ) ;
  assign n9275 = n5153 | n5951 ;
  assign n9276 = n3386 & n7111 ;
  assign n9277 = n6722 ^ n4729 ^ 1'b0 ;
  assign n9278 = n5229 & n9277 ;
  assign n9279 = n533 | n3797 ;
  assign n9281 = ( n558 & n1639 ) | ( n558 & ~n3354 ) | ( n1639 & ~n3354 ) ;
  assign n9280 = n2589 & n5582 ;
  assign n9282 = n9281 ^ n9280 ^ 1'b0 ;
  assign n9283 = ( ~n8403 & n9279 ) | ( ~n8403 & n9282 ) | ( n9279 & n9282 ) ;
  assign n9284 = n5119 | n5915 ;
  assign n9287 = n7328 ^ n2001 ^ 1'b0 ;
  assign n9288 = n8349 & n9287 ;
  assign n9289 = n6851 & n9288 ;
  assign n9290 = n8188 & n9289 ;
  assign n9285 = ~n276 & n971 ;
  assign n9286 = n5700 & n9285 ;
  assign n9291 = n9290 ^ n9286 ^ 1'b0 ;
  assign n9292 = n4216 | n9291 ;
  assign n9293 = n4134 | n9292 ;
  assign n9294 = n342 | n871 ;
  assign n9295 = n61 & ~n9294 ;
  assign n9296 = n1361 & ~n9295 ;
  assign n9297 = n9296 ^ n6011 ^ 1'b0 ;
  assign n9298 = n3563 & ~n9297 ;
  assign n9299 = ( ~n4549 & n5602 ) | ( ~n4549 & n9298 ) | ( n5602 & n9298 ) ;
  assign n9302 = n309 & n7047 ;
  assign n9303 = n9302 ^ n764 ^ 1'b0 ;
  assign n9300 = ( ~n360 & n2561 ) | ( ~n360 & n5563 ) | ( n2561 & n5563 ) ;
  assign n9301 = ~n961 & n9300 ;
  assign n9304 = n9303 ^ n9301 ^ 1'b0 ;
  assign n9305 = n4341 ^ n2596 ^ 1'b0 ;
  assign n9306 = n5831 | n9305 ;
  assign n9307 = ~n1209 & n3909 ;
  assign n9308 = n4047 ^ n1716 ^ n570 ;
  assign n9309 = n9308 ^ n8145 ^ n1370 ;
  assign n9310 = ~n9307 & n9309 ;
  assign n9311 = n5164 & n9310 ;
  assign n9312 = n1348 | n6008 ;
  assign n9313 = n2367 | n3447 ;
  assign n9314 = n7844 ^ n7113 ^ 1'b0 ;
  assign n9315 = n9314 ^ n8826 ^ 1'b0 ;
  assign n9317 = n2676 ^ n882 ^ 1'b0 ;
  assign n9316 = ~n5178 & n7237 ;
  assign n9318 = n9317 ^ n9316 ^ 1'b0 ;
  assign n9319 = n3699 | n9318 ;
  assign n9320 = n7254 | n9319 ;
  assign n9321 = n2326 ^ n1796 ^ 1'b0 ;
  assign n9322 = n9321 ^ n1748 ^ 1'b0 ;
  assign n9323 = ( n368 & n7234 ) | ( n368 & n9322 ) | ( n7234 & n9322 ) ;
  assign n9324 = n7657 ^ n6977 ^ n6414 ;
  assign n9325 = n1176 | n5572 ;
  assign n9326 = n6720 ^ n4767 ^ 1'b0 ;
  assign n9327 = n4719 & n7116 ;
  assign n9328 = n9327 ^ n240 ^ 1'b0 ;
  assign n9329 = ~n4489 & n5806 ;
  assign n9330 = ~n203 & n9329 ;
  assign n9331 = ~n621 & n9330 ;
  assign n9332 = ~n968 & n3373 ;
  assign n9333 = n6833 & n9332 ;
  assign n9334 = ( n4158 & ~n6524 ) | ( n4158 & n9179 ) | ( ~n6524 & n9179 ) ;
  assign n9335 = n1461 ^ n1026 ^ n650 ;
  assign n9336 = ( n2513 & ~n6122 ) | ( n2513 & n9335 ) | ( ~n6122 & n9335 ) ;
  assign n9337 = n9336 ^ n4291 ^ 1'b0 ;
  assign n9338 = n1861 ^ n691 ^ 1'b0 ;
  assign n9339 = n3174 & ~n9338 ;
  assign n9340 = n2464 & ~n9339 ;
  assign n9343 = n1988 ^ n137 ^ 1'b0 ;
  assign n9344 = n1137 | n9343 ;
  assign n9345 = n9344 ^ n2019 ^ n139 ;
  assign n9346 = ~n8906 & n9345 ;
  assign n9341 = n9246 ^ n8894 ^ 1'b0 ;
  assign n9342 = n403 & ~n9341 ;
  assign n9347 = n9346 ^ n9342 ^ 1'b0 ;
  assign n9349 = n2365 | n4502 ;
  assign n9350 = n9349 ^ n6389 ^ 1'b0 ;
  assign n9348 = ~n411 & n1746 ;
  assign n9351 = n9350 ^ n9348 ^ 1'b0 ;
  assign n9352 = n6862 ^ n4704 ^ n4024 ;
  assign n9353 = n9352 ^ n5571 ^ 1'b0 ;
  assign n9354 = ( n1875 & n3367 ) | ( n1875 & ~n5896 ) | ( n3367 & ~n5896 ) ;
  assign n9355 = n3923 ^ n3384 ^ 1'b0 ;
  assign n9356 = n3443 ^ n170 ^ 1'b0 ;
  assign n9357 = ~n6495 & n9356 ;
  assign n9358 = n3452 & ~n4927 ;
  assign n9359 = n2653 | n9358 ;
  assign n9360 = n9359 ^ n3345 ^ 1'b0 ;
  assign n9361 = n4253 & n9360 ;
  assign n9362 = ( n1787 & n1791 ) | ( n1787 & n5877 ) | ( n1791 & n5877 ) ;
  assign n9363 = ~n3564 & n9362 ;
  assign n9364 = n1412 | n4390 ;
  assign n9365 = n9364 ^ n884 ^ 1'b0 ;
  assign n9366 = n2825 | n9365 ;
  assign n9367 = n9366 ^ n8251 ^ 1'b0 ;
  assign n9368 = ~n1126 & n6100 ;
  assign n9369 = n9368 ^ n7457 ^ 1'b0 ;
  assign n9370 = n4701 & ~n6475 ;
  assign n9371 = n9369 & n9370 ;
  assign n9372 = n8961 ^ n7940 ^ n4345 ;
  assign n9373 = n1463 ^ n41 ^ 1'b0 ;
  assign n9374 = n9373 ^ n4334 ^ 1'b0 ;
  assign n9375 = n3432 & ~n6972 ;
  assign n9376 = ~n1169 & n9375 ;
  assign n9377 = n3967 | n6960 ;
  assign n9378 = ( n1737 & n9376 ) | ( n1737 & n9377 ) | ( n9376 & n9377 ) ;
  assign n9379 = ( n8188 & n9374 ) | ( n8188 & ~n9378 ) | ( n9374 & ~n9378 ) ;
  assign n9380 = ~n5200 & n5520 ;
  assign n9381 = n7558 ^ n6297 ^ 1'b0 ;
  assign n9382 = n3392 | n9381 ;
  assign n9383 = n9380 | n9382 ;
  assign n9384 = n9383 ^ n8911 ^ 1'b0 ;
  assign n9385 = n1235 & n1699 ;
  assign n9386 = ( ~n942 & n2258 ) | ( ~n942 & n9385 ) | ( n2258 & n9385 ) ;
  assign n9387 = n3088 & n9245 ;
  assign n9388 = n9387 ^ n1238 ^ 1'b0 ;
  assign n9389 = n5522 & n6756 ;
  assign n9390 = ~n9388 & n9389 ;
  assign n9391 = n9390 ^ n4645 ^ 1'b0 ;
  assign n9392 = n8049 ^ n3383 ^ 1'b0 ;
  assign n9393 = n5052 ^ n1238 ^ 1'b0 ;
  assign n9394 = ~n6330 & n9393 ;
  assign n9395 = n9394 ^ n9216 ^ 1'b0 ;
  assign n9396 = n32 & ~n4477 ;
  assign n9397 = n916 & n9396 ;
  assign n9398 = n2216 & ~n9397 ;
  assign n9399 = ~n2918 & n9398 ;
  assign n9400 = n668 | n4730 ;
  assign n9401 = n9400 ^ n3131 ^ 1'b0 ;
  assign n9402 = n5227 ^ n4568 ^ 1'b0 ;
  assign n9403 = ~n3983 & n6115 ;
  assign n9404 = n6761 & n9403 ;
  assign n9405 = n5948 | n9404 ;
  assign n9406 = n9405 ^ n4723 ^ 1'b0 ;
  assign n9407 = n1595 & n2510 ;
  assign n9408 = n9407 ^ n2226 ^ 1'b0 ;
  assign n9409 = ( n695 & n9406 ) | ( n695 & n9408 ) | ( n9406 & n9408 ) ;
  assign n9414 = n4971 ^ n1691 ^ 1'b0 ;
  assign n9410 = n1339 ^ n1109 ^ 1'b0 ;
  assign n9411 = n3324 | n9410 ;
  assign n9412 = n1262 & ~n9411 ;
  assign n9413 = n2348 & n9412 ;
  assign n9415 = n9414 ^ n9413 ^ 1'b0 ;
  assign n9416 = n1367 ^ n1094 ^ n905 ;
  assign n9417 = n4084 & n9416 ;
  assign n9418 = ( n1237 & ~n1553 ) | ( n1237 & n9417 ) | ( ~n1553 & n9417 ) ;
  assign n9419 = n5848 ^ n5809 ^ n5285 ;
  assign n9420 = n9419 ^ n4260 ^ n2592 ;
  assign n9421 = n9420 ^ n8551 ^ 1'b0 ;
  assign n9422 = n381 & ~n9421 ;
  assign n9423 = n5353 & n7941 ;
  assign n9424 = n6128 ^ n2374 ^ 1'b0 ;
  assign n9425 = n8208 ^ n3948 ^ n968 ;
  assign n9426 = n3838 ^ n1852 ^ 1'b0 ;
  assign n9427 = n6564 & ~n8756 ;
  assign n9428 = n1310 & n9427 ;
  assign n9429 = n9426 | n9428 ;
  assign n9430 = n1627 | n9429 ;
  assign n9431 = ~n1346 & n9131 ;
  assign n9432 = n9431 ^ n2451 ^ 1'b0 ;
  assign n9433 = n6051 ^ n2807 ^ n514 ;
  assign n9434 = n1564 ^ n401 ^ 1'b0 ;
  assign n9435 = n9433 & ~n9434 ;
  assign n9436 = n929 & n5372 ;
  assign n9437 = n2623 & ~n5361 ;
  assign n9438 = n563 & n9437 ;
  assign n9439 = n2871 & ~n3500 ;
  assign n9440 = n1380 ^ n1289 ^ n819 ;
  assign n9441 = n9440 ^ n8673 ^ 1'b0 ;
  assign n9442 = n845 ^ n826 ^ 1'b0 ;
  assign n9443 = n4939 & ~n9442 ;
  assign n9445 = n263 & n2125 ;
  assign n9446 = n9445 ^ n7956 ^ 1'b0 ;
  assign n9447 = n9446 ^ n2879 ^ 1'b0 ;
  assign n9448 = n4889 | n9447 ;
  assign n9444 = n4972 ^ n1274 ^ 1'b0 ;
  assign n9449 = n9448 ^ n9444 ^ 1'b0 ;
  assign n9450 = n5913 ^ n910 ^ 1'b0 ;
  assign n9451 = ( n3059 & ~n8158 ) | ( n3059 & n9450 ) | ( ~n8158 & n9450 ) ;
  assign n9452 = n8555 ^ n5481 ^ n1221 ;
  assign n9453 = n734 & n6520 ;
  assign n9454 = ( n7049 & n9452 ) | ( n7049 & ~n9453 ) | ( n9452 & ~n9453 ) ;
  assign n9455 = n3745 ^ n629 ^ 1'b0 ;
  assign n9456 = n5392 ^ n1220 ^ 1'b0 ;
  assign n9457 = ~n9455 & n9456 ;
  assign n9458 = n1777 | n8960 ;
  assign n9459 = n7275 | n9458 ;
  assign n9460 = n3521 & n9459 ;
  assign n9464 = n5377 ^ n1043 ^ 1'b0 ;
  assign n9465 = ~n7057 & n9464 ;
  assign n9461 = n1919 & ~n3891 ;
  assign n9462 = ~n7374 & n9461 ;
  assign n9463 = ~n471 & n9462 ;
  assign n9466 = n9465 ^ n9463 ^ 1'b0 ;
  assign n9467 = n697 & n9466 ;
  assign n9468 = ( n1893 & ~n5346 ) | ( n1893 & n8713 ) | ( ~n5346 & n8713 ) ;
  assign n9469 = n9468 ^ n3334 ^ 1'b0 ;
  assign n9470 = n4311 & ~n9469 ;
  assign n9471 = n1465 ^ n1411 ^ n1387 ;
  assign n9472 = n3157 & ~n9471 ;
  assign n9473 = n9472 ^ n2184 ^ 1'b0 ;
  assign n9474 = n9473 ^ n2790 ^ 1'b0 ;
  assign n9475 = ~n5236 & n5599 ;
  assign n9476 = n9475 ^ x7 ^ 1'b0 ;
  assign n9477 = n9474 | n9476 ;
  assign n9478 = n9470 | n9477 ;
  assign n9479 = n9220 ^ n6852 ^ 1'b0 ;
  assign n9480 = n9479 ^ n736 ^ 1'b0 ;
  assign n9481 = n2913 | n9480 ;
  assign n9482 = ~n545 & n2845 ;
  assign n9483 = n9482 ^ n2077 ^ 1'b0 ;
  assign n9484 = n2421 ^ n326 ^ 1'b0 ;
  assign n9485 = n2925 & n2976 ;
  assign n9488 = n6024 & n8234 ;
  assign n9489 = n9488 ^ n5831 ^ 1'b0 ;
  assign n9490 = n9489 ^ n5490 ^ n164 ;
  assign n9491 = n1737 & n5822 ;
  assign n9492 = n9490 & n9491 ;
  assign n9486 = ( n3045 & n5295 ) | ( n3045 & n6996 ) | ( n5295 & n6996 ) ;
  assign n9487 = n5102 | n9486 ;
  assign n9493 = n9492 ^ n9487 ^ n7216 ;
  assign n9494 = n4552 ^ n2906 ^ n1167 ;
  assign n9495 = n9494 ^ n3294 ^ n42 ;
  assign n9496 = ( n1661 & n6860 ) | ( n1661 & n9495 ) | ( n6860 & n9495 ) ;
  assign n9497 = n3926 ^ n2321 ^ 1'b0 ;
  assign n9498 = n2081 & ~n9497 ;
  assign n9499 = n9498 ^ n2791 ^ 1'b0 ;
  assign n9500 = n9496 & ~n9499 ;
  assign n9501 = n1665 | n9500 ;
  assign n9502 = n5069 & ~n8035 ;
  assign n9503 = n976 & n9502 ;
  assign n9504 = n8131 ^ n1406 ^ 1'b0 ;
  assign n9505 = ~n730 & n4869 ;
  assign n9506 = n9505 ^ n1842 ^ 1'b0 ;
  assign n9507 = ~n299 & n2009 ;
  assign n9508 = n1439 | n9507 ;
  assign n9509 = n1176 & ~n9508 ;
  assign n9510 = n1303 & n3406 ;
  assign n9511 = n8970 & n9510 ;
  assign n9512 = n4150 & ~n9511 ;
  assign n9513 = n9512 ^ n329 ^ 1'b0 ;
  assign n9514 = n9509 | n9513 ;
  assign n9515 = n2297 | n4226 ;
  assign n9516 = n9515 ^ n2552 ^ 1'b0 ;
  assign n9517 = n1548 ^ n234 ^ 1'b0 ;
  assign n9518 = n9516 & n9517 ;
  assign n9519 = n4214 & n9518 ;
  assign n9520 = n9519 ^ n3377 ^ n3294 ;
  assign n9521 = n3454 & n9520 ;
  assign n9522 = n9514 & n9521 ;
  assign n9523 = ~n3092 & n7418 ;
  assign n9524 = n7094 & n9523 ;
  assign n9525 = n916 & ~n9524 ;
  assign n9526 = n9525 ^ n1775 ^ 1'b0 ;
  assign n9527 = n1674 & n6264 ;
  assign n9528 = n744 | n6869 ;
  assign n9529 = n2897 | n3592 ;
  assign n9530 = n5364 & ~n8958 ;
  assign n9531 = n8329 ^ n580 ^ 1'b0 ;
  assign n9532 = n3309 & ~n9531 ;
  assign n9533 = n9532 ^ n7650 ^ 1'b0 ;
  assign n9534 = ~n3892 & n3934 ;
  assign n9535 = n9534 ^ n8558 ^ 1'b0 ;
  assign n9536 = n9535 ^ n1600 ^ 1'b0 ;
  assign n9537 = n1302 ^ n957 ^ 1'b0 ;
  assign n9538 = n3739 & ~n9537 ;
  assign n9539 = ( n563 & ~n856 ) | ( n563 & n9538 ) | ( ~n856 & n9538 ) ;
  assign n9540 = n9539 ^ n8234 ^ 1'b0 ;
  assign n9541 = n2045 & ~n9540 ;
  assign n9542 = n9541 ^ n1746 ^ 1'b0 ;
  assign n9543 = ~n9536 & n9542 ;
  assign n9544 = n7218 | n8692 ;
  assign n9545 = n6978 & n9544 ;
  assign n9546 = n9250 ^ n5637 ^ 1'b0 ;
  assign n9547 = n1156 & ~n9546 ;
  assign n9548 = n1294 & n9547 ;
  assign n9549 = n7675 ^ x10 ^ 1'b0 ;
  assign n9550 = n33 & ~n3850 ;
  assign n9551 = n1026 & ~n5512 ;
  assign n9552 = ~n3057 & n9551 ;
  assign n9553 = ( ~n9549 & n9550 ) | ( ~n9549 & n9552 ) | ( n9550 & n9552 ) ;
  assign n9554 = n6566 ^ n1526 ^ 1'b0 ;
  assign n9555 = n6276 & n9554 ;
  assign n9556 = ~n321 & n9555 ;
  assign n9557 = n9556 ^ n9148 ^ 1'b0 ;
  assign n9558 = n2280 & ~n5861 ;
  assign n9559 = n3426 | n9558 ;
  assign n9560 = n9559 ^ n4541 ^ 1'b0 ;
  assign n9561 = n7417 & n9560 ;
  assign n9562 = n2454 & n9561 ;
  assign n9563 = n5197 ^ n887 ^ 1'b0 ;
  assign n9564 = ( n5284 & n5572 ) | ( n5284 & ~n6396 ) | ( n5572 & ~n6396 ) ;
  assign n9565 = ~n1701 & n9564 ;
  assign n9566 = n536 & n1302 ;
  assign n9567 = n9566 ^ n1103 ^ 1'b0 ;
  assign n9568 = ~n9565 & n9567 ;
  assign n9575 = n2966 ^ n833 ^ 1'b0 ;
  assign n9576 = n2190 & n9575 ;
  assign n9572 = n4121 ^ n2340 ^ 1'b0 ;
  assign n9573 = n756 | n9572 ;
  assign n9574 = n3524 & ~n9573 ;
  assign n9577 = n9576 ^ n9574 ^ 1'b0 ;
  assign n9569 = n7541 ^ n7163 ^ 1'b0 ;
  assign n9570 = n5625 & n9569 ;
  assign n9571 = ( n230 & n4058 ) | ( n230 & n9570 ) | ( n4058 & n9570 ) ;
  assign n9578 = n9577 ^ n9571 ^ n4562 ;
  assign n9582 = n8980 ^ n3569 ^ 1'b0 ;
  assign n9583 = n246 & n9582 ;
  assign n9579 = n839 & ~n7490 ;
  assign n9580 = n4009 & n9579 ;
  assign n9581 = n7893 | n9580 ;
  assign n9584 = n9583 ^ n9581 ^ 1'b0 ;
  assign n9585 = n3214 ^ n383 ^ 1'b0 ;
  assign n9586 = ~n5663 & n9585 ;
  assign n9587 = ~n1296 & n6288 ;
  assign n9588 = n9587 ^ n2004 ^ 1'b0 ;
  assign n9589 = n9588 ^ n3660 ^ n3266 ;
  assign n9590 = n6909 ^ n923 ^ 1'b0 ;
  assign n9591 = n1360 | n9590 ;
  assign n9592 = n3564 & ~n9591 ;
  assign n9593 = ~n2172 & n9592 ;
  assign n9594 = n9593 ^ n1405 ^ 1'b0 ;
  assign n9595 = ~n1723 & n3872 ;
  assign n9596 = n4001 & n9595 ;
  assign n9597 = ~n4099 & n7186 ;
  assign n9598 = n7939 ^ n3082 ^ 1'b0 ;
  assign n9599 = n6456 ^ n4894 ^ 1'b0 ;
  assign n9600 = n7563 & ~n9599 ;
  assign n9601 = ( n1561 & n3904 ) | ( n1561 & n4208 ) | ( n3904 & n4208 ) ;
  assign n9602 = n9601 ^ n5072 ^ 1'b0 ;
  assign n9603 = n247 & n9602 ;
  assign n9604 = n9603 ^ n41 ^ 1'b0 ;
  assign n9605 = n9446 & n9604 ;
  assign n9607 = n4653 ^ n1827 ^ 1'b0 ;
  assign n9608 = n7650 & n9607 ;
  assign n9609 = n3940 | n4390 ;
  assign n9610 = n1490 | n9609 ;
  assign n9611 = n9610 ^ n6225 ^ 1'b0 ;
  assign n9612 = n9608 & ~n9611 ;
  assign n9606 = n8210 ^ n2231 ^ n416 ;
  assign n9613 = n9612 ^ n9606 ^ 1'b0 ;
  assign n9614 = ~n4002 & n7852 ;
  assign n9615 = ~n1173 & n7284 ;
  assign n9616 = n9615 ^ n6667 ^ 1'b0 ;
  assign n9617 = n406 & ~n3116 ;
  assign n9618 = n9617 ^ n1664 ^ 1'b0 ;
  assign n9619 = ~n7878 & n9618 ;
  assign n9622 = n3772 ^ n2991 ^ 1'b0 ;
  assign n9623 = n563 & ~n9622 ;
  assign n9624 = n9623 ^ n5183 ^ n1853 ;
  assign n9620 = ( n6793 & n7886 ) | ( n6793 & ~n8784 ) | ( n7886 & ~n8784 ) ;
  assign n9621 = n9620 ^ n4319 ^ n3034 ;
  assign n9625 = n9624 ^ n9621 ^ 1'b0 ;
  assign n9626 = n922 | n2889 ;
  assign n9627 = n2164 | n3312 ;
  assign n9628 = n1801 & n3886 ;
  assign n9629 = n1854 ^ n44 ^ 1'b0 ;
  assign n9630 = n1888 & n9629 ;
  assign n9631 = n5754 | n9630 ;
  assign n9632 = ~n9628 & n9631 ;
  assign n9633 = n5876 & n9632 ;
  assign n9634 = ( n517 & n5179 ) | ( n517 & n6614 ) | ( n5179 & n6614 ) ;
  assign n9635 = n2140 | n3645 ;
  assign n9636 = n865 & n9635 ;
  assign n9637 = n2599 | n6253 ;
  assign n9638 = n1980 & ~n9637 ;
  assign n9639 = n2745 | n9638 ;
  assign n9640 = n668 & n5172 ;
  assign n9641 = n4364 & ~n9012 ;
  assign n9642 = n9641 ^ n9233 ^ 1'b0 ;
  assign n9643 = n9642 ^ n962 ^ 1'b0 ;
  assign n9644 = n5848 & ~n7365 ;
  assign n9645 = n5209 ^ n5147 ^ n2377 ;
  assign n9646 = ( n1114 & ~n1622 ) | ( n1114 & n6877 ) | ( ~n1622 & n6877 ) ;
  assign n9647 = ~n2025 & n5902 ;
  assign n9648 = n518 | n2152 ;
  assign n9649 = n2294 & ~n9648 ;
  assign n9650 = n7773 & ~n9649 ;
  assign n9651 = n9650 ^ n6868 ^ 1'b0 ;
  assign n9652 = n2514 | n9651 ;
  assign n9653 = ~n987 & n4363 ;
  assign n9654 = n1063 & ~n7099 ;
  assign n9655 = n8793 & n9654 ;
  assign n9656 = n9655 ^ n7977 ^ 1'b0 ;
  assign n9657 = n1693 | n6426 ;
  assign n9658 = n91 | n9657 ;
  assign n9659 = n1272 & n3345 ;
  assign n9660 = n9658 & n9659 ;
  assign n9661 = n9660 ^ n3677 ^ 1'b0 ;
  assign n9662 = x6 & n7144 ;
  assign n9663 = ~n3882 & n9662 ;
  assign n9664 = n8493 ^ n6381 ^ 1'b0 ;
  assign n9665 = n735 & ~n3922 ;
  assign n9666 = n9665 ^ n424 ^ 1'b0 ;
  assign n9667 = n9666 ^ n5502 ^ n2818 ;
  assign n9668 = n725 & n1260 ;
  assign n9669 = n9667 & n9668 ;
  assign n9670 = ( n2098 & n3737 ) | ( n2098 & ~n8282 ) | ( n3737 & ~n8282 ) ;
  assign n9671 = n6223 & ~n9670 ;
  assign n9672 = n2853 | n9671 ;
  assign n9673 = n957 & ~n9672 ;
  assign n9674 = n6560 ^ n3914 ^ 1'b0 ;
  assign n9675 = n9189 ^ n8664 ^ 1'b0 ;
  assign n9676 = ~n9674 & n9675 ;
  assign n9677 = n2804 ^ n228 ^ 1'b0 ;
  assign n9678 = n9471 | n9677 ;
  assign n9679 = ~n2145 & n9678 ;
  assign n9680 = n6996 ^ n6376 ^ 1'b0 ;
  assign n9681 = n8857 ^ n3221 ^ 1'b0 ;
  assign n9682 = n2686 & n3838 ;
  assign n9683 = n769 & n9682 ;
  assign n9684 = ~n3541 & n4743 ;
  assign n9685 = n9684 ^ n927 ^ 1'b0 ;
  assign n9686 = ( ~n7523 & n9683 ) | ( ~n7523 & n9685 ) | ( n9683 & n9685 ) ;
  assign n9687 = n9603 ^ n5934 ^ n400 ;
  assign n9688 = n7844 ^ n6140 ^ n2824 ;
  assign n9689 = ~n1114 & n6874 ;
  assign n9690 = n9615 & n9689 ;
  assign n9691 = n9690 ^ n6810 ^ 1'b0 ;
  assign n9692 = n9688 & ~n9691 ;
  assign n9693 = n3079 & n9692 ;
  assign n9694 = n9693 ^ n9628 ^ 1'b0 ;
  assign n9695 = n8633 ^ n4430 ^ 1'b0 ;
  assign n9696 = n9052 & n9695 ;
  assign n9697 = n811 | n9208 ;
  assign n9698 = n9696 | n9697 ;
  assign n9699 = ( n7645 & n8580 ) | ( n7645 & ~n9628 ) | ( n8580 & ~n9628 ) ;
  assign n9700 = n5759 & ~n9402 ;
  assign n9702 = n4602 ^ n2966 ^ n865 ;
  assign n9701 = n2720 & ~n8406 ;
  assign n9703 = n9702 ^ n9701 ^ 1'b0 ;
  assign n9704 = ~n1450 & n3016 ;
  assign n9705 = n9704 ^ n5122 ^ 1'b0 ;
  assign n9706 = ( n1148 & n5261 ) | ( n1148 & n8066 ) | ( n5261 & n8066 ) ;
  assign n9707 = n774 & ~n4922 ;
  assign n9708 = n5788 | n9707 ;
  assign n9709 = n1596 | n9708 ;
  assign n9710 = n9709 ^ n3401 ^ 1'b0 ;
  assign n9711 = ~n8657 & n9710 ;
  assign n9712 = n9711 ^ n6167 ^ 1'b0 ;
  assign n9713 = n190 | n394 ;
  assign n9714 = ( ~n3680 & n4048 ) | ( ~n3680 & n9713 ) | ( n4048 & n9713 ) ;
  assign n9715 = n9714 ^ n9538 ^ 1'b0 ;
  assign n9716 = ~n2284 & n7019 ;
  assign n9720 = ~n1105 & n8595 ;
  assign n9721 = n9720 ^ n6976 ^ 1'b0 ;
  assign n9717 = n9115 ^ n8750 ^ 1'b0 ;
  assign n9718 = n6481 ^ n2582 ^ 1'b0 ;
  assign n9719 = ~n9717 & n9718 ;
  assign n9722 = n9721 ^ n9719 ^ 1'b0 ;
  assign n9723 = ( n1238 & ~n1539 ) | ( n1238 & n9265 ) | ( ~n1539 & n9265 ) ;
  assign n9724 = ~n2447 & n4536 ;
  assign n9725 = n5234 ^ n350 ^ 1'b0 ;
  assign n9726 = ~n3753 & n9725 ;
  assign n9727 = ~n5537 & n9726 ;
  assign n9728 = n4330 & ~n9727 ;
  assign n9729 = n9728 ^ n9357 ^ 1'b0 ;
  assign n9730 = n9290 | n9605 ;
  assign n9731 = n324 & ~n423 ;
  assign n9732 = ~n578 & n9731 ;
  assign n9733 = ( x9 & n6490 ) | ( x9 & n9732 ) | ( n6490 & n9732 ) ;
  assign n9734 = n272 & n9733 ;
  assign n9735 = n9734 ^ n740 ^ 1'b0 ;
  assign n9736 = ~n2534 & n9735 ;
  assign n9737 = n9736 ^ n9108 ^ n4542 ;
  assign n9738 = n3923 & ~n4880 ;
  assign n9739 = ~n2570 & n9738 ;
  assign n9740 = n9739 ^ n8024 ^ 1'b0 ;
  assign n9741 = n9740 ^ n736 ^ n298 ;
  assign n9742 = n718 | n3790 ;
  assign n9743 = n9742 ^ n3614 ^ 1'b0 ;
  assign n9744 = n9743 ^ n1535 ^ 1'b0 ;
  assign n9745 = n2187 | n9744 ;
  assign n9746 = ( ~n6426 & n7278 ) | ( ~n6426 & n9745 ) | ( n7278 & n9745 ) ;
  assign n9747 = n6638 ^ n336 ^ 1'b0 ;
  assign n9748 = ~n8016 & n9747 ;
  assign n9749 = n2539 ^ n420 ^ 1'b0 ;
  assign n9750 = n9748 & n9749 ;
  assign n9757 = n3384 & n3899 ;
  assign n9758 = ( n108 & n434 ) | ( n108 & ~n9757 ) | ( n434 & ~n9757 ) ;
  assign n9759 = n5233 & n9758 ;
  assign n9751 = n3224 ^ n760 ^ 1'b0 ;
  assign n9753 = n5585 ^ n1076 ^ 1'b0 ;
  assign n9752 = n8630 ^ n6026 ^ 1'b0 ;
  assign n9754 = n9753 ^ n9752 ^ 1'b0 ;
  assign n9755 = n5661 & n9754 ;
  assign n9756 = n9751 & n9755 ;
  assign n9760 = n9759 ^ n9756 ^ 1'b0 ;
  assign n9761 = n8856 ^ n3789 ^ 1'b0 ;
  assign n9762 = n7917 ^ n1680 ^ 1'b0 ;
  assign n9763 = n8195 | n9762 ;
  assign n9764 = ( n4647 & ~n5161 ) | ( n4647 & n9763 ) | ( ~n5161 & n9763 ) ;
  assign n9765 = ~n2930 & n5867 ;
  assign n9766 = ~n7495 & n9765 ;
  assign n9767 = ~n3085 & n6879 ;
  assign n9768 = n9767 ^ n5186 ^ 1'b0 ;
  assign n9769 = ~n1835 & n2551 ;
  assign n9770 = ( n2070 & n4574 ) | ( n2070 & n9769 ) | ( n4574 & n9769 ) ;
  assign n9771 = n7542 & n8799 ;
  assign n9772 = ~n9770 & n9771 ;
  assign n9773 = n5700 ^ n2580 ^ 1'b0 ;
  assign n9774 = n1206 | n9773 ;
  assign n9775 = n2553 | n5028 ;
  assign n9776 = n9775 ^ n4422 ^ 1'b0 ;
  assign n9777 = n9774 & n9776 ;
  assign n9778 = ~n2541 & n9777 ;
  assign n9779 = ~n2403 & n9778 ;
  assign n9780 = ( n5570 & n7332 ) | ( n5570 & n7757 ) | ( n7332 & n7757 ) ;
  assign n9781 = n8232 ^ n8164 ^ n572 ;
  assign n9782 = n9781 ^ n5519 ^ n2645 ;
  assign n9785 = n4382 ^ n1153 ^ n966 ;
  assign n9786 = n9785 ^ n1126 ^ 1'b0 ;
  assign n9787 = n2943 | n9786 ;
  assign n9783 = ( n418 & n1661 ) | ( n418 & ~n2211 ) | ( n1661 & ~n2211 ) ;
  assign n9784 = n9467 & n9783 ;
  assign n9788 = n9787 ^ n9784 ^ 1'b0 ;
  assign n9789 = n9788 ^ n7478 ^ 1'b0 ;
  assign n9790 = n6738 | n7087 ;
  assign n9791 = n7996 ^ n2395 ^ 1'b0 ;
  assign n9792 = n2049 & n9791 ;
  assign n9793 = n7697 | n9792 ;
  assign n9794 = n8625 ^ n769 ^ 1'b0 ;
  assign n9795 = n9704 ^ n4105 ^ 1'b0 ;
  assign n9796 = n3238 | n5353 ;
  assign n9797 = n9796 ^ n624 ^ 1'b0 ;
  assign n9798 = n9795 & n9797 ;
  assign n9799 = n309 & n4034 ;
  assign n9800 = n9799 ^ n5725 ^ 1'b0 ;
  assign n9801 = n9800 ^ n866 ^ 1'b0 ;
  assign n9802 = n7952 ^ n259 ^ 1'b0 ;
  assign n9803 = n260 & n3248 ;
  assign n9804 = n9803 ^ n7917 ^ 1'b0 ;
  assign n9805 = n3148 & n4230 ;
  assign n9806 = n8539 ^ n2094 ^ n1412 ;
  assign n9807 = n893 | n7493 ;
  assign n9808 = n3060 | n9807 ;
  assign n9809 = ~n1472 & n9716 ;
  assign n9810 = ~n319 & n8077 ;
  assign n9811 = n9810 ^ n3260 ^ 1'b0 ;
  assign n9812 = ~n9809 & n9811 ;
  assign n9813 = n9812 ^ n4187 ^ 1'b0 ;
  assign n9814 = n4216 & n6810 ;
  assign n9815 = n9814 ^ n448 ^ n260 ;
  assign n9816 = ( n3941 & n4365 ) | ( n3941 & ~n9815 ) | ( n4365 & ~n9815 ) ;
  assign n9817 = n1891 & n9816 ;
  assign n9818 = n5820 ^ n780 ^ 1'b0 ;
  assign n9819 = n672 & ~n5380 ;
  assign n9820 = n889 ^ n73 ^ 1'b0 ;
  assign n9821 = n4825 | n6289 ;
  assign n9822 = n9821 ^ n6474 ^ 1'b0 ;
  assign n9823 = n4639 & n9822 ;
  assign n9824 = ~n811 & n1247 ;
  assign n9825 = n9824 ^ n4308 ^ 1'b0 ;
  assign n9826 = n1630 | n9825 ;
  assign n9827 = n1943 & n4788 ;
  assign n9828 = ( n1200 & n3526 ) | ( n1200 & ~n3608 ) | ( n3526 & ~n3608 ) ;
  assign n9829 = n6115 & ~n9828 ;
  assign n9830 = n7641 ^ n777 ^ 1'b0 ;
  assign n9832 = n5276 | n9713 ;
  assign n9831 = ~n147 & n2497 ;
  assign n9833 = n9832 ^ n9831 ^ 1'b0 ;
  assign n9834 = ~n3463 & n9833 ;
  assign n9835 = n9834 ^ n7002 ^ 1'b0 ;
  assign n9836 = n9271 | n9835 ;
  assign n9837 = n9836 ^ n2836 ^ 1'b0 ;
  assign n9838 = n4328 | n9837 ;
  assign n9839 = ( n2890 & n3043 ) | ( n2890 & n5732 ) | ( n3043 & n5732 ) ;
  assign n9840 = ( n1135 & n1628 ) | ( n1135 & ~n9839 ) | ( n1628 & ~n9839 ) ;
  assign n9841 = n23 & ~n9840 ;
  assign n9842 = n4114 & n6066 ;
  assign n9843 = n523 & n9842 ;
  assign n9844 = n6917 & n8355 ;
  assign n9845 = ~n2754 & n9844 ;
  assign n9846 = n9845 ^ n4700 ^ 1'b0 ;
  assign n9847 = n9843 | n9846 ;
  assign n9852 = n496 ^ n411 ^ n318 ;
  assign n9853 = n1341 & ~n9852 ;
  assign n9849 = n3361 & ~n5406 ;
  assign n9848 = ~n7348 & n8474 ;
  assign n9850 = n9849 ^ n9848 ^ 1'b0 ;
  assign n9851 = ~n2696 & n9850 ;
  assign n9854 = n9853 ^ n9851 ^ 1'b0 ;
  assign n9855 = n5222 & n9854 ;
  assign n9856 = ~n989 & n5353 ;
  assign n9857 = ~n2461 & n9856 ;
  assign n9858 = ( n99 & ~n6289 ) | ( n99 & n9857 ) | ( ~n6289 & n9857 ) ;
  assign n9859 = n1983 | n9858 ;
  assign n9860 = n4239 & ~n9859 ;
  assign n9861 = n9855 & n9860 ;
  assign n9862 = n9861 ^ n8032 ^ 1'b0 ;
  assign n9863 = n1182 & n8639 ;
  assign n9864 = n3162 ^ n2362 ^ 1'b0 ;
  assign n9865 = ~n45 & n4733 ;
  assign n9866 = ~n2199 & n9865 ;
  assign n9867 = n2539 & ~n9866 ;
  assign n9868 = n9864 & n9867 ;
  assign n9869 = n9868 ^ n8110 ^ n7970 ;
  assign n9871 = n3679 & n4431 ;
  assign n9872 = n9871 ^ n1812 ^ 1'b0 ;
  assign n9873 = n9872 ^ n6412 ^ 1'b0 ;
  assign n9874 = n7929 & n9873 ;
  assign n9870 = ~n3798 & n8775 ;
  assign n9875 = n9874 ^ n9870 ^ 1'b0 ;
  assign n9878 = ~n6191 & n7120 ;
  assign n9879 = n9878 ^ n905 ^ 1'b0 ;
  assign n9876 = n837 | n2667 ;
  assign n9877 = n3359 | n9876 ;
  assign n9880 = n9879 ^ n9877 ^ n1431 ;
  assign n9881 = ~n4187 & n7633 ;
  assign n9882 = n9881 ^ n3893 ^ 1'b0 ;
  assign n9883 = n328 & ~n2137 ;
  assign n9884 = n1515 & n9883 ;
  assign n9885 = n8729 ^ n5519 ^ n3756 ;
  assign n9886 = n9885 ^ n2500 ^ n2195 ;
  assign n9887 = n134 & ~n3229 ;
  assign n9888 = n4116 ^ n1666 ^ 1'b0 ;
  assign n9889 = n887 & ~n9888 ;
  assign n9890 = n9889 ^ n704 ^ 1'b0 ;
  assign n9891 = n9887 & ~n9890 ;
  assign n9892 = n9886 & n9891 ;
  assign n9893 = n9892 ^ n1561 ^ 1'b0 ;
  assign n9894 = n3107 ^ n2172 ^ 1'b0 ;
  assign n9895 = n2214 ^ n637 ^ 1'b0 ;
  assign n9896 = ~n2804 & n9895 ;
  assign n9897 = n441 & n2206 ;
  assign n9898 = n9897 ^ n41 ^ 1'b0 ;
  assign n9899 = n191 | n1890 ;
  assign n9900 = ~n9898 & n9899 ;
  assign n9901 = n9900 ^ n2588 ^ 1'b0 ;
  assign n9902 = n9901 ^ n619 ^ n156 ;
  assign n9903 = n9902 ^ n44 ^ 1'b0 ;
  assign n9904 = n9903 ^ n4263 ^ n3899 ;
  assign n9905 = n4847 ^ n2666 ^ 1'b0 ;
  assign n9906 = n9792 ^ n1387 ^ 1'b0 ;
  assign n9907 = n9404 | n9906 ;
  assign n9909 = ( n142 & n962 ) | ( n142 & ~n1441 ) | ( n962 & ~n1441 ) ;
  assign n9910 = ( ~n169 & n5166 ) | ( ~n169 & n9909 ) | ( n5166 & n9909 ) ;
  assign n9908 = n9263 ^ n8754 ^ n5540 ;
  assign n9911 = n9910 ^ n9908 ^ 1'b0 ;
  assign n9912 = ~n2770 & n7541 ;
  assign n9913 = n9912 ^ n1996 ^ 1'b0 ;
  assign n9914 = n3786 & n9913 ;
  assign n9915 = n2234 & ~n9914 ;
  assign n9916 = ~n1052 & n1105 ;
  assign n9917 = n3512 & n9916 ;
  assign n9918 = n1103 | n2286 ;
  assign n9919 = ( n780 & n3709 ) | ( n780 & n9918 ) | ( n3709 & n9918 ) ;
  assign n9920 = ~n8630 & n9919 ;
  assign n9921 = ( n4348 & n4424 ) | ( n4348 & ~n7445 ) | ( n4424 & ~n7445 ) ;
  assign n9922 = n2149 & ~n9921 ;
  assign n9923 = n9922 ^ n6131 ^ 1'b0 ;
  assign n9924 = n7391 ^ n1091 ^ 1'b0 ;
  assign n9925 = n5708 & ~n9924 ;
  assign n9926 = ~n9923 & n9925 ;
  assign n9927 = ( n2831 & n7880 ) | ( n2831 & n9378 ) | ( n7880 & n9378 ) ;
  assign n9928 = n2622 & n4204 ;
  assign n9929 = n9714 & n9928 ;
  assign n9930 = ( ~n937 & n9927 ) | ( ~n937 & n9929 ) | ( n9927 & n9929 ) ;
  assign n9931 = n2025 | n9930 ;
  assign n9932 = n1823 & ~n9931 ;
  assign n9933 = n1741 ^ n927 ^ 1'b0 ;
  assign n9934 = n9933 ^ n3888 ^ 1'b0 ;
  assign n9935 = n2531 ^ n2146 ^ 1'b0 ;
  assign n9936 = n9935 ^ n1798 ^ 1'b0 ;
  assign n9937 = n9936 ^ n5047 ^ 1'b0 ;
  assign n9938 = n4892 ^ n3259 ^ 1'b0 ;
  assign n9939 = n8398 ^ n2211 ^ 1'b0 ;
  assign n9940 = n710 | n5955 ;
  assign n9941 = n2148 | n9940 ;
  assign n9942 = n9939 & n9941 ;
  assign n9943 = n8552 ^ n2892 ^ 1'b0 ;
  assign n9944 = ~n6009 & n9943 ;
  assign n9945 = ~n4021 & n9944 ;
  assign n9946 = n9945 ^ n2911 ^ 1'b0 ;
  assign n9947 = ( n4887 & ~n9463 ) | ( n4887 & n9946 ) | ( ~n9463 & n9946 ) ;
  assign n9948 = n9947 ^ n6630 ^ 1'b0 ;
  assign n9949 = n2485 | n9384 ;
  assign n9950 = n9949 ^ n8743 ^ 1'b0 ;
  assign n9951 = n966 & ~n4897 ;
  assign n9952 = n8813 | n9951 ;
  assign n9953 = ~n3170 & n4310 ;
  assign n9954 = ~n9952 & n9953 ;
  assign n9955 = ( n532 & n3181 ) | ( n532 & ~n7516 ) | ( n3181 & ~n7516 ) ;
  assign n9956 = ( n448 & ~n6475 ) | ( n448 & n9955 ) | ( ~n6475 & n9955 ) ;
  assign n9957 = n9956 ^ n6695 ^ 1'b0 ;
  assign n9958 = n3916 & n9957 ;
  assign n9959 = n6083 ^ n2573 ^ n1142 ;
  assign n9960 = n9959 ^ n2445 ^ 1'b0 ;
  assign n9961 = n7960 | n9960 ;
  assign n9962 = ~n806 & n1003 ;
  assign n9963 = ~n718 & n1167 ;
  assign n9964 = n9962 & n9963 ;
  assign n9965 = n1346 ^ n1045 ^ 1'b0 ;
  assign n9966 = n9965 ^ n1082 ^ 1'b0 ;
  assign n9967 = n9434 ^ n8889 ^ n411 ;
  assign n9968 = ( n3816 & ~n4228 ) | ( n3816 & n9967 ) | ( ~n4228 & n9967 ) ;
  assign n9969 = n2307 | n7364 ;
  assign n9970 = n1688 | n4490 ;
  assign n9971 = n9970 ^ n6136 ^ 1'b0 ;
  assign n9972 = n9969 | n9971 ;
  assign n9973 = ~n2081 & n3638 ;
  assign n9974 = ~n455 & n2484 ;
  assign n9975 = n9974 ^ n3622 ^ 1'b0 ;
  assign n9976 = n9973 | n9975 ;
  assign n9977 = n2876 | n9976 ;
  assign n9978 = n9977 ^ n3579 ^ 1'b0 ;
  assign n9979 = n1967 & ~n9978 ;
  assign n9980 = n524 & n5533 ;
  assign n9981 = n9980 ^ x8 ^ 1'b0 ;
  assign n9982 = ~n5312 & n9981 ;
  assign n9983 = n1105 & n6296 ;
  assign n9984 = n2544 ^ n2114 ^ 1'b0 ;
  assign n9985 = n5954 & n7197 ;
  assign n9986 = n7655 | n9414 ;
  assign n9987 = ( n9984 & n9985 ) | ( n9984 & ~n9986 ) | ( n9985 & ~n9986 ) ;
  assign n9988 = n2373 ^ n1889 ^ 1'b0 ;
  assign n9989 = ~n2469 & n9988 ;
  assign n9990 = ~n2680 & n9989 ;
  assign n9991 = n9990 ^ n4618 ^ 1'b0 ;
  assign n9992 = n1251 | n1545 ;
  assign n9993 = n318 | n9992 ;
  assign n9994 = ~n3372 & n9993 ;
  assign n9995 = n9994 ^ n794 ^ 1'b0 ;
  assign n9996 = n8030 ^ n4381 ^ n1848 ;
  assign n9997 = n816 | n2291 ;
  assign n9998 = n9997 ^ n7663 ^ n2794 ;
  assign n10002 = n351 & n2399 ;
  assign n10000 = n1167 & ~n8911 ;
  assign n10001 = ~n3481 & n10000 ;
  assign n9999 = n6437 ^ n2937 ^ n2851 ;
  assign n10003 = n10002 ^ n10001 ^ n9999 ;
  assign n10004 = ~n3918 & n6991 ;
  assign n10005 = n7240 & ~n10004 ;
  assign n10006 = n37 & n6261 ;
  assign n10007 = n5961 & n10006 ;
  assign n10008 = n1360 | n3777 ;
  assign n10009 = n10008 ^ n3044 ^ 1'b0 ;
  assign n10010 = ~n10007 & n10009 ;
  assign n10011 = n5954 & ~n7796 ;
  assign n10012 = n10011 ^ n3694 ^ 1'b0 ;
  assign n10013 = ~n202 & n10012 ;
  assign n10014 = ~n7279 & n10013 ;
  assign n10017 = n2316 & ~n7366 ;
  assign n10015 = n8119 ^ n5569 ^ 1'b0 ;
  assign n10016 = n2836 | n10015 ;
  assign n10018 = n10017 ^ n10016 ^ 1'b0 ;
  assign n10019 = n223 & ~n10018 ;
  assign n10020 = ~n2818 & n10019 ;
  assign n10021 = n156 | n4936 ;
  assign n10022 = n4711 & n7099 ;
  assign n10023 = ~n2591 & n10022 ;
  assign n10024 = n4502 | n10023 ;
  assign n10025 = n4093 | n10024 ;
  assign n10026 = n10025 ^ n5773 ^ 1'b0 ;
  assign n10027 = n10026 ^ n9481 ^ 1'b0 ;
  assign n10028 = n1485 | n3488 ;
  assign n10029 = n10028 ^ n2039 ^ 1'b0 ;
  assign n10030 = n9196 ^ n2595 ^ 1'b0 ;
  assign n10031 = n10029 & n10030 ;
  assign n10032 = n6050 ^ n2298 ^ 1'b0 ;
  assign n10033 = ~n3946 & n10032 ;
  assign n10035 = ~n2039 & n4544 ;
  assign n10034 = n4459 ^ n2691 ^ 1'b0 ;
  assign n10036 = n10035 ^ n10034 ^ 1'b0 ;
  assign n10037 = n3128 & n10036 ;
  assign n10038 = ~n2149 & n4724 ;
  assign n10039 = n4719 ^ n641 ^ 1'b0 ;
  assign n10040 = n582 & ~n10039 ;
  assign n10041 = n4039 & n10040 ;
  assign n10042 = ~n9008 & n10041 ;
  assign n10043 = n10038 & ~n10042 ;
  assign n10044 = ~n6360 & n10043 ;
  assign n10045 = n1518 ^ n698 ^ 1'b0 ;
  assign n10046 = n1623 & n10045 ;
  assign n10047 = n10046 ^ n6455 ^ 1'b0 ;
  assign n10048 = ~n10044 & n10047 ;
  assign n10049 = n9619 ^ n8334 ^ n8115 ;
  assign n10050 = ( n360 & ~n4368 ) | ( n360 & n9571 ) | ( ~n4368 & n9571 ) ;
  assign n10051 = n1771 | n6692 ;
  assign n10053 = n1167 ^ n1164 ^ n421 ;
  assign n10054 = n1630 & n10053 ;
  assign n10052 = n7053 ^ n5870 ^ 1'b0 ;
  assign n10055 = n10054 ^ n10052 ^ 1'b0 ;
  assign n10056 = n8001 | n8686 ;
  assign n10057 = ( n747 & n926 ) | ( n747 & n4100 ) | ( n926 & n4100 ) ;
  assign n10058 = n397 & n10057 ;
  assign n10059 = n2004 ^ n1869 ^ 1'b0 ;
  assign n10060 = n4937 | n8408 ;
  assign n10061 = ~n1135 & n7989 ;
  assign n10062 = ~n5484 & n10061 ;
  assign n10063 = ( n2885 & ~n10060 ) | ( n2885 & n10062 ) | ( ~n10060 & n10062 ) ;
  assign n10064 = n3680 & n4330 ;
  assign n10065 = n10064 ^ n2258 ^ 1'b0 ;
  assign n10066 = n10065 ^ n2316 ^ 1'b0 ;
  assign n10067 = n3268 & n4252 ;
  assign n10068 = n10067 ^ n6607 ^ 1'b0 ;
  assign n10069 = n10068 ^ n5262 ^ 1'b0 ;
  assign n10070 = n4823 & n10069 ;
  assign n10071 = n10070 ^ n2475 ^ 1'b0 ;
  assign n10072 = n10071 ^ n6380 ^ n4283 ;
  assign n10073 = n2443 ^ n2084 ^ n1403 ;
  assign n10074 = n10073 ^ n3709 ^ n104 ;
  assign n10075 = n1053 & ~n4201 ;
  assign n10076 = n5085 & n10075 ;
  assign n10077 = ( n6622 & n8912 ) | ( n6622 & ~n10076 ) | ( n8912 & ~n10076 ) ;
  assign n10078 = n1679 & ~n5106 ;
  assign n10079 = n1429 ^ n915 ^ 1'b0 ;
  assign n10080 = n6197 ^ n2098 ^ n1178 ;
  assign n10081 = n10080 ^ n8314 ^ 1'b0 ;
  assign n10082 = n10079 | n10081 ;
  assign n10083 = n2657 & n7029 ;
  assign n10084 = ~n9245 & n10083 ;
  assign n10085 = n987 & ~n10084 ;
  assign n10086 = n1784 & n4671 ;
  assign n10087 = n4111 & n8097 ;
  assign n10088 = n2145 ^ n263 ^ 1'b0 ;
  assign n10089 = n846 & ~n9162 ;
  assign n10090 = ~n10088 & n10089 ;
  assign n10091 = n10090 ^ n7483 ^ n1560 ;
  assign n10092 = n2880 & ~n4025 ;
  assign n10093 = n9717 & n10092 ;
  assign n10094 = n10093 ^ n5717 ^ n2544 ;
  assign n10095 = n2111 | n7657 ;
  assign n10096 = n9406 | n10095 ;
  assign n10097 = n4041 & n6289 ;
  assign n10098 = ~n411 & n10097 ;
  assign n10099 = n5080 & ~n10098 ;
  assign n10100 = n10099 ^ n6140 ^ 1'b0 ;
  assign n10101 = n10100 ^ n5954 ^ 1'b0 ;
  assign n10102 = n10101 ^ n923 ^ 1'b0 ;
  assign n10104 = n2853 ^ n687 ^ 1'b0 ;
  assign n10105 = n7596 | n10104 ;
  assign n10103 = n4214 & n8546 ;
  assign n10106 = n10105 ^ n10103 ^ 1'b0 ;
  assign n10107 = n650 & n4966 ;
  assign n10108 = n4862 & n10107 ;
  assign n10109 = n2719 & n7457 ;
  assign n10110 = ~n5931 & n10109 ;
  assign n10111 = ( ~n9490 & n10108 ) | ( ~n9490 & n10110 ) | ( n10108 & n10110 ) ;
  assign n10112 = n283 ^ n72 ^ 1'b0 ;
  assign n10113 = n7168 & ~n10112 ;
  assign n10114 = n10113 ^ n1585 ^ 1'b0 ;
  assign n10115 = n10114 ^ n5732 ^ n3819 ;
  assign n10118 = ( n2622 & n3354 ) | ( n2622 & ~n4443 ) | ( n3354 & ~n4443 ) ;
  assign n10119 = ~n7393 & n10118 ;
  assign n10120 = ~n2772 & n10119 ;
  assign n10116 = n1595 & ~n7441 ;
  assign n10117 = n10116 ^ n5725 ^ 1'b0 ;
  assign n10121 = n10120 ^ n10117 ^ 1'b0 ;
  assign n10122 = n799 | n10121 ;
  assign n10124 = n5045 | n10053 ;
  assign n10123 = n4674 | n7587 ;
  assign n10125 = n10124 ^ n10123 ^ 1'b0 ;
  assign n10126 = n177 & n5304 ;
  assign n10127 = n10126 ^ n4784 ^ 1'b0 ;
  assign n10128 = n10127 ^ n6707 ^ 1'b0 ;
  assign n10129 = n5982 & n10128 ;
  assign n10130 = ~n10125 & n10129 ;
  assign n10131 = n4099 ^ n1804 ^ 1'b0 ;
  assign n10132 = n1231 & n10131 ;
  assign n10133 = ~n962 & n10132 ;
  assign n10134 = n927 & ~n10133 ;
  assign n10135 = n10134 ^ n7698 ^ 1'b0 ;
  assign n10136 = n13 & ~n598 ;
  assign n10137 = n5268 ^ n2261 ^ 1'b0 ;
  assign n10138 = n1322 | n10137 ;
  assign n10139 = ( n7009 & n10136 ) | ( n7009 & n10138 ) | ( n10136 & n10138 ) ;
  assign n10140 = n10139 ^ n6544 ^ 1'b0 ;
  assign n10141 = n4977 ^ n1610 ^ 1'b0 ;
  assign n10142 = n1744 & n10141 ;
  assign n10143 = ~n911 & n10142 ;
  assign n10144 = n7813 ^ n3415 ^ 1'b0 ;
  assign n10145 = n3211 | n10144 ;
  assign n10146 = n7752 ^ n2867 ^ 1'b0 ;
  assign n10147 = ~n3772 & n10146 ;
  assign n10148 = n10147 ^ n6890 ^ 1'b0 ;
  assign n10149 = n7374 & n10148 ;
  assign n10150 = ~n10145 & n10149 ;
  assign n10151 = n10150 ^ n6520 ^ 1'b0 ;
  assign n10152 = n4635 | n6842 ;
  assign n10153 = n2840 & ~n10152 ;
  assign n10154 = n7435 ^ n5986 ^ 1'b0 ;
  assign n10156 = n3750 ^ n2146 ^ 1'b0 ;
  assign n10157 = ~n1250 & n10156 ;
  assign n10155 = ( n205 & n2888 ) | ( n205 & n4062 ) | ( n2888 & n4062 ) ;
  assign n10158 = n10157 ^ n10155 ^ 1'b0 ;
  assign n10159 = n8747 | n10158 ;
  assign n10160 = n10159 ^ n191 ^ 1'b0 ;
  assign n10161 = ~n6643 & n10160 ;
  assign n10162 = n3877 ^ n2447 ^ 1'b0 ;
  assign n10163 = n2918 & ~n10162 ;
  assign n10164 = n10163 ^ n1875 ^ n1603 ;
  assign n10165 = n7418 ^ n2939 ^ n2811 ;
  assign n10166 = ~n875 & n3801 ;
  assign n10167 = ~n10165 & n10166 ;
  assign n10168 = n10164 | n10167 ;
  assign n10169 = n10168 ^ n7141 ^ 1'b0 ;
  assign n10170 = n1371 & ~n5022 ;
  assign n10171 = ~n3131 & n10170 ;
  assign n10172 = n4992 & n10171 ;
  assign n10173 = n10172 ^ n7140 ^ 1'b0 ;
  assign n10175 = n353 & ~n3988 ;
  assign n10176 = n10175 ^ n3144 ^ 1'b0 ;
  assign n10174 = n3135 | n7033 ;
  assign n10177 = n10176 ^ n10174 ^ 1'b0 ;
  assign n10178 = n1572 | n7898 ;
  assign n10179 = n1713 & n4310 ;
  assign n10180 = ~n1642 & n10179 ;
  assign n10181 = n10180 ^ n1482 ^ n886 ;
  assign n10182 = n10127 ^ n7060 ^ 1'b0 ;
  assign n10183 = n10181 | n10182 ;
  assign n10184 = ~n3192 & n7405 ;
  assign n10185 = n3926 & n10184 ;
  assign n10186 = n2056 & n10185 ;
  assign n10187 = n172 | n221 ;
  assign n10188 = n9433 & n9901 ;
  assign n10189 = ~n10187 & n10188 ;
  assign n10190 = ~n4097 & n10189 ;
  assign n10191 = n5988 ^ n3027 ^ 1'b0 ;
  assign n10192 = n4540 | n10191 ;
  assign n10193 = n3835 & ~n10192 ;
  assign n10194 = n1636 & n10193 ;
  assign n10195 = n1407 | n10194 ;
  assign n10196 = n8633 | n8929 ;
  assign n10197 = n2060 ^ n875 ^ 1'b0 ;
  assign n10198 = n448 ^ n40 ^ 1'b0 ;
  assign n10199 = n1381 | n10198 ;
  assign n10200 = ( n306 & ~n5036 ) | ( n306 & n5155 ) | ( ~n5036 & n5155 ) ;
  assign n10201 = n10200 ^ n688 ^ 1'b0 ;
  assign n10202 = ~n9973 & n10201 ;
  assign n10203 = ~n10199 & n10202 ;
  assign n10204 = n10197 & n10203 ;
  assign n10207 = n3575 | n5050 ;
  assign n10205 = n153 & n1312 ;
  assign n10206 = n10205 ^ n6139 ^ 1'b0 ;
  assign n10208 = n10207 ^ n10206 ^ 1'b0 ;
  assign n10209 = n7004 | n10208 ;
  assign n10210 = n7267 ^ n5442 ^ n811 ;
  assign n10211 = n5471 ^ n4212 ^ 1'b0 ;
  assign n10212 = ( n6149 & n8885 ) | ( n6149 & ~n10211 ) | ( n8885 & ~n10211 ) ;
  assign n10213 = ~n1709 & n4580 ;
  assign n10214 = n246 & ~n5414 ;
  assign n10215 = n710 & n10214 ;
  assign n10216 = n8604 | n10215 ;
  assign n10217 = n2180 | n10216 ;
  assign n10218 = n4990 ^ n729 ^ 1'b0 ;
  assign n10219 = n8289 ^ n3408 ^ 1'b0 ;
  assign n10220 = n4422 & n10219 ;
  assign n10221 = n10220 ^ n6601 ^ n6181 ;
  assign n10222 = n10136 ^ n3402 ^ 1'b0 ;
  assign n10223 = n6067 ^ n2416 ^ 1'b0 ;
  assign n10224 = n10223 ^ n6614 ^ 1'b0 ;
  assign n10225 = n1078 & ~n10224 ;
  assign n10226 = n10222 & n10225 ;
  assign n10227 = ( ~n864 & n2565 ) | ( ~n864 & n6917 ) | ( n2565 & n6917 ) ;
  assign n10228 = n10227 ^ n110 ^ 1'b0 ;
  assign n10229 = n3000 & n4025 ;
  assign n10230 = ( n319 & ~n2935 ) | ( n319 & n10229 ) | ( ~n2935 & n10229 ) ;
  assign n10231 = n3145 & ~n9804 ;
  assign n10232 = n2940 ^ n1728 ^ 1'b0 ;
  assign n10233 = ( n5361 & n5517 ) | ( n5361 & n9952 ) | ( n5517 & n9952 ) ;
  assign n10234 = n3825 ^ n940 ^ 1'b0 ;
  assign n10235 = ( n2387 & ~n3635 ) | ( n2387 & n10234 ) | ( ~n3635 & n10234 ) ;
  assign n10236 = n1247 | n10235 ;
  assign n10237 = n4185 & n6736 ;
  assign n10238 = ~n4356 & n10237 ;
  assign n10240 = n139 | n7402 ;
  assign n10239 = ~n962 & n1213 ;
  assign n10241 = n10240 ^ n10239 ^ n5738 ;
  assign n10242 = n10241 ^ n7633 ^ 1'b0 ;
  assign n10243 = ~n4765 & n10242 ;
  assign n10244 = ~n2754 & n10243 ;
  assign n10245 = n2885 & n4626 ;
  assign n10246 = n6044 ^ n4696 ^ 1'b0 ;
  assign n10247 = n4954 & n10246 ;
  assign n10248 = n8851 ^ n795 ^ 1'b0 ;
  assign n10249 = n3909 & n10248 ;
  assign n10250 = n614 & ~n771 ;
  assign n10251 = n7568 ^ n6188 ^ 1'b0 ;
  assign n10252 = ~n10250 & n10251 ;
  assign n10253 = n63 & ~n4971 ;
  assign n10254 = ( n8154 & n9457 ) | ( n8154 & ~n10253 ) | ( n9457 & ~n10253 ) ;
  assign n10255 = n7815 ^ n2100 ^ 1'b0 ;
  assign n10256 = n10255 ^ n9469 ^ n3603 ;
  assign n10257 = ~n16 & n10086 ;
  assign n10258 = ~n5144 & n10257 ;
  assign n10259 = n1472 & ~n9444 ;
  assign n10260 = n10259 ^ n8177 ^ 1'b0 ;
  assign n10261 = n10260 ^ n3874 ^ 1'b0 ;
  assign n10262 = n1625 ^ n396 ^ 1'b0 ;
  assign n10263 = ~n1982 & n10262 ;
  assign n10264 = ( n654 & n2025 ) | ( n654 & ~n10263 ) | ( n2025 & ~n10263 ) ;
  assign n10265 = n10264 ^ n9437 ^ n285 ;
  assign n10266 = n3528 | n10265 ;
  assign n10267 = n1032 ^ n809 ^ 1'b0 ;
  assign n10268 = n10267 ^ n8751 ^ 1'b0 ;
  assign n10269 = n8094 & n10268 ;
  assign n10270 = ( n293 & ~n3571 ) | ( n293 & n5072 ) | ( ~n3571 & n5072 ) ;
  assign n10271 = ( n3904 & ~n6024 ) | ( n3904 & n7522 ) | ( ~n6024 & n7522 ) ;
  assign n10272 = n3615 | n10271 ;
  assign n10273 = n8903 ^ n7812 ^ n2839 ;
  assign n10274 = ( n245 & ~n6234 ) | ( n245 & n6784 ) | ( ~n6234 & n6784 ) ;
  assign n10275 = ~n3482 & n4763 ;
  assign n10276 = ~n3784 & n10275 ;
  assign n10277 = n4663 ^ n4045 ^ n1871 ;
  assign n10278 = n10277 ^ n4588 ^ 1'b0 ;
  assign n10279 = n194 & n10278 ;
  assign n10280 = n6140 ^ n2732 ^ n46 ;
  assign n10281 = n1261 & ~n2776 ;
  assign n10282 = n10281 ^ n4440 ^ 1'b0 ;
  assign n10288 = n2940 | n8046 ;
  assign n10283 = n6064 & ~n6351 ;
  assign n10284 = n10283 ^ n4368 ^ 1'b0 ;
  assign n10285 = n1907 & n8047 ;
  assign n10286 = n10284 & n10285 ;
  assign n10287 = n10286 ^ n2986 ^ 1'b0 ;
  assign n10289 = n10288 ^ n10287 ^ 1'b0 ;
  assign n10290 = n10282 | n10289 ;
  assign n10291 = ( n4067 & ~n4403 ) | ( n4067 & n6210 ) | ( ~n4403 & n6210 ) ;
  assign n10292 = ( ~n10280 & n10290 ) | ( ~n10280 & n10291 ) | ( n10290 & n10291 ) ;
  assign n10293 = n1650 & ~n8425 ;
  assign n10294 = n10293 ^ n8168 ^ 1'b0 ;
  assign n10295 = ~n213 & n254 ;
  assign n10296 = n3501 | n10295 ;
  assign n10297 = n10296 ^ n6466 ^ n5568 ;
  assign n10298 = n44 & n5916 ;
  assign n10299 = n10298 ^ n408 ^ 1'b0 ;
  assign n10300 = n9669 ^ n2058 ^ 1'b0 ;
  assign n10301 = ~n10299 & n10300 ;
  assign n10302 = n814 & ~n1467 ;
  assign n10303 = n1924 & n10302 ;
  assign n10304 = n10303 ^ n3114 ^ n1937 ;
  assign n10305 = n10304 ^ n1094 ^ 1'b0 ;
  assign n10306 = n3306 & ~n9084 ;
  assign n10307 = n9994 & n10306 ;
  assign n10308 = n10307 ^ n4896 ^ 1'b0 ;
  assign n10309 = n661 & ~n4114 ;
  assign n10310 = n452 & n7169 ;
  assign n10311 = n10309 & n10310 ;
  assign n10312 = n7307 & n7868 ;
  assign n10313 = n9595 ^ n2421 ^ 1'b0 ;
  assign n10316 = n4818 ^ n2907 ^ n32 ;
  assign n10314 = n1309 ^ n953 ^ 1'b0 ;
  assign n10315 = ~n9821 & n10314 ;
  assign n10317 = n10316 ^ n10315 ^ 1'b0 ;
  assign n10318 = n10313 | n10317 ;
  assign n10319 = ( n1189 & n3189 ) | ( n1189 & ~n7600 ) | ( n3189 & ~n7600 ) ;
  assign n10320 = n1213 & ~n7657 ;
  assign n10321 = n10319 | n10320 ;
  assign n10322 = n4779 & n10321 ;
  assign n10323 = n3874 ^ n2510 ^ 1'b0 ;
  assign n10324 = n1201 | n10323 ;
  assign n10325 = n10324 ^ n2294 ^ 1'b0 ;
  assign n10326 = n5700 ^ n2544 ^ n376 ;
  assign n10327 = ~n4450 & n10326 ;
  assign n10328 = n4077 & n10327 ;
  assign n10329 = n8472 & ~n10328 ;
  assign n10330 = n3780 ^ n205 ^ 1'b0 ;
  assign n10331 = n4078 ^ n85 ^ 1'b0 ;
  assign n10332 = n2374 ^ n1419 ^ 1'b0 ;
  assign n10333 = n8408 & n10332 ;
  assign n10334 = n10333 ^ n1897 ^ 1'b0 ;
  assign n10335 = ~n10331 & n10334 ;
  assign n10336 = n6261 ^ n6050 ^ 1'b0 ;
  assign n10337 = n7956 | n10336 ;
  assign n10338 = n46 & ~n10296 ;
  assign n10339 = ~n1531 & n10338 ;
  assign n10340 = n6893 | n10339 ;
  assign n10341 = n7872 ^ n2207 ^ 1'b0 ;
  assign n10342 = n7872 & n10341 ;
  assign n10343 = n4534 ^ n1545 ^ 1'b0 ;
  assign n10344 = n5481 ^ n4016 ^ n1728 ;
  assign n10345 = ~n1517 & n5229 ;
  assign n10346 = n8539 ^ n2617 ^ 1'b0 ;
  assign n10347 = n4356 ^ n3650 ^ n811 ;
  assign n10348 = n1343 ^ n1334 ^ n1041 ;
  assign n10349 = n2770 & n10348 ;
  assign n10350 = ~n4579 & n10349 ;
  assign n10351 = n10350 ^ n518 ^ 1'b0 ;
  assign n10352 = n1436 & ~n10351 ;
  assign n10359 = n1155 & ~n8168 ;
  assign n10360 = n10017 & n10359 ;
  assign n10356 = ~n3563 & n5227 ;
  assign n10357 = ( n4452 & n5961 ) | ( n4452 & ~n10356 ) | ( n5961 & ~n10356 ) ;
  assign n10353 = n3486 ^ n697 ^ 1'b0 ;
  assign n10354 = n6034 | n10353 ;
  assign n10355 = n1213 & ~n10354 ;
  assign n10358 = n10357 ^ n10355 ^ 1'b0 ;
  assign n10361 = n10360 ^ n10358 ^ 1'b0 ;
  assign n10362 = ~n1118 & n2705 ;
  assign n10363 = ~n499 & n10362 ;
  assign n10364 = ~n3354 & n10363 ;
  assign n10365 = n4319 ^ n2775 ^ 1'b0 ;
  assign n10366 = n1061 & n10365 ;
  assign n10367 = n6157 & n10366 ;
  assign n10368 = n10364 & n10367 ;
  assign n10369 = ~n234 & n6759 ;
  assign n10370 = n3560 & n10369 ;
  assign n10371 = n9653 & n10370 ;
  assign n10372 = n6353 ^ n2113 ^ 1'b0 ;
  assign n10373 = ~n769 & n8354 ;
  assign n10374 = n1777 & ~n7698 ;
  assign n10375 = n10374 ^ n5258 ^ n3739 ;
  assign n10376 = n6646 ^ n142 ^ 1'b0 ;
  assign n10377 = n10376 ^ n5335 ^ n846 ;
  assign n10378 = ( n5758 & n7196 ) | ( n5758 & n10377 ) | ( n7196 & n10377 ) ;
  assign n10379 = n108 & n523 ;
  assign n10380 = n10379 ^ n3365 ^ n1023 ;
  assign n10381 = n10380 ^ n1877 ^ 1'b0 ;
  assign n10382 = n32 & ~n2177 ;
  assign n10383 = ~n6947 & n10382 ;
  assign n10384 = n478 & n3019 ;
  assign n10385 = n2662 & n4215 ;
  assign n10386 = n5376 & n10385 ;
  assign n10387 = n5038 | n10386 ;
  assign n10388 = n3183 & n5888 ;
  assign n10389 = n44 & ~n2889 ;
  assign n10390 = n10389 ^ n10200 ^ 1'b0 ;
  assign n10391 = n10390 ^ n5955 ^ 1'b0 ;
  assign n10392 = n10388 & ~n10391 ;
  assign n10393 = n1647 & ~n2128 ;
  assign n10394 = n782 & ~n5554 ;
  assign n10395 = ~n1810 & n4968 ;
  assign n10396 = n4683 | n8895 ;
  assign n10397 = ( n1201 & n6105 ) | ( n1201 & n7638 ) | ( n6105 & n7638 ) ;
  assign n10398 = n10397 ^ n1484 ^ 1'b0 ;
  assign n10399 = ( n1666 & ~n5794 ) | ( n1666 & n6641 ) | ( ~n5794 & n6641 ) ;
  assign n10400 = n10271 | n10399 ;
  assign n10402 = n1410 & ~n5255 ;
  assign n10401 = n853 & n2887 ;
  assign n10403 = n10402 ^ n10401 ^ 1'b0 ;
  assign n10404 = n739 | n10403 ;
  assign n10405 = n8890 ^ n4536 ^ n3281 ;
  assign n10406 = n10405 ^ n4320 ^ 1'b0 ;
  assign n10410 = n2804 & n5033 ;
  assign n10411 = ~n3456 & n10410 ;
  assign n10412 = n10411 ^ n6571 ^ n2801 ;
  assign n10413 = n1526 & ~n5501 ;
  assign n10414 = n184 & n10413 ;
  assign n10415 = ( n5591 & ~n10412 ) | ( n5591 & n10414 ) | ( ~n10412 & n10414 ) ;
  assign n10407 = n5110 ^ n4605 ^ n3244 ;
  assign n10408 = n10407 ^ n3362 ^ 1'b0 ;
  assign n10409 = n4648 | n10408 ;
  assign n10416 = n10415 ^ n10409 ^ 1'b0 ;
  assign n10417 = n741 & n7508 ;
  assign n10418 = n2454 & n7303 ;
  assign n10419 = n3659 & n5108 ;
  assign n10420 = n10419 ^ n9027 ^ 1'b0 ;
  assign n10421 = n10420 ^ n6276 ^ n2168 ;
  assign n10422 = n2213 ^ n2051 ^ 1'b0 ;
  assign n10423 = n6005 & ~n10422 ;
  assign n10426 = n2490 ^ n2421 ^ 1'b0 ;
  assign n10424 = ~n322 & n5070 ;
  assign n10425 = n4880 | n10424 ;
  assign n10427 = n10426 ^ n10425 ^ n4427 ;
  assign n10428 = n5061 ^ n1787 ^ 1'b0 ;
  assign n10429 = n1650 & n10428 ;
  assign n10430 = n3661 & n10429 ;
  assign n10431 = n8024 | n10430 ;
  assign n10432 = n10427 | n10431 ;
  assign n10433 = ( n1412 & n2206 ) | ( n1412 & n4325 ) | ( n2206 & n4325 ) ;
  assign n10434 = ~n7282 & n10229 ;
  assign n10435 = n10434 ^ n3082 ^ 1'b0 ;
  assign n10436 = n7649 ^ n4951 ^ n1463 ;
  assign n10437 = n6101 | n9361 ;
  assign n10438 = n185 & ~n10437 ;
  assign n10439 = n10436 | n10438 ;
  assign n10440 = n10439 ^ n5578 ^ 1'b0 ;
  assign n10442 = n968 & ~n4325 ;
  assign n10441 = ( n126 & n1238 ) | ( n126 & ~n4574 ) | ( n1238 & ~n4574 ) ;
  assign n10443 = n10442 ^ n10441 ^ 1'b0 ;
  assign n10444 = ( ~n1035 & n2687 ) | ( ~n1035 & n2807 ) | ( n2687 & n2807 ) ;
  assign n10445 = n3964 & n9615 ;
  assign n10446 = n10444 & ~n10445 ;
  assign n10447 = n5626 | n6144 ;
  assign n10448 = n10447 ^ n1416 ^ 1'b0 ;
  assign n10449 = n10118 ^ n166 ^ 1'b0 ;
  assign n10450 = n10449 ^ n6632 ^ 1'b0 ;
  assign n10451 = n953 & n3844 ;
  assign n10452 = n3542 | n10451 ;
  assign n10453 = n4702 & n10452 ;
  assign n10454 = n10453 ^ n2569 ^ 1'b0 ;
  assign n10455 = n299 & n9021 ;
  assign n10456 = n10454 & n10455 ;
  assign n10457 = n1345 & ~n10456 ;
  assign n10458 = ~n383 & n2177 ;
  assign n10459 = n10458 ^ n3698 ^ 1'b0 ;
  assign n10460 = ~n4412 & n10459 ;
  assign n10461 = n7672 & n10460 ;
  assign n10462 = n5406 ^ n2863 ^ 1'b0 ;
  assign n10463 = n5673 ^ n3390 ^ 1'b0 ;
  assign n10464 = ~n10462 & n10463 ;
  assign n10465 = n9295 ^ n3166 ^ 1'b0 ;
  assign n10466 = n3634 ^ n1686 ^ 1'b0 ;
  assign n10467 = ~n2869 & n10466 ;
  assign n10468 = ( ~n9018 & n10465 ) | ( ~n9018 & n10467 ) | ( n10465 & n10467 ) ;
  assign n10469 = n10468 ^ n209 ^ 1'b0 ;
  assign n10470 = n10469 ^ n2902 ^ n2718 ;
  assign n10471 = n250 & n10470 ;
  assign n10472 = n9930 & n10471 ;
  assign n10473 = n2379 & ~n7927 ;
  assign n10476 = n299 & n7348 ;
  assign n10477 = n10476 ^ n3998 ^ 1'b0 ;
  assign n10474 = n30 | n5373 ;
  assign n10475 = n850 | n10474 ;
  assign n10478 = n10477 ^ n10475 ^ 1'b0 ;
  assign n10479 = n2262 ^ n1679 ^ 1'b0 ;
  assign n10480 = ( n3897 & ~n4064 ) | ( n3897 & n10479 ) | ( ~n4064 & n10479 ) ;
  assign n10481 = n8398 ^ n4914 ^ 1'b0 ;
  assign n10482 = n1241 & ~n10481 ;
  assign n10483 = ~n826 & n4837 ;
  assign n10484 = ( n2106 & ~n7514 ) | ( n2106 & n10483 ) | ( ~n7514 & n10483 ) ;
  assign n10485 = ~n395 & n4345 ;
  assign n10486 = n141 & n10485 ;
  assign n10487 = n125 & n10486 ;
  assign n10488 = n1145 & ~n6022 ;
  assign n10489 = n7164 ^ n4102 ^ 1'b0 ;
  assign n10490 = n10488 & ~n10489 ;
  assign n10491 = n7069 ^ n5182 ^ n2999 ;
  assign n10492 = n624 & ~n6813 ;
  assign n10493 = n6380 ^ n3679 ^ n139 ;
  assign n10494 = n1794 | n10493 ;
  assign n10495 = n5725 | n10494 ;
  assign n10496 = n10495 ^ n8241 ^ 1'b0 ;
  assign n10497 = n3709 | n4263 ;
  assign n10498 = n10497 ^ n6924 ^ 1'b0 ;
  assign n10499 = ( n4044 & n4147 ) | ( n4044 & n4285 ) | ( n4147 & n4285 ) ;
  assign n10500 = ~n1980 & n3620 ;
  assign n10501 = n5361 & n9000 ;
  assign n10502 = n961 | n6339 ;
  assign n10503 = n10502 ^ n1279 ^ 1'b0 ;
  assign n10507 = n1684 & n1700 ;
  assign n10508 = ~n7106 & n10507 ;
  assign n10509 = n2783 & n10508 ;
  assign n10510 = n10509 ^ n1290 ^ 1'b0 ;
  assign n10511 = n431 & n10510 ;
  assign n10504 = n2330 | n5219 ;
  assign n10505 = n10504 ^ n1484 ^ 1'b0 ;
  assign n10506 = n935 & ~n10505 ;
  assign n10512 = n10511 ^ n10506 ^ n188 ;
  assign n10513 = n2051 ^ n1079 ^ 1'b0 ;
  assign n10514 = n10512 | n10513 ;
  assign n10516 = n4475 ^ n1277 ^ n1058 ;
  assign n10515 = ~n434 & n6874 ;
  assign n10517 = n10516 ^ n10515 ^ 1'b0 ;
  assign n10518 = n10517 ^ n668 ^ 1'b0 ;
  assign n10519 = n3578 | n10518 ;
  assign n10520 = n23 | n6585 ;
  assign n10521 = ( n879 & n10519 ) | ( n879 & ~n10520 ) | ( n10519 & ~n10520 ) ;
  assign n10522 = ~n3107 & n4171 ;
  assign n10523 = ~n3792 & n10522 ;
  assign n10525 = n6245 ^ n3938 ^ 1'b0 ;
  assign n10526 = n3858 & ~n10525 ;
  assign n10524 = n7618 ^ n7500 ^ n4959 ;
  assign n10527 = n10526 ^ n10524 ^ 1'b0 ;
  assign n10528 = n169 & n10527 ;
  assign n10529 = n1824 ^ n1295 ^ 1'b0 ;
  assign n10530 = ~n496 & n10529 ;
  assign n10531 = n10530 ^ n6450 ^ 1'b0 ;
  assign n10532 = n10531 ^ n3566 ^ 1'b0 ;
  assign n10533 = n3077 ^ n1415 ^ 1'b0 ;
  assign n10534 = ~n4311 & n10533 ;
  assign n10535 = n7462 ^ n1225 ^ 1'b0 ;
  assign n10536 = n5879 & n10535 ;
  assign n10537 = ~n10534 & n10536 ;
  assign n10538 = n10391 | n10537 ;
  assign n10539 = n8154 & ~n10538 ;
  assign n10549 = n3650 | n5078 ;
  assign n10540 = n6995 ^ n6470 ^ n3080 ;
  assign n10541 = n5724 & n10540 ;
  assign n10542 = n8595 & ~n10541 ;
  assign n10543 = n10542 ^ n261 ^ 1'b0 ;
  assign n10544 = ~n156 & n10543 ;
  assign n10545 = ~n867 & n1793 ;
  assign n10546 = n2372 & n10545 ;
  assign n10547 = n10544 & ~n10546 ;
  assign n10548 = n8223 & n10547 ;
  assign n10550 = n10549 ^ n10548 ^ 1'b0 ;
  assign n10551 = ( n2864 & ~n3537 ) | ( n2864 & n5724 ) | ( ~n3537 & n5724 ) ;
  assign n10552 = n5673 ^ n1558 ^ 1'b0 ;
  assign n10553 = n3379 & ~n10552 ;
  assign n10554 = ~n2192 & n8766 ;
  assign n10555 = n10554 ^ n44 ^ 1'b0 ;
  assign n10556 = ( ~n10551 & n10553 ) | ( ~n10551 & n10555 ) | ( n10553 & n10555 ) ;
  assign n10557 = ( n3694 & n7428 ) | ( n3694 & ~n10556 ) | ( n7428 & ~n10556 ) ;
  assign n10558 = ~n3914 & n10301 ;
  assign n10559 = ~n8676 & n10558 ;
  assign n10560 = n126 & ~n1391 ;
  assign n10561 = n10390 ^ n1400 ^ 1'b0 ;
  assign n10562 = ~n10560 & n10561 ;
  assign n10563 = n6353 ^ n3040 ^ 1'b0 ;
  assign n10564 = n1773 | n3832 ;
  assign n10565 = ( n7699 & ~n10563 ) | ( n7699 & n10564 ) | ( ~n10563 & n10564 ) ;
  assign n10566 = n4083 & n7965 ;
  assign n10567 = n769 & n10566 ;
  assign n10568 = n5854 & n8707 ;
  assign n10569 = n1189 ^ n624 ^ 1'b0 ;
  assign n10570 = n3929 ^ n598 ^ 1'b0 ;
  assign n10571 = n10569 & n10570 ;
  assign n10572 = n10571 ^ n9732 ^ n3741 ;
  assign n10573 = n4508 ^ n1250 ^ 1'b0 ;
  assign n10574 = n7045 | n10573 ;
  assign n10575 = n299 & ~n2058 ;
  assign n10576 = n10574 & ~n10575 ;
  assign n10577 = n10576 ^ n1736 ^ 1'b0 ;
  assign n10578 = n4830 ^ n2954 ^ 1'b0 ;
  assign n10579 = n3774 | n8325 ;
  assign n10580 = n10579 ^ n2180 ^ 1'b0 ;
  assign n10581 = n10578 & n10580 ;
  assign n10582 = n6430 & n10581 ;
  assign n10583 = n1260 & ~n6868 ;
  assign n10584 = n1480 ^ n169 ^ 1'b0 ;
  assign n10585 = ~n10583 & n10584 ;
  assign n10586 = n10018 ^ n4024 ^ 1'b0 ;
  assign n10587 = n5088 ^ n3214 ^ 1'b0 ;
  assign n10588 = n4432 & ~n10587 ;
  assign n10589 = n8281 ^ n8135 ^ 1'b0 ;
  assign n10590 = n8383 & n10589 ;
  assign n10591 = n10590 ^ n3802 ^ 1'b0 ;
  assign n10592 = n6142 ^ n3912 ^ n3585 ;
  assign n10593 = n1561 | n3951 ;
  assign n10594 = n9914 ^ n4994 ^ n2556 ;
  assign n10595 = n863 & n4204 ;
  assign n10596 = n6514 & n10595 ;
  assign n10597 = n10054 ^ n2483 ^ n102 ;
  assign n10598 = n10597 ^ n9388 ^ n1279 ;
  assign n10599 = n10598 ^ n7653 ^ 1'b0 ;
  assign n10600 = n236 & n8807 ;
  assign n10601 = n8031 ^ n7996 ^ n5312 ;
  assign n10602 = n57 & ~n117 ;
  assign n10603 = n117 & n10602 ;
  assign n10604 = n168 & ~n10603 ;
  assign n10605 = ~n168 & n10604 ;
  assign n10606 = x10 & ~n10605 ;
  assign n10607 = ~x10 & n10606 ;
  assign n10608 = n1094 & n10607 ;
  assign n10609 = n1309 & ~n1395 ;
  assign n10610 = n10608 & n10609 ;
  assign n10611 = n868 | n1148 ;
  assign n10612 = n868 & ~n10611 ;
  assign n10613 = n401 | n10612 ;
  assign n10614 = n10610 & ~n10613 ;
  assign n10615 = n2422 | n3214 ;
  assign n10616 = n3214 & ~n10615 ;
  assign n10617 = ~n260 & n2305 ;
  assign n10618 = ~n10616 & n10617 ;
  assign n10619 = n10614 & n10618 ;
  assign n10620 = n10619 ^ n9864 ^ 1'b0 ;
  assign n10621 = n10601 & n10620 ;
  assign n10622 = n5697 | n6844 ;
  assign n10623 = n10622 ^ n8251 ^ 1'b0 ;
  assign n10624 = n7182 ^ n5261 ^ n830 ;
  assign n10625 = n2382 ^ n465 ^ 1'b0 ;
  assign n10626 = n10625 ^ n755 ^ 1'b0 ;
  assign n10627 = n10626 ^ n3570 ^ 1'b0 ;
  assign n10628 = ~n2885 & n10627 ;
  assign n10629 = ~n744 & n10628 ;
  assign n10630 = ~n8463 & n10629 ;
  assign n10631 = n1138 | n4399 ;
  assign n10632 = n312 & n3581 ;
  assign n10633 = n10632 ^ n3879 ^ n3692 ;
  assign n10634 = n5570 ^ n4757 ^ 1'b0 ;
  assign n10635 = n10633 | n10634 ;
  assign n10637 = ~n63 & n2168 ;
  assign n10638 = n10637 ^ n1459 ^ 1'b0 ;
  assign n10636 = n4036 | n10393 ;
  assign n10639 = n10638 ^ n10636 ^ 1'b0 ;
  assign n10640 = n7617 ^ n4350 ^ 1'b0 ;
  assign n10641 = ~n6965 & n10640 ;
  assign n10642 = n10641 ^ n493 ^ 1'b0 ;
  assign n10643 = ~n10639 & n10642 ;
  assign n10644 = ( n2111 & n2586 ) | ( n2111 & ~n3814 ) | ( n2586 & ~n3814 ) ;
  assign n10645 = n759 | n10598 ;
  assign n10646 = n10644 | n10645 ;
  assign n10647 = n609 & n1079 ;
  assign n10648 = ( n7878 & ~n8348 ) | ( n7878 & n10647 ) | ( ~n8348 & n10647 ) ;
  assign n10649 = ( ~n829 & n3342 ) | ( ~n829 & n10456 ) | ( n3342 & n10456 ) ;
  assign n10650 = ( n2635 & n10161 ) | ( n2635 & n10649 ) | ( n10161 & n10649 ) ;
  assign n10651 = ~n191 & n9700 ;
  assign n10652 = n10651 ^ n1455 ^ 1'b0 ;
  assign n10653 = n5011 & ~n10652 ;
  assign n10654 = n8929 & n10653 ;
  assign n10655 = n1350 ^ n467 ^ 1'b0 ;
  assign n10656 = n201 & n10655 ;
  assign n10657 = n5684 ^ n972 ^ 1'b0 ;
  assign n10658 = n10656 & n10657 ;
  assign n10659 = ( n1090 & n4888 ) | ( n1090 & n5172 ) | ( n4888 & n5172 ) ;
  assign n10660 = n10659 ^ n550 ^ 1'b0 ;
  assign n10661 = n3533 & ~n4247 ;
  assign n10662 = n10660 & n10661 ;
  assign n10663 = n7371 ^ n5802 ^ 1'b0 ;
  assign n10664 = ~n10662 & n10663 ;
  assign n10665 = n7269 ^ n2214 ^ 1'b0 ;
  assign n10666 = n761 & ~n1652 ;
  assign n10667 = n10666 ^ n6156 ^ 1'b0 ;
  assign n10668 = n9950 ^ n74 ^ 1'b0 ;
  assign n10669 = n2911 | n6855 ;
  assign n10670 = n10669 ^ n5066 ^ 1'b0 ;
  assign n10672 = ~n1979 & n10430 ;
  assign n10671 = n84 | n4028 ;
  assign n10673 = n10672 ^ n10671 ^ 1'b0 ;
  assign n10674 = n1182 ^ n582 ^ 1'b0 ;
  assign n10675 = n10674 ^ n3931 ^ 1'b0 ;
  assign n10676 = ~n4531 & n10029 ;
  assign n10677 = n10676 ^ n5047 ^ n4000 ;
  assign n10680 = n2644 ^ n2177 ^ 1'b0 ;
  assign n10681 = n2644 & n10680 ;
  assign n10682 = n10681 ^ n5845 ^ 1'b0 ;
  assign n10678 = n1280 ^ n773 ^ 1'b0 ;
  assign n10679 = n2861 | n10678 ;
  assign n10683 = n10682 ^ n10679 ^ 1'b0 ;
  assign n10684 = ~n8591 & n10683 ;
  assign n10685 = n7666 ^ n1650 ^ 1'b0 ;
  assign n10686 = n6987 ^ n2076 ^ n1865 ;
  assign n10687 = n10686 ^ n2671 ^ 1'b0 ;
  assign n10688 = n7721 | n10687 ;
  assign n10694 = n1407 & n1848 ;
  assign n10695 = ~n2573 & n10694 ;
  assign n10696 = n10695 ^ n162 ^ 1'b0 ;
  assign n10697 = n1303 & n10696 ;
  assign n10698 = ~n4515 & n10697 ;
  assign n10699 = n10698 ^ n511 ^ 1'b0 ;
  assign n10690 = ~n4662 & n4796 ;
  assign n10691 = n4703 ^ n2433 ^ 1'b0 ;
  assign n10692 = ~n10690 & n10691 ;
  assign n10693 = n8500 & n10692 ;
  assign n10700 = n10699 ^ n10693 ^ 1'b0 ;
  assign n10701 = n10700 ^ n3593 ^ 1'b0 ;
  assign n10702 = n7293 & n10701 ;
  assign n10703 = n10702 ^ n8537 ^ 1'b0 ;
  assign n10704 = ~n1665 & n8823 ;
  assign n10705 = n10704 ^ n5891 ^ 1'b0 ;
  assign n10706 = ~n6796 & n10705 ;
  assign n10707 = n10703 & n10706 ;
  assign n10689 = n759 & n1234 ;
  assign n10708 = n10707 ^ n10689 ^ x3 ;
  assign n10709 = n532 & n1695 ;
  assign n10710 = n4667 ^ n1283 ^ 1'b0 ;
  assign n10711 = ~n10709 & n10710 ;
  assign n10712 = n10711 ^ n10485 ^ 1'b0 ;
  assign n10715 = n3062 | n8542 ;
  assign n10713 = ~n1485 & n4966 ;
  assign n10714 = n10713 ^ n2028 ^ 1'b0 ;
  assign n10716 = n10715 ^ n10714 ^ n2986 ;
  assign n10717 = n6695 & n10716 ;
  assign n10718 = n4144 & n6085 ;
  assign n10719 = n1575 & n10718 ;
  assign n10720 = n496 | n10719 ;
  assign n10721 = n6972 ^ n100 ^ 1'b0 ;
  assign n10722 = n10721 ^ n5696 ^ n1650 ;
  assign n10723 = n8789 ^ n2972 ^ 1'b0 ;
  assign n10724 = ~n6363 & n10723 ;
  assign n10725 = ~n2942 & n3187 ;
  assign n10726 = n2623 & ~n10725 ;
  assign n10727 = ( n168 & n3027 ) | ( n168 & ~n3170 ) | ( n3027 & ~n3170 ) ;
  assign n10728 = ~n1633 & n10727 ;
  assign n10729 = n668 & n10728 ;
  assign n10730 = n10729 ^ n5482 ^ 1'b0 ;
  assign n10731 = n3680 & ~n10730 ;
  assign n10732 = n10731 ^ n6899 ^ 1'b0 ;
  assign n10733 = ~n6304 & n10732 ;
  assign n10734 = n7026 ^ n2906 ^ 1'b0 ;
  assign n10736 = n2549 ^ n1457 ^ 1'b0 ;
  assign n10737 = n304 & ~n10736 ;
  assign n10735 = n3256 & ~n3698 ;
  assign n10738 = n10737 ^ n10735 ^ 1'b0 ;
  assign n10739 = n1001 | n10738 ;
  assign n10740 = n4399 & n10739 ;
  assign n10741 = ~n10734 & n10740 ;
  assign n10742 = n1201 | n10741 ;
  assign n10743 = n10742 ^ n5848 ^ 1'b0 ;
  assign n10744 = n3305 ^ n729 ^ 1'b0 ;
  assign n10745 = n5134 | n10744 ;
  assign n10746 = n10743 & ~n10745 ;
  assign n10747 = n10746 ^ n3329 ^ 1'b0 ;
  assign n10748 = n2612 | n3263 ;
  assign n10749 = ~n6097 & n6704 ;
  assign n10750 = n220 & n5707 ;
  assign n10751 = n9816 & n10750 ;
  assign n10752 = n4000 ^ n3938 ^ n1120 ;
  assign n10753 = ( n395 & ~n1409 ) | ( n395 & n10752 ) | ( ~n1409 & n10752 ) ;
  assign n10754 = n8355 ^ n2241 ^ 1'b0 ;
  assign n10755 = n4986 ^ n2787 ^ 1'b0 ;
  assign n10756 = n10755 ^ n530 ^ 1'b0 ;
  assign n10758 = n4686 ^ n2974 ^ 1'b0 ;
  assign n10759 = n628 | n5732 ;
  assign n10760 = n10758 & ~n10759 ;
  assign n10761 = n9244 | n10760 ;
  assign n10757 = ~n3691 & n6222 ;
  assign n10762 = n10761 ^ n10757 ^ 1'b0 ;
  assign n10763 = n2494 | n10762 ;
  assign n10764 = n2485 & ~n10763 ;
  assign n10765 = n2816 | n8421 ;
  assign n10766 = n187 | n3526 ;
  assign n10767 = n10766 ^ n3318 ^ 1'b0 ;
  assign n10768 = n946 | n10767 ;
  assign n10769 = n10768 ^ n7844 ^ n7213 ;
  assign n10770 = n631 | n888 ;
  assign n10771 = n3246 & ~n10770 ;
  assign n10772 = n10771 ^ n5351 ^ n3606 ;
  assign n10773 = n3260 & n4693 ;
  assign n10774 = n10234 ^ n5942 ^ n1185 ;
  assign n10775 = n10774 ^ n5078 ^ 1'b0 ;
  assign n10776 = n312 & n5520 ;
  assign n10777 = n10776 ^ n1167 ^ 1'b0 ;
  assign n10778 = n10777 ^ n6931 ^ 1'b0 ;
  assign n10779 = ~n6332 & n10778 ;
  assign n10780 = n7082 | n10779 ;
  assign n10781 = ( ~n7645 & n10223 ) | ( ~n7645 & n10780 ) | ( n10223 & n10780 ) ;
  assign n10782 = n452 & ~n645 ;
  assign n10783 = n10782 ^ n4135 ^ 1'b0 ;
  assign n10784 = ( n1289 & n2345 ) | ( n1289 & n3170 ) | ( n2345 & n3170 ) ;
  assign n10785 = n5488 ^ n99 ^ 1'b0 ;
  assign n10786 = n7236 & ~n10785 ;
  assign n10787 = n10784 & n10786 ;
  assign n10788 = n10787 ^ n2954 ^ 1'b0 ;
  assign n10789 = n46 & ~n10788 ;
  assign n10790 = n10789 ^ n2621 ^ 1'b0 ;
  assign n10791 = n6470 | n10790 ;
  assign n10792 = n9879 & ~n10450 ;
  assign n10793 = ( ~n1546 & n1640 ) | ( ~n1546 & n6692 ) | ( n1640 & n6692 ) ;
  assign n10794 = n10793 ^ n4082 ^ n267 ;
  assign n10795 = n10794 ^ n1583 ^ 1'b0 ;
  assign n10796 = ~n38 & n3784 ;
  assign n10797 = n10796 ^ n1436 ^ 1'b0 ;
  assign n10798 = n2870 | n3473 ;
  assign n10799 = ( n4455 & ~n5748 ) | ( n4455 & n10798 ) | ( ~n5748 & n10798 ) ;
  assign n10800 = ( n1993 & n6277 ) | ( n1993 & ~n8490 ) | ( n6277 & ~n8490 ) ;
  assign n10801 = n10799 & n10800 ;
  assign n10802 = n10801 ^ n4114 ^ 1'b0 ;
  assign n10803 = n8030 & ~n9562 ;
  assign n10804 = ( n6030 & n7977 ) | ( n6030 & ~n9839 ) | ( n7977 & ~n9839 ) ;
  assign n10805 = n10804 ^ n177 ^ 1'b0 ;
  assign n10806 = n2836 & ~n10805 ;
  assign n10807 = ~n1461 & n10806 ;
  assign n10808 = n115 & n3304 ;
  assign n10809 = ~n23 & n10808 ;
  assign n10810 = n6451 ^ n1300 ^ 1'b0 ;
  assign n10811 = ( n2922 & n8899 ) | ( n2922 & ~n10810 ) | ( n8899 & ~n10810 ) ;
  assign n10812 = ( n51 & n201 ) | ( n51 & n1006 ) | ( n201 & n1006 ) ;
  assign n10813 = n10812 ^ n3802 ^ 1'b0 ;
  assign n10814 = n10813 ^ n372 ^ 1'b0 ;
  assign n10815 = n10814 ^ n7450 ^ 1'b0 ;
  assign n10816 = n1826 & ~n5800 ;
  assign n10817 = n10816 ^ n5091 ^ n375 ;
  assign n10818 = n5195 ^ n532 ^ 1'b0 ;
  assign n10819 = n2039 & n10818 ;
  assign n10820 = n2999 & n3765 ;
  assign n10821 = n5425 & ~n10820 ;
  assign n10822 = n1387 | n10821 ;
  assign n10823 = n5450 | n8277 ;
  assign n10824 = n10823 ^ n5585 ^ 1'b0 ;
  assign n10825 = n2036 ^ n1307 ^ n500 ;
  assign n10826 = n10825 ^ n2831 ^ 1'b0 ;
  assign n10827 = ~n5037 & n10826 ;
  assign n10831 = ~n1511 & n6154 ;
  assign n10832 = n10831 ^ n496 ^ 1'b0 ;
  assign n10828 = n57 & ~n6774 ;
  assign n10829 = n10828 ^ n5189 ^ 1'b0 ;
  assign n10830 = n10738 | n10829 ;
  assign n10833 = n10832 ^ n10830 ^ 1'b0 ;
  assign n10834 = n8566 ^ n883 ^ 1'b0 ;
  assign n10835 = n7516 & n10834 ;
  assign n10836 = n1312 & ~n10835 ;
  assign n10840 = ~n2640 & n10786 ;
  assign n10841 = n10840 ^ n1640 ^ 1'b0 ;
  assign n10839 = n447 & ~n3185 ;
  assign n10837 = n1031 | n10197 ;
  assign n10838 = n5657 & ~n10837 ;
  assign n10842 = n10841 ^ n10839 ^ n10838 ;
  assign n10843 = n2573 | n3608 ;
  assign n10844 = n4048 | n10843 ;
  assign n10845 = n1072 ^ n1045 ^ 1'b0 ;
  assign n10846 = n10845 ^ n5137 ^ 1'b0 ;
  assign n10847 = n10846 ^ n5851 ^ 1'b0 ;
  assign n10848 = n10844 & n10847 ;
  assign n10849 = n4093 & n7409 ;
  assign n10850 = n3548 ^ n2871 ^ 1'b0 ;
  assign n10851 = n1727 & ~n6620 ;
  assign n10852 = ( n4345 & n10850 ) | ( n4345 & n10851 ) | ( n10850 & n10851 ) ;
  assign n10853 = n961 | n10852 ;
  assign n10854 = n10853 ^ n6220 ^ 1'b0 ;
  assign n10855 = n779 & ~n10854 ;
  assign n10856 = n4796 & n10855 ;
  assign n10857 = ( ~n436 & n10849 ) | ( ~n436 & n10856 ) | ( n10849 & n10856 ) ;
  assign n10858 = n2873 ^ n2678 ^ 1'b0 ;
  assign n10859 = ~n9832 & n10858 ;
  assign n10860 = n8149 & ~n9255 ;
  assign n10861 = ~n7469 & n10860 ;
  assign n10862 = n3737 & ~n4445 ;
  assign n10863 = ~n5554 & n10862 ;
  assign n10864 = n1482 ^ n882 ^ 1'b0 ;
  assign n10865 = n430 & ~n10864 ;
  assign n10866 = n4129 | n8714 ;
  assign n10867 = n10865 | n10866 ;
  assign n10868 = n4428 & ~n10719 ;
  assign n10869 = n10868 ^ n10012 ^ 1'b0 ;
  assign n10870 = n10867 & ~n10869 ;
  assign n10871 = n5470 ^ n2258 ^ 1'b0 ;
  assign n10872 = ~n5040 & n10871 ;
  assign n10873 = ~n1196 & n7715 ;
  assign n10876 = n3238 & n6821 ;
  assign n10874 = n6309 | n7701 ;
  assign n10875 = n10874 ^ n9416 ^ n5219 ;
  assign n10877 = n10876 ^ n10875 ^ 1'b0 ;
  assign n10878 = n5223 & n10877 ;
  assign n10884 = ( ~n235 & n2471 ) | ( ~n235 & n7443 ) | ( n2471 & n7443 ) ;
  assign n10885 = n4186 & n10884 ;
  assign n10879 = n6259 | n10008 ;
  assign n10880 = n7759 ^ n4665 ^ 1'b0 ;
  assign n10881 = ~n694 & n10880 ;
  assign n10882 = n10879 & n10881 ;
  assign n10883 = n10882 ^ n6695 ^ 1'b0 ;
  assign n10886 = n10885 ^ n10883 ^ n4652 ;
  assign n10892 = n2917 ^ n2428 ^ 1'b0 ;
  assign n10887 = ~n1841 & n2982 ;
  assign n10888 = n3741 | n10887 ;
  assign n10889 = n10888 ^ n7535 ^ 1'b0 ;
  assign n10890 = n8254 & ~n10889 ;
  assign n10891 = ~n255 & n10890 ;
  assign n10893 = n10892 ^ n10891 ^ 1'b0 ;
  assign n10894 = n10893 ^ n1742 ^ 1'b0 ;
  assign n10895 = n647 & ~n7927 ;
  assign n10896 = ~n3409 & n5039 ;
  assign n10897 = ~n10895 & n10896 ;
  assign n10898 = n7228 ^ n301 ^ 1'b0 ;
  assign n10899 = n1003 & ~n2088 ;
  assign n10900 = n7815 ^ n7004 ^ 1'b0 ;
  assign n10901 = n10180 ^ n176 ^ 1'b0 ;
  assign n10902 = ~n3198 & n10901 ;
  assign n10903 = n2088 | n8048 ;
  assign n10904 = ~n9011 & n10903 ;
  assign n10905 = n5488 & n10904 ;
  assign n10906 = n852 | n10905 ;
  assign n10907 = n10906 ^ n749 ^ 1'b0 ;
  assign n10908 = n1407 & ~n5313 ;
  assign n10909 = n10908 ^ n1940 ^ 1'b0 ;
  assign n10910 = ( n46 & n3138 ) | ( n46 & n7019 ) | ( n3138 & n7019 ) ;
  assign n10911 = ~n1206 & n6607 ;
  assign n10912 = n10910 & ~n10911 ;
  assign n10913 = ~n10909 & n10912 ;
  assign n10914 = n3648 ^ n3175 ^ 1'b0 ;
  assign n10915 = ~n3528 & n10914 ;
  assign n10916 = n283 & ~n7888 ;
  assign n10917 = ~n8110 & n10916 ;
  assign n10918 = n6449 & ~n10917 ;
  assign n10919 = ~n10915 & n10918 ;
  assign n10920 = n10919 ^ n1622 ^ n994 ;
  assign n10921 = ~n809 & n1597 ;
  assign n10922 = n10921 ^ n644 ^ 1'b0 ;
  assign n10923 = n135 & ~n10922 ;
  assign n10924 = ~n477 & n10923 ;
  assign n10925 = n469 & ~n6866 ;
  assign n10926 = ~n1886 & n10925 ;
  assign n10927 = n3539 & n5438 ;
  assign n10928 = n10926 & n10927 ;
  assign n10929 = n4221 ^ n1927 ^ 1'b0 ;
  assign n10930 = n6150 | n10929 ;
  assign n10931 = n9792 ^ n8019 ^ 1'b0 ;
  assign n10932 = ~n6424 & n10931 ;
  assign n10933 = n10932 ^ n9436 ^ 1'b0 ;
  assign n10934 = ~n3051 & n8516 ;
  assign n10935 = n2745 & n5006 ;
  assign n10936 = ~n1226 & n8683 ;
  assign n10937 = n3398 & n4536 ;
  assign n10938 = n10936 & n10937 ;
  assign n10939 = ( n3676 & ~n8262 ) | ( n3676 & n9273 ) | ( ~n8262 & n9273 ) ;
  assign n10940 = ( ~n1960 & n3027 ) | ( ~n1960 & n10939 ) | ( n3027 & n10939 ) ;
  assign n10941 = ( n1243 & n7287 ) | ( n1243 & n10919 ) | ( n7287 & n10919 ) ;
  assign n10942 = n3630 ^ n1263 ^ 1'b0 ;
  assign n10943 = ( n577 & n2276 ) | ( n577 & ~n7183 ) | ( n2276 & ~n7183 ) ;
  assign n10944 = ~n2840 & n10943 ;
  assign n10945 = ~n2089 & n10944 ;
  assign n10946 = ( n7094 & n10942 ) | ( n7094 & ~n10945 ) | ( n10942 & ~n10945 ) ;
  assign n10947 = n6071 ^ n2106 ^ 1'b0 ;
  assign n10948 = n10946 | n10947 ;
  assign n10949 = n23 | n3817 ;
  assign n10950 = n1030 & ~n10949 ;
  assign n10951 = n8721 ^ n5228 ^ 1'b0 ;
  assign n10952 = n10951 ^ n3137 ^ n1728 ;
  assign n10953 = n8106 & ~n10952 ;
  assign n10954 = n10953 ^ n98 ^ 1'b0 ;
  assign n10955 = n5384 | n10954 ;
  assign n10956 = n8470 | n10955 ;
  assign n10957 = n10950 | n10956 ;
  assign n10958 = n1770 ^ n1642 ^ 1'b0 ;
  assign n10959 = n993 & ~n5816 ;
  assign n10960 = n4719 | n9378 ;
  assign n10961 = n5202 & n10960 ;
  assign n10962 = ~n3620 & n10961 ;
  assign n10963 = n10962 ^ n7600 ^ 1'b0 ;
  assign n10964 = n8447 ^ n4890 ^ 1'b0 ;
  assign n10965 = ~n3170 & n10964 ;
  assign n10966 = n6150 & n10965 ;
  assign n10967 = n5331 ^ n4914 ^ 1'b0 ;
  assign n10968 = n9470 ^ n6927 ^ n3563 ;
  assign n10969 = n10968 ^ n10598 ^ n6844 ;
  assign n10970 = ~n694 & n5572 ;
  assign n10971 = n10970 ^ n2745 ^ 1'b0 ;
  assign n10972 = n6168 | n10949 ;
  assign n10973 = n10972 ^ n104 ^ 1'b0 ;
  assign n10974 = n8015 ^ n441 ^ 1'b0 ;
  assign n10975 = ~n4397 & n4542 ;
  assign n10976 = n7988 | n10420 ;
  assign n10977 = n5931 ^ n2460 ^ 1'b0 ;
  assign n10978 = n6144 | n10808 ;
  assign n10979 = n5521 ^ n4023 ^ 1'b0 ;
  assign n10980 = n5314 | n10979 ;
  assign n10981 = ~n3647 & n10980 ;
  assign n10982 = n8994 ^ n6078 ^ 1'b0 ;
  assign n10983 = n1265 | n4533 ;
  assign n10984 = n10983 ^ n10451 ^ 1'b0 ;
  assign n10985 = n891 & n10984 ;
  assign n10986 = n10985 ^ n8636 ^ 1'b0 ;
  assign n10987 = n4142 & ~n4366 ;
  assign n10988 = n2859 | n4586 ;
  assign n10989 = n5676 | n10988 ;
  assign n10990 = ( n3456 & n7867 ) | ( n3456 & ~n10989 ) | ( n7867 & ~n10989 ) ;
  assign n10993 = n6302 & ~n8105 ;
  assign n10991 = n2216 & n2368 ;
  assign n10992 = n5879 | n10991 ;
  assign n10994 = n10993 ^ n10992 ^ 1'b0 ;
  assign n10995 = n676 & ~n10994 ;
  assign n10996 = n2108 | n10007 ;
  assign n10997 = n10996 ^ n9956 ^ 1'b0 ;
  assign n11001 = n1047 | n2128 ;
  assign n11002 = n6142 | n11001 ;
  assign n10998 = n57 & ~n4058 ;
  assign n10999 = ( ~n5377 & n7272 ) | ( ~n5377 & n10998 ) | ( n7272 & n10998 ) ;
  assign n11000 = ~n4863 & n10999 ;
  assign n11003 = n11002 ^ n11000 ^ n26 ;
  assign n11004 = ~n740 & n2710 ;
  assign n11005 = n7494 | n10396 ;
  assign n11006 = n11005 ^ n5128 ^ 1'b0 ;
  assign n11007 = ~n2196 & n9426 ;
  assign n11008 = n4327 ^ n4233 ^ 1'b0 ;
  assign n11009 = n1023 & ~n11008 ;
  assign n11015 = n10709 ^ n7276 ^ n4330 ;
  assign n11010 = n2696 ^ n1287 ^ 1'b0 ;
  assign n11011 = n11010 ^ n3330 ^ 1'b0 ;
  assign n11012 = n604 | n11011 ;
  assign n11013 = n4240 & ~n11012 ;
  assign n11014 = n11013 ^ n9722 ^ n1723 ;
  assign n11016 = n11015 ^ n11014 ^ 1'b0 ;
  assign n11017 = ~n6071 & n11016 ;
  assign n11018 = ( n11007 & n11009 ) | ( n11007 & ~n11017 ) | ( n11009 & ~n11017 ) ;
  assign n11021 = ( ~n177 & n183 ) | ( ~n177 & n530 ) | ( n183 & n530 ) ;
  assign n11019 = n2414 & n3759 ;
  assign n11020 = n3773 & ~n11019 ;
  assign n11022 = n11021 ^ n11020 ^ 1'b0 ;
  assign n11023 = n2449 | n3607 ;
  assign n11024 = n4383 ^ n563 ^ 1'b0 ;
  assign n11025 = n5661 & n11024 ;
  assign n11026 = ~n6554 & n11025 ;
  assign n11027 = n11023 & n11026 ;
  assign n11028 = n11027 ^ n1520 ^ 1'b0 ;
  assign n11029 = n7226 ^ n4608 ^ 1'b0 ;
  assign n11030 = n1869 ^ n806 ^ 1'b0 ;
  assign n11031 = ~n10884 & n11030 ;
  assign n11032 = n11031 ^ n7306 ^ 1'b0 ;
  assign n11033 = n6616 | n11032 ;
  assign n11036 = n4536 ^ n4105 ^ 1'b0 ;
  assign n11034 = n3923 & n8889 ;
  assign n11035 = n11034 ^ n7090 ^ 1'b0 ;
  assign n11037 = n11036 ^ n11035 ^ 1'b0 ;
  assign n11038 = n3207 | n9519 ;
  assign n11039 = n4469 & n7641 ;
  assign n11040 = ~n1577 & n11039 ;
  assign n11041 = ( n1255 & n4809 ) | ( n1255 & ~n11040 ) | ( n4809 & ~n11040 ) ;
  assign n11042 = n9576 ^ n3358 ^ n2397 ;
  assign n11043 = n301 & n6357 ;
  assign n11044 = n11043 ^ n7123 ^ 1'b0 ;
  assign n11045 = ( n10931 & ~n11042 ) | ( n10931 & n11044 ) | ( ~n11042 & n11044 ) ;
  assign n11046 = n2581 & ~n2797 ;
  assign n11047 = n289 & ~n8542 ;
  assign n11048 = ~n11046 & n11047 ;
  assign n11049 = ~n1198 & n1281 ;
  assign n11050 = n3811 & n11049 ;
  assign n11051 = n2985 ^ n1944 ^ 1'b0 ;
  assign n11052 = n971 | n11051 ;
  assign n11053 = n1849 ^ n1590 ^ 1'b0 ;
  assign n11054 = ~n4678 & n6059 ;
  assign n11055 = ~n11053 & n11054 ;
  assign n11056 = n842 & n11055 ;
  assign n11057 = n11056 ^ n2577 ^ 1'b0 ;
  assign n11068 = n54 | n263 ;
  assign n11069 = n11068 ^ n4815 ^ 1'b0 ;
  assign n11070 = n59 & ~n11069 ;
  assign n11058 = n6759 ^ n4424 ^ 1'b0 ;
  assign n11059 = ~n1149 & n4458 ;
  assign n11060 = n11059 ^ n2935 ^ n36 ;
  assign n11061 = ~n8006 & n11060 ;
  assign n11062 = n11058 & n11061 ;
  assign n11063 = n11062 ^ n5596 ^ 1'b0 ;
  assign n11064 = n6205 ^ n1302 ^ 1'b0 ;
  assign n11065 = n2606 & n8258 ;
  assign n11066 = n11064 & n11065 ;
  assign n11067 = n11063 & ~n11066 ;
  assign n11071 = n11070 ^ n11067 ^ 1'b0 ;
  assign n11072 = ~n3081 & n10088 ;
  assign n11073 = ( ~n4890 & n8472 ) | ( ~n4890 & n11072 ) | ( n8472 & n11072 ) ;
  assign n11074 = n10753 ^ n5324 ^ 1'b0 ;
  assign n11075 = n9103 ^ n4247 ^ 1'b0 ;
  assign n11076 = n962 & ~n11075 ;
  assign n11077 = n7325 ^ n6076 ^ n3113 ;
  assign n11078 = ( ~n4237 & n4704 ) | ( ~n4237 & n11077 ) | ( n4704 & n11077 ) ;
  assign n11081 = n7713 ^ n5640 ^ 1'b0 ;
  assign n11079 = ( n1022 & n4012 ) | ( n1022 & n10046 ) | ( n4012 & n10046 ) ;
  assign n11080 = n5114 & ~n11079 ;
  assign n11082 = n11081 ^ n11080 ^ 1'b0 ;
  assign n11083 = ( ~n5229 & n7706 ) | ( ~n5229 & n10002 ) | ( n7706 & n10002 ) ;
  assign n11084 = n11083 ^ n607 ^ 1'b0 ;
  assign n11085 = n11082 & n11084 ;
  assign n11086 = ~n5893 & n11085 ;
  assign n11090 = ( n1010 & ~n5511 ) | ( n1010 & n7025 ) | ( ~n5511 & n7025 ) ;
  assign n11087 = n2132 & ~n3449 ;
  assign n11088 = n11087 ^ n9459 ^ 1'b0 ;
  assign n11089 = n303 | n11088 ;
  assign n11091 = n11090 ^ n11089 ^ 1'b0 ;
  assign n11092 = n1822 & n11002 ;
  assign n11093 = n8659 & n11092 ;
  assign n11094 = ( n59 & n1606 ) | ( n59 & n11093 ) | ( n1606 & n11093 ) ;
  assign n11095 = n666 & ~n4712 ;
  assign n11096 = n134 & ~n3848 ;
  assign n11097 = n11096 ^ n9558 ^ 1'b0 ;
  assign n11098 = ~n11095 & n11097 ;
  assign n11099 = n1495 & ~n5667 ;
  assign n11100 = ~n3842 & n11099 ;
  assign n11101 = n7318 | n11100 ;
  assign n11102 = n3575 | n9371 ;
  assign n11103 = n505 & ~n11102 ;
  assign n11104 = n11103 ^ n8442 ^ n3357 ;
  assign n11106 = ~n228 & n2188 ;
  assign n11107 = n11106 ^ n4632 ^ 1'b0 ;
  assign n11108 = n11107 ^ n5571 ^ 1'b0 ;
  assign n11109 = n11108 ^ n6343 ^ 1'b0 ;
  assign n11110 = n6174 ^ n4287 ^ 1'b0 ;
  assign n11111 = n7362 | n11110 ;
  assign n11112 = n4014 & ~n11111 ;
  assign n11113 = n11112 ^ n5118 ^ 1'b0 ;
  assign n11114 = n11109 & n11113 ;
  assign n11105 = ~n617 & n8043 ;
  assign n11115 = n11114 ^ n11105 ^ 1'b0 ;
  assign n11116 = n7655 ^ n352 ^ 1'b0 ;
  assign n11117 = n2481 ^ n477 ^ 1'b0 ;
  assign n11118 = ( ~n2154 & n2190 ) | ( ~n2154 & n11117 ) | ( n2190 & n11117 ) ;
  assign n11119 = n4877 | n5481 ;
  assign n11120 = ( ~n7754 & n8866 ) | ( ~n7754 & n10379 ) | ( n8866 & n10379 ) ;
  assign n11121 = n11120 ^ n4832 ^ 1'b0 ;
  assign n11122 = ~n1318 & n11121 ;
  assign n11123 = ~n6485 & n11122 ;
  assign n11124 = n10223 | n11123 ;
  assign n11125 = n2034 ^ n1643 ^ 1'b0 ;
  assign n11126 = ~n2601 & n11125 ;
  assign n11127 = n2728 & n11126 ;
  assign n11128 = n11127 ^ n2664 ^ 1'b0 ;
  assign n11129 = ( n6326 & n7055 ) | ( n6326 & n11128 ) | ( n7055 & n11128 ) ;
  assign n11130 = n2089 ^ n209 ^ 1'b0 ;
  assign n11131 = n1079 & ~n3105 ;
  assign n11132 = n11131 ^ n7836 ^ n7773 ;
  assign n11133 = n11132 ^ n9197 ^ 1'b0 ;
  assign n11134 = n11130 | n11133 ;
  assign n11135 = n1602 & ~n2304 ;
  assign n11136 = n624 & n11135 ;
  assign n11137 = n8978 ^ n3018 ^ 1'b0 ;
  assign n11138 = n4115 ^ n863 ^ 1'b0 ;
  assign n11139 = ~n1612 & n7763 ;
  assign n11140 = n11139 ^ n3775 ^ 1'b0 ;
  assign n11141 = n1170 ^ n446 ^ 1'b0 ;
  assign n11142 = n11140 | n11141 ;
  assign n11143 = ( ~n2422 & n4769 ) | ( ~n2422 & n11142 ) | ( n4769 & n11142 ) ;
  assign n11144 = ~n11138 & n11143 ;
  assign n11145 = ( n2135 & ~n11137 ) | ( n2135 & n11144 ) | ( ~n11137 & n11144 ) ;
  assign n11146 = n10978 ^ n10850 ^ 1'b0 ;
  assign n11147 = ~n8754 & n11146 ;
  assign n11152 = n5062 ^ n734 ^ 1'b0 ;
  assign n11148 = n121 & n2173 ;
  assign n11149 = n11148 ^ n1368 ^ 1'b0 ;
  assign n11150 = n11149 ^ n10393 ^ n6919 ;
  assign n11151 = n1063 & ~n11150 ;
  assign n11153 = n11152 ^ n11151 ^ 1'b0 ;
  assign n11154 = ( n799 & n9066 ) | ( n799 & n9208 ) | ( n9066 & n9208 ) ;
  assign n11155 = n1170 & n4846 ;
  assign n11156 = n11155 ^ n3970 ^ 1'b0 ;
  assign n11157 = ~n11154 & n11156 ;
  assign n11158 = ~n6451 & n9528 ;
  assign n11159 = n11158 ^ n496 ^ 1'b0 ;
  assign n11160 = n4590 ^ n607 ^ 1'b0 ;
  assign n11161 = n4311 & n11160 ;
  assign n11162 = ( n467 & n1368 ) | ( n467 & ~n11161 ) | ( n1368 & ~n11161 ) ;
  assign n11163 = ~n5110 & n11162 ;
  assign n11164 = n1134 ^ n381 ^ 1'b0 ;
  assign n11165 = n2064 | n4366 ;
  assign n11166 = n11165 ^ n3009 ^ 1'b0 ;
  assign n11167 = n42 | n11166 ;
  assign n11168 = ~n11164 & n11167 ;
  assign n11169 = n1527 & n11168 ;
  assign n11170 = ( n1767 & n2538 ) | ( n1767 & n4002 ) | ( n2538 & n4002 ) ;
  assign n11171 = n10204 & n11170 ;
  assign n11172 = n777 & ~n5160 ;
  assign n11173 = n1728 & n5878 ;
  assign n11175 = n332 | n9535 ;
  assign n11176 = n8091 ^ n4961 ^ 1'b0 ;
  assign n11177 = ~n11175 & n11176 ;
  assign n11174 = n3364 | n9045 ;
  assign n11178 = n11177 ^ n11174 ^ 1'b0 ;
  assign n11179 = n4483 ^ n455 ^ 1'b0 ;
  assign n11180 = n5109 & n11179 ;
  assign n11181 = n6858 ^ n85 ^ 1'b0 ;
  assign n11182 = n698 | n11181 ;
  assign n11183 = n3660 & ~n11182 ;
  assign n11184 = n11183 ^ n6732 ^ 1'b0 ;
  assign n11185 = n10163 ^ n2584 ^ 1'b0 ;
  assign n11186 = ~n5370 & n11185 ;
  assign n11187 = n11186 ^ n1835 ^ 1'b0 ;
  assign n11188 = ~n2181 & n9849 ;
  assign n11189 = n9548 ^ n6129 ^ 1'b0 ;
  assign n11191 = n5583 | n7721 ;
  assign n11192 = n9245 | n11191 ;
  assign n11193 = n8047 ^ n940 ^ 1'b0 ;
  assign n11194 = n11192 & n11193 ;
  assign n11190 = ( ~n2373 & n3761 ) | ( ~n2373 & n5338 ) | ( n3761 & n5338 ) ;
  assign n11195 = n11194 ^ n11190 ^ 1'b0 ;
  assign n11196 = n2083 & ~n5323 ;
  assign n11197 = n11196 ^ n830 ^ 1'b0 ;
  assign n11198 = n5856 | n11197 ;
  assign n11199 = n11195 | n11198 ;
  assign n11200 = n63 | n2389 ;
  assign n11201 = n1326 & ~n11200 ;
  assign n11202 = n285 | n11201 ;
  assign n11203 = n324 & ~n1465 ;
  assign n11204 = n11203 ^ n1938 ^ 1'b0 ;
  assign n11205 = n11204 ^ n6951 ^ 1'b0 ;
  assign n11206 = n4706 | n11205 ;
  assign n11207 = n349 & ~n11206 ;
  assign n11208 = n4447 ^ n919 ^ 1'b0 ;
  assign n11209 = ~n11207 & n11208 ;
  assign n11210 = ~n607 & n11209 ;
  assign n11211 = n11202 & ~n11210 ;
  assign n11212 = n2456 & n4364 ;
  assign n11213 = n11212 ^ n3855 ^ 1'b0 ;
  assign n11214 = n1188 & n5171 ;
  assign n11215 = ~n11213 & n11214 ;
  assign n11216 = n11215 ^ n2633 ^ 1'b0 ;
  assign n11217 = n4844 & ~n6660 ;
  assign n11218 = ~n3264 & n11217 ;
  assign n11219 = n3241 ^ n2158 ^ 1'b0 ;
  assign n11220 = n11219 ^ n6833 ^ n1412 ;
  assign n11221 = n5107 ^ n3141 ^ 1'b0 ;
  assign n11222 = n2696 & ~n7659 ;
  assign n11223 = n4708 ^ n779 ^ 1'b0 ;
  assign n11224 = ~n4815 & n11223 ;
  assign n11225 = n11224 ^ n4211 ^ 1'b0 ;
  assign n11226 = ~n2617 & n11225 ;
  assign n11227 = n9330 ^ n1439 ^ n1426 ;
  assign n11228 = n11227 ^ n548 ^ 1'b0 ;
  assign n11229 = n3737 | n11228 ;
  assign n11230 = n6199 & ~n7126 ;
  assign n11231 = n9713 ^ n4674 ^ n1461 ;
  assign n11232 = n7058 ^ n3322 ^ 1'b0 ;
  assign n11233 = n4576 & n11232 ;
  assign n11234 = n411 & n10136 ;
  assign n11235 = ( n4355 & n6942 ) | ( n4355 & n11234 ) | ( n6942 & n11234 ) ;
  assign n11236 = ~n1934 & n8793 ;
  assign n11237 = n11236 ^ n2309 ^ 1'b0 ;
  assign n11238 = n5090 & ~n11237 ;
  assign n11239 = n8179 ^ n291 ^ 1'b0 ;
  assign n11247 = ( ~n3049 & n4480 ) | ( ~n3049 & n8113 ) | ( n4480 & n8113 ) ;
  assign n11248 = n740 | n5084 ;
  assign n11249 = n11247 & ~n11248 ;
  assign n11240 = n5011 & n5509 ;
  assign n11241 = n1003 & n11240 ;
  assign n11242 = n2271 & ~n2732 ;
  assign n11243 = n11242 ^ n2934 ^ 1'b0 ;
  assign n11244 = n1737 & n4962 ;
  assign n11245 = ( n1346 & n11243 ) | ( n1346 & ~n11244 ) | ( n11243 & ~n11244 ) ;
  assign n11246 = n11241 | n11245 ;
  assign n11250 = n11249 ^ n11246 ^ 1'b0 ;
  assign n11251 = n6204 ^ n2784 ^ 1'b0 ;
  assign n11252 = ~n1068 & n4637 ;
  assign n11253 = n2218 & n11252 ;
  assign n11254 = n11253 ^ n10263 ^ n1373 ;
  assign n11255 = ( n2431 & ~n6792 ) | ( n2431 & n10062 ) | ( ~n6792 & n10062 ) ;
  assign n11256 = ~n11254 & n11255 ;
  assign n11257 = n1492 ^ n131 ^ 1'b0 ;
  assign n11258 = n567 & n11257 ;
  assign n11259 = n11258 ^ n7929 ^ 1'b0 ;
  assign n11260 = ~n8267 & n11259 ;
  assign n11261 = n1832 & ~n2627 ;
  assign n11262 = n11261 ^ n4345 ^ 1'b0 ;
  assign n11263 = n2549 | n11262 ;
  assign n11264 = n256 | n11263 ;
  assign n11265 = ~n9420 & n11264 ;
  assign n11266 = n11265 ^ n586 ^ 1'b0 ;
  assign n11267 = n11260 & ~n11266 ;
  assign n11268 = n11267 ^ n4992 ^ 1'b0 ;
  assign n11269 = ~n2818 & n11268 ;
  assign n11271 = n4704 ^ n4091 ^ 1'b0 ;
  assign n11270 = n6616 & ~n6653 ;
  assign n11272 = n11271 ^ n11270 ^ 1'b0 ;
  assign n11273 = n6579 & ~n11272 ;
  assign n11274 = n10980 ^ n324 ^ 1'b0 ;
  assign n11275 = n7387 ^ n1262 ^ 1'b0 ;
  assign n11277 = ( n3385 & n4696 ) | ( n3385 & n4906 ) | ( n4696 & n4906 ) ;
  assign n11276 = n197 & n230 ;
  assign n11278 = n11277 ^ n11276 ^ 1'b0 ;
  assign n11279 = n4336 & ~n11278 ;
  assign n11281 = n7231 ^ n3024 ^ 1'b0 ;
  assign n11280 = ~n4588 & n6480 ;
  assign n11282 = n11281 ^ n11280 ^ 1'b0 ;
  assign n11285 = ( n2177 & n4477 ) | ( n2177 & n5661 ) | ( n4477 & n5661 ) ;
  assign n11283 = n3437 ^ n2278 ^ n1898 ;
  assign n11284 = ~n1502 & n11283 ;
  assign n11286 = n11285 ^ n11284 ^ 1'b0 ;
  assign n11287 = n1456 & ~n11286 ;
  assign n11288 = n11287 ^ n4573 ^ 1'b0 ;
  assign n11289 = n11288 ^ n747 ^ 1'b0 ;
  assign n11290 = n9073 | n11289 ;
  assign n11291 = n5891 ^ n1095 ^ 1'b0 ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11293 = n8145 & ~n9395 ;
  assign n11294 = n498 & n11293 ;
  assign n11295 = n3894 ^ n2568 ^ 1'b0 ;
  assign n11296 = n5068 ^ n3923 ^ 1'b0 ;
  assign n11298 = n1972 & n4932 ;
  assign n11299 = n5946 | n11298 ;
  assign n11300 = n11299 ^ n5352 ^ 1'b0 ;
  assign n11297 = n3223 & ~n5854 ;
  assign n11301 = n11300 ^ n11297 ^ 1'b0 ;
  assign n11302 = n2552 ^ n1546 ^ 1'b0 ;
  assign n11303 = n2337 | n11302 ;
  assign n11304 = n11303 ^ n6977 ^ 1'b0 ;
  assign n11305 = n3784 & n8515 ;
  assign n11306 = n5853 | n8635 ;
  assign n11307 = n9792 | n11306 ;
  assign n11308 = n315 | n890 ;
  assign n11309 = n11308 ^ n9206 ^ 1'b0 ;
  assign n11310 = n1336 & ~n11309 ;
  assign n11311 = ~n4439 & n11310 ;
  assign n11312 = n5526 ^ n5374 ^ 1'b0 ;
  assign n11313 = n1151 & n3049 ;
  assign n11314 = n11313 ^ n8153 ^ 1'b0 ;
  assign n11315 = n498 | n11314 ;
  assign n11316 = n7831 | n11315 ;
  assign n11317 = n11204 ^ n1830 ^ 1'b0 ;
  assign n11318 = ~n2650 & n11317 ;
  assign n11319 = n8325 ^ n1274 ^ 1'b0 ;
  assign n11320 = n11318 & n11319 ;
  assign n11322 = n9688 ^ n1340 ^ 1'b0 ;
  assign n11321 = n3619 & n7832 ;
  assign n11323 = n11322 ^ n11321 ^ 1'b0 ;
  assign n11324 = ~n4830 & n7975 ;
  assign n11325 = n11324 ^ n4304 ^ 1'b0 ;
  assign n11326 = n4008 | n4688 ;
  assign n11327 = n7153 & ~n11326 ;
  assign n11331 = ~n2989 & n10349 ;
  assign n11328 = n2381 | n5529 ;
  assign n11329 = n5957 | n11328 ;
  assign n11330 = n11329 ^ n2086 ^ 1'b0 ;
  assign n11332 = n11331 ^ n11330 ^ 1'b0 ;
  assign n11333 = n1376 | n11091 ;
  assign n11334 = ( ~n1186 & n3908 ) | ( ~n1186 & n4590 ) | ( n3908 & n4590 ) ;
  assign n11335 = n11334 ^ n6555 ^ n2740 ;
  assign n11336 = n8018 | n11335 ;
  assign n11337 = n11336 ^ n4114 ^ 1'b0 ;
  assign n11338 = n8083 ^ n1032 ^ 1'b0 ;
  assign n11339 = n4430 & ~n11338 ;
  assign n11340 = n11339 ^ n183 ^ 1'b0 ;
  assign n11341 = n5653 & n8362 ;
  assign n11343 = n4465 & ~n5985 ;
  assign n11344 = n6352 & n11343 ;
  assign n11342 = ~n1875 & n3878 ;
  assign n11345 = n11344 ^ n11342 ^ 1'b0 ;
  assign n11346 = n11341 & ~n11345 ;
  assign n11347 = ( n41 & ~n2500 ) | ( n41 & n5562 ) | ( ~n2500 & n5562 ) ;
  assign n11348 = n11347 ^ n3745 ^ 1'b0 ;
  assign n11349 = n1233 | n11348 ;
  assign n11350 = n11349 ^ n5656 ^ n3790 ;
  assign n11351 = n5793 ^ n1400 ^ 1'b0 ;
  assign n11352 = n11350 & n11351 ;
  assign n11353 = n10200 ^ n7078 ^ 1'b0 ;
  assign n11354 = n6265 ^ n5751 ^ 1'b0 ;
  assign n11355 = n209 & n11354 ;
  assign n11356 = n11344 ^ n5007 ^ 1'b0 ;
  assign n11357 = ( ~n2324 & n5090 ) | ( ~n2324 & n11356 ) | ( n5090 & n11356 ) ;
  assign n11358 = ~n7186 & n9549 ;
  assign n11359 = ~n2098 & n11358 ;
  assign n11360 = n11359 ^ n5651 ^ 1'b0 ;
  assign n11361 = n1538 | n4880 ;
  assign n11362 = n11361 ^ n463 ^ 1'b0 ;
  assign n11363 = n11360 & n11362 ;
  assign n11364 = n2620 & ~n8285 ;
  assign n11365 = n10079 & n11364 ;
  assign n11366 = n8735 & n11365 ;
  assign n11367 = ( n7547 & n11363 ) | ( n7547 & n11366 ) | ( n11363 & n11366 ) ;
  assign n11368 = n1209 & n2436 ;
  assign n11369 = n654 & n11368 ;
  assign n11370 = n11369 ^ n3633 ^ 1'b0 ;
  assign n11371 = ~n2768 & n11370 ;
  assign n11372 = n11371 ^ n9745 ^ 1'b0 ;
  assign n11373 = n11372 ^ n9615 ^ n9104 ;
  assign n11374 = n2313 & ~n2896 ;
  assign n11375 = n1209 & n11374 ;
  assign n11376 = n11375 ^ n6868 ^ 1'b0 ;
  assign n11377 = n156 | n11376 ;
  assign n11378 = n2991 | n11377 ;
  assign n11379 = n8049 & ~n11378 ;
  assign n11380 = n9128 ^ n6802 ^ 1'b0 ;
  assign n11381 = n2493 & n11380 ;
  assign n11382 = n6049 & ~n10269 ;
  assign n11383 = ( n717 & n5823 ) | ( n717 & ~n8099 ) | ( n5823 & ~n8099 ) ;
  assign n11384 = n962 & ~n11383 ;
  assign n11385 = n11384 ^ n4536 ^ 1'b0 ;
  assign n11386 = n2416 ^ n2254 ^ 1'b0 ;
  assign n11387 = n1520 | n5423 ;
  assign n11388 = n1807 & ~n11387 ;
  assign n11389 = n11388 ^ n4054 ^ 1'b0 ;
  assign n11390 = n11389 ^ n1063 ^ 1'b0 ;
  assign n11391 = ~n3285 & n11390 ;
  assign n11392 = n5099 ^ n2173 ^ 1'b0 ;
  assign n11393 = n1210 & ~n11392 ;
  assign n11394 = n178 & ~n2583 ;
  assign n11395 = ~n728 & n11394 ;
  assign n11396 = n11395 ^ n5113 ^ 1'b0 ;
  assign n11397 = n11393 & ~n11396 ;
  assign n11398 = n11397 ^ n8094 ^ 1'b0 ;
  assign n11399 = ( n2330 & n11391 ) | ( n2330 & ~n11398 ) | ( n11391 & ~n11398 ) ;
  assign n11400 = n3773 & n5315 ;
  assign n11401 = ~n1079 & n11400 ;
  assign n11402 = n11401 ^ n619 ^ n62 ;
  assign n11403 = n6693 & ~n6775 ;
  assign n11404 = ( n1499 & n2330 ) | ( n1499 & n4188 ) | ( n2330 & n4188 ) ;
  assign n11405 = n7463 ^ n1138 ^ 1'b0 ;
  assign n11406 = n11404 & n11405 ;
  assign n11407 = n4462 & ~n8257 ;
  assign n11408 = ~n8622 & n11407 ;
  assign n11409 = n2194 | n11408 ;
  assign n11410 = ~n2752 & n11409 ;
  assign n11411 = n2245 ^ n1444 ^ 1'b0 ;
  assign n11412 = n1718 | n11411 ;
  assign n11413 = n1875 & ~n11412 ;
  assign n11414 = n691 | n3700 ;
  assign n11415 = n7645 | n11414 ;
  assign n11416 = n2896 | n11415 ;
  assign n11417 = n5101 | n11416 ;
  assign n11418 = n8608 | n11417 ;
  assign n11419 = n5082 | n9965 ;
  assign n11420 = n9746 ^ n91 ^ 1'b0 ;
  assign n11421 = n10140 ^ n6278 ^ 1'b0 ;
  assign n11422 = n8693 & ~n11421 ;
  assign n11432 = n6572 ^ n5972 ^ 1'b0 ;
  assign n11429 = n1604 & n6908 ;
  assign n11427 = ( ~n3020 & n4135 ) | ( ~n3020 & n4227 ) | ( n4135 & n4227 ) ;
  assign n11428 = n2064 & n11427 ;
  assign n11423 = n63 | n3676 ;
  assign n11424 = n11423 ^ n1613 ^ 1'b0 ;
  assign n11425 = ~n3593 & n11424 ;
  assign n11426 = n11425 ^ n10500 ^ 1'b0 ;
  assign n11430 = n11429 ^ n11428 ^ n11426 ;
  assign n11431 = n8298 & n11430 ;
  assign n11433 = n11432 ^ n11431 ^ 1'b0 ;
  assign n11437 = n3807 ^ n1583 ^ 1'b0 ;
  assign n11434 = n7443 ^ n3234 ^ 1'b0 ;
  assign n11435 = n5094 & ~n11434 ;
  assign n11436 = n2492 & n11435 ;
  assign n11438 = n11437 ^ n11436 ^ 1'b0 ;
  assign n11439 = n4339 ^ n842 ^ 1'b0 ;
  assign n11440 = n11439 ^ n5234 ^ 1'b0 ;
  assign n11441 = n11440 ^ n991 ^ 1'b0 ;
  assign n11442 = ~n11438 & n11441 ;
  assign n11443 = n6636 ^ n4873 ^ 1'b0 ;
  assign n11444 = n648 ^ n63 ^ 1'b0 ;
  assign n11445 = n100 & n11444 ;
  assign n11446 = ~n4205 & n11445 ;
  assign n11449 = n8398 ^ n7325 ^ 1'b0 ;
  assign n11450 = ~n942 & n11449 ;
  assign n11451 = n2154 & n3299 ;
  assign n11452 = n6466 & n11451 ;
  assign n11453 = ~n11450 & n11452 ;
  assign n11448 = ~n473 & n4604 ;
  assign n11447 = n2218 & n10841 ;
  assign n11454 = n11453 ^ n11448 ^ n11447 ;
  assign n11455 = n11454 ^ n2943 ^ 1'b0 ;
  assign n11456 = n10900 & ~n11455 ;
  assign n11457 = n9127 ^ n2657 ^ 1'b0 ;
  assign n11458 = ~n2453 & n11457 ;
  assign n11459 = ~n2933 & n7308 ;
  assign n11460 = ( ~n2633 & n2801 ) | ( ~n2633 & n3227 ) | ( n2801 & n3227 ) ;
  assign n11461 = n2350 | n11460 ;
  assign n11462 = n11459 & ~n11461 ;
  assign n11465 = ( ~n427 & n2874 ) | ( ~n427 & n6213 ) | ( n2874 & n6213 ) ;
  assign n11463 = n1231 & ~n3232 ;
  assign n11464 = n11463 ^ n2282 ^ 1'b0 ;
  assign n11466 = n11465 ^ n11464 ^ x6 ;
  assign n11467 = n11466 ^ n7935 ^ 1'b0 ;
  assign n11468 = n4512 & ~n5044 ;
  assign n11469 = n11468 ^ n3301 ^ 1'b0 ;
  assign n11470 = ( ~n3183 & n7297 ) | ( ~n3183 & n9764 ) | ( n7297 & n9764 ) ;
  assign n11471 = n4147 & ~n4371 ;
  assign n11472 = n11471 ^ n1523 ^ 1'b0 ;
  assign n11473 = n11363 ^ n6713 ^ n4006 ;
  assign n11474 = n6191 | n11473 ;
  assign n11475 = n4518 & ~n11474 ;
  assign n11477 = n6000 & ~n8657 ;
  assign n11478 = n11477 ^ n386 ^ 1'b0 ;
  assign n11479 = ( n5535 & ~n7988 ) | ( n5535 & n11478 ) | ( ~n7988 & n11478 ) ;
  assign n11480 = n994 & n5280 ;
  assign n11481 = ~n8148 & n11480 ;
  assign n11482 = n11479 & n11481 ;
  assign n11476 = n7729 & n8055 ;
  assign n11483 = n11482 ^ n11476 ^ 1'b0 ;
  assign n11484 = n2195 ^ n816 ^ 1'b0 ;
  assign n11485 = ~n1232 & n11484 ;
  assign n11486 = n11485 ^ n8590 ^ 1'b0 ;
  assign n11487 = ( n2926 & n5534 ) | ( n2926 & ~n11486 ) | ( n5534 & ~n11486 ) ;
  assign n11488 = n11487 ^ n2992 ^ 1'b0 ;
  assign n11489 = n11055 ^ n10353 ^ 1'b0 ;
  assign n11490 = ~n11488 & n11489 ;
  assign n11491 = ~n6157 & n9104 ;
  assign n11492 = n4661 ^ n3254 ^ 1'b0 ;
  assign n11493 = n2939 & ~n11492 ;
  assign n11494 = ~n5841 & n11493 ;
  assign n11495 = n1641 & n11007 ;
  assign n11496 = n2736 & ~n11495 ;
  assign n11497 = n11496 ^ n11256 ^ 1'b0 ;
  assign n11498 = ( n982 & n6178 ) | ( n982 & ~n6789 ) | ( n6178 & ~n6789 ) ;
  assign n11499 = n366 & ~n3341 ;
  assign n11500 = ~n8052 & n11499 ;
  assign n11501 = n3560 & ~n8582 ;
  assign n11502 = n11500 & n11501 ;
  assign n11503 = n8730 ^ n7873 ^ n6590 ;
  assign n11504 = n985 & ~n6246 ;
  assign n11505 = ~n4056 & n11504 ;
  assign n11506 = n5368 & n10249 ;
  assign n11507 = n6535 & n11506 ;
  assign n11509 = ~n1521 & n3679 ;
  assign n11510 = n7652 & n11509 ;
  assign n11508 = ( ~n607 & n1249 ) | ( ~n607 & n6528 ) | ( n1249 & n6528 ) ;
  assign n11511 = n11510 ^ n11508 ^ 1'b0 ;
  assign n11512 = n1772 | n3686 ;
  assign n11513 = n3799 | n11512 ;
  assign n11514 = n10303 ^ n987 ^ 1'b0 ;
  assign n11516 = n9961 ^ n209 ^ 1'b0 ;
  assign n11515 = n1612 & ~n3255 ;
  assign n11517 = n11516 ^ n11515 ^ 1'b0 ;
  assign n11518 = n150 | n5116 ;
  assign n11519 = n8335 ^ n2561 ^ 1'b0 ;
  assign n11520 = n11518 | n11519 ;
  assign n11521 = n11520 ^ n5110 ^ 1'b0 ;
  assign n11522 = n1013 | n9404 ;
  assign n11523 = n1103 & ~n11522 ;
  assign n11524 = ( n5766 & n6802 ) | ( n5766 & n7935 ) | ( n6802 & n7935 ) ;
  assign n11525 = ~n3823 & n3950 ;
  assign n11526 = n11525 ^ n1505 ^ 1'b0 ;
  assign n11527 = n11526 ^ n135 ^ 1'b0 ;
  assign n11528 = ( ~n5543 & n11524 ) | ( ~n5543 & n11527 ) | ( n11524 & n11527 ) ;
  assign n11529 = n2547 ^ n2132 ^ 1'b0 ;
  assign n11530 = ~n1840 & n2925 ;
  assign n11531 = ~n22 & n11530 ;
  assign n11532 = n5722 ^ n5395 ^ n1889 ;
  assign n11533 = n1866 & ~n11532 ;
  assign n11534 = n11531 & n11533 ;
  assign n11535 = ( n1234 & n3581 ) | ( n1234 & n11534 ) | ( n3581 & n11534 ) ;
  assign n11536 = n9621 ^ n414 ^ n332 ;
  assign n11537 = n2049 & ~n10361 ;
  assign n11538 = n3824 & n11537 ;
  assign n11539 = n1982 | n10514 ;
  assign n11540 = n9798 | n11539 ;
  assign n11541 = n3749 & ~n9625 ;
  assign n11542 = n11541 ^ n4460 ^ 1'b0 ;
  assign n11543 = n6827 ^ n6275 ^ 1'b0 ;
  assign n11544 = ~n3363 & n5903 ;
  assign n11545 = n11544 ^ n7847 ^ n4195 ;
  assign n11546 = n11545 ^ n2588 ^ 1'b0 ;
  assign n11547 = n629 | n10108 ;
  assign n11548 = ~n1295 & n11547 ;
  assign n11549 = n11548 ^ n7818 ^ 1'b0 ;
  assign n11550 = n3486 & ~n11123 ;
  assign n11551 = ~n7013 & n11550 ;
  assign n11552 = n5649 ^ n1382 ^ n243 ;
  assign n11553 = n4728 & n11552 ;
  assign n11554 = n8061 & n11553 ;
  assign n11557 = n687 & ~n3043 ;
  assign n11558 = ~n5570 & n11557 ;
  assign n11555 = ~n799 & n5874 ;
  assign n11556 = ~n9130 & n11555 ;
  assign n11559 = n11558 ^ n11556 ^ 1'b0 ;
  assign n11560 = n6983 ^ n3949 ^ 1'b0 ;
  assign n11561 = ~n1542 & n6097 ;
  assign n11562 = ( n10791 & n11560 ) | ( n10791 & n11561 ) | ( n11560 & n11561 ) ;
  assign n11563 = n3560 ^ n156 ^ 1'b0 ;
  assign n11564 = ( n2432 & n7535 ) | ( n2432 & ~n11563 ) | ( n7535 & ~n11563 ) ;
  assign n11565 = n5524 ^ n934 ^ 1'b0 ;
  assign n11566 = n11565 ^ n9815 ^ 1'b0 ;
  assign n11567 = n3094 ^ n2182 ^ 1'b0 ;
  assign n11568 = n3100 | n9704 ;
  assign n11569 = n3577 | n10948 ;
  assign n11570 = n8486 ^ n2951 ^ n2544 ;
  assign n11571 = n9479 ^ n6790 ^ 1'b0 ;
  assign n11572 = n11570 & ~n11571 ;
  assign n11573 = n5986 ^ n448 ^ 1'b0 ;
  assign n11574 = n344 & n4376 ;
  assign n11581 = n11356 ^ n3412 ^ 1'b0 ;
  assign n11580 = n887 & ~n8193 ;
  assign n11582 = n11581 ^ n11580 ^ 1'b0 ;
  assign n11575 = ( n3656 & n3851 ) | ( n3656 & ~n6143 ) | ( n3851 & ~n6143 ) ;
  assign n11576 = n11376 | n11575 ;
  assign n11577 = n11576 ^ n77 ^ 1'b0 ;
  assign n11578 = n8651 ^ n5793 ^ 1'b0 ;
  assign n11579 = n11577 & n11578 ;
  assign n11583 = n11582 ^ n11579 ^ 1'b0 ;
  assign n11584 = n3769 ^ n1694 ^ 1'b0 ;
  assign n11585 = n944 & ~n11584 ;
  assign n11586 = n7670 ^ n3959 ^ 1'b0 ;
  assign n11587 = n3373 & n11586 ;
  assign n11588 = n11587 ^ n6352 ^ 1'b0 ;
  assign n11589 = n2926 | n11588 ;
  assign n11590 = n11585 & ~n11589 ;
  assign n11591 = n11590 ^ n6422 ^ 1'b0 ;
  assign n11592 = n4008 ^ n1368 ^ 1'b0 ;
  assign n11593 = n2966 | n11592 ;
  assign n11594 = n3371 | n6462 ;
  assign n11595 = n5891 ^ n2896 ^ 1'b0 ;
  assign n11596 = n1364 & n1712 ;
  assign n11597 = n11596 ^ n4670 ^ n2758 ;
  assign n11598 = n3104 | n5986 ;
  assign n11599 = n2983 | n11598 ;
  assign n11600 = n1654 | n2649 ;
  assign n11601 = n7271 & ~n11600 ;
  assign n11602 = n11601 ^ n5008 ^ 1'b0 ;
  assign n11603 = n8306 ^ n714 ^ 1'b0 ;
  assign n11604 = n4142 & ~n11603 ;
  assign n11605 = n11604 ^ n3584 ^ 1'b0 ;
  assign n11606 = n11605 ^ n2745 ^ n381 ;
  assign n11607 = n7903 & n9363 ;
  assign n11608 = n4817 & ~n5301 ;
  assign n11609 = n6322 & n11608 ;
  assign n11610 = n2384 ^ n1516 ^ n514 ;
  assign n11611 = n11610 ^ n2953 ^ 1'b0 ;
  assign n11612 = n998 & n11611 ;
  assign n11613 = n3406 & ~n6866 ;
  assign n11614 = n11613 ^ n2390 ^ 1'b0 ;
  assign n11615 = n8265 ^ n7904 ^ 1'b0 ;
  assign n11616 = n9911 | n11615 ;
  assign n11617 = n3898 | n11616 ;
  assign n11619 = n6949 ^ n753 ^ n180 ;
  assign n11618 = n6844 ^ n4114 ^ 1'b0 ;
  assign n11620 = n11619 ^ n11618 ^ n3075 ;
  assign n11621 = n1964 | n4216 ;
  assign n11622 = n11621 ^ n2752 ^ 1'b0 ;
  assign n11623 = n8756 ^ n4694 ^ 1'b0 ;
  assign n11624 = n9002 | n11623 ;
  assign n11626 = n2994 ^ n839 ^ n514 ;
  assign n11627 = n6398 & ~n9885 ;
  assign n11628 = n11627 ^ n2857 ^ 1'b0 ;
  assign n11629 = n11626 & ~n11628 ;
  assign n11630 = ~n7211 & n11629 ;
  assign n11625 = ~n4406 & n10267 ;
  assign n11631 = n11630 ^ n11625 ^ 1'b0 ;
  assign n11632 = ( ~n405 & n963 ) | ( ~n405 & n5628 ) | ( n963 & n5628 ) ;
  assign n11633 = n2687 & ~n6933 ;
  assign n11634 = ( ~n9674 & n11202 ) | ( ~n9674 & n11633 ) | ( n11202 & n11633 ) ;
  assign n11635 = n1175 & ~n5578 ;
  assign n11636 = n2014 & n3599 ;
  assign n11637 = n9766 | n11636 ;
  assign n11638 = n11635 & ~n11637 ;
  assign n11639 = n11634 | n11638 ;
  assign n11640 = n11632 & ~n11639 ;
  assign n11641 = n65 | n745 ;
  assign n11642 = n3229 & ~n11641 ;
  assign n11643 = n11642 ^ n4429 ^ n3054 ;
  assign n11644 = ( ~n908 & n2005 ) | ( ~n908 & n6763 ) | ( n2005 & n6763 ) ;
  assign n11645 = ~n2385 & n4981 ;
  assign n11646 = n6620 & n11645 ;
  assign n11647 = n1120 & ~n11646 ;
  assign n11648 = n11647 ^ n3542 ^ 1'b0 ;
  assign n11649 = n11648 ^ n10224 ^ 1'b0 ;
  assign n11650 = n8043 & ~n11649 ;
  assign n11651 = n3357 ^ n3232 ^ 1'b0 ;
  assign n11652 = n983 & ~n11651 ;
  assign n11654 = n2271 & n7870 ;
  assign n11655 = n11654 ^ n2524 ^ 1'b0 ;
  assign n11656 = ( n2860 & n6064 ) | ( n2860 & n11655 ) | ( n6064 & n11655 ) ;
  assign n11653 = n5008 ^ n2328 ^ n191 ;
  assign n11657 = n11656 ^ n11653 ^ n5740 ;
  assign n11658 = n3038 ^ n216 ^ 1'b0 ;
  assign n11659 = ~n4990 & n11658 ;
  assign n11660 = n6159 & n11659 ;
  assign n11661 = ~n2986 & n8310 ;
  assign n11662 = n11660 & n11661 ;
  assign n11663 = n7017 ^ n1684 ^ 1'b0 ;
  assign n11664 = n3421 | n11663 ;
  assign n11665 = n2588 ^ n1064 ^ 1'b0 ;
  assign n11666 = n11664 | n11665 ;
  assign n11669 = n756 | n6814 ;
  assign n11670 = n11669 ^ n8630 ^ 1'b0 ;
  assign n11667 = ( n223 & n4264 ) | ( n223 & ~n7640 ) | ( n4264 & ~n7640 ) ;
  assign n11668 = n11667 ^ n5663 ^ 1'b0 ;
  assign n11671 = n11670 ^ n11668 ^ 1'b0 ;
  assign n11672 = n4515 ^ n1506 ^ 1'b0 ;
  assign n11673 = n7678 ^ n1980 ^ 1'b0 ;
  assign n11674 = ( ~n115 & n7697 ) | ( ~n115 & n11673 ) | ( n7697 & n11673 ) ;
  assign n11675 = n11672 & ~n11674 ;
  assign n11676 = n9839 & n11675 ;
  assign n11677 = n11671 | n11676 ;
  assign n11678 = n5684 & ~n11677 ;
  assign n11679 = n1726 & ~n9800 ;
  assign n11680 = ~n5953 & n11679 ;
  assign n11681 = n2980 ^ n1990 ^ 1'b0 ;
  assign n11682 = n150 & n11681 ;
  assign n11683 = n95 & n3319 ;
  assign n11684 = n6956 & n11683 ;
  assign n11685 = ~n11682 & n11684 ;
  assign n11686 = n11685 ^ n2050 ^ 1'b0 ;
  assign n11687 = n11680 | n11686 ;
  assign n11688 = n11687 ^ n2756 ^ 1'b0 ;
  assign n11689 = n3998 & n11688 ;
  assign n11690 = ~n809 & n9444 ;
  assign n11691 = n11690 ^ n5958 ^ 1'b0 ;
  assign n11692 = ~n1579 & n5272 ;
  assign n11693 = ( ~n811 & n4085 ) | ( ~n811 & n4647 ) | ( n4085 & n4647 ) ;
  assign n11694 = n2787 & ~n3988 ;
  assign n11695 = n7051 & n11694 ;
  assign n11696 = ( n4285 & n11693 ) | ( n4285 & ~n11695 ) | ( n11693 & ~n11695 ) ;
  assign n11697 = ~n11692 & n11696 ;
  assign n11698 = n6062 ^ n5942 ^ 1'b0 ;
  assign n11699 = n3568 ^ n3544 ^ 1'b0 ;
  assign n11700 = n7681 & n11699 ;
  assign n11701 = ( n1094 & n1877 ) | ( n1094 & n3310 ) | ( n1877 & n3310 ) ;
  assign n11702 = n11701 ^ n960 ^ 1'b0 ;
  assign n11703 = n475 & n11702 ;
  assign n11704 = n11703 ^ n6269 ^ 1'b0 ;
  assign n11705 = n9271 ^ n7411 ^ 1'b0 ;
  assign n11706 = ~n2667 & n11705 ;
  assign n11707 = n11706 ^ n3379 ^ 1'b0 ;
  assign n11708 = ~n2577 & n10942 ;
  assign n11709 = n6238 & n8551 ;
  assign n11710 = n2666 & n11709 ;
  assign n11711 = ~n11708 & n11710 ;
  assign n11712 = n10684 ^ n8585 ^ 1'b0 ;
  assign n11713 = ( n2289 & ~n4309 ) | ( n2289 & n5145 ) | ( ~n4309 & n5145 ) ;
  assign n11714 = n2539 & ~n9099 ;
  assign n11715 = n4961 & n11714 ;
  assign n11716 = n7265 ^ n951 ^ 1'b0 ;
  assign n11717 = n11716 ^ n156 ^ 1'b0 ;
  assign n11718 = n2832 ^ n271 ^ 1'b0 ;
  assign n11719 = n11718 ^ n7977 ^ 1'b0 ;
  assign n11720 = ~n4691 & n11719 ;
  assign n11722 = n2783 & n3245 ;
  assign n11721 = n913 & ~n10296 ;
  assign n11723 = n11722 ^ n11721 ^ 1'b0 ;
  assign n11724 = n434 | n4775 ;
  assign n11725 = n11408 & ~n11724 ;
  assign n11726 = ~n9765 & n11725 ;
  assign n11727 = n11726 ^ n10821 ^ 1'b0 ;
  assign n11728 = n856 & n7701 ;
  assign n11729 = ~n4218 & n11728 ;
  assign n11730 = n2525 ^ n696 ^ 1'b0 ;
  assign n11731 = n11730 ^ n8476 ^ 1'b0 ;
  assign n11732 = n2952 & ~n6855 ;
  assign n11733 = n11732 ^ n216 ^ 1'b0 ;
  assign n11734 = n3327 ^ n2196 ^ 1'b0 ;
  assign n11735 = n8274 ^ n4735 ^ n3307 ;
  assign n11737 = n2642 ^ n1770 ^ n1258 ;
  assign n11736 = n990 | n1076 ;
  assign n11738 = n11737 ^ n11736 ^ n3310 ;
  assign n11740 = n9843 ^ n2791 ^ n1960 ;
  assign n11739 = n1359 | n4291 ;
  assign n11741 = n11740 ^ n11739 ^ 1'b0 ;
  assign n11742 = n953 & ~n11680 ;
  assign n11743 = n11741 & n11742 ;
  assign n11744 = n9549 ^ n8783 ^ 1'b0 ;
  assign n11745 = n4100 & ~n4365 ;
  assign n11746 = n11745 ^ n5915 ^ n2798 ;
  assign n11747 = ~n1964 & n2374 ;
  assign n11748 = n10555 & n11747 ;
  assign n11749 = ( n2146 & n6073 ) | ( n2146 & ~n11748 ) | ( n6073 & ~n11748 ) ;
  assign n11750 = n4417 & n11749 ;
  assign n11751 = n7630 ^ n3084 ^ 1'b0 ;
  assign n11752 = n11751 ^ n7055 ^ 1'b0 ;
  assign n11753 = n2114 | n11670 ;
  assign n11754 = n534 ^ n312 ^ 1'b0 ;
  assign n11755 = n255 | n11754 ;
  assign n11756 = n73 & ~n11755 ;
  assign n11757 = n9727 ^ n5965 ^ 1'b0 ;
  assign n11758 = n9893 & n11757 ;
  assign n11759 = n11756 & n11758 ;
  assign n11760 = n1142 & ~n1913 ;
  assign n11761 = ~n5282 & n11760 ;
  assign n11762 = ~n11759 & n11761 ;
  assign n11763 = ( n882 & ~n948 ) | ( n882 & n1926 ) | ( ~n948 & n1926 ) ;
  assign n11765 = n8799 ^ n1871 ^ 1'b0 ;
  assign n11766 = n6361 & ~n11765 ;
  assign n11764 = ( n4134 & n4803 ) | ( n4134 & n9055 ) | ( n4803 & n9055 ) ;
  assign n11767 = n11766 ^ n11764 ^ 1'b0 ;
  assign n11768 = ~n11763 & n11767 ;
  assign n11769 = n6493 ^ n2037 ^ 1'b0 ;
  assign n11770 = n11769 ^ n8622 ^ 1'b0 ;
  assign n11771 = n11768 & ~n11770 ;
  assign n11772 = n6272 | n11771 ;
  assign n11773 = ~n3046 & n11772 ;
  assign n11776 = n2040 | n3526 ;
  assign n11777 = n6125 | n11776 ;
  assign n11774 = ~n2953 & n4715 ;
  assign n11775 = n954 | n11774 ;
  assign n11778 = n11777 ^ n11775 ^ 1'b0 ;
  assign n11779 = ~n603 & n3168 ;
  assign n11780 = n1556 & n11779 ;
  assign n11781 = n6431 ^ n4770 ^ n3861 ;
  assign n11782 = n11781 ^ n101 ^ 1'b0 ;
  assign n11783 = n4278 ^ n1513 ^ 1'b0 ;
  assign n11784 = n11782 & ~n11783 ;
  assign n11785 = n11784 ^ n400 ^ 1'b0 ;
  assign n11786 = n11785 ^ n2350 ^ n1221 ;
  assign n11787 = n4436 | n11786 ;
  assign n11788 = n2662 | n11787 ;
  assign n11789 = ( n2335 & ~n7545 ) | ( n2335 & n8398 ) | ( ~n7545 & n8398 ) ;
  assign n11790 = ( n1444 & n6614 ) | ( n1444 & ~n7642 ) | ( n6614 & ~n7642 ) ;
  assign n11791 = ~n11789 & n11790 ;
  assign n11792 = n3574 & n11791 ;
  assign n11793 = n9513 ^ n3770 ^ 1'b0 ;
  assign n11794 = n3566 & n11793 ;
  assign n11795 = n7457 ^ n7009 ^ 1'b0 ;
  assign n11796 = n11795 ^ n157 ^ 1'b0 ;
  assign n11797 = ~n3234 & n11796 ;
  assign n11798 = n11797 ^ n135 ^ 1'b0 ;
  assign n11800 = n276 ^ n91 ^ 1'b0 ;
  assign n11801 = n1055 & n11800 ;
  assign n11802 = ~n1812 & n11801 ;
  assign n11799 = n1170 & n4954 ;
  assign n11803 = n11802 ^ n11799 ^ 1'b0 ;
  assign n11804 = n3555 | n9643 ;
  assign n11805 = ~n7584 & n11804 ;
  assign n11806 = n2606 & ~n6350 ;
  assign n11807 = n11806 ^ n478 ^ 1'b0 ;
  assign n11808 = n6745 & ~n11807 ;
  assign n11809 = n408 & ~n6765 ;
  assign n11810 = n11809 ^ n5100 ^ 1'b0 ;
  assign n11811 = n11810 ^ n10442 ^ n9872 ;
  assign n11812 = n7201 & n11811 ;
  assign n11813 = n7300 ^ n2425 ^ 1'b0 ;
  assign n11814 = ~n93 & n1209 ;
  assign n11815 = n11814 ^ n870 ^ 1'b0 ;
  assign n11816 = n5338 & n8833 ;
  assign n11817 = n11816 ^ n536 ^ 1'b0 ;
  assign n11818 = n11815 & n11817 ;
  assign n11819 = n3248 & ~n10079 ;
  assign n11820 = n11819 ^ n1096 ^ 1'b0 ;
  assign n11822 = n2414 & n4011 ;
  assign n11823 = n11822 ^ n3094 ^ 1'b0 ;
  assign n11821 = n641 | n7482 ;
  assign n11824 = n11823 ^ n11821 ^ 1'b0 ;
  assign n11825 = ~n2851 & n11824 ;
  assign n11832 = ~n2449 & n8423 ;
  assign n11833 = n11832 ^ n1632 ^ n1334 ;
  assign n11826 = n3414 ^ n2660 ^ n177 ;
  assign n11827 = ~n5424 & n11826 ;
  assign n11828 = ~n203 & n7815 ;
  assign n11829 = n11828 ^ n8707 ^ 1'b0 ;
  assign n11830 = n11829 ^ n10054 ^ 1'b0 ;
  assign n11831 = n11827 & n11830 ;
  assign n11834 = n11833 ^ n11831 ^ 1'b0 ;
  assign n11835 = n2759 ^ n1633 ^ 1'b0 ;
  assign n11836 = ~n8287 & n11835 ;
  assign n11837 = ( n601 & ~n911 ) | ( n601 & n9014 ) | ( ~n911 & n9014 ) ;
  assign n11838 = n8741 ^ n8037 ^ 1'b0 ;
  assign n11839 = n7366 & ~n11838 ;
  assign n11840 = ~n11837 & n11839 ;
  assign n11841 = n11840 ^ n1184 ^ 1'b0 ;
  assign n11844 = ( n1114 & n3807 ) | ( n1114 & n3899 ) | ( n3807 & n3899 ) ;
  assign n11842 = n5276 & n8371 ;
  assign n11843 = n63 & n11842 ;
  assign n11845 = n11844 ^ n11843 ^ 1'b0 ;
  assign n11846 = ~n11355 & n11845 ;
  assign n11847 = n8208 ^ n1628 ^ n772 ;
  assign n11848 = n4371 | n8989 ;
  assign n11849 = n4258 & ~n7506 ;
  assign n11850 = n11849 ^ n10305 ^ 1'b0 ;
  assign n11852 = n5281 ^ n1135 ^ 1'b0 ;
  assign n11851 = n7862 ^ n5893 ^ 1'b0 ;
  assign n11853 = n11852 ^ n11851 ^ 1'b0 ;
  assign n11854 = n6535 ^ n4696 ^ 1'b0 ;
  assign n11858 = n400 | n2550 ;
  assign n11859 = n10493 & ~n11858 ;
  assign n11856 = ~n965 & n4231 ;
  assign n11857 = n9253 & n11856 ;
  assign n11860 = n11859 ^ n11857 ^ 1'b0 ;
  assign n11861 = n1841 & n11860 ;
  assign n11855 = n1155 & ~n2350 ;
  assign n11862 = n11861 ^ n11855 ^ 1'b0 ;
  assign n11863 = n3248 ^ n839 ^ 1'b0 ;
  assign n11864 = ~n1532 & n11863 ;
  assign n11865 = n10488 ^ n7467 ^ 1'b0 ;
  assign n11866 = ( ~n826 & n1061 ) | ( ~n826 & n4153 ) | ( n1061 & n4153 ) ;
  assign n11867 = n5327 ^ n3876 ^ 1'b0 ;
  assign n11868 = ( n5018 & ~n8292 ) | ( n5018 & n11867 ) | ( ~n8292 & n11867 ) ;
  assign n11869 = n11866 & ~n11868 ;
  assign n11870 = n11869 ^ n11354 ^ 1'b0 ;
  assign n11871 = n11870 ^ n637 ^ 1'b0 ;
  assign n11872 = n11871 ^ n5400 ^ 1'b0 ;
  assign n11873 = n1545 & n6557 ;
  assign n11874 = n5543 & ~n9902 ;
  assign n11875 = n11874 ^ n5747 ^ 1'b0 ;
  assign n11876 = ~n191 & n3597 ;
  assign n11877 = n11875 & ~n11876 ;
  assign n11878 = n11314 ^ n2051 ^ 1'b0 ;
  assign n11879 = n11470 & ~n11878 ;
  assign n11880 = n7070 | n11445 ;
  assign n11881 = n7718 ^ n466 ^ 1'b0 ;
  assign n11882 = n2274 | n5880 ;
  assign n11883 = n55 & ~n4846 ;
  assign n11884 = ( ~n4460 & n6166 ) | ( ~n4460 & n11883 ) | ( n6166 & n11883 ) ;
  assign n11885 = ~n11882 & n11884 ;
  assign n11886 = n11885 ^ n8489 ^ 1'b0 ;
  assign n11887 = ~n11401 & n11852 ;
  assign n11888 = ~n808 & n11887 ;
  assign n11889 = n8530 & ~n11888 ;
  assign n11890 = ~n11886 & n11889 ;
  assign n11891 = n650 | n4723 ;
  assign n11892 = n11891 ^ n2582 ^ 1'b0 ;
  assign n11893 = ( ~n951 & n7506 ) | ( ~n951 & n11892 ) | ( n7506 & n11892 ) ;
  assign n11894 = n2558 & ~n5667 ;
  assign n11895 = n2939 & ~n3450 ;
  assign n11896 = n11895 ^ n2493 ^ 1'b0 ;
  assign n11897 = n10017 & ~n11896 ;
  assign n11898 = ~n4105 & n11897 ;
  assign n11899 = n4896 & ~n5607 ;
  assign n11900 = n11899 ^ n1093 ^ 1'b0 ;
  assign n11901 = n8389 & ~n11900 ;
  assign n11903 = n1179 & ~n10223 ;
  assign n11904 = n11903 ^ n3190 ^ 1'b0 ;
  assign n11902 = ~n5872 & n11764 ;
  assign n11905 = n11904 ^ n11902 ^ 1'b0 ;
  assign n11906 = n7343 ^ n5424 ^ n2211 ;
  assign n11907 = n11906 ^ n5146 ^ n4543 ;
  assign n11908 = n8953 & ~n11907 ;
  assign n11909 = n11905 & ~n11908 ;
  assign n11910 = n4264 & n11909 ;
  assign n11911 = n11901 & n11910 ;
  assign n11912 = n1316 & n2045 ;
  assign n11913 = ~n6134 & n11166 ;
  assign n11914 = n11913 ^ n2076 ^ 1'b0 ;
  assign n11915 = n11914 ^ n7813 ^ 1'b0 ;
  assign n11916 = ( n9128 & n11912 ) | ( n9128 & n11915 ) | ( n11912 & n11915 ) ;
  assign n11917 = n10171 ^ n10008 ^ 1'b0 ;
  assign n11918 = n9236 | n11917 ;
  assign n11919 = n11918 ^ n3997 ^ 1'b0 ;
  assign n11921 = n4461 ^ n580 ^ n303 ;
  assign n11922 = ( ~n2754 & n5563 ) | ( ~n2754 & n11570 ) | ( n5563 & n11570 ) ;
  assign n11924 = n7233 ^ n3205 ^ 1'b0 ;
  assign n11923 = n1849 & n10563 ;
  assign n11925 = n11924 ^ n11923 ^ 1'b0 ;
  assign n11926 = ~n11922 & n11925 ;
  assign n11927 = n11921 & n11926 ;
  assign n11920 = ~n5578 & n8285 ;
  assign n11928 = n11927 ^ n11920 ^ 1'b0 ;
  assign n11931 = n4801 ^ n3229 ^ 1'b0 ;
  assign n11932 = n11931 ^ n4171 ^ 1'b0 ;
  assign n11933 = n1010 | n3951 ;
  assign n11934 = n11932 | n11933 ;
  assign n11935 = n5881 ^ n5732 ^ 1'b0 ;
  assign n11936 = n11934 & n11935 ;
  assign n11929 = n11843 ^ n4287 ^ 1'b0 ;
  assign n11930 = n10886 & n11929 ;
  assign n11937 = n11936 ^ n11930 ^ 1'b0 ;
  assign n11938 = n5667 | n11937 ;
  assign n11939 = n65 | n321 ;
  assign n11940 = n1339 | n11939 ;
  assign n11941 = ( n525 & n3503 ) | ( n525 & n11940 ) | ( n3503 & n11940 ) ;
  assign n11942 = n8919 ^ n1311 ^ 1'b0 ;
  assign n11943 = n11942 ^ n9314 ^ n368 ;
  assign n11947 = ~n2622 & n5352 ;
  assign n11948 = n2023 & n11947 ;
  assign n11944 = ~n548 & n784 ;
  assign n11945 = n6004 & n11944 ;
  assign n11946 = n2576 & n11945 ;
  assign n11949 = n11948 ^ n11946 ^ n2357 ;
  assign n11950 = n11069 ^ n5186 ^ 1'b0 ;
  assign n11951 = ~n4326 & n6304 ;
  assign n11952 = n11951 ^ n471 ^ 1'b0 ;
  assign n11953 = n11952 ^ n9118 ^ 1'b0 ;
  assign n11954 = ~n1658 & n11953 ;
  assign n11955 = n3973 ^ n72 ^ 1'b0 ;
  assign n11956 = n6446 ^ n6082 ^ n4685 ;
  assign n11957 = n1188 & ~n11956 ;
  assign n11959 = ~n157 & n2270 ;
  assign n11960 = ~n1251 & n11959 ;
  assign n11961 = n1964 & n11960 ;
  assign n11962 = n11961 ^ n7525 ^ 1'b0 ;
  assign n11958 = n5852 ^ n127 ^ 1'b0 ;
  assign n11963 = n11962 ^ n11958 ^ 1'b0 ;
  assign n11964 = n9522 ^ n3365 ^ 1'b0 ;
  assign n11965 = n5837 ^ n2815 ^ 1'b0 ;
  assign n11966 = n11965 ^ n6278 ^ n817 ;
  assign n11967 = ( n6660 & n7435 ) | ( n6660 & n9337 ) | ( n7435 & n9337 ) ;
  assign n11968 = ~n3542 & n9483 ;
  assign n11969 = n5797 & n8888 ;
  assign n11970 = n11969 ^ n9137 ^ 1'b0 ;
  assign n11971 = ~n4382 & n11970 ;
  assign n11972 = n6745 & ~n11266 ;
  assign n11973 = ~n2876 & n11972 ;
  assign n11974 = n3517 ^ n1134 ^ 1'b0 ;
  assign n11975 = ( n2866 & ~n5101 ) | ( n2866 & n11974 ) | ( ~n5101 & n11974 ) ;
  assign n11976 = n10999 & n11975 ;
  assign n11977 = n467 & ~n4066 ;
  assign n11978 = n11977 ^ n10509 ^ 1'b0 ;
  assign n11979 = n11976 | n11978 ;
  assign n11980 = n9169 | n11979 ;
  assign n11981 = n6322 & ~n9678 ;
  assign n11982 = n11981 ^ n8332 ^ 1'b0 ;
  assign n11983 = n1456 & n3346 ;
  assign n11984 = n11982 & ~n11983 ;
  assign n11985 = n9546 | n11984 ;
  assign n11986 = n1232 & ~n11985 ;
  assign n11987 = n3359 & ~n11986 ;
  assign n11988 = n7365 & n7374 ;
  assign n11989 = n2682 & ~n6696 ;
  assign n11990 = n11989 ^ n3248 ^ 1'b0 ;
  assign n11991 = n777 & ~n11990 ;
  assign n11992 = n4120 ^ n951 ^ 1'b0 ;
  assign n11993 = n2773 & ~n11992 ;
  assign n11994 = n11993 ^ n9886 ^ 1'b0 ;
  assign n11995 = n11991 & ~n11994 ;
  assign n11996 = n11995 ^ n3911 ^ 1'b0 ;
  assign n11997 = ~n4925 & n11777 ;
  assign n11998 = n9189 ^ n5543 ^ n5114 ;
  assign n11999 = ( ~n2502 & n2648 ) | ( ~n2502 & n5479 ) | ( n2648 & n5479 ) ;
  assign n12000 = ( ~n405 & n771 ) | ( ~n405 & n11999 ) | ( n771 & n11999 ) ;
  assign n12003 = n1427 ^ n263 ^ 1'b0 ;
  assign n12001 = n4140 | n10444 ;
  assign n12002 = n331 & ~n12001 ;
  assign n12004 = n12003 ^ n12002 ^ n8655 ;
  assign n12005 = ~n1395 & n3443 ;
  assign n12006 = ( n4383 & n8251 ) | ( n4383 & n8521 ) | ( n8251 & n8521 ) ;
  assign n12007 = n3755 | n12006 ;
  assign n12008 = ~n8830 & n12007 ;
  assign n12009 = ~n4004 & n6807 ;
  assign n12010 = n12009 ^ n7130 ^ 1'b0 ;
  assign n12011 = ~n3744 & n10176 ;
  assign n12012 = n12011 ^ n2354 ^ 1'b0 ;
  assign n12013 = ~n1435 & n12012 ;
  assign n12014 = n12013 ^ n10930 ^ 1'b0 ;
  assign n12015 = n4304 & ~n5459 ;
  assign n12016 = n12015 ^ n1826 ^ 1'b0 ;
  assign n12017 = n1032 | n1666 ;
  assign n12018 = n2129 | n12017 ;
  assign n12019 = n1522 ^ n1240 ^ 1'b0 ;
  assign n12020 = n12018 & n12019 ;
  assign n12021 = n12020 ^ n5344 ^ 1'b0 ;
  assign n12022 = n2292 ^ n1437 ^ 1'b0 ;
  assign n12024 = ( ~n2542 & n5881 ) | ( ~n2542 & n6495 ) | ( n5881 & n6495 ) ;
  assign n12023 = n809 | n3945 ;
  assign n12025 = n12024 ^ n12023 ^ 1'b0 ;
  assign n12026 = n536 | n2214 ;
  assign n12027 = n9634 ^ n2992 ^ 1'b0 ;
  assign n12028 = n12026 & ~n12027 ;
  assign n12029 = n6363 ^ n4920 ^ 1'b0 ;
  assign n12030 = ~n6634 & n12029 ;
  assign n12031 = n12030 ^ n11283 ^ 1'b0 ;
  assign n12032 = n2164 & n12031 ;
  assign n12033 = n12032 ^ n5615 ^ 1'b0 ;
  assign n12034 = n513 & ~n12033 ;
  assign n12035 = n2271 & n3957 ;
  assign n12036 = ~n1355 & n12035 ;
  assign n12037 = ( n1932 & n3198 ) | ( n1932 & ~n12036 ) | ( n3198 & ~n12036 ) ;
  assign n12038 = n11365 & ~n12037 ;
  assign n12040 = ~n529 & n1102 ;
  assign n12039 = n1600 & n4998 ;
  assign n12041 = n12040 ^ n12039 ^ 1'b0 ;
  assign n12042 = n835 & n12041 ;
  assign n12043 = n1547 & n3655 ;
  assign n12044 = n951 & n12043 ;
  assign n12045 = n2321 | n12044 ;
  assign n12046 = n12045 ^ n1109 ^ 1'b0 ;
  assign n12047 = n12042 & ~n12046 ;
  assign n12048 = ~n5806 & n12047 ;
  assign n12049 = n1157 | n3786 ;
  assign n12050 = n12049 ^ n7925 ^ n3595 ;
  assign n12051 = ~n4604 & n12050 ;
  assign n12056 = n2568 ^ n808 ^ n115 ;
  assign n12054 = n7322 ^ n1206 ^ n434 ;
  assign n12052 = n1658 ^ n108 ^ 1'b0 ;
  assign n12053 = n3870 & ~n12052 ;
  assign n12055 = n12054 ^ n12053 ^ n3336 ;
  assign n12057 = n12056 ^ n12055 ^ n3308 ;
  assign n12058 = ( n1370 & n3486 ) | ( n1370 & ~n3593 ) | ( n3486 & ~n3593 ) ;
  assign n12059 = n11464 ^ n6949 ^ n4275 ;
  assign n12060 = ~n6104 & n12059 ;
  assign n12061 = n124 & n12060 ;
  assign n12062 = n4693 | n11544 ;
  assign n12063 = n5420 & ~n6929 ;
  assign n12064 = n5891 | n11366 ;
  assign n12065 = n2733 & ~n12064 ;
  assign n12066 = ( n2876 & n2963 ) | ( n2876 & n4756 ) | ( n2963 & n4756 ) ;
  assign n12067 = n1129 | n12066 ;
  assign n12068 = n12067 ^ n5337 ^ 1'b0 ;
  assign n12069 = ~n2874 & n3401 ;
  assign n12070 = ~n4741 & n12069 ;
  assign n12071 = n378 & ~n2322 ;
  assign n12072 = n5776 & ~n9454 ;
  assign n12073 = n12071 & n12072 ;
  assign n12075 = n3741 & ~n10108 ;
  assign n12074 = ~n5615 & n8157 ;
  assign n12076 = n12075 ^ n12074 ^ 1'b0 ;
  assign n12077 = n2727 & n9330 ;
  assign n12078 = n4869 & ~n10825 ;
  assign n12079 = n12078 ^ n3158 ^ 1'b0 ;
  assign n12080 = n12077 | n12079 ;
  assign n12081 = ( ~n259 & n2412 ) | ( ~n259 & n5120 ) | ( n2412 & n5120 ) ;
  assign n12082 = n12081 ^ n2213 ^ n1426 ;
  assign n12084 = n5533 ^ n2583 ^ 1'b0 ;
  assign n12083 = n2497 & n10804 ;
  assign n12085 = n12084 ^ n12083 ^ 1'b0 ;
  assign n12086 = ~n9406 & n12085 ;
  assign n12087 = ~n2798 & n4337 ;
  assign n12088 = n12087 ^ n1343 ^ 1'b0 ;
  assign n12089 = n3383 ^ n1645 ^ 1'b0 ;
  assign n12090 = n3312 | n12089 ;
  assign n12091 = n4343 ^ n501 ^ 1'b0 ;
  assign n12092 = n12091 ^ n1768 ^ 1'b0 ;
  assign n12093 = n1891 & ~n12092 ;
  assign n12094 = n12093 ^ n3269 ^ 1'b0 ;
  assign n12095 = n12090 | n12094 ;
  assign n12096 = n7215 & n8751 ;
  assign n12097 = n12096 ^ n3312 ^ 1'b0 ;
  assign n12098 = ~n6287 & n12097 ;
  assign n12099 = n10850 & n12098 ;
  assign n12100 = n7033 ^ n4212 ^ 1'b0 ;
  assign n12101 = ~n6212 & n6837 ;
  assign n12102 = n1407 & n2196 ;
  assign n12103 = n4217 ^ n1120 ^ 1'b0 ;
  assign n12104 = n830 | n7195 ;
  assign n12105 = n12104 ^ n545 ^ 1'b0 ;
  assign n12106 = n12103 & n12105 ;
  assign n12107 = n6317 ^ n771 ^ 1'b0 ;
  assign n12108 = n7057 ^ n201 ^ 1'b0 ;
  assign n12110 = n1361 & n4452 ;
  assign n12111 = ~n1520 & n12110 ;
  assign n12109 = n448 | n9866 ;
  assign n12112 = n12111 ^ n12109 ^ 1'b0 ;
  assign n12113 = n994 ^ n780 ^ 1'b0 ;
  assign n12114 = ~n4975 & n12113 ;
  assign n12115 = ~n5244 & n12114 ;
  assign n12116 = ( n1484 & n7737 ) | ( n1484 & ~n7987 ) | ( n7737 & ~n7987 ) ;
  assign n12121 = n4430 ^ n3882 ^ 1'b0 ;
  assign n12118 = n5538 ^ n4275 ^ 1'b0 ;
  assign n12119 = n9253 & n12118 ;
  assign n12117 = n4863 | n10079 ;
  assign n12120 = n12119 ^ n12117 ^ 1'b0 ;
  assign n12122 = n12121 ^ n12120 ^ 1'b0 ;
  assign n12123 = n310 & ~n12122 ;
  assign n12124 = n8371 & ~n12123 ;
  assign n12126 = ( n1542 & n5149 ) | ( n1542 & n6808 ) | ( n5149 & n6808 ) ;
  assign n12127 = n12126 ^ n2786 ^ 1'b0 ;
  assign n12125 = n1523 & ~n3870 ;
  assign n12128 = n12127 ^ n12125 ^ 1'b0 ;
  assign n12130 = n8101 ^ n8024 ^ 1'b0 ;
  assign n12131 = n5066 & n12130 ;
  assign n12129 = n7588 ^ n350 ^ 1'b0 ;
  assign n12132 = n12131 ^ n12129 ^ 1'b0 ;
  assign n12133 = n9956 | n12132 ;
  assign n12134 = n8748 ^ n1582 ^ 1'b0 ;
  assign n12135 = ~n6060 & n12134 ;
  assign n12136 = n11359 ^ n8822 ^ 1'b0 ;
  assign n12137 = n9724 ^ n8072 ^ 1'b0 ;
  assign n12138 = n12136 & ~n12137 ;
  assign n12139 = n8424 ^ n5937 ^ 1'b0 ;
  assign n12140 = ( n647 & n919 ) | ( n647 & ~n6024 ) | ( n919 & ~n6024 ) ;
  assign n12141 = n12140 ^ n3551 ^ 1'b0 ;
  assign n12142 = n12139 & ~n12141 ;
  assign n12143 = n10288 ^ n4143 ^ 1'b0 ;
  assign n12146 = n4951 ^ n3769 ^ n1082 ;
  assign n12144 = n9833 ^ n1710 ^ 1'b0 ;
  assign n12145 = ~n8289 & n12144 ;
  assign n12147 = n12146 ^ n12145 ^ 1'b0 ;
  assign n12148 = n3658 | n12147 ;
  assign n12149 = n12143 | n12148 ;
  assign n12150 = ~n3742 & n12149 ;
  assign n12151 = n3212 & ~n4552 ;
  assign n12152 = n6129 ^ n3185 ^ 1'b0 ;
  assign n12153 = n2124 & n12152 ;
  assign n12158 = ~n2390 & n3353 ;
  assign n12159 = n12158 ^ n1050 ^ 1'b0 ;
  assign n12160 = n10779 ^ n7558 ^ 1'b0 ;
  assign n12161 = n12159 & ~n12160 ;
  assign n12154 = n9539 | n9740 ;
  assign n12155 = n7523 & ~n12154 ;
  assign n12156 = n1460 & ~n12056 ;
  assign n12157 = ~n12155 & n12156 ;
  assign n12162 = n12161 ^ n12157 ^ 1'b0 ;
  assign n12163 = n3067 ^ n3043 ^ 1'b0 ;
  assign n12164 = n12163 ^ n7567 ^ 1'b0 ;
  assign n12165 = ( n2733 & ~n3257 ) | ( n2733 & n4235 ) | ( ~n3257 & n4235 ) ;
  assign n12166 = n3112 & ~n5457 ;
  assign n12167 = n3662 & n6953 ;
  assign n12168 = n12167 ^ n6304 ^ n2876 ;
  assign n12169 = n12166 | n12168 ;
  assign n12170 = n12165 & n12169 ;
  assign n12171 = n6016 & n12170 ;
  assign n12172 = n2945 & n7187 ;
  assign n12173 = n1695 & n12172 ;
  assign n12174 = n8740 & ~n10329 ;
  assign n12175 = ~n838 & n6683 ;
  assign n12176 = n11508 & n12175 ;
  assign n12177 = n12176 ^ n5172 ^ 1'b0 ;
  assign n12178 = n5241 ^ n1554 ^ 1'b0 ;
  assign n12179 = n710 | n3343 ;
  assign n12180 = n12179 ^ n5713 ^ 1'b0 ;
  assign n12181 = n1585 | n3106 ;
  assign n12182 = n11723 & ~n12181 ;
  assign n12183 = n12182 ^ n6562 ^ 1'b0 ;
  assign n12184 = n10500 ^ n5389 ^ n1589 ;
  assign n12185 = n12184 ^ n4402 ^ n3517 ;
  assign n12186 = n12185 ^ n44 ^ 1'b0 ;
  assign n12187 = n7908 | n9951 ;
  assign n12188 = n3644 | n8651 ;
  assign n12189 = n11658 ^ n1603 ^ 1'b0 ;
  assign n12190 = n12188 & ~n12189 ;
  assign n12191 = n4371 ^ n2561 ^ n42 ;
  assign n12192 = n310 & ~n12191 ;
  assign n12193 = n5796 ^ n3971 ^ 1'b0 ;
  assign n12194 = ~n1823 & n12193 ;
  assign n12195 = n2334 ^ n1770 ^ 1'b0 ;
  assign n12196 = n7489 & n12195 ;
  assign n12198 = n12040 ^ n9140 ^ n3779 ;
  assign n12197 = n7915 ^ n383 ^ 1'b0 ;
  assign n12199 = n12198 ^ n12197 ^ 1'b0 ;
  assign n12200 = n8232 & n10374 ;
  assign n12201 = ~n3167 & n3918 ;
  assign n12202 = ~n3898 & n12201 ;
  assign n12203 = n11628 & ~n12202 ;
  assign n12204 = ~n7228 & n12203 ;
  assign n12205 = n9126 ^ n8260 ^ n2535 ;
  assign n12206 = n5130 & ~n9201 ;
  assign n12207 = n4150 & ~n12206 ;
  assign n12208 = ~n12205 & n12207 ;
  assign n12209 = n10051 ^ n2055 ^ 1'b0 ;
  assign n12210 = n8148 | n12209 ;
  assign n12211 = n12210 ^ n9917 ^ 1'b0 ;
  assign n12212 = n3303 & ~n7937 ;
  assign n12213 = n4428 ^ n1376 ^ 1'b0 ;
  assign n12214 = n2713 & n7251 ;
  assign n12215 = ~n7768 & n12214 ;
  assign n12216 = n12215 ^ n837 ^ 1'b0 ;
  assign n12217 = n12216 ^ n8223 ^ n4054 ;
  assign n12218 = n3096 & ~n3871 ;
  assign n12219 = n12218 ^ n8597 ^ 1'b0 ;
  assign n12220 = n3339 ^ n1064 ^ 1'b0 ;
  assign n12221 = n5912 ^ n1843 ^ 1'b0 ;
  assign n12222 = ( n26 & n953 ) | ( n26 & n12221 ) | ( n953 & n12221 ) ;
  assign n12223 = n12222 ^ n1563 ^ 1'b0 ;
  assign n12224 = n12220 & n12223 ;
  assign n12225 = n6149 & ~n8618 ;
  assign n12226 = n11934 ^ n4207 ^ 1'b0 ;
  assign n12227 = n9217 | n12226 ;
  assign n12228 = n10597 | n12227 ;
  assign n12229 = n12228 ^ n7550 ^ 1'b0 ;
  assign n12230 = n526 ^ n352 ^ 1'b0 ;
  assign n12231 = n2756 & ~n12230 ;
  assign n12232 = n5446 & ~n8821 ;
  assign n12233 = ~n157 & n12232 ;
  assign n12234 = n6602 ^ n3898 ^ n740 ;
  assign n12235 = n3826 ^ n2251 ^ 1'b0 ;
  assign n12236 = n3224 ^ n1278 ^ 1'b0 ;
  assign n12237 = n1721 & ~n12236 ;
  assign n12238 = ~n125 & n12237 ;
  assign n12239 = n3984 & n12238 ;
  assign n12240 = n2012 & ~n12239 ;
  assign n12241 = n11132 & n12240 ;
  assign n12242 = n12241 ^ n3519 ^ 1'b0 ;
  assign n12243 = n11391 & n12242 ;
  assign n12244 = n137 & n7022 ;
  assign n12245 = n12244 ^ n8259 ^ 1'b0 ;
  assign n12246 = ~n59 & n2276 ;
  assign n12247 = n12246 ^ n1221 ^ 1'b0 ;
  assign n12248 = n10196 | n12247 ;
  assign n12249 = ( n1149 & n5836 ) | ( n1149 & ~n12248 ) | ( n5836 & ~n12248 ) ;
  assign n12250 = ~n1135 & n2496 ;
  assign n12251 = n12250 ^ n3332 ^ 1'b0 ;
  assign n12252 = ~n7782 & n12251 ;
  assign n12253 = n9221 & n12252 ;
  assign n12254 = n6136 & ~n11459 ;
  assign n12255 = n12254 ^ n2645 ^ 1'b0 ;
  assign n12256 = n4326 ^ n3926 ^ 1'b0 ;
  assign n12257 = n12255 & n12256 ;
  assign n12258 = n650 & n9326 ;
  assign n12259 = n473 & n2471 ;
  assign n12260 = n12259 ^ n3245 ^ 1'b0 ;
  assign n12261 = n8998 ^ n1976 ^ n488 ;
  assign n12262 = ( ~n4366 & n12260 ) | ( ~n4366 & n12261 ) | ( n12260 & n12261 ) ;
  assign n12263 = ( ~n2745 & n7583 ) | ( ~n2745 & n7601 ) | ( n7583 & n7601 ) ;
  assign n12264 = n12263 ^ n3844 ^ 1'b0 ;
  assign n12265 = ~x10 & n12264 ;
  assign n12266 = n12265 ^ n510 ^ 1'b0 ;
  assign n12267 = n6280 | n12266 ;
  assign n12268 = n1682 & ~n4667 ;
  assign n12269 = n2113 | n12268 ;
  assign n12270 = n600 & ~n1368 ;
  assign n12271 = n12270 ^ n5254 ^ 1'b0 ;
  assign n12273 = n4690 ^ n2745 ^ n797 ;
  assign n12274 = n3957 & n12273 ;
  assign n12275 = n76 & n12274 ;
  assign n12272 = n6758 & n7025 ;
  assign n12276 = n12275 ^ n12272 ^ 1'b0 ;
  assign n12277 = n7236 ^ n4043 ^ 1'b0 ;
  assign n12278 = n12277 ^ n2934 ^ 1'b0 ;
  assign n12279 = n5673 & ~n12278 ;
  assign n12280 = n1281 & ~n4884 ;
  assign n12281 = n7392 & n12280 ;
  assign n12282 = n3943 & n12281 ;
  assign n12283 = n12282 ^ n8841 ^ 1'b0 ;
  assign n12284 = n863 | n1138 ;
  assign n12285 = n7198 ^ n5309 ^ 1'b0 ;
  assign n12286 = n2595 & n2880 ;
  assign n12287 = n12285 & n12286 ;
  assign n12288 = n7245 ^ n3222 ^ 1'b0 ;
  assign n12289 = n8934 ^ n8594 ^ 1'b0 ;
  assign n12290 = ~n2992 & n5016 ;
  assign n12291 = ( n1704 & n8947 ) | ( n1704 & ~n12290 ) | ( n8947 & ~n12290 ) ;
  assign n12292 = n101 & ~n12291 ;
  assign n12293 = ( ~n8509 & n12289 ) | ( ~n8509 & n12292 ) | ( n12289 & n12292 ) ;
  assign n12294 = n6020 | n8065 ;
  assign n12295 = n5616 & ~n12294 ;
  assign n12296 = n1731 & ~n12295 ;
  assign n12297 = n6746 ^ n492 ^ 1'b0 ;
  assign n12298 = n1419 & ~n12297 ;
  assign n12299 = n5095 & n10228 ;
  assign n12300 = ~n12298 & n12299 ;
  assign n12301 = n12300 ^ n4607 ^ 1'b0 ;
  assign n12304 = n2110 ^ n301 ^ 1'b0 ;
  assign n12302 = ( n523 & n4134 ) | ( n523 & n7176 ) | ( n4134 & n7176 ) ;
  assign n12303 = ( n203 & n11682 ) | ( n203 & n12302 ) | ( n11682 & n12302 ) ;
  assign n12305 = n12304 ^ n12303 ^ 1'b0 ;
  assign n12310 = ~n1926 & n8735 ;
  assign n12311 = ( n4165 & n6161 ) | ( n4165 & ~n12310 ) | ( n6161 & ~n12310 ) ;
  assign n12306 = n3202 ^ n1489 ^ 1'b0 ;
  assign n12307 = ~n944 & n12306 ;
  assign n12308 = n12307 ^ n7859 ^ 1'b0 ;
  assign n12309 = n10903 & ~n12308 ;
  assign n12312 = n12311 ^ n12309 ^ 1'b0 ;
  assign n12313 = n1645 & ~n12312 ;
  assign n12317 = n965 & ~n8406 ;
  assign n12318 = n11756 ^ n1197 ^ 1'b0 ;
  assign n12319 = n12317 & n12318 ;
  assign n12314 = n4521 ^ n2190 ^ 1'b0 ;
  assign n12315 = n4507 & ~n10385 ;
  assign n12316 = n12314 | n12315 ;
  assign n12320 = n12319 ^ n12316 ^ 1'b0 ;
  assign n12321 = n172 & ~n332 ;
  assign n12322 = n4471 | n9584 ;
  assign n12323 = n4121 | n5684 ;
  assign n12324 = ( n6442 & n6611 ) | ( n6442 & ~n8009 ) | ( n6611 & ~n8009 ) ;
  assign n12325 = n3579 ^ n3522 ^ n2205 ;
  assign n12326 = n12325 ^ n5881 ^ 1'b0 ;
  assign n12327 = n12324 & n12326 ;
  assign n12328 = ( ~n3426 & n12323 ) | ( ~n3426 & n12327 ) | ( n12323 & n12327 ) ;
  assign n12332 = n2528 & n10171 ;
  assign n12329 = n4287 & n11162 ;
  assign n12330 = ~n134 & n12329 ;
  assign n12331 = n6497 & ~n12330 ;
  assign n12333 = n12332 ^ n12331 ^ 1'b0 ;
  assign n12334 = ~n1162 & n2319 ;
  assign n12335 = n4531 & n12334 ;
  assign n12336 = n11356 & ~n12335 ;
  assign n12337 = n12336 ^ n4976 ^ 1'b0 ;
  assign n12338 = n12337 ^ n7653 ^ 1'b0 ;
  assign n12339 = n3342 & ~n12338 ;
  assign n12340 = n9981 & n12339 ;
  assign n12341 = ~n3362 & n4736 ;
  assign n12342 = n12197 & n12341 ;
  assign n12343 = n1315 & ~n8153 ;
  assign n12345 = ~n3138 & n11283 ;
  assign n12346 = n12345 ^ n177 ^ 1'b0 ;
  assign n12344 = n1700 & n1880 ;
  assign n12347 = n12346 ^ n12344 ^ 1'b0 ;
  assign n12348 = n12220 & ~n12347 ;
  assign n12349 = n12348 ^ n6797 ^ 1'b0 ;
  assign n12350 = n6899 ^ n3570 ^ 1'b0 ;
  assign n12351 = ~n957 & n12350 ;
  assign n12352 = n5862 ^ n98 ^ 1'b0 ;
  assign n12353 = n4104 & n12352 ;
  assign n12359 = n3969 & ~n11190 ;
  assign n12360 = n6101 & n12359 ;
  assign n12354 = n1800 & ~n2693 ;
  assign n12355 = n12354 ^ n6180 ^ 1'b0 ;
  assign n12356 = ~n4413 & n12355 ;
  assign n12357 = n5519 & n12356 ;
  assign n12358 = n12357 ^ n7868 ^ n7213 ;
  assign n12361 = n12360 ^ n12358 ^ 1'b0 ;
  assign n12362 = n12353 & ~n12361 ;
  assign n12363 = n11888 ^ n8678 ^ 1'b0 ;
  assign n12364 = n6139 & ~n6424 ;
  assign n12365 = ~n299 & n2524 ;
  assign n12366 = n8574 & n12365 ;
  assign n12367 = n5706 & n8555 ;
  assign n12368 = ~n3868 & n12367 ;
  assign n12369 = n12368 ^ n10163 ^ n5718 ;
  assign n12370 = n534 & n12369 ;
  assign n12371 = n12370 ^ n4405 ^ 1'b0 ;
  assign n12372 = ~n11538 & n12371 ;
  assign n12373 = n6880 ^ n6091 ^ 1'b0 ;
  assign n12374 = n12373 ^ n5813 ^ n1006 ;
  assign n12377 = n1179 & ~n1525 ;
  assign n12375 = n3459 | n8889 ;
  assign n12376 = n115 & n12375 ;
  assign n12378 = n12377 ^ n12376 ^ 1'b0 ;
  assign n12379 = ~n3463 & n7126 ;
  assign n12381 = n5599 & ~n9414 ;
  assign n12382 = n4730 & n12381 ;
  assign n12380 = n1727 & n10816 ;
  assign n12383 = n12382 ^ n12380 ^ 1'b0 ;
  assign n12384 = n6702 | n12383 ;
  assign n12385 = n3855 & ~n10827 ;
  assign n12386 = n1122 & ~n2805 ;
  assign n12387 = ~n4704 & n12386 ;
  assign n12388 = n12387 ^ n654 ^ 1'b0 ;
  assign n12389 = n5354 & ~n6574 ;
  assign n12390 = n12389 ^ n2801 ^ 1'b0 ;
  assign n12391 = n8133 & n12097 ;
  assign n12392 = n4890 | n5657 ;
  assign n12393 = n10017 & ~n12392 ;
  assign n12394 = n12393 ^ n4805 ^ 1'b0 ;
  assign n12395 = n12394 ^ n8183 ^ n1285 ;
  assign n12396 = n10715 ^ n837 ^ 1'b0 ;
  assign n12397 = ~n276 & n12396 ;
  assign n12398 = n6481 & n8625 ;
  assign n12399 = n12397 & n12398 ;
  assign n12400 = n7133 ^ n592 ^ 1'b0 ;
  assign n12401 = n6855 | n7026 ;
  assign n12402 = n11260 ^ n6850 ^ 1'b0 ;
  assign n12403 = ( n3919 & n12401 ) | ( n3919 & ~n12402 ) | ( n12401 & ~n12402 ) ;
  assign n12404 = n3060 & n6293 ;
  assign n12405 = n2036 & n12404 ;
  assign n12406 = n349 | n8304 ;
  assign n12408 = n4405 & n6756 ;
  assign n12409 = ~n3983 & n12408 ;
  assign n12407 = n6299 ^ n1032 ^ 1'b0 ;
  assign n12410 = n12409 ^ n12407 ^ n4084 ;
  assign n12411 = n10843 ^ n4055 ^ 1'b0 ;
  assign n12412 = n3717 ^ n656 ^ 1'b0 ;
  assign n12413 = n3057 & n12412 ;
  assign n12414 = n12411 & n12413 ;
  assign n12415 = n10046 & ~n10679 ;
  assign n12416 = n12415 ^ n3426 ^ n2524 ;
  assign n12417 = n6879 & n12089 ;
  assign n12418 = n2495 & n12417 ;
  assign n12419 = n3312 ^ n1467 ^ 1'b0 ;
  assign n12420 = ~n11042 & n12419 ;
  assign n12421 = n12420 ^ n4316 ^ 1'b0 ;
  assign n12422 = n12418 & ~n12421 ;
  assign n12423 = n3104 ^ n903 ^ n794 ;
  assign n12424 = n2001 & n7801 ;
  assign n12425 = n12424 ^ n2277 ^ 1'b0 ;
  assign n12426 = n2198 ^ n1248 ^ n205 ;
  assign n12427 = n3557 & n12426 ;
  assign n12428 = n12425 & n12427 ;
  assign n12429 = n6929 ^ n803 ^ 1'b0 ;
  assign n12430 = n12428 | n12429 ;
  assign n12431 = n12423 & n12430 ;
  assign n12432 = n12431 ^ n9819 ^ n9036 ;
  assign n12433 = n2562 ^ n49 ^ 1'b0 ;
  assign n12434 = ~n271 & n960 ;
  assign n12435 = n12434 ^ n3920 ^ 1'b0 ;
  assign n12436 = n7140 | n12435 ;
  assign n12437 = n12436 ^ n6477 ^ 1'b0 ;
  assign n12438 = n7374 ^ n5091 ^ 1'b0 ;
  assign n12439 = n4210 & ~n12438 ;
  assign n12440 = ~x10 & n3151 ;
  assign n12441 = n8911 | n12440 ;
  assign n12442 = n12441 ^ n5145 ^ n1060 ;
  assign n12443 = n2878 ^ n816 ^ 1'b0 ;
  assign n12444 = n12443 ^ n3575 ^ n417 ;
  assign n12445 = n1322 ^ n352 ^ n82 ;
  assign n12446 = ~n3696 & n12445 ;
  assign n12447 = n12446 ^ n12025 ^ 1'b0 ;
  assign n12448 = n6169 ^ n4667 ^ 1'b0 ;
  assign n12449 = n5946 | n12448 ;
  assign n12450 = n7791 ^ n3060 ^ 1'b0 ;
  assign n12451 = ~n12449 & n12450 ;
  assign n12452 = n12451 ^ n10202 ^ n7585 ;
  assign n12453 = n378 | n5130 ;
  assign n12454 = n5020 | n12453 ;
  assign n12455 = n1880 & n12454 ;
  assign n12456 = n12455 ^ n3923 ^ 1'b0 ;
  assign n12457 = ( n137 & ~n4965 ) | ( n137 & n12456 ) | ( ~n4965 & n12456 ) ;
  assign n12458 = n11235 | n12457 ;
  assign n12459 = n12458 ^ n1007 ^ 1'b0 ;
  assign n12460 = ~n4427 & n10155 ;
  assign n12461 = ~n1412 & n1431 ;
  assign n12462 = n12461 ^ n1922 ^ 1'b0 ;
  assign n12463 = n12460 | n12462 ;
  assign n12464 = n2476 ^ n1509 ^ 1'b0 ;
  assign n12465 = n2623 & n12464 ;
  assign n12466 = ( ~n169 & n1672 ) | ( ~n169 & n12454 ) | ( n1672 & n12454 ) ;
  assign n12467 = n12466 ^ n11286 ^ 1'b0 ;
  assign n12468 = n5517 | n12467 ;
  assign n12469 = n12468 ^ n6623 ^ 1'b0 ;
  assign n12470 = ~n2287 & n12469 ;
  assign n12471 = ~n4237 & n12470 ;
  assign n12472 = n12471 ^ n8012 ^ 1'b0 ;
  assign n12473 = n1698 | n5162 ;
  assign n12474 = ~n903 & n12473 ;
  assign n12475 = n12474 ^ n1599 ^ 1'b0 ;
  assign n12476 = ( n6578 & ~n12472 ) | ( n6578 & n12475 ) | ( ~n12472 & n12475 ) ;
  assign n12477 = ( n8455 & n10153 ) | ( n8455 & n12476 ) | ( n10153 & n12476 ) ;
  assign n12478 = n797 ^ n777 ^ 1'b0 ;
  assign n12479 = n7040 & ~n7886 ;
  assign n12480 = n293 | n12479 ;
  assign n12481 = n3061 & ~n3443 ;
  assign n12482 = n10709 ^ n8522 ^ 1'b0 ;
  assign n12483 = n8323 ^ n6213 ^ n4618 ;
  assign n12484 = n6661 & n9494 ;
  assign n12485 = n12484 ^ n2745 ^ 1'b0 ;
  assign n12486 = n4221 & ~n12485 ;
  assign n12487 = ~n12483 & n12486 ;
  assign n12488 = n3179 & ~n6073 ;
  assign n12489 = n816 & n1353 ;
  assign n12490 = n1124 ^ n471 ^ 1'b0 ;
  assign n12491 = n7773 ^ n2168 ^ n1022 ;
  assign n12492 = n12491 ^ n3564 ^ 1'b0 ;
  assign n12493 = n2230 & ~n12492 ;
  assign n12494 = n12493 ^ n1634 ^ 1'b0 ;
  assign n12495 = n12494 ^ n9286 ^ n3918 ;
  assign n12496 = n10705 ^ n5494 ^ 1'b0 ;
  assign n12497 = n1578 & ~n12496 ;
  assign n12500 = n1527 ^ n1018 ^ n383 ;
  assign n12499 = n211 | n666 ;
  assign n12501 = n12500 ^ n12499 ^ 1'b0 ;
  assign n12502 = ~n7008 & n12501 ;
  assign n12503 = ( n4394 & ~n8099 ) | ( n4394 & n12502 ) | ( ~n8099 & n12502 ) ;
  assign n12498 = n9511 ^ n704 ^ 1'b0 ;
  assign n12504 = n12503 ^ n12498 ^ 1'b0 ;
  assign n12505 = ~n445 & n4927 ;
  assign n12506 = n5292 ^ n4175 ^ 1'b0 ;
  assign n12507 = ( n12275 & ~n12505 ) | ( n12275 & n12506 ) | ( ~n12505 & n12506 ) ;
  assign n12508 = n797 & ~n7441 ;
  assign n12509 = n12508 ^ n8207 ^ 1'b0 ;
  assign n12510 = ~n12507 & n12509 ;
  assign n12511 = n9519 | n10942 ;
  assign n12512 = n12511 ^ n12314 ^ 1'b0 ;
  assign n12513 = n12512 ^ n12260 ^ 1'b0 ;
  assign n12514 = ~n2387 & n12513 ;
  assign n12520 = n10163 ^ n547 ^ 1'b0 ;
  assign n12521 = ~n5169 & n6970 ;
  assign n12522 = ~n1153 & n12521 ;
  assign n12523 = n1611 & ~n12522 ;
  assign n12524 = ~n12520 & n12523 ;
  assign n12515 = ( n361 & n3762 ) | ( n361 & n6890 ) | ( n3762 & n6890 ) ;
  assign n12516 = n2058 | n12515 ;
  assign n12517 = n12516 ^ n4996 ^ 1'b0 ;
  assign n12518 = n12517 ^ n8976 ^ 1'b0 ;
  assign n12519 = n10171 & ~n12518 ;
  assign n12525 = n12524 ^ n12519 ^ n8436 ;
  assign n12530 = ~n366 & n5486 ;
  assign n12526 = n5954 ^ n4741 ^ 1'b0 ;
  assign n12527 = n2064 & n12526 ;
  assign n12528 = ~n6942 & n12527 ;
  assign n12529 = n1290 & n12528 ;
  assign n12531 = n12530 ^ n12529 ^ 1'b0 ;
  assign n12532 = n5596 & ~n10835 ;
  assign n12533 = n12532 ^ n160 ^ 1'b0 ;
  assign n12534 = n1105 | n12533 ;
  assign n12535 = n10832 | n12534 ;
  assign n12536 = ~n3070 & n6763 ;
  assign n12537 = n12536 ^ n7836 ^ 1'b0 ;
  assign n12538 = ~n5897 & n8673 ;
  assign n12539 = n12538 ^ n2521 ^ 1'b0 ;
  assign n12540 = n1296 | n6550 ;
  assign n12541 = n1885 & n2456 ;
  assign n12542 = n966 & ~n12541 ;
  assign n12543 = n12542 ^ n1562 ^ 1'b0 ;
  assign n12544 = n12543 ^ n2172 ^ 1'b0 ;
  assign n12545 = ~n8140 & n12544 ;
  assign n12546 = n7583 ^ n3112 ^ 1'b0 ;
  assign n12547 = n2682 & ~n12546 ;
  assign n12548 = n12547 ^ n6305 ^ n991 ;
  assign n12549 = n145 & ~n12548 ;
  assign n12550 = n3092 | n11786 ;
  assign n12551 = n12550 ^ n2220 ^ 1'b0 ;
  assign n12552 = n1202 & n1531 ;
  assign n12553 = n12552 ^ n4720 ^ 1'b0 ;
  assign n12554 = n12553 ^ n1517 ^ 1'b0 ;
  assign n12555 = n6948 ^ n3439 ^ 1'b0 ;
  assign n12556 = n6362 | n12555 ;
  assign n12557 = n2156 & ~n2825 ;
  assign n12558 = n1820 ^ n947 ^ 1'b0 ;
  assign n12559 = n3433 ^ n2489 ^ 1'b0 ;
  assign n12560 = n12558 | n12559 ;
  assign n12561 = n1890 ^ n1185 ^ 1'b0 ;
  assign n12562 = n698 | n12561 ;
  assign n12563 = n5886 | n12562 ;
  assign n12564 = n12560 & ~n12563 ;
  assign n12566 = n1712 | n11984 ;
  assign n12567 = n10390 | n12566 ;
  assign n12565 = n3893 & n7707 ;
  assign n12568 = n12567 ^ n12565 ^ 1'b0 ;
  assign n12569 = n1013 | n1832 ;
  assign n12570 = n3751 & ~n12569 ;
  assign n12571 = n4767 ^ n1633 ^ 1'b0 ;
  assign n12572 = n12570 | n12571 ;
  assign n12573 = n12572 ^ n11832 ^ 1'b0 ;
  assign n12574 = n1859 | n7103 ;
  assign n12575 = n4121 & ~n12574 ;
  assign n12576 = n6388 & ~n6802 ;
  assign n12577 = n2304 ^ n401 ^ 1'b0 ;
  assign n12578 = n4897 & ~n12577 ;
  assign n12579 = n12578 ^ n11929 ^ 1'b0 ;
  assign n12580 = n12576 & n12579 ;
  assign n12581 = ~n2281 & n12580 ;
  assign n12582 = n7956 ^ n6648 ^ n3466 ;
  assign n12583 = n12582 ^ n11598 ^ 1'b0 ;
  assign n12584 = n850 & n12583 ;
  assign n12585 = n5704 & n12584 ;
  assign n12586 = n12382 ^ n5837 ^ 1'b0 ;
  assign n12587 = n12586 ^ n11931 ^ n9417 ;
  assign n12588 = n6119 ^ n4461 ^ 1'b0 ;
  assign n12589 = ( ~n3312 & n8314 ) | ( ~n3312 & n12588 ) | ( n8314 & n12588 ) ;
  assign n12590 = n12589 ^ n3636 ^ 1'b0 ;
  assign n12591 = n1592 & ~n3730 ;
  assign n12592 = n12591 ^ n1110 ^ 1'b0 ;
  assign n12593 = n1822 & n12592 ;
  assign n12594 = n5519 ^ n2880 ^ 1'b0 ;
  assign n12595 = n10308 & ~n12594 ;
  assign n12596 = n12595 ^ n11419 ^ 1'b0 ;
  assign n12597 = ~n11931 & n12596 ;
  assign n12598 = n1904 & ~n3532 ;
  assign n12599 = n1330 & n12598 ;
  assign n12600 = n7348 & ~n12599 ;
  assign n12601 = n1927 & ~n1952 ;
  assign n12602 = n521 | n9140 ;
  assign n12603 = n12602 ^ n5016 ^ 1'b0 ;
  assign n12604 = n5039 & n12603 ;
  assign n12605 = ~n257 & n767 ;
  assign n12606 = n5688 & n12605 ;
  assign n12607 = n6960 | n12606 ;
  assign n12608 = ( n4377 & n6667 ) | ( n4377 & n9260 ) | ( n6667 & n9260 ) ;
  assign n12609 = n353 & ~n12051 ;
  assign n12610 = n12609 ^ n11161 ^ 1'b0 ;
  assign n12611 = n11745 ^ n6976 ^ n3620 ;
  assign n12612 = ( n1279 & ~n9008 ) | ( n1279 & n10958 ) | ( ~n9008 & n10958 ) ;
  assign n12613 = n3812 | n12612 ;
  assign n12614 = n12611 | n12613 ;
  assign n12615 = n12614 ^ n8089 ^ 1'b0 ;
  assign n12616 = n8770 | n12615 ;
  assign n12617 = n11334 ^ n6638 ^ 1'b0 ;
  assign n12618 = n790 ^ n551 ^ 1'b0 ;
  assign n12619 = n2370 & n4113 ;
  assign n12620 = n12619 ^ n245 ^ 1'b0 ;
  assign n12621 = n12620 ^ n4424 ^ 1'b0 ;
  assign n12622 = n7011 | n12621 ;
  assign n12623 = n3521 | n12622 ;
  assign n12624 = n5683 & n6785 ;
  assign n12625 = n12624 ^ n3800 ^ 1'b0 ;
  assign n12626 = n12625 ^ n1476 ^ 1'b0 ;
  assign n12627 = n777 | n4471 ;
  assign n12628 = ~n3914 & n12627 ;
  assign n12629 = n12626 & n12628 ;
  assign n12630 = n6455 & ~n11931 ;
  assign n12631 = n2230 ^ n334 ^ 1'b0 ;
  assign n12632 = n12631 ^ n10371 ^ n3770 ;
  assign n12633 = n10229 & n12632 ;
  assign n12634 = n5053 | n5861 ;
  assign n12635 = n8340 ^ n887 ^ 1'b0 ;
  assign n12636 = n12635 ^ n6358 ^ 1'b0 ;
  assign n12637 = n12634 & ~n12636 ;
  assign n12638 = n10917 ^ n10376 ^ 1'b0 ;
  assign n12639 = ~n5013 & n8049 ;
  assign n12640 = n271 | n6014 ;
  assign n12641 = n12640 ^ n3170 ^ 1'b0 ;
  assign n12642 = n12641 ^ n10532 ^ n1767 ;
  assign n12643 = ~n1676 & n10349 ;
  assign n12644 = n12643 ^ n8372 ^ 1'b0 ;
  assign n12645 = ( n3176 & n9045 ) | ( n3176 & n12644 ) | ( n9045 & n12644 ) ;
  assign n12646 = ~n4410 & n7150 ;
  assign n12647 = ~n7150 & n12646 ;
  assign n12648 = n4154 | n4690 ;
  assign n12649 = n12647 & ~n12648 ;
  assign n12650 = n12649 ^ n5914 ^ 1'b0 ;
  assign n12651 = n8373 & n12650 ;
  assign n12652 = ~n10656 & n12651 ;
  assign n12653 = n4454 | n5370 ;
  assign n12654 = n8608 | n12653 ;
  assign n12655 = n6938 | n9201 ;
  assign n12656 = ~n11051 & n12655 ;
  assign n12657 = ~n575 & n12656 ;
  assign n12658 = ( ~n778 & n853 ) | ( ~n778 & n2966 ) | ( n853 & n2966 ) ;
  assign n12659 = n12658 ^ n1330 ^ n1079 ;
  assign n12660 = n3379 & n8920 ;
  assign n12661 = n12660 ^ n299 ^ 1'b0 ;
  assign n12662 = n1167 ^ n496 ^ n40 ;
  assign n12663 = n3636 | n6585 ;
  assign n12664 = ( n2764 & ~n12662 ) | ( n2764 & n12663 ) | ( ~n12662 & n12663 ) ;
  assign n12665 = n3848 | n12664 ;
  assign n12666 = ~n287 & n7561 ;
  assign n12667 = ~n813 & n12666 ;
  assign n12668 = ~n10775 & n12667 ;
  assign n12669 = n11044 ^ n2745 ^ 1'b0 ;
  assign n12670 = n10180 | n12669 ;
  assign n12671 = n12668 & n12670 ;
  assign n12672 = ( x11 & n608 ) | ( x11 & n5277 ) | ( n608 & n5277 ) ;
  assign n12673 = n12672 ^ n4959 ^ 1'b0 ;
  assign n12674 = n6866 & ~n12673 ;
  assign n12675 = ( n3128 & n3413 ) | ( n3128 & ~n9251 ) | ( n3413 & ~n9251 ) ;
  assign n12676 = n12675 ^ n5145 ^ 1'b0 ;
  assign n12677 = n2818 & ~n12676 ;
  assign n12678 = n12677 ^ n3236 ^ 1'b0 ;
  assign n12679 = n11514 ^ n5039 ^ 1'b0 ;
  assign n12680 = n184 | n5047 ;
  assign n12681 = n95 | n6107 ;
  assign n12682 = n12681 ^ n8614 ^ 1'b0 ;
  assign n12683 = ~n10065 & n12682 ;
  assign n12684 = n281 | n3439 ;
  assign n12685 = n11443 ^ n8777 ^ 1'b0 ;
  assign n12686 = n6660 ^ n446 ^ 1'b0 ;
  assign n12687 = n221 | n12686 ;
  assign n12688 = n6511 & n7006 ;
  assign n12689 = ~n4454 & n5128 ;
  assign n12690 = n12689 ^ n7641 ^ 1'b0 ;
  assign n12691 = n12690 ^ n7875 ^ n4629 ;
  assign n12692 = n3495 ^ n1151 ^ 1'b0 ;
  assign n12693 = n12692 ^ n2345 ^ 1'b0 ;
  assign n12694 = ( n1303 & n2078 ) | ( n1303 & n12693 ) | ( n2078 & n12693 ) ;
  assign n12695 = n2385 ^ n1891 ^ 1'b0 ;
  assign n12696 = n2081 & ~n5101 ;
  assign n12697 = n12696 ^ n5595 ^ 1'b0 ;
  assign n12698 = n6357 & n12411 ;
  assign n12699 = n168 & ~n7361 ;
  assign n12700 = n12699 ^ n12425 ^ 1'b0 ;
  assign n12701 = n12700 ^ n12385 ^ n2490 ;
  assign n12702 = ( ~n2646 & n4632 ) | ( ~n2646 & n12055 ) | ( n4632 & n12055 ) ;
  assign n12706 = n112 | n3579 ;
  assign n12707 = n2841 & ~n12706 ;
  assign n12704 = n9550 ^ n5356 ^ n2454 ;
  assign n12705 = n12704 ^ n3951 ^ n2521 ;
  assign n12708 = n12707 ^ n12705 ^ 1'b0 ;
  assign n12703 = n8793 ^ n6888 ^ 1'b0 ;
  assign n12709 = n12708 ^ n12703 ^ n11318 ;
  assign n12711 = n600 & ~n1295 ;
  assign n12710 = n1363 | n1991 ;
  assign n12712 = n12711 ^ n12710 ^ 1'b0 ;
  assign n12713 = n6787 ^ n1791 ^ 1'b0 ;
  assign n12714 = n2556 & n4142 ;
  assign n12715 = n12714 ^ n7958 ^ 1'b0 ;
  assign n12716 = n7380 & ~n9628 ;
  assign n12717 = ~n12715 & n12716 ;
  assign n12718 = ~n2228 & n8829 ;
  assign n12719 = n9937 ^ n6729 ^ 1'b0 ;
  assign n12720 = ~n4617 & n12719 ;
  assign n12721 = ~n9118 & n12720 ;
  assign n12722 = n5380 & n12721 ;
  assign n12723 = ( ~n3203 & n7795 ) | ( ~n3203 & n11941 ) | ( n7795 & n11941 ) ;
  assign n12724 = n102 & ~n4667 ;
  assign n12725 = n12724 ^ n494 ^ 1'b0 ;
  assign n12726 = n12725 ^ n7535 ^ 1'b0 ;
  assign n12727 = n5174 & ~n12726 ;
  assign n12728 = n7870 ^ n7034 ^ 1'b0 ;
  assign n12729 = n12728 ^ n3773 ^ 1'b0 ;
  assign n12730 = n2606 & ~n12729 ;
  assign n12731 = n9245 ^ n1238 ^ 1'b0 ;
  assign n12732 = ~n4419 & n12731 ;
  assign n12735 = n3122 | n6129 ;
  assign n12736 = n1149 | n12735 ;
  assign n12733 = n3387 | n7864 ;
  assign n12734 = n5058 | n12733 ;
  assign n12737 = n12736 ^ n12734 ^ n709 ;
  assign n12738 = n1851 | n5740 ;
  assign n12739 = n4525 | n12738 ;
  assign n12740 = n12739 ^ n7398 ^ 1'b0 ;
  assign n12741 = n4009 & n12740 ;
  assign n12742 = n5107 ^ n822 ^ 1'b0 ;
  assign n12743 = n12742 ^ n2432 ^ 1'b0 ;
  assign n12744 = ~n12741 & n12743 ;
  assign n12745 = ~n395 & n4548 ;
  assign n12746 = n1446 | n4740 ;
  assign n12747 = ( n714 & n7049 ) | ( n714 & ~n7974 ) | ( n7049 & ~n7974 ) ;
  assign n12748 = n4720 ^ n3377 ^ n514 ;
  assign n12749 = ~n1053 & n12748 ;
  assign n12750 = n3713 | n12749 ;
  assign n12751 = n10560 ^ n9147 ^ n2405 ;
  assign n12752 = n12751 ^ n12196 ^ 1'b0 ;
  assign n12753 = ( n305 & ~n4574 ) | ( n305 & n6712 ) | ( ~n4574 & n6712 ) ;
  assign n12754 = n12753 ^ n11815 ^ 1'b0 ;
  assign n12755 = n12754 ^ n8319 ^ n2440 ;
  assign n12756 = ~n4230 & n5169 ;
  assign n12757 = n9619 | n12756 ;
  assign n12758 = n12757 ^ n5137 ^ 1'b0 ;
  assign n12759 = ~n2025 & n6899 ;
  assign n12765 = ~n84 & n2211 ;
  assign n12766 = n12765 ^ n3912 ^ 1'b0 ;
  assign n12767 = n2837 | n12766 ;
  assign n12760 = n4627 ^ n3542 ^ n1075 ;
  assign n12761 = n11143 | n12760 ;
  assign n12762 = n451 | n12761 ;
  assign n12763 = n8414 | n12762 ;
  assign n12764 = n4693 & ~n12763 ;
  assign n12768 = n12767 ^ n12764 ^ n1484 ;
  assign n12769 = n108 & ~n4577 ;
  assign n12770 = n12769 ^ n761 ^ 1'b0 ;
  assign n12771 = n12770 ^ n12548 ^ n7802 ;
  assign n12772 = ( n6221 & ~n10679 ) | ( n6221 & n12771 ) | ( ~n10679 & n12771 ) ;
  assign n12773 = n12772 ^ n3010 ^ 1'b0 ;
  assign n12774 = n7842 ^ n3833 ^ 1'b0 ;
  assign n12775 = n1029 & n12774 ;
  assign n12776 = ~n1000 & n12775 ;
  assign n12777 = n12773 & n12776 ;
  assign n12778 = n4465 ^ n739 ^ 1'b0 ;
  assign n12779 = n101 | n12778 ;
  assign n12780 = n2113 & ~n3119 ;
  assign n12781 = n12272 ^ n4567 ^ 1'b0 ;
  assign n12782 = ~n12780 & n12781 ;
  assign n12783 = ~n1201 & n12782 ;
  assign n12784 = n12783 ^ n9126 ^ 1'b0 ;
  assign n12785 = n12784 ^ n8823 ^ n2019 ;
  assign n12786 = n12779 | n12785 ;
  assign n12787 = n6406 | n12786 ;
  assign n12788 = n12718 ^ n6616 ^ 1'b0 ;
  assign n12789 = n3962 ^ n2492 ^ 1'b0 ;
  assign n12790 = n2173 & n9245 ;
  assign n12791 = ~n12789 & n12790 ;
  assign n12792 = n12791 ^ n8029 ^ 1'b0 ;
  assign n12793 = n5866 & ~n12792 ;
  assign n12794 = n1295 & n1442 ;
  assign n12795 = n10707 ^ n771 ^ 1'b0 ;
  assign n12796 = n12794 | n12795 ;
  assign n12797 = n12796 ^ n12502 ^ 1'b0 ;
  assign n12798 = n2434 ^ n601 ^ 1'b0 ;
  assign n12799 = ( n1459 & ~n7831 ) | ( n1459 & n12798 ) | ( ~n7831 & n12798 ) ;
  assign n12800 = n9624 & n12799 ;
  assign n12801 = n11594 ^ n10311 ^ 1'b0 ;
  assign n12802 = n10254 | n12801 ;
  assign n12803 = ( ~n68 & n2452 ) | ( ~n68 & n6914 ) | ( n2452 & n6914 ) ;
  assign n12804 = ~n8465 & n12803 ;
  assign n12805 = n12804 ^ n10340 ^ 1'b0 ;
  assign n12806 = n657 | n4541 ;
  assign n12807 = ~n2995 & n12806 ;
  assign n12808 = n7828 ^ n5307 ^ 1'b0 ;
  assign n12809 = n5284 ^ n544 ^ 1'b0 ;
  assign n12810 = n195 & n12809 ;
  assign n12815 = n5471 & n8030 ;
  assign n12814 = n8395 ^ n5580 ^ n481 ;
  assign n12811 = ~n7056 & n7383 ;
  assign n12812 = n12811 ^ n6379 ^ 1'b0 ;
  assign n12813 = ~n1591 & n12812 ;
  assign n12816 = n12815 ^ n12814 ^ n12813 ;
  assign n12817 = ~n12810 & n12816 ;
  assign n12818 = ( ~n607 & n1723 ) | ( ~n607 & n10712 ) | ( n1723 & n10712 ) ;
  assign n12819 = n10038 ^ n9140 ^ n1706 ;
  assign n12820 = n3479 & ~n12819 ;
  assign n12821 = n8170 ^ n578 ^ 1'b0 ;
  assign n12822 = n12821 ^ n11216 ^ 1'b0 ;
  assign n12823 = n3951 & n10113 ;
  assign n12825 = ~n1168 & n3133 ;
  assign n12826 = n12825 ^ n3469 ^ 1'b0 ;
  assign n12827 = n12826 ^ n2651 ^ n1386 ;
  assign n12824 = ~n9765 & n10349 ;
  assign n12828 = n12827 ^ n12824 ^ 1'b0 ;
  assign n12829 = n1623 & ~n6420 ;
  assign n12830 = n6381 & n12829 ;
  assign n12831 = n12830 ^ n3784 ^ n645 ;
  assign n12832 = ~n5748 & n12831 ;
  assign n12833 = ~n9146 & n12832 ;
  assign n12834 = n3558 ^ n710 ^ 1'b0 ;
  assign n12835 = n3692 & ~n12834 ;
  assign n12836 = n12835 ^ n11771 ^ 1'b0 ;
  assign n12837 = n3098 & ~n7290 ;
  assign n12838 = ( n3825 & n8462 ) | ( n3825 & ~n12837 ) | ( n8462 & ~n12837 ) ;
  assign n12839 = n12838 ^ n9282 ^ n332 ;
  assign n12840 = n1182 & ~n2944 ;
  assign n12841 = n5713 | n7208 ;
  assign n12842 = n12841 ^ n1563 ^ 1'b0 ;
  assign n12843 = ~n4518 & n7975 ;
  assign n12844 = ~n12842 & n12843 ;
  assign n12845 = ~n12840 & n12844 ;
  assign n12846 = n3332 & n7147 ;
  assign n12847 = n12846 ^ n7588 ^ 1'b0 ;
  assign n12848 = n9530 ^ n2888 ^ 1'b0 ;
  assign n12849 = n6383 | n12848 ;
  assign n12850 = n5645 | n12849 ;
  assign n12851 = n5457 ^ n442 ^ 1'b0 ;
  assign n12852 = n8792 ^ n799 ^ 1'b0 ;
  assign n12853 = n8700 & ~n12852 ;
  assign n12854 = n4728 ^ n59 ^ 1'b0 ;
  assign n12855 = n12854 ^ n8647 ^ 1'b0 ;
  assign n12856 = ( ~n9809 & n12853 ) | ( ~n9809 & n12855 ) | ( n12853 & n12855 ) ;
  assign n12857 = n12856 ^ n8912 ^ 1'b0 ;
  assign n12858 = ~n1632 & n1940 ;
  assign n12859 = n11508 & n12858 ;
  assign n12860 = n12859 ^ n9558 ^ 1'b0 ;
  assign n12861 = n11010 ^ n8070 ^ n4053 ;
  assign n12862 = ~n3769 & n12861 ;
  assign n12863 = n12862 ^ n11531 ^ 1'b0 ;
  assign n12864 = n12863 ^ n11729 ^ 1'b0 ;
  assign n12865 = n4728 & n8975 ;
  assign n12866 = n12865 ^ n417 ^ 1'b0 ;
  assign n12867 = n5377 & n7989 ;
  assign n12868 = n12867 ^ n12010 ^ 1'b0 ;
  assign n12869 = n12866 | n12868 ;
  assign n12870 = n6047 & ~n12869 ;
  assign n12871 = ~n3691 & n9903 ;
  assign n12872 = n3296 & n12871 ;
  assign n12873 = n12872 ^ n11754 ^ n7690 ;
  assign n12874 = n3105 | n3614 ;
  assign n12875 = ( ~n1856 & n2397 ) | ( ~n1856 & n7440 ) | ( n2397 & n7440 ) ;
  assign n12876 = n3112 ^ n35 ^ 1'b0 ;
  assign n12877 = ~n32 & n12876 ;
  assign n12878 = n1075 & ~n12877 ;
  assign n12879 = n951 & ~n11756 ;
  assign n12880 = n6513 ^ n492 ^ 1'b0 ;
  assign n12881 = n10922 ^ n5233 ^ 1'b0 ;
  assign n12882 = ~n12880 & n12881 ;
  assign n12883 = n12879 & n12882 ;
  assign n12884 = n1428 & ~n12883 ;
  assign n12885 = n5538 ^ n4735 ^ 1'b0 ;
  assign n12886 = n12885 ^ n5806 ^ 1'b0 ;
  assign n12887 = n11771 ^ n3602 ^ 1'b0 ;
  assign n12888 = n12887 ^ n897 ^ 1'b0 ;
  assign n12889 = ~n12854 & n12888 ;
  assign n12890 = n2328 ^ n960 ^ 1'b0 ;
  assign n12891 = n8498 ^ n6583 ^ 1'b0 ;
  assign n12892 = n3870 & ~n12891 ;
  assign n12893 = ~n12890 & n12892 ;
  assign n12895 = n1825 & ~n3413 ;
  assign n12896 = n6044 & n12895 ;
  assign n12897 = n772 & ~n12896 ;
  assign n12898 = ~n2277 & n12897 ;
  assign n12894 = n7405 ^ n2242 ^ 1'b0 ;
  assign n12899 = n12898 ^ n12894 ^ n4346 ;
  assign n12902 = ~n7312 & n10816 ;
  assign n12903 = n12902 ^ n118 ^ 1'b0 ;
  assign n12904 = n12903 ^ n601 ^ 1'b0 ;
  assign n12900 = ~n5032 & n11035 ;
  assign n12901 = n12900 ^ n5883 ^ 1'b0 ;
  assign n12905 = n12904 ^ n12901 ^ 1'b0 ;
  assign n12906 = n12899 & ~n12905 ;
  assign n12907 = n3252 | n10054 ;
  assign n12908 = n12907 ^ n10563 ^ 1'b0 ;
  assign n12909 = n2254 & n12908 ;
  assign n12911 = n324 & ~n2418 ;
  assign n12912 = ~n18 & n12911 ;
  assign n12913 = n1470 & ~n2817 ;
  assign n12914 = n12912 & n12913 ;
  assign n12915 = ~n7003 & n12914 ;
  assign n12910 = ~n4325 & n7847 ;
  assign n12916 = n12915 ^ n12910 ^ 1'b0 ;
  assign n12917 = ~n3669 & n5059 ;
  assign n12918 = n12917 ^ n797 ^ 1'b0 ;
  assign n12919 = n12918 ^ n7406 ^ 1'b0 ;
  assign n12920 = n12916 & n12919 ;
  assign n12921 = n5614 & n6564 ;
  assign n12922 = n9860 ^ n1447 ^ 1'b0 ;
  assign n12923 = n9388 & ~n12922 ;
  assign n12924 = n11339 & n12923 ;
  assign n12925 = n5007 & n12924 ;
  assign n12926 = ~n4079 & n5295 ;
  assign n12927 = n12926 ^ n8068 ^ n6438 ;
  assign n12928 = n859 | n12026 ;
  assign n12929 = n289 & n500 ;
  assign n12931 = ~n2631 & n7087 ;
  assign n12930 = n51 | n2580 ;
  assign n12932 = n12931 ^ n12930 ^ 1'b0 ;
  assign n12933 = ~n2303 & n7844 ;
  assign n12934 = n7017 | n12933 ;
  assign n12935 = ( ~n1173 & n1360 ) | ( ~n1173 & n3218 ) | ( n1360 & n3218 ) ;
  assign n12936 = n12935 ^ n2258 ^ 1'b0 ;
  assign n12937 = n1391 & ~n12936 ;
  assign n12938 = n12937 ^ n10329 ^ n2330 ;
  assign n12939 = ( n2158 & n3466 ) | ( n2158 & ~n6262 ) | ( n3466 & ~n6262 ) ;
  assign n12940 = n12939 ^ n914 ^ 1'b0 ;
  assign n12941 = n12940 ^ n4728 ^ 1'b0 ;
  assign n12942 = ( n2488 & n11944 ) | ( n2488 & n12941 ) | ( n11944 & n12941 ) ;
  assign n12943 = n4251 ^ n1232 ^ 1'b0 ;
  assign n12944 = n2431 & n5231 ;
  assign n12945 = ~n443 & n12944 ;
  assign n12946 = n4387 & n12945 ;
  assign n12947 = n12946 ^ n727 ^ 1'b0 ;
  assign n12948 = n7010 & n8281 ;
  assign n12949 = n12947 & n12948 ;
  assign n12950 = n5650 | n12949 ;
  assign n12951 = n1082 & ~n1779 ;
  assign n12952 = n6093 ^ n2330 ^ n723 ;
  assign n12953 = ~n7208 & n12952 ;
  assign n12954 = n12953 ^ n3119 ^ 1'b0 ;
  assign n12955 = ( n5697 & n12951 ) | ( n5697 & n12954 ) | ( n12951 & n12954 ) ;
  assign n12956 = ( n1050 & n7507 ) | ( n1050 & ~n12955 ) | ( n7507 & ~n12955 ) ;
  assign n12957 = n12150 ^ n5811 ^ 1'b0 ;
  assign n12958 = n3734 ^ n881 ^ 1'b0 ;
  assign n12959 = ( n5102 & ~n6109 ) | ( n5102 & n12958 ) | ( ~n6109 & n12958 ) ;
  assign n12960 = n11404 & ~n12959 ;
  assign n12961 = n8058 ^ n5256 ^ 1'b0 ;
  assign n12962 = n12961 ^ n7852 ^ 1'b0 ;
  assign n12963 = n4439 & ~n12962 ;
  assign n12964 = n2922 ^ n72 ^ 1'b0 ;
  assign n12965 = n8316 & n12964 ;
  assign n12966 = ( ~n1135 & n4060 ) | ( ~n1135 & n4563 ) | ( n4060 & n4563 ) ;
  assign n12967 = n12966 ^ n11602 ^ n4555 ;
  assign n12968 = n2819 & n3333 ;
  assign n12969 = ~n6166 & n12968 ;
  assign n12970 = n12969 ^ n8480 ^ 1'b0 ;
  assign n12971 = n4434 & ~n12970 ;
  assign n12972 = ~n2677 & n12971 ;
  assign n12973 = n12972 ^ n1727 ^ 1'b0 ;
  assign n12974 = ~n2561 & n12973 ;
  assign n12975 = n11558 & ~n12974 ;
  assign n12978 = n1461 & ~n3307 ;
  assign n12979 = n12978 ^ n10393 ^ 1'b0 ;
  assign n12976 = n5124 ^ n2581 ^ 1'b0 ;
  assign n12977 = ~n8267 & n12976 ;
  assign n12980 = n12979 ^ n12977 ^ 1'b0 ;
  assign n12981 = ( n2714 & ~n5788 ) | ( n2714 & n10323 ) | ( ~n5788 & n10323 ) ;
  assign n12982 = ~n4340 & n12981 ;
  assign n12983 = n7751 & n12982 ;
  assign n12984 = n461 | n9524 ;
  assign n12985 = n3761 & ~n12984 ;
  assign n12986 = n12481 ^ n11411 ^ 1'b0 ;
  assign n12987 = n104 & n3195 ;
  assign n12988 = n12987 ^ n1272 ^ 1'b0 ;
  assign n12989 = n11042 ^ n7348 ^ 1'b0 ;
  assign n12990 = ~n157 & n2836 ;
  assign n12991 = n12990 ^ n7634 ^ 1'b0 ;
  assign n12992 = n8115 & n12991 ;
  assign n12997 = n977 & n6229 ;
  assign n12993 = n5986 & n7366 ;
  assign n12994 = n12993 ^ n4849 ^ 1'b0 ;
  assign n12995 = n8775 & ~n12994 ;
  assign n12996 = n3593 | n12995 ;
  assign n12998 = n12997 ^ n12996 ^ 1'b0 ;
  assign n12999 = n10990 ^ n7269 ^ 1'b0 ;
  assign n13000 = n3387 & n9032 ;
  assign n13001 = n13000 ^ x4 ^ 1'b0 ;
  assign n13003 = ~n2922 & n4584 ;
  assign n13004 = n3568 & n13003 ;
  assign n13002 = n4886 | n10424 ;
  assign n13005 = n13004 ^ n13002 ^ 1'b0 ;
  assign n13006 = ~n13001 & n13005 ;
  assign n13007 = ( n3916 & ~n5623 ) | ( n3916 & n10527 ) | ( ~n5623 & n10527 ) ;
  assign n13008 = n9197 & n13007 ;
  assign n13009 = n13008 ^ n9578 ^ 1'b0 ;
  assign n13010 = n6776 | n13009 ;
  assign n13011 = n10352 ^ n9795 ^ 1'b0 ;
  assign n13012 = n5089 ^ n545 ^ 1'b0 ;
  assign n13013 = n8303 | n13012 ;
  assign n13014 = n3463 | n11302 ;
  assign n13015 = n644 | n13014 ;
  assign n13016 = ~n13013 & n13015 ;
  assign n13017 = ~n11454 & n13016 ;
  assign n13018 = ~n269 & n1507 ;
  assign n13019 = n888 | n13018 ;
  assign n13020 = n55 | n4071 ;
  assign n13021 = n13020 ^ n8103 ^ n4330 ;
  assign n13022 = n1612 & n12500 ;
  assign n13023 = n13022 ^ n687 ^ 1'b0 ;
  assign n13024 = n7236 ^ n6546 ^ 1'b0 ;
  assign n13025 = ~n3654 & n13024 ;
  assign n13026 = n3459 ^ n2070 ^ 1'b0 ;
  assign n13027 = n5620 & ~n13026 ;
  assign n13028 = ~n13025 & n13027 ;
  assign n13034 = ( ~n2382 & n5569 ) | ( ~n2382 & n10723 ) | ( n5569 & n10723 ) ;
  assign n13032 = n1380 & n6368 ;
  assign n13029 = n289 & ~n3469 ;
  assign n13030 = n5722 & n13029 ;
  assign n13031 = n3926 & ~n13030 ;
  assign n13033 = n13032 ^ n13031 ^ n8879 ;
  assign n13035 = n13034 ^ n13033 ^ 1'b0 ;
  assign n13036 = n657 | n895 ;
  assign n13037 = n13036 ^ n1768 ^ 1'b0 ;
  assign n13038 = n13037 ^ n6051 ^ n842 ;
  assign n13041 = n5280 & ~n8150 ;
  assign n13039 = n6692 ^ n5557 ^ 1'b0 ;
  assign n13040 = n484 | n13039 ;
  assign n13042 = n13041 ^ n13040 ^ 1'b0 ;
  assign n13044 = n3201 ^ n889 ^ 1'b0 ;
  assign n13045 = n4368 | n13044 ;
  assign n13046 = n13045 ^ n544 ^ 1'b0 ;
  assign n13043 = n5359 & n6725 ;
  assign n13047 = n13046 ^ n13043 ^ 1'b0 ;
  assign n13048 = n2149 ^ n881 ^ 1'b0 ;
  assign n13049 = ~n1164 & n13048 ;
  assign n13050 = n13049 ^ n8453 ^ n2346 ;
  assign n13051 = n13050 ^ n4364 ^ n1064 ;
  assign n13060 = n5453 ^ n5292 ^ n4847 ;
  assign n13061 = n5481 ^ n2152 ^ 1'b0 ;
  assign n13062 = n13060 & ~n13061 ;
  assign n13052 = n8703 ^ n6675 ^ 1'b0 ;
  assign n13053 = n2403 | n6091 ;
  assign n13054 = n4866 | n13053 ;
  assign n13055 = ~n42 & n13054 ;
  assign n13056 = n13055 ^ n2666 ^ 1'b0 ;
  assign n13057 = ( n3214 & n10115 ) | ( n3214 & ~n13056 ) | ( n10115 & ~n13056 ) ;
  assign n13058 = n13052 | n13057 ;
  assign n13059 = n13058 ^ n10267 ^ 1'b0 ;
  assign n13063 = n13062 ^ n13059 ^ 1'b0 ;
  assign n13064 = n8801 ^ n7483 ^ 1'b0 ;
  assign n13065 = ( n3709 & n8404 ) | ( n3709 & n10741 ) | ( n8404 & n10741 ) ;
  assign n13066 = n11019 | n13065 ;
  assign n13067 = n13066 ^ n740 ^ 1'b0 ;
  assign n13068 = n13067 ^ n12509 ^ n10133 ;
  assign n13069 = n2048 & n13068 ;
  assign n13070 = n5522 & n12319 ;
  assign n13071 = ~n13069 & n13070 ;
  assign n13072 = n3392 ^ n228 ^ 1'b0 ;
  assign n13073 = ( n4660 & n5352 ) | ( n4660 & ~n13072 ) | ( n5352 & ~n13072 ) ;
  assign n13074 = ~n1917 & n8790 ;
  assign n13075 = n13074 ^ n1200 ^ 1'b0 ;
  assign n13076 = n13075 ^ n6614 ^ 1'b0 ;
  assign n13077 = n2147 | n13076 ;
  assign n13078 = n577 & ~n13077 ;
  assign n13079 = n13078 ^ n2684 ^ 1'b0 ;
  assign n13080 = ( n4965 & n13073 ) | ( n4965 & ~n13079 ) | ( n13073 & ~n13079 ) ;
  assign n13081 = n545 & n11007 ;
  assign n13082 = ( n5132 & ~n5720 ) | ( n5132 & n13081 ) | ( ~n5720 & n13081 ) ;
  assign n13083 = ~n2755 & n13082 ;
  assign n13084 = n13083 ^ n6888 ^ 1'b0 ;
  assign n13085 = n2177 ^ n1619 ^ 1'b0 ;
  assign n13086 = n6590 & ~n13085 ;
  assign n13087 = ~n968 & n4576 ;
  assign n13088 = ~n13086 & n13087 ;
  assign n13089 = n13088 ^ n9490 ^ 1'b0 ;
  assign n13090 = ~n362 & n10034 ;
  assign n13091 = n4204 ^ n3955 ^ 1'b0 ;
  assign n13092 = n647 & ~n13091 ;
  assign n13093 = n13092 ^ n8199 ^ 1'b0 ;
  assign n13094 = n1017 & ~n4784 ;
  assign n13095 = n4201 | n13094 ;
  assign n13096 = n13095 ^ n3387 ^ 1'b0 ;
  assign n13097 = n3564 ^ n1147 ^ 1'b0 ;
  assign n13103 = n2721 | n3225 ;
  assign n13098 = n11002 ^ n3061 ^ 1'b0 ;
  assign n13099 = ~n888 & n13098 ;
  assign n13100 = n13099 ^ n12423 ^ 1'b0 ;
  assign n13101 = n6614 & n13100 ;
  assign n13102 = n13101 ^ n1465 ^ 1'b0 ;
  assign n13104 = n13103 ^ n13102 ^ n6541 ;
  assign n13105 = n11180 & ~n13104 ;
  assign n13106 = n11527 & n13105 ;
  assign n13107 = n5909 ^ n3022 ^ 1'b0 ;
  assign n13108 = ~n13073 & n13107 ;
  assign n13109 = n9155 ^ n2277 ^ 1'b0 ;
  assign n13110 = n13109 ^ n11253 ^ 1'b0 ;
  assign n13111 = n1820 ^ n893 ^ 1'b0 ;
  assign n13112 = ( n4617 & ~n10528 ) | ( n4617 & n13111 ) | ( ~n10528 & n13111 ) ;
  assign n13113 = n13112 ^ n1096 ^ 1'b0 ;
  assign n13114 = ( n5515 & ~n7944 ) | ( n5515 & n13113 ) | ( ~n7944 & n13113 ) ;
  assign n13115 = n10632 & n12319 ;
  assign n13116 = n13115 ^ n6533 ^ 1'b0 ;
  assign n13117 = n6219 ^ n2738 ^ 1'b0 ;
  assign n13118 = ~n3588 & n9610 ;
  assign n13119 = n13118 ^ n6656 ^ 1'b0 ;
  assign n13120 = n9702 ^ n7867 ^ 1'b0 ;
  assign n13121 = n3319 & n13120 ;
  assign n13122 = n13121 ^ n8199 ^ n4264 ;
  assign n13124 = n2580 ^ n1041 ^ 1'b0 ;
  assign n13123 = n4006 ^ n3135 ^ n471 ;
  assign n13125 = n13124 ^ n13123 ^ 1'b0 ;
  assign n13126 = ~n8448 & n9919 ;
  assign n13127 = ~n13125 & n13126 ;
  assign n13128 = ~n965 & n1409 ;
  assign n13129 = n13128 ^ n2650 ^ 1'b0 ;
  assign n13136 = n3167 & ~n9681 ;
  assign n13130 = n8540 ^ n5898 ^ 1'b0 ;
  assign n13131 = n3847 | n13130 ;
  assign n13132 = n13131 ^ n1506 ^ 1'b0 ;
  assign n13133 = n5809 & ~n13132 ;
  assign n13134 = n8374 ^ n228 ^ 1'b0 ;
  assign n13135 = n13133 & ~n13134 ;
  assign n13137 = n13136 ^ n13135 ^ 1'b0 ;
  assign n13138 = n11201 ^ n10034 ^ 1'b0 ;
  assign n13139 = n1636 | n5175 ;
  assign n13140 = n4371 ^ n2428 ^ 1'b0 ;
  assign n13141 = n11544 & n13140 ;
  assign n13142 = n3159 & n6810 ;
  assign n13143 = ( n141 & ~n7468 ) | ( n141 & n13142 ) | ( ~n7468 & n13142 ) ;
  assign n13144 = n6638 & ~n13143 ;
  assign n13145 = n13144 ^ n13038 ^ 1'b0 ;
  assign n13146 = ~n4668 & n7097 ;
  assign n13147 = n13146 ^ n134 ^ 1'b0 ;
  assign n13148 = ( x10 & ~n310 ) | ( x10 & n10588 ) | ( ~n310 & n10588 ) ;
  assign n13149 = n2214 & n3639 ;
  assign n13150 = n727 & ~n5050 ;
  assign n13151 = ~n3897 & n13150 ;
  assign n13152 = n6546 & ~n13151 ;
  assign n13153 = ~n649 & n13152 ;
  assign n13154 = n13153 ^ n11226 ^ 1'b0 ;
  assign n13155 = ( n2118 & n3495 ) | ( n2118 & n5092 ) | ( n3495 & n5092 ) ;
  assign n13156 = n411 | n498 ;
  assign n13157 = n13155 | n13156 ;
  assign n13158 = n9372 & n13157 ;
  assign n13159 = n4728 ^ n1262 ^ 1'b0 ;
  assign n13160 = n13159 ^ n3214 ^ n2885 ;
  assign n13161 = n6504 ^ n1340 ^ 1'b0 ;
  assign n13162 = ~n63 & n13161 ;
  assign n13163 = ~n7718 & n12684 ;
  assign n13164 = n9377 & n13163 ;
  assign n13166 = n2937 & n4322 ;
  assign n13167 = n13166 ^ n1830 ^ 1'b0 ;
  assign n13168 = ~n183 & n13167 ;
  assign n13169 = n13168 ^ n1628 ^ 1'b0 ;
  assign n13165 = ~n10366 & n11867 ;
  assign n13170 = n13169 ^ n13165 ^ n10711 ;
  assign n13171 = n1138 | n1506 ;
  assign n13172 = n13171 ^ n3027 ^ 1'b0 ;
  assign n13173 = n2569 & n10247 ;
  assign n13174 = n13172 & n13173 ;
  assign n13175 = n2980 ^ n408 ^ 1'b0 ;
  assign n13176 = n736 | n887 ;
  assign n13177 = ( ~n10263 & n13175 ) | ( ~n10263 & n13176 ) | ( n13175 & n13176 ) ;
  assign n13178 = ( n6790 & n7985 ) | ( n6790 & n13177 ) | ( n7985 & n13177 ) ;
  assign n13179 = n3263 & n13178 ;
  assign n13180 = ~n5167 & n7130 ;
  assign n13181 = n4640 ^ n3906 ^ 1'b0 ;
  assign n13182 = n13180 | n13181 ;
  assign n13190 = ~n4454 & n12827 ;
  assign n13191 = n4153 & n13190 ;
  assign n13187 = ~n3252 & n6504 ;
  assign n13188 = n2783 & n13187 ;
  assign n13189 = n316 & ~n13188 ;
  assign n13192 = n13191 ^ n13189 ^ 1'b0 ;
  assign n13183 = n8198 ^ n1701 ^ 1'b0 ;
  assign n13184 = n2569 ^ n1898 ^ 1'b0 ;
  assign n13185 = n13184 ^ n2584 ^ 1'b0 ;
  assign n13186 = ~n13183 & n13185 ;
  assign n13193 = n13192 ^ n13186 ^ n4982 ;
  assign n13194 = ~n1934 & n4273 ;
  assign n13195 = n13194 ^ n9341 ^ 1'b0 ;
  assign n13196 = n2674 ^ n1760 ^ 1'b0 ;
  assign n13197 = n8842 ^ n3159 ^ n2784 ;
  assign n13198 = n6235 ^ n448 ^ 1'b0 ;
  assign n13199 = ( n6110 & ~n9250 ) | ( n6110 & n13198 ) | ( ~n9250 & n13198 ) ;
  assign n13200 = n694 & n12321 ;
  assign n13201 = n271 & n13200 ;
  assign n13202 = n11131 ^ n7017 ^ n4393 ;
  assign n13204 = n1684 & ~n6078 ;
  assign n13205 = n13204 ^ n1063 ^ 1'b0 ;
  assign n13206 = n11518 ^ n8067 ^ n4842 ;
  assign n13207 = ~n13205 & n13206 ;
  assign n13203 = n1988 | n4054 ;
  assign n13208 = n13207 ^ n13203 ^ 1'b0 ;
  assign n13210 = n5242 ^ n1628 ^ 1'b0 ;
  assign n13209 = n1984 ^ n532 ^ 1'b0 ;
  assign n13211 = n13210 ^ n13209 ^ 1'b0 ;
  assign n13212 = n1374 | n12543 ;
  assign n13213 = n13212 ^ n9634 ^ 1'b0 ;
  assign n13216 = ( x10 & ~n5106 ) | ( x10 & n9241 ) | ( ~n5106 & n9241 ) ;
  assign n13214 = ~n247 & n2597 ;
  assign n13215 = ~n3750 & n13214 ;
  assign n13217 = n13216 ^ n13215 ^ n7087 ;
  assign n13220 = n11636 ^ n9566 ^ n3166 ;
  assign n13221 = ( n401 & ~n10163 ) | ( n401 & n13220 ) | ( ~n10163 & n13220 ) ;
  assign n13222 = n13221 ^ n11626 ^ 1'b0 ;
  assign n13218 = n11243 ^ n5970 ^ n799 ;
  assign n13219 = ~n1991 & n13218 ;
  assign n13223 = n13222 ^ n13219 ^ 1'b0 ;
  assign n13224 = ( n5178 & n5344 ) | ( n5178 & n8165 ) | ( n5344 & n8165 ) ;
  assign n13225 = n2627 | n5066 ;
  assign n13226 = ( n2130 & ~n8350 ) | ( n2130 & n12644 ) | ( ~n8350 & n12644 ) ;
  assign n13227 = n10070 ^ n4723 ^ 1'b0 ;
  assign n13228 = n13226 & ~n13227 ;
  assign n13229 = n13225 & n13228 ;
  assign n13230 = ~n386 & n13229 ;
  assign n13231 = ( n96 & n13224 ) | ( n96 & n13230 ) | ( n13224 & n13230 ) ;
  assign n13232 = n3421 & ~n12227 ;
  assign n13233 = n10252 ^ n7021 ^ 1'b0 ;
  assign n13234 = n893 & n6941 ;
  assign n13235 = n13234 ^ n1033 ^ 1'b0 ;
  assign n13236 = n13235 ^ n5229 ^ 1'b0 ;
  assign n13237 = ~n13233 & n13236 ;
  assign n13238 = n9597 ^ n132 ^ 1'b0 ;
  assign n13239 = ~n3440 & n5724 ;
  assign n13240 = n2225 ^ n1664 ^ 1'b0 ;
  assign n13241 = ~n7052 & n13240 ;
  assign n13242 = ~n13239 & n13241 ;
  assign n13243 = n1571 ^ n682 ^ n383 ;
  assign n13244 = n462 & ~n13243 ;
  assign n13245 = ~n6781 & n13244 ;
  assign n13246 = n6475 & ~n13245 ;
  assign n13247 = ( n4070 & n4948 ) | ( n4070 & n13246 ) | ( n4948 & n13246 ) ;
  assign n13248 = n12081 ^ n3244 ^ 1'b0 ;
  assign n13249 = n13248 ^ n7072 ^ 1'b0 ;
  assign n13250 = ( n6096 & ~n8127 ) | ( n6096 & n9887 ) | ( ~n8127 & n9887 ) ;
  assign n13251 = ( n1138 & ~n4493 ) | ( n1138 & n13250 ) | ( ~n4493 & n13250 ) ;
  assign n13255 = n4239 | n9378 ;
  assign n13256 = n13255 ^ n5495 ^ 1'b0 ;
  assign n13257 = n7425 ^ n4105 ^ n3890 ;
  assign n13258 = n340 & n7238 ;
  assign n13259 = n13257 & ~n13258 ;
  assign n13260 = n13256 & n13259 ;
  assign n13252 = n3030 ^ n44 ^ 1'b0 ;
  assign n13253 = n11065 | n13252 ;
  assign n13254 = ~n10723 & n13253 ;
  assign n13261 = n13260 ^ n13254 ^ 1'b0 ;
  assign n13262 = ( n6616 & ~n12630 ) | ( n6616 & n12637 ) | ( ~n12630 & n12637 ) ;
  assign n13265 = ( n230 & ~n1622 ) | ( n230 & n4249 ) | ( ~n1622 & n4249 ) ;
  assign n13263 = n7323 ^ n3288 ^ n977 ;
  assign n13264 = n154 & n13263 ;
  assign n13266 = n13265 ^ n13264 ^ 1'b0 ;
  assign n13267 = n9104 & n9857 ;
  assign n13268 = n11239 & n13267 ;
  assign n13269 = n3510 & n4702 ;
  assign n13270 = n13269 ^ n5748 ^ 1'b0 ;
  assign n13271 = n13270 ^ n1509 ^ 1'b0 ;
  assign n13272 = n564 & ~n13271 ;
  assign n13273 = n469 & n10176 ;
  assign n13274 = n13273 ^ n11137 ^ 1'b0 ;
  assign n13275 = n301 & ~n1415 ;
  assign n13276 = n13275 ^ n3691 ^ 1'b0 ;
  assign n13277 = n2750 & ~n13276 ;
  assign n13278 = n8057 & n13277 ;
  assign n13279 = n13278 ^ n7945 ^ 1'b0 ;
  assign n13280 = n13274 | n13279 ;
  assign n13281 = n4084 ^ n2309 ^ 1'b0 ;
  assign n13282 = ~n147 & n13281 ;
  assign n13283 = n3387 ^ n3151 ^ n1207 ;
  assign n13284 = n13283 ^ n4462 ^ n2370 ;
  assign n13285 = ( n10546 & n12109 ) | ( n10546 & n13284 ) | ( n12109 & n13284 ) ;
  assign n13286 = n2976 & ~n7262 ;
  assign n13287 = n11249 & ~n13286 ;
  assign n13288 = n426 | n13287 ;
  assign n13289 = n4128 & ~n13288 ;
  assign n13290 = n3816 ^ n3684 ^ 1'b0 ;
  assign n13291 = n5307 & ~n13290 ;
  assign n13292 = n13291 ^ n1811 ^ 1'b0 ;
  assign n13293 = ~n2982 & n13292 ;
  assign n13294 = n1660 ^ n953 ^ 1'b0 ;
  assign n13295 = n4123 | n13294 ;
  assign n13296 = n7228 & ~n10654 ;
  assign n13297 = ( ~n8975 & n13295 ) | ( ~n8975 & n13296 ) | ( n13295 & n13296 ) ;
  assign n13298 = n10282 | n13297 ;
  assign n13299 = n2502 & ~n13298 ;
  assign n13300 = n13299 ^ n11965 ^ 1'b0 ;
  assign n13301 = ~n16 & n4488 ;
  assign n13302 = n10829 | n13301 ;
  assign n13303 = n13301 & ~n13302 ;
  assign n13305 = n8463 ^ n1823 ^ 1'b0 ;
  assign n13306 = n10371 | n13305 ;
  assign n13304 = n9808 & n12960 ;
  assign n13307 = n13306 ^ n13304 ^ 1'b0 ;
  assign n13308 = ~n1045 & n5470 ;
  assign n13310 = n2661 & ~n7223 ;
  assign n13311 = n13310 ^ n7699 ^ 1'b0 ;
  assign n13309 = n1596 & n10568 ;
  assign n13312 = n13311 ^ n13309 ^ 1'b0 ;
  assign n13313 = n996 | n2832 ;
  assign n13314 = n1569 & ~n13313 ;
  assign n13315 = n13172 & ~n13314 ;
  assign n13316 = n13315 ^ n13277 ^ n926 ;
  assign n13317 = n10719 & ~n13316 ;
  assign n13318 = n2379 & n4014 ;
  assign n13319 = ~n2379 & n13318 ;
  assign n13320 = n8271 & ~n13319 ;
  assign n13321 = n12882 & n13320 ;
  assign n13322 = n6995 & n13321 ;
  assign n13324 = n3665 & ~n4490 ;
  assign n13325 = n6727 & n13324 ;
  assign n13326 = n6866 & ~n13325 ;
  assign n13323 = n4278 & n4357 ;
  assign n13327 = n13326 ^ n13323 ^ 1'b0 ;
  assign n13328 = n8730 & n8912 ;
  assign n13329 = ~n953 & n13328 ;
  assign n13330 = n3127 & n3486 ;
  assign n13331 = ( n5259 & ~n7046 ) | ( n5259 & n13330 ) | ( ~n7046 & n13330 ) ;
  assign n13332 = ( ~n98 & n13329 ) | ( ~n98 & n13331 ) | ( n13329 & n13331 ) ;
  assign n13333 = n1784 ^ n1298 ^ 1'b0 ;
  assign n13334 = n10794 & ~n13333 ;
  assign n13335 = n13334 ^ n11170 ^ n5394 ;
  assign n13336 = n8210 ^ x10 ^ 1'b0 ;
  assign n13337 = ~n1103 & n13336 ;
  assign n13338 = n4751 ^ n499 ^ 1'b0 ;
  assign n13339 = n2932 & ~n13338 ;
  assign n13340 = n13339 ^ n10883 ^ 1'b0 ;
  assign n13341 = ~n5594 & n12383 ;
  assign n13342 = n13341 ^ n101 ^ 1'b0 ;
  assign n13343 = n3884 & n4840 ;
  assign n13344 = n10031 ^ n6205 ^ 1'b0 ;
  assign n13345 = ~n2362 & n12979 ;
  assign n13346 = n13345 ^ n11007 ^ n2971 ;
  assign n13347 = n11827 & ~n13346 ;
  assign n13348 = n13344 & n13347 ;
  assign n13349 = n2674 & ~n3318 ;
  assign n13350 = n13349 ^ n12599 ^ 1'b0 ;
  assign n13351 = n13350 ^ n12053 ^ n10057 ;
  assign n13352 = ( ~n1960 & n10200 ) | ( ~n1960 & n13351 ) | ( n10200 & n13351 ) ;
  assign n13353 = n1155 & ~n7136 ;
  assign n13354 = ~n4711 & n13353 ;
  assign n13360 = n5590 ^ n4045 ^ 1'b0 ;
  assign n13361 = n2025 | n13360 ;
  assign n13362 = n13361 ^ n12441 ^ 1'b0 ;
  assign n13356 = n2733 ^ n32 ^ 1'b0 ;
  assign n13357 = n809 ^ n652 ^ 1'b0 ;
  assign n13358 = ~n2944 & n13357 ;
  assign n13359 = ~n13356 & n13358 ;
  assign n13363 = n13362 ^ n13359 ^ n4296 ;
  assign n13355 = ~n6873 & n13182 ;
  assign n13364 = n13363 ^ n13355 ^ 1'b0 ;
  assign n13365 = n12198 ^ n10568 ^ n5873 ;
  assign n13366 = n884 & n5103 ;
  assign n13367 = n13366 ^ n750 ^ 1'b0 ;
  assign n13368 = n12281 | n13367 ;
  assign n13369 = n938 | n1789 ;
  assign n13370 = n13368 & ~n13369 ;
  assign n13371 = ~n4949 & n8695 ;
  assign n13372 = n4326 & ~n13371 ;
  assign n13373 = n923 | n4579 ;
  assign n13374 = n12530 & ~n13373 ;
  assign n13375 = n205 | n10073 ;
  assign n13376 = n4607 & ~n13375 ;
  assign n13377 = n13376 ^ n4849 ^ 1'b0 ;
  assign n13378 = n13377 ^ n1409 ^ 1'b0 ;
  assign n13379 = ~n13374 & n13378 ;
  assign n13380 = n13379 ^ n3797 ^ 1'b0 ;
  assign n13381 = ~n44 & n122 ;
  assign n13382 = n13381 ^ n1777 ^ 1'b0 ;
  assign n13383 = n1389 | n13382 ;
  assign n13384 = n5761 & ~n13383 ;
  assign n13385 = ( n3211 & n11064 ) | ( n3211 & ~n13384 ) | ( n11064 & ~n13384 ) ;
  assign n13386 = n1623 & n11949 ;
  assign n13387 = ~n7657 & n13386 ;
  assign n13388 = ( n11331 & n12441 ) | ( n11331 & ~n13387 ) | ( n12441 & ~n13387 ) ;
  assign n13389 = n366 & n6909 ;
  assign n13390 = n13389 ^ n10564 ^ 1'b0 ;
  assign n13391 = n3969 ^ n1220 ^ 1'b0 ;
  assign n13392 = n4976 ^ n2065 ^ 1'b0 ;
  assign n13393 = ~n13391 & n13392 ;
  assign n13394 = n688 & ~n6239 ;
  assign n13395 = n876 & n9146 ;
  assign n13396 = n13395 ^ n5753 ^ 1'b0 ;
  assign n13397 = n1681 ^ n543 ^ 1'b0 ;
  assign n13398 = n13396 & n13397 ;
  assign n13399 = ~n4638 & n13398 ;
  assign n13400 = n2083 & ~n4074 ;
  assign n13401 = n12440 & ~n13400 ;
  assign n13402 = ~n197 & n13401 ;
  assign n13403 = n2461 & ~n3811 ;
  assign n13404 = n6700 & n13403 ;
  assign n13405 = n13402 | n13404 ;
  assign n13406 = n7554 & ~n13405 ;
  assign n13407 = n13406 ^ n6422 ^ 1'b0 ;
  assign n13408 = n8264 ^ n5033 ^ 1'b0 ;
  assign n13409 = n5484 & n6457 ;
  assign n13410 = n13409 ^ n7207 ^ 1'b0 ;
  assign n13411 = n12780 ^ n11137 ^ 1'b0 ;
  assign n13412 = n13410 & ~n13411 ;
  assign n13413 = n13412 ^ n1350 ^ 1'b0 ;
  assign n13416 = n2502 & n8097 ;
  assign n13417 = ~n6746 & n13416 ;
  assign n13414 = n9126 ^ n8474 ^ 1'b0 ;
  assign n13415 = n1783 | n13414 ;
  assign n13418 = n13417 ^ n13415 ^ n3306 ;
  assign n13419 = n10263 & ~n11409 ;
  assign n13420 = ~n6664 & n13419 ;
  assign n13421 = n13420 ^ n98 ^ 1'b0 ;
  assign n13422 = n13421 ^ n12593 ^ n10838 ;
  assign n13424 = ~n1166 & n8707 ;
  assign n13425 = n1052 & n13424 ;
  assign n13423 = ~n5147 & n6790 ;
  assign n13426 = n13425 ^ n13423 ^ n8955 ;
  assign n13427 = n11159 ^ n3593 ^ 1'b0 ;
  assign n13428 = ~n2999 & n10227 ;
  assign n13429 = ( n3801 & n6161 ) | ( n3801 & ~n13331 ) | ( n6161 & ~n13331 ) ;
  assign n13430 = n3567 & n13429 ;
  assign n13431 = n93 | n6370 ;
  assign n13432 = n13430 | n13431 ;
  assign n13433 = n9924 & n10136 ;
  assign n13434 = ~n1783 & n2790 ;
  assign n13435 = n3104 & n13434 ;
  assign n13436 = n7891 ^ n7481 ^ n5026 ;
  assign n13437 = n1569 & n1611 ;
  assign n13438 = n13437 ^ n10390 ^ n2997 ;
  assign n13439 = n2897 | n4100 ;
  assign n13440 = ( n6885 & ~n11374 ) | ( n6885 & n13439 ) | ( ~n11374 & n13439 ) ;
  assign n13441 = n13438 & n13440 ;
  assign n13442 = n13436 & n13441 ;
  assign n13443 = n9292 ^ n5897 ^ 1'b0 ;
  assign n13444 = n4104 ^ n3131 ^ 1'b0 ;
  assign n13445 = ( ~n3823 & n11701 ) | ( ~n3823 & n13444 ) | ( n11701 & n13444 ) ;
  assign n13446 = n6736 ^ n3619 ^ n3470 ;
  assign n13447 = n826 | n3384 ;
  assign n13448 = n816 & ~n13447 ;
  assign n13449 = n13446 & ~n13448 ;
  assign n13450 = n550 & n5535 ;
  assign n13451 = n13450 ^ n6304 ^ 1'b0 ;
  assign n13452 = n6027 & n9226 ;
  assign n13453 = ~n6821 & n13452 ;
  assign n13454 = ~n3003 & n13363 ;
  assign n13455 = n13454 ^ n8518 ^ 1'b0 ;
  assign n13456 = ( n3481 & n6930 ) | ( n3481 & n13455 ) | ( n6930 & n13455 ) ;
  assign n13457 = n890 | n2032 ;
  assign n13458 = n589 & ~n1772 ;
  assign n13459 = n13458 ^ n2616 ^ 1'b0 ;
  assign n13460 = n5253 & n6591 ;
  assign n13461 = n13460 ^ n9393 ^ 1'b0 ;
  assign n13462 = ( n2391 & n2403 ) | ( n2391 & ~n3687 ) | ( n2403 & ~n3687 ) ;
  assign n13463 = n4645 | n5610 ;
  assign n13464 = n10807 & n13463 ;
  assign n13465 = n13464 ^ n11073 ^ n1381 ;
  assign n13466 = n5940 & n9120 ;
  assign n13467 = n11538 & n13466 ;
  assign n13468 = n8539 ^ n5128 ^ 1'b0 ;
  assign n13469 = n947 & n13468 ;
  assign n13470 = n13469 ^ n4578 ^ 1'b0 ;
  assign n13473 = n1195 | n3571 ;
  assign n13471 = n236 & ~n9050 ;
  assign n13472 = n6657 & n13471 ;
  assign n13474 = n13473 ^ n13472 ^ 1'b0 ;
  assign n13475 = ~n11771 & n13474 ;
  assign n13476 = n352 & n5377 ;
  assign n13477 = n13476 ^ n1087 ^ n878 ;
  assign n13478 = n6533 ^ n5965 ^ n5123 ;
  assign n13479 = n6474 & ~n13478 ;
  assign n13480 = ~n5447 & n13479 ;
  assign n13481 = n13480 ^ n1348 ^ 1'b0 ;
  assign n13482 = ~n13477 & n13481 ;
  assign n13483 = ~n4818 & n13482 ;
  assign n13484 = n9217 | n13483 ;
  assign n13485 = n6647 & ~n13484 ;
  assign n13486 = n5569 | n13485 ;
  assign n13487 = n2307 | n3216 ;
  assign n13488 = n11116 & ~n13487 ;
  assign n13489 = n8362 ^ n317 ^ 1'b0 ;
  assign n13490 = n8107 ^ n7598 ^ 1'b0 ;
  assign n13495 = n1348 & ~n3636 ;
  assign n13496 = n13495 ^ n3906 ^ 1'b0 ;
  assign n13497 = ( n1645 & n7921 ) | ( n1645 & ~n13496 ) | ( n7921 & ~n13496 ) ;
  assign n13491 = n5933 ^ n2374 ^ n154 ;
  assign n13492 = ~n10073 & n13491 ;
  assign n13493 = n13492 ^ n11626 ^ 1'b0 ;
  assign n13494 = n13051 | n13493 ;
  assign n13498 = n13497 ^ n13494 ^ 1'b0 ;
  assign n13499 = n108 & n2995 ;
  assign n13500 = ~n3084 & n13499 ;
  assign n13501 = n4536 & n7599 ;
  assign n13502 = ~n7269 & n13501 ;
  assign n13503 = n9676 & ~n13502 ;
  assign n13504 = ( ~n2438 & n13500 ) | ( ~n2438 & n13503 ) | ( n13500 & n13503 ) ;
  assign n13505 = ( n44 & n1554 ) | ( n44 & n2919 ) | ( n1554 & n2919 ) ;
  assign n13506 = n3749 & n13356 ;
  assign n13507 = n6481 & n13506 ;
  assign n13508 = n13505 & ~n13507 ;
  assign n13509 = n3867 & n13507 ;
  assign n13510 = n13426 & n13509 ;
  assign n13511 = ~n10380 & n13510 ;
  assign n13512 = n13511 ^ n13335 ^ 1'b0 ;
  assign n13513 = ~n12761 & n13512 ;
  assign n13514 = n1820 ^ n523 ^ 1'b0 ;
  assign n13515 = n13514 ^ n2343 ^ 1'b0 ;
  assign n13516 = n7974 & n13515 ;
  assign n13517 = n9258 & ~n12401 ;
  assign n13518 = n1235 & n11292 ;
  assign n13519 = n13518 ^ n4465 ^ 1'b0 ;
  assign n13520 = n5997 & ~n13519 ;
  assign n13521 = n12750 ^ n6188 ^ n63 ;
  assign n13522 = n5957 ^ n4742 ^ n3120 ;
  assign n13523 = n5494 ^ n2825 ^ 1'b0 ;
  assign n13524 = n13522 & n13523 ;
  assign n13525 = n1233 | n7032 ;
  assign n13526 = n13525 ^ n10950 ^ 1'b0 ;
  assign n13527 = n1264 & n1974 ;
  assign n13528 = n13527 ^ n8007 ^ 1'b0 ;
  assign n13529 = n6052 | n13528 ;
  assign n13530 = ( n245 & ~n12821 ) | ( n245 & n13529 ) | ( ~n12821 & n13529 ) ;
  assign n13531 = ~n788 & n3637 ;
  assign n13532 = n13531 ^ n1861 ^ 1'b0 ;
  assign n13533 = n13532 ^ n9595 ^ n1507 ;
  assign n13536 = n1784 & n3116 ;
  assign n13537 = n13536 ^ n969 ^ 1'b0 ;
  assign n13534 = n704 | n6551 ;
  assign n13535 = ~n7315 & n13534 ;
  assign n13538 = n13537 ^ n13535 ^ n2476 ;
  assign n13539 = n40 & ~n2418 ;
  assign n13540 = ( ~n216 & n570 ) | ( ~n216 & n13539 ) | ( n570 & n13539 ) ;
  assign n13541 = n13540 ^ n5359 ^ 1'b0 ;
  assign n13542 = ~n645 & n6014 ;
  assign n13543 = n612 & ~n6149 ;
  assign n13544 = n13543 ^ n11345 ^ n1623 ;
  assign n13545 = n8869 ^ n3973 ^ 1'b0 ;
  assign n13546 = n1822 & ~n3964 ;
  assign n13547 = ~n7787 & n13546 ;
  assign n13548 = n7101 | n11172 ;
  assign n13549 = n306 & n7499 ;
  assign n13550 = ( n754 & n1616 ) | ( n754 & ~n1813 ) | ( n1616 & ~n1813 ) ;
  assign n13551 = n800 & ~n6641 ;
  assign n13552 = n13550 & n13551 ;
  assign n13553 = n6144 & n10934 ;
  assign n13554 = ~n7153 & n13553 ;
  assign n13555 = n4854 & ~n5122 ;
  assign n13556 = n10658 | n13555 ;
  assign n13557 = n12317 ^ n2902 ^ 1'b0 ;
  assign n13558 = ~n7931 & n11741 ;
  assign n13559 = n13558 ^ n5521 ^ 1'b0 ;
  assign n13560 = n13559 ^ n6105 ^ 1'b0 ;
  assign n13561 = n1661 | n3105 ;
  assign n13562 = n6345 & ~n13248 ;
  assign n13563 = n13562 ^ n543 ^ 1'b0 ;
  assign n13564 = n9194 & ~n10838 ;
  assign n13565 = n13564 ^ n9779 ^ 1'b0 ;
  assign n13566 = n177 & ~n7270 ;
  assign n13567 = n117 & n2457 ;
  assign n13568 = ( ~n864 & n13075 ) | ( ~n864 & n13567 ) | ( n13075 & n13567 ) ;
  assign n13569 = n13566 | n13568 ;
  assign n13570 = n6040 & n9781 ;
  assign n13571 = n3575 & n13570 ;
  assign n13572 = n13571 ^ n10481 ^ 1'b0 ;
  assign n13573 = n4377 ^ n411 ^ 1'b0 ;
  assign n13574 = n3898 & ~n13573 ;
  assign n13577 = n4877 | n7010 ;
  assign n13575 = n1209 & ~n1527 ;
  assign n13576 = n13575 ^ n12020 ^ 1'b0 ;
  assign n13578 = n13577 ^ n13576 ^ n6699 ;
  assign n13579 = n11680 ^ n1722 ^ 1'b0 ;
  assign n13580 = n6332 ^ n5852 ^ 1'b0 ;
  assign n13581 = n1784 & ~n13580 ;
  assign n13582 = ~n13579 & n13581 ;
  assign n13583 = n236 & n10031 ;
  assign n13584 = n1435 | n2815 ;
  assign n13585 = ( n1129 & ~n10130 ) | ( n1129 & n13584 ) | ( ~n10130 & n13584 ) ;
  assign n13586 = n10594 ^ n8073 ^ 1'b0 ;
  assign n13587 = n443 ^ n37 ^ 1'b0 ;
  assign n13588 = n596 | n4077 ;
  assign n13589 = n682 | n13588 ;
  assign n13590 = ~n7780 & n13589 ;
  assign n13591 = n13590 ^ n2330 ^ 1'b0 ;
  assign n13592 = ~n272 & n13591 ;
  assign n13593 = n13587 & n13592 ;
  assign n13594 = n10323 & n11114 ;
  assign n13595 = n151 & n13594 ;
  assign n13596 = n263 | n2337 ;
  assign n13597 = n13596 ^ n1874 ^ 1'b0 ;
  assign n13598 = n2352 ^ n1489 ^ 1'b0 ;
  assign n13599 = ~n1944 & n13598 ;
  assign n13600 = n11505 & n13599 ;
  assign n13601 = n4761 & ~n13600 ;
  assign n13602 = ~n8242 & n13601 ;
  assign n13603 = n13602 ^ n13387 ^ n1135 ;
  assign n13604 = n696 & ~n946 ;
  assign n13605 = n3850 & n13604 ;
  assign n13606 = n3148 & n4803 ;
  assign n13607 = n13605 & n13606 ;
  assign n13608 = n11782 ^ n2769 ^ 1'b0 ;
  assign n13609 = n8919 ^ n2558 ^ 1'b0 ;
  assign n13610 = n5847 ^ n1721 ^ n611 ;
  assign n13611 = ~n5667 & n13610 ;
  assign n13612 = n6549 ^ n3304 ^ 1'b0 ;
  assign n13613 = n8099 & n13612 ;
  assign n13614 = ~n13611 & n13613 ;
  assign n13615 = ~n7026 & n7254 ;
  assign n13616 = ~n3020 & n13615 ;
  assign n13617 = n2756 & ~n13616 ;
  assign n13618 = n10361 ^ n6336 ^ 1'b0 ;
  assign n13619 = n1026 & ~n13618 ;
  assign n13620 = n1563 & ~n7094 ;
  assign n13621 = ~n1560 & n5265 ;
  assign n13622 = n9849 & ~n13621 ;
  assign n13623 = ~n5436 & n13622 ;
  assign n13624 = n13623 ^ n12379 ^ 1'b0 ;
  assign n13625 = n13620 | n13624 ;
  assign n13626 = n9546 ^ n4305 ^ 1'b0 ;
  assign n13627 = ( n1155 & n3087 ) | ( n1155 & ~n9993 ) | ( n3087 & ~n9993 ) ;
  assign n13628 = n11923 & ~n13627 ;
  assign n13629 = n13628 ^ n13558 ^ 1'b0 ;
  assign n13630 = n9448 ^ n2588 ^ 1'b0 ;
  assign n13631 = ~n1389 & n13630 ;
  assign n13632 = n13631 ^ n13315 ^ 1'b0 ;
  assign n13633 = n13632 ^ n13155 ^ 1'b0 ;
  assign n13634 = n4717 | n13633 ;
  assign n13635 = n2092 & n5128 ;
  assign n13636 = ~n1210 & n13635 ;
  assign n13637 = n9308 & n13636 ;
  assign n13638 = n4131 & n8626 ;
  assign n13639 = n318 & ~n13638 ;
  assign n13640 = n13639 ^ n1285 ^ 1'b0 ;
  assign n13641 = n9924 ^ n3531 ^ 1'b0 ;
  assign n13642 = n13640 & ~n13641 ;
  assign n13643 = n3638 ^ n2250 ^ 1'b0 ;
  assign n13644 = n13643 ^ n3307 ^ n2517 ;
  assign n13645 = ( n7536 & ~n8560 ) | ( n7536 & n12826 ) | ( ~n8560 & n12826 ) ;
  assign n13646 = ( n588 & ~n6041 ) | ( n588 & n13645 ) | ( ~n6041 & n13645 ) ;
  assign n13647 = ~n13644 & n13646 ;
  assign n13648 = n13647 ^ n11633 ^ 1'b0 ;
  assign n13649 = ( n4678 & n5444 ) | ( n4678 & n7790 ) | ( n5444 & n7790 ) ;
  assign n13650 = n3884 | n5734 ;
  assign n13651 = n13650 ^ n11233 ^ n5327 ;
  assign n13652 = n3221 ^ n2694 ^ 1'b0 ;
  assign n13653 = n4260 & n13652 ;
  assign n13654 = n356 & ~n13653 ;
  assign n13655 = n6670 & ~n11113 ;
  assign n13656 = n13655 ^ n8697 ^ 1'b0 ;
  assign n13657 = n3183 & n13656 ;
  assign n13658 = n13657 ^ n12220 ^ 1'b0 ;
  assign n13659 = n1294 ^ n583 ^ 1'b0 ;
  assign n13660 = n6280 | n13659 ;
  assign n13661 = n5626 & n9432 ;
  assign n13663 = n7917 ^ n1650 ^ n1305 ;
  assign n13664 = n7927 | n13663 ;
  assign n13662 = ~n4404 & n4654 ;
  assign n13665 = n13664 ^ n13662 ^ 1'b0 ;
  assign n13666 = n11779 ^ n7373 ^ 1'b0 ;
  assign n13667 = n1475 & n13666 ;
  assign n13668 = n7432 ^ n3256 ^ 1'b0 ;
  assign n13670 = n7380 ^ n6346 ^ n350 ;
  assign n13669 = n7047 & ~n12211 ;
  assign n13671 = n13670 ^ n13669 ^ 1'b0 ;
  assign n13672 = ( n2594 & ~n5803 ) | ( n2594 & n8768 ) | ( ~n5803 & n8768 ) ;
  assign n13673 = n13672 ^ n10010 ^ 1'b0 ;
  assign n13675 = ~n3541 & n7584 ;
  assign n13676 = n13675 ^ n1068 ^ 1'b0 ;
  assign n13674 = n9688 & ~n11635 ;
  assign n13677 = n13676 ^ n13674 ^ 1'b0 ;
  assign n13678 = n13677 ^ n13298 ^ 1'b0 ;
  assign n13679 = n1409 & ~n1533 ;
  assign n13680 = ~n3242 & n7150 ;
  assign n13681 = ~n7089 & n13680 ;
  assign n13682 = n13681 ^ n2568 ^ 1'b0 ;
  assign n13683 = n13682 ^ n4679 ^ 1'b0 ;
  assign n13684 = n13683 ^ n3784 ^ n2084 ;
  assign n13685 = n1745 & ~n5691 ;
  assign n13686 = n13685 ^ n6811 ^ 1'b0 ;
  assign n13687 = n13686 ^ n594 ^ 1'b0 ;
  assign n13688 = n13684 & ~n13687 ;
  assign n13689 = n3715 ^ n1213 ^ 1'b0 ;
  assign n13690 = ~n1895 & n4818 ;
  assign n13691 = n13690 ^ n209 ^ 1'b0 ;
  assign n13692 = ~n13689 & n13691 ;
  assign n13693 = n1319 & ~n4345 ;
  assign n13694 = n13692 & ~n13693 ;
  assign n13697 = n2425 ^ n1979 ^ 1'b0 ;
  assign n13695 = ( ~n905 & n2605 ) | ( ~n905 & n11921 ) | ( n2605 & n11921 ) ;
  assign n13696 = n126 & ~n13695 ;
  assign n13698 = n13697 ^ n13696 ^ 1'b0 ;
  assign n13699 = n7788 ^ n3482 ^ 1'b0 ;
  assign n13700 = n5151 ^ n534 ^ 1'b0 ;
  assign n13701 = n13161 & ~n13700 ;
  assign n13702 = ~n4769 & n13701 ;
  assign n13703 = n6513 ^ n4163 ^ n3124 ;
  assign n13704 = n2648 & ~n13703 ;
  assign n13705 = n13704 ^ n272 ^ 1'b0 ;
  assign n13706 = ( ~n462 & n9235 ) | ( ~n462 & n13705 ) | ( n9235 & n13705 ) ;
  assign n13711 = n8145 & n12435 ;
  assign n13712 = n713 & n13711 ;
  assign n13707 = n4923 | n9026 ;
  assign n13708 = ( n1625 & n6684 ) | ( n1625 & n13707 ) | ( n6684 & n13707 ) ;
  assign n13709 = n2497 & ~n13708 ;
  assign n13710 = n8655 & n13709 ;
  assign n13713 = n13712 ^ n13710 ^ n9501 ;
  assign n13714 = ~n8171 & n11009 ;
  assign n13716 = n1170 & n7495 ;
  assign n13715 = ( n1368 & n7400 ) | ( n1368 & ~n11859 ) | ( n7400 & ~n11859 ) ;
  assign n13717 = n13716 ^ n13715 ^ 1'b0 ;
  assign n13718 = n13717 ^ n7242 ^ 1'b0 ;
  assign n13719 = ~n6088 & n13718 ;
  assign n13720 = n734 | n13516 ;
  assign n13724 = n4168 | n5312 ;
  assign n13725 = n4640 | n13724 ;
  assign n13726 = ~n10579 & n13725 ;
  assign n13721 = n5970 & ~n8919 ;
  assign n13722 = n1744 | n2549 ;
  assign n13723 = n13721 | n13722 ;
  assign n13727 = n13726 ^ n13723 ^ 1'b0 ;
  assign n13728 = n59 | n893 ;
  assign n13729 = n228 & ~n13728 ;
  assign n13730 = n607 | n2695 ;
  assign n13731 = ~n13729 & n13730 ;
  assign n13732 = n13731 ^ n5866 ^ 1'b0 ;
  assign n13733 = n13732 ^ n6947 ^ 1'b0 ;
  assign n13734 = ~n2339 & n6142 ;
  assign n13735 = n13734 ^ n11458 ^ 1'b0 ;
  assign n13736 = ( n74 & n3635 ) | ( n74 & ~n3846 ) | ( n3635 & ~n3846 ) ;
  assign n13740 = ~n8047 & n8537 ;
  assign n13737 = n9011 ^ n4068 ^ n921 ;
  assign n13738 = ~n2129 & n13737 ;
  assign n13739 = n13738 ^ n2740 ^ 1'b0 ;
  assign n13741 = n13740 ^ n13739 ^ 1'b0 ;
  assign n13742 = ~n6805 & n13546 ;
  assign n13743 = n13742 ^ n5841 ^ 1'b0 ;
  assign n13744 = n1025 & ~n6411 ;
  assign n13745 = n13744 ^ n411 ^ 1'b0 ;
  assign n13746 = n13745 ^ n1374 ^ 1'b0 ;
  assign n13747 = n13743 | n13746 ;
  assign n13748 = n10375 ^ n2375 ^ 1'b0 ;
  assign n13749 = n5804 ^ n4264 ^ 1'b0 ;
  assign n13750 = n5389 & n10715 ;
  assign n13751 = n5180 & n13750 ;
  assign n13754 = ~n2101 & n9029 ;
  assign n13752 = n2416 & n5951 ;
  assign n13753 = n881 & n13752 ;
  assign n13755 = n13754 ^ n13753 ^ 1'b0 ;
  assign n13756 = n13751 | n13755 ;
  assign n13757 = n11660 & ~n13756 ;
  assign n13758 = n3263 & ~n8166 ;
  assign n13759 = n8198 | n13758 ;
  assign n13760 = n11057 | n13759 ;
  assign n13761 = n5438 ^ n2115 ^ 1'b0 ;
  assign n13762 = ~n2831 & n10388 ;
  assign n13763 = n216 & ~n3271 ;
  assign n13764 = n13151 ^ n6156 ^ n4105 ;
  assign n13765 = n6805 & ~n13764 ;
  assign n13766 = n13763 & n13765 ;
  assign n13767 = n2712 | n13766 ;
  assign n13768 = n13767 ^ n6895 ^ 1'b0 ;
  assign n13769 = n4457 & n13496 ;
  assign n13770 = n13769 ^ n10534 ^ n7807 ;
  assign n13771 = n977 & ~n4078 ;
  assign n13772 = n9702 ^ n4250 ^ n38 ;
  assign n13773 = n209 & n7954 ;
  assign n13774 = n13772 & n13773 ;
  assign n13775 = n13771 | n13774 ;
  assign n13776 = n9779 ^ n250 ^ 1'b0 ;
  assign n13777 = n10072 & n13776 ;
  assign n13778 = n174 | n2147 ;
  assign n13779 = n8070 ^ n1572 ^ 1'b0 ;
  assign n13780 = n1351 | n13779 ;
  assign n13781 = n7254 & ~n13780 ;
  assign n13782 = ~n13086 & n13781 ;
  assign n13783 = ( n4356 & n13778 ) | ( n4356 & ~n13782 ) | ( n13778 & ~n13782 ) ;
  assign n13784 = n12658 ^ n1809 ^ 1'b0 ;
  assign n13785 = n985 & ~n13784 ;
  assign n13786 = n2537 ^ n20 ^ 1'b0 ;
  assign n13787 = ~n2650 & n13786 ;
  assign n13788 = n12163 & n13787 ;
  assign n13789 = ~n10068 & n13788 ;
  assign n13790 = n7035 & ~n13789 ;
  assign n13791 = ~n1177 & n13790 ;
  assign n13803 = n833 | n8218 ;
  assign n13804 = n10206 & ~n13803 ;
  assign n13792 = n4216 | n5258 ;
  assign n13795 = n3708 & ~n7842 ;
  assign n13794 = n958 & n3508 ;
  assign n13796 = n13795 ^ n13794 ^ 1'b0 ;
  assign n13793 = n834 | n3571 ;
  assign n13797 = n13796 ^ n13793 ^ 1'b0 ;
  assign n13798 = n7338 & n13797 ;
  assign n13799 = ~n987 & n7245 ;
  assign n13800 = n13799 ^ n8177 ^ 1'b0 ;
  assign n13801 = ~n13798 & n13800 ;
  assign n13802 = n13792 & n13801 ;
  assign n13805 = n13804 ^ n13802 ^ 1'b0 ;
  assign n13806 = ~n13791 & n13805 ;
  assign n13807 = ~n10124 & n13737 ;
  assign n13808 = n13807 ^ n11302 ^ 1'b0 ;
  assign n13809 = ~n7115 & n8347 ;
  assign n13810 = n13809 ^ n1695 ^ 1'b0 ;
  assign n13811 = n63 & ~n4612 ;
  assign n13812 = n13811 ^ n7069 ^ n780 ;
  assign n13813 = n3666 & n10719 ;
  assign n13814 = n11135 ^ n1319 ^ 1'b0 ;
  assign n13815 = n13814 ^ n2058 ^ 1'b0 ;
  assign n13816 = n8655 | n13815 ;
  assign n13817 = n3336 | n13816 ;
  assign n13818 = n9156 ^ n4116 ^ 1'b0 ;
  assign n13819 = ~n5129 & n5740 ;
  assign n13820 = n2226 & ~n7284 ;
  assign n13821 = n13820 ^ n12541 ^ 1'b0 ;
  assign n13822 = n576 | n1653 ;
  assign n13823 = n13822 ^ n5062 ^ 1'b0 ;
  assign n13824 = n1029 ^ n276 ^ 1'b0 ;
  assign n13825 = n13823 | n13824 ;
  assign n13826 = n13825 ^ n4376 ^ 1'b0 ;
  assign n13827 = n2432 & ~n13826 ;
  assign n13828 = n13827 ^ n3357 ^ 1'b0 ;
  assign n13829 = n13821 & n13828 ;
  assign n13831 = n7378 & ~n9734 ;
  assign n13832 = ~n1153 & n13831 ;
  assign n13833 = n11646 ^ n5635 ^ 1'b0 ;
  assign n13834 = n13832 | n13833 ;
  assign n13835 = n3530 ^ n2159 ^ 1'b0 ;
  assign n13836 = n3688 | n13835 ;
  assign n13837 = n13836 ^ n1848 ^ 1'b0 ;
  assign n13838 = n11223 & ~n13837 ;
  assign n13839 = n2515 & n13838 ;
  assign n13840 = ~n3303 & n13839 ;
  assign n13841 = n13834 & n13840 ;
  assign n13830 = ~n2761 & n8551 ;
  assign n13842 = n13841 ^ n13830 ^ 1'b0 ;
  assign n13844 = n5350 ^ x10 ^ 1'b0 ;
  assign n13843 = n1586 & n4469 ;
  assign n13845 = n13844 ^ n13843 ^ 1'b0 ;
  assign n13846 = ~n1248 & n5766 ;
  assign n13847 = n2745 & n4290 ;
  assign n13848 = n13847 ^ n2070 ^ 1'b0 ;
  assign n13849 = n13848 ^ n13845 ^ n11385 ;
  assign n13850 = n4693 | n9074 ;
  assign n13851 = n3051 | n5093 ;
  assign n13852 = n13851 ^ n1668 ^ 1'b0 ;
  assign n13853 = n6039 | n13852 ;
  assign n13854 = n63 | n2041 ;
  assign n13855 = n8907 ^ n3214 ^ n1082 ;
  assign n13856 = n12403 ^ n3069 ^ 1'b0 ;
  assign n13857 = ~n13855 & n13856 ;
  assign n13858 = ~n13854 & n13857 ;
  assign n13859 = n13125 ^ n1151 ^ 1'b0 ;
  assign n13860 = ( n4976 & n5915 ) | ( n4976 & n7133 ) | ( n5915 & n7133 ) ;
  assign n13861 = n4743 & ~n13860 ;
  assign n13862 = n13861 ^ n5251 ^ 1'b0 ;
  assign n13863 = n3542 ^ n2556 ^ 1'b0 ;
  assign n13864 = n6477 & n7746 ;
  assign n13865 = ~n13863 & n13864 ;
  assign n13866 = n8441 ^ n2213 ^ 1'b0 ;
  assign n13867 = n13865 | n13866 ;
  assign n13868 = n13867 ^ n8727 ^ 1'b0 ;
  assign n13869 = n8906 ^ n922 ^ 1'b0 ;
  assign n13870 = n13868 & ~n13869 ;
  assign n13871 = n9361 ^ n8882 ^ n7790 ;
  assign n13872 = n2925 & n8157 ;
  assign n13873 = ~n13871 & n13872 ;
  assign n13874 = n596 & n2412 ;
  assign n13875 = ~n2412 & n13874 ;
  assign n13876 = ( n933 & n7190 ) | ( n933 & ~n10008 ) | ( n7190 & ~n10008 ) ;
  assign n13877 = n13875 & ~n13876 ;
  assign n13878 = ~n6526 & n13877 ;
  assign n13879 = n2118 & ~n10054 ;
  assign n13880 = n6965 ^ n3027 ^ 1'b0 ;
  assign n13881 = n13879 & n13880 ;
  assign n13882 = n13881 ^ n3040 ^ 1'b0 ;
  assign n13883 = n543 & ~n13882 ;
  assign n13884 = ~n10362 & n13883 ;
  assign n13885 = n10433 & n12748 ;
  assign n13886 = n13885 ^ n12509 ^ 1'b0 ;
  assign n13887 = n43 | n13886 ;
  assign n13888 = n4186 | n8382 ;
  assign n13889 = n13888 ^ n2992 ^ 1'b0 ;
  assign n13890 = n13889 ^ n1865 ^ 1'b0 ;
  assign n13891 = n13890 ^ n8741 ^ 1'b0 ;
  assign n13892 = n4743 & n11458 ;
  assign n13893 = n13891 & n13892 ;
  assign n13894 = n2441 & ~n13893 ;
  assign n13895 = n13894 ^ n12305 ^ 1'b0 ;
  assign n13897 = n2036 | n3603 ;
  assign n13898 = n3603 & ~n13897 ;
  assign n13899 = n13898 ^ n8465 ^ n7358 ;
  assign n13896 = ( n79 & ~n6924 ) | ( n79 & n11249 ) | ( ~n6924 & n11249 ) ;
  assign n13900 = n13899 ^ n13896 ^ n1766 ;
  assign n13901 = ~n3869 & n12056 ;
  assign n13902 = n13901 ^ n11044 ^ 1'b0 ;
  assign n13903 = n37 & n7128 ;
  assign n13904 = n13751 ^ n2321 ^ 1'b0 ;
  assign n13905 = n5453 ^ n2226 ^ 1'b0 ;
  assign n13906 = n13905 ^ n4477 ^ 1'b0 ;
  assign n13907 = n13904 & n13906 ;
  assign n13908 = n3205 & ~n4503 ;
  assign n13909 = n2143 & n13908 ;
  assign n13910 = n5606 | n13909 ;
  assign n13911 = n260 & ~n13910 ;
  assign n13912 = n7028 | n13911 ;
  assign n13913 = n13912 ^ n3916 ^ 1'b0 ;
  assign n13914 = n2125 ^ n916 ^ 1'b0 ;
  assign n13915 = n159 | n8205 ;
  assign n13916 = n9484 & ~n13915 ;
  assign n13917 = n4741 | n6036 ;
  assign n13918 = ( n4896 & n7147 ) | ( n4896 & ~n10062 ) | ( n7147 & ~n10062 ) ;
  assign n13919 = ( ~n3465 & n13917 ) | ( ~n3465 & n13918 ) | ( n13917 & n13918 ) ;
  assign n13920 = n8076 | n13919 ;
  assign n13925 = n1838 | n8404 ;
  assign n13926 = n13925 ^ n4060 ^ 1'b0 ;
  assign n13927 = n3975 ^ n3600 ^ 1'b0 ;
  assign n13928 = n13926 & ~n13927 ;
  assign n13929 = n1856 | n13928 ;
  assign n13930 = n13929 ^ n517 ^ 1'b0 ;
  assign n13921 = ( n3361 & n5750 ) | ( n3361 & n7638 ) | ( n5750 & n7638 ) ;
  assign n13922 = n13921 ^ n1340 ^ 1'b0 ;
  assign n13923 = ~x10 & n13922 ;
  assign n13924 = n7052 | n13923 ;
  assign n13931 = n13930 ^ n13924 ^ 1'b0 ;
  assign n13932 = n7646 ^ n2804 ^ n37 ;
  assign n13933 = n13932 ^ n2060 ^ 1'b0 ;
  assign n13934 = n13933 ^ n12476 ^ 1'b0 ;
  assign n13939 = n5584 ^ n5457 ^ 1'b0 ;
  assign n13940 = ( ~n6809 & n10263 ) | ( ~n6809 & n13939 ) | ( n10263 & n13939 ) ;
  assign n13935 = n9015 ^ x3 ^ 1'b0 ;
  assign n13936 = n2348 & ~n13935 ;
  assign n13937 = ( n1307 & n7636 ) | ( n1307 & ~n13936 ) | ( n7636 & ~n13936 ) ;
  assign n13938 = n13937 ^ n2270 ^ 1'b0 ;
  assign n13941 = n13940 ^ n13938 ^ n2414 ;
  assign n13942 = ( n4169 & n4273 ) | ( n4169 & n11899 ) | ( n4273 & n11899 ) ;
  assign n13943 = ( n906 & ~n3029 ) | ( n906 & n3886 ) | ( ~n3029 & n3886 ) ;
  assign n13944 = n13943 ^ n7294 ^ 1'b0 ;
  assign n13945 = ~n1690 & n13944 ;
  assign n13946 = n13945 ^ n5197 ^ n3717 ;
  assign n13947 = n1579 & ~n3968 ;
  assign n13948 = n3097 | n6514 ;
  assign n13949 = n7449 | n13948 ;
  assign n13950 = ( ~n3221 & n13947 ) | ( ~n3221 & n13949 ) | ( n13947 & n13949 ) ;
  assign n13951 = ( n7067 & n13946 ) | ( n7067 & n13950 ) | ( n13946 & n13950 ) ;
  assign n13952 = n10597 ^ n4495 ^ n250 ;
  assign n13953 = ( n1463 & n9238 ) | ( n1463 & n13952 ) | ( n9238 & n13952 ) ;
  assign n13954 = n2330 | n13953 ;
  assign n13955 = n7716 ^ n2679 ^ 1'b0 ;
  assign n13956 = n7880 | n13955 ;
  assign n13957 = n9093 | n13956 ;
  assign n13958 = n3201 ^ n2785 ^ 1'b0 ;
  assign n13959 = n3897 & n13958 ;
  assign n13960 = n13959 ^ n5986 ^ 1'b0 ;
  assign n13961 = n3603 | n13960 ;
  assign n13962 = n13957 | n13961 ;
  assign n13963 = ~n3189 & n9267 ;
  assign n13964 = n368 & n3811 ;
  assign n13965 = n1686 | n13964 ;
  assign n13967 = n3622 & n4059 ;
  assign n13968 = n13967 ^ n5423 ^ 1'b0 ;
  assign n13966 = n4495 & n8083 ;
  assign n13969 = n13968 ^ n13966 ^ 1'b0 ;
  assign n13970 = n13969 ^ n12833 ^ n9666 ;
  assign n13971 = n8117 ^ n5418 ^ 1'b0 ;
  assign n13972 = ~n923 & n13971 ;
  assign n13973 = ( n4780 & ~n12237 ) | ( n4780 & n13972 ) | ( ~n12237 & n13972 ) ;
  assign n13974 = n7335 ^ n1264 ^ 1'b0 ;
  assign n13975 = n13974 ^ n6394 ^ 1'b0 ;
  assign n13976 = n13973 & n13975 ;
  assign n13977 = n11331 ^ n5977 ^ n3423 ;
  assign n13978 = n13977 ^ n5937 ^ 1'b0 ;
  assign n13979 = ~n13976 & n13978 ;
  assign n13980 = n4113 ^ n2435 ^ 1'b0 ;
  assign n13981 = ~n4151 & n13980 ;
  assign n13982 = n13981 ^ n10543 ^ 1'b0 ;
  assign n13983 = n2810 & n6221 ;
  assign n13984 = n13983 ^ n6541 ^ 1'b0 ;
  assign n13985 = ~n2549 & n13984 ;
  assign n13986 = n13985 ^ n10451 ^ 1'b0 ;
  assign n13987 = n6052 | n11445 ;
  assign n13988 = n13986 | n13987 ;
  assign n13989 = n4177 & ~n13988 ;
  assign n13990 = ~n11321 & n13989 ;
  assign n13991 = n9563 ^ n374 ^ 1'b0 ;
  assign n13992 = n7895 ^ n5506 ^ n1909 ;
  assign n13993 = ( n4948 & n6352 ) | ( n4948 & n13992 ) | ( n6352 & n13992 ) ;
  assign n13994 = n4569 & n4685 ;
  assign n13995 = n13993 & n13994 ;
  assign n13996 = n8953 ^ n1542 ^ 1'b0 ;
  assign n13997 = n6682 & n13996 ;
  assign n13998 = n13997 ^ n5100 ^ 1'b0 ;
  assign n13999 = ~n12087 & n13998 ;
  assign n14000 = n6241 ^ n5607 ^ 1'b0 ;
  assign n14001 = n390 & n14000 ;
  assign n14002 = n6620 ^ n2048 ^ n1478 ;
  assign n14003 = n1096 & n2053 ;
  assign n14004 = n14002 & n14003 ;
  assign n14005 = n14004 ^ n11664 ^ 1'b0 ;
  assign n14006 = n9168 ^ n7314 ^ 1'b0 ;
  assign n14007 = n1418 & n14006 ;
  assign n14008 = n1091 & ~n2631 ;
  assign n14009 = n14008 ^ n5214 ^ 1'b0 ;
  assign n14010 = n1276 ^ n93 ^ 1'b0 ;
  assign n14011 = n14010 ^ n9853 ^ n2476 ;
  assign n14012 = n14011 ^ n8133 ^ 1'b0 ;
  assign n14013 = n3457 & ~n14012 ;
  assign n14014 = n14013 ^ n6212 ^ 1'b0 ;
  assign n14016 = n7055 ^ n1436 ^ 1'b0 ;
  assign n14015 = ~n7140 & n10806 ;
  assign n14017 = n14016 ^ n14015 ^ 1'b0 ;
  assign n14018 = n8912 & ~n14017 ;
  assign n14019 = n12761 & n14018 ;
  assign n14022 = n8842 & n11777 ;
  assign n14020 = n2322 | n3093 ;
  assign n14021 = n10192 | n14020 ;
  assign n14023 = n14022 ^ n14021 ^ 1'b0 ;
  assign n14024 = ( n7039 & n10329 ) | ( n7039 & n14023 ) | ( n10329 & n14023 ) ;
  assign n14030 = n4263 ^ n1721 ^ 1'b0 ;
  assign n14031 = n3333 ^ n2497 ^ 1'b0 ;
  assign n14032 = ~n14030 & n14031 ;
  assign n14028 = n1400 & n6102 ;
  assign n14029 = n5124 & n14028 ;
  assign n14025 = n711 & ~n6275 ;
  assign n14026 = n14025 ^ n4688 ^ 1'b0 ;
  assign n14027 = ~n12736 & n14026 ;
  assign n14033 = n14032 ^ n14029 ^ n14027 ;
  assign n14034 = n6808 | n13710 ;
  assign n14035 = n14033 & ~n14034 ;
  assign n14036 = n6993 ^ n4159 ^ 1'b0 ;
  assign n14037 = n203 & n14036 ;
  assign n14039 = n4380 & ~n4541 ;
  assign n14040 = n14039 ^ n5374 ^ 1'b0 ;
  assign n14041 = n14040 ^ n4430 ^ 1'b0 ;
  assign n14042 = n3923 & n14041 ;
  assign n14038 = n145 & ~n5017 ;
  assign n14043 = n14042 ^ n14038 ^ 1'b0 ;
  assign n14044 = n5511 ^ n4728 ^ 1'b0 ;
  assign n14045 = n7016 & ~n14044 ;
  assign n14046 = n6229 ^ n4186 ^ 1'b0 ;
  assign n14047 = n14045 & ~n14046 ;
  assign n14048 = ( n1883 & n8552 ) | ( n1883 & ~n9339 ) | ( n8552 & ~n9339 ) ;
  assign n14049 = n14039 ^ n4109 ^ n790 ;
  assign n14052 = ( n961 & n5055 ) | ( n961 & ~n5725 ) | ( n5055 & ~n5725 ) ;
  assign n14050 = n8389 & n11347 ;
  assign n14051 = n14050 ^ n1138 ^ 1'b0 ;
  assign n14053 = n14052 ^ n14051 ^ 1'b0 ;
  assign n14054 = n14049 | n14053 ;
  assign n14055 = ( n5632 & n8074 ) | ( n5632 & ~n11796 ) | ( n8074 & ~n11796 ) ;
  assign n14056 = ~n733 & n3750 ;
  assign n14057 = n14056 ^ n2813 ^ 1'b0 ;
  assign n14058 = n1000 & ~n5234 ;
  assign n14059 = n14057 & n14058 ;
  assign n14060 = n656 | n14059 ;
  assign n14061 = n14060 ^ n3761 ^ 1'b0 ;
  assign n14062 = n13780 | n14061 ;
  assign n14063 = n14055 | n14062 ;
  assign n14064 = n3634 ^ n2108 ^ n502 ;
  assign n14065 = ~n8108 & n14064 ;
  assign n14066 = ( n451 & n5273 ) | ( n451 & n8555 ) | ( n5273 & n8555 ) ;
  assign n14067 = n3720 & ~n6205 ;
  assign n14068 = ( n8815 & n14066 ) | ( n8815 & n14067 ) | ( n14066 & n14067 ) ;
  assign n14077 = n4769 ^ n2712 ^ 1'b0 ;
  assign n14069 = n1383 & ~n1921 ;
  assign n14070 = n2324 ^ n484 ^ 1'b0 ;
  assign n14071 = n1089 & ~n14070 ;
  assign n14072 = n6120 & n14071 ;
  assign n14073 = ~n14069 & n14072 ;
  assign n14074 = n12140 ^ n890 ^ 1'b0 ;
  assign n14075 = ( n4028 & ~n14073 ) | ( n4028 & n14074 ) | ( ~n14073 & n14074 ) ;
  assign n14076 = n9318 | n14075 ;
  assign n14078 = n14077 ^ n14076 ^ n4696 ;
  assign n14079 = n6976 & n14078 ;
  assign n14080 = n14079 ^ n13111 ^ 1'b0 ;
  assign n14082 = n6745 ^ n2745 ^ n321 ;
  assign n14083 = n14082 ^ n8369 ^ 1'b0 ;
  assign n14081 = ~n4892 & n7530 ;
  assign n14084 = n14083 ^ n14081 ^ 1'b0 ;
  assign n14085 = n2422 | n9210 ;
  assign n14086 = n14085 ^ n4503 ^ 1'b0 ;
  assign n14087 = n14084 | n14086 ;
  assign n14088 = n9110 | n14087 ;
  assign n14089 = n10657 ^ n6510 ^ 1'b0 ;
  assign n14090 = n4271 ^ n2223 ^ 1'b0 ;
  assign n14091 = n14089 & n14090 ;
  assign n14092 = n2807 | n3984 ;
  assign n14093 = n6308 & ~n14092 ;
  assign n14094 = n5656 & ~n14093 ;
  assign n14097 = n5162 ^ n4222 ^ n3282 ;
  assign n14095 = n3824 & ~n10044 ;
  assign n14096 = ~n13953 & n14095 ;
  assign n14098 = n14097 ^ n14096 ^ 1'b0 ;
  assign n14099 = ( n9713 & n11341 ) | ( n9713 & ~n12371 ) | ( n11341 & ~n12371 ) ;
  assign n14100 = n14099 ^ n13762 ^ 1'b0 ;
  assign n14102 = n1156 & ~n2864 ;
  assign n14101 = n569 & n3255 ;
  assign n14103 = n14102 ^ n14101 ^ n13987 ;
  assign n14104 = n8901 | n14103 ;
  assign n14105 = n3406 ^ n1841 ^ 1'b0 ;
  assign n14106 = n4599 & ~n14105 ;
  assign n14107 = n14106 ^ n403 ^ 1'b0 ;
  assign n14108 = n1384 & n1817 ;
  assign n14109 = ~n14107 & n14108 ;
  assign n14110 = n6272 & ~n12124 ;
  assign n14111 = ~n1081 & n2830 ;
  assign n14112 = ~n2569 & n14111 ;
  assign n14117 = n3833 ^ n572 ^ 1'b0 ;
  assign n14118 = n3330 & ~n14117 ;
  assign n14119 = n14118 ^ n962 ^ 1'b0 ;
  assign n14113 = n7186 ^ n6475 ^ 1'b0 ;
  assign n14114 = n2289 & ~n14113 ;
  assign n14115 = n7920 & n14114 ;
  assign n14116 = n14115 ^ n6189 ^ 1'b0 ;
  assign n14120 = n14119 ^ n14116 ^ 1'b0 ;
  assign n14121 = n14112 & ~n14120 ;
  assign n14123 = ~n8330 & n10711 ;
  assign n14124 = n12357 & n14123 ;
  assign n14122 = n3632 | n4096 ;
  assign n14125 = n14124 ^ n14122 ^ 1'b0 ;
  assign n14126 = n1036 & ~n8683 ;
  assign n14127 = n10018 & ~n14126 ;
  assign n14130 = n590 & n2582 ;
  assign n14131 = n2418 & n14130 ;
  assign n14132 = n6187 | n14131 ;
  assign n14133 = n14132 ^ n2165 ^ 1'b0 ;
  assign n14134 = n3876 & n14133 ;
  assign n14128 = n7778 & ~n9374 ;
  assign n14129 = ~n12383 & n14128 ;
  assign n14135 = n14134 ^ n14129 ^ n41 ;
  assign n14136 = n740 & n2020 ;
  assign n14137 = n12119 ^ n8530 ^ n7189 ;
  assign n14138 = n14137 ^ n7380 ^ 1'b0 ;
  assign n14139 = n14136 & n14138 ;
  assign n14142 = n13950 ^ n9649 ^ 1'b0 ;
  assign n14143 = n2483 & ~n14142 ;
  assign n14140 = n12971 ^ n10219 ^ 1'b0 ;
  assign n14141 = n4212 & n14140 ;
  assign n14144 = n14143 ^ n14141 ^ 1'b0 ;
  assign n14145 = ( ~n2605 & n5890 ) | ( ~n2605 & n8409 ) | ( n5890 & n8409 ) ;
  assign n14146 = n14145 ^ n3607 ^ n3069 ;
  assign n14147 = n14146 ^ n9232 ^ 1'b0 ;
  assign n14148 = n8417 & ~n14147 ;
  assign n14149 = ~n835 & n11345 ;
  assign n14150 = ~n14148 & n14149 ;
  assign n14151 = ( n4114 & ~n4608 ) | ( n4114 & n11418 ) | ( ~n4608 & n11418 ) ;
  assign n14152 = n5968 ^ n4488 ^ 1'b0 ;
  assign n14153 = ~n3810 & n5108 ;
  assign n14154 = n13188 ^ n7298 ^ n5313 ;
  assign n14155 = n5693 & ~n14154 ;
  assign n14156 = n14155 ^ n3151 ^ 1'b0 ;
  assign n14157 = n14156 ^ n5648 ^ 1'b0 ;
  assign n14158 = n5086 | n5657 ;
  assign n14159 = n12127 ^ n5089 ^ 1'b0 ;
  assign n14160 = n6076 | n7757 ;
  assign n14161 = n2217 | n14160 ;
  assign n14162 = n261 | n2186 ;
  assign n14163 = ( n1228 & ~n1334 ) | ( n1228 & n3322 ) | ( ~n1334 & n3322 ) ;
  assign n14164 = n6725 & n14163 ;
  assign n14165 = n3450 | n9428 ;
  assign n14166 = n14165 ^ n9103 ^ 1'b0 ;
  assign n14167 = ( n5808 & n10553 ) | ( n5808 & n12317 ) | ( n10553 & n12317 ) ;
  assign n14168 = n9298 & n14167 ;
  assign n14169 = n8960 ^ n8706 ^ n8130 ;
  assign n14170 = ( ~n4002 & n6506 ) | ( ~n4002 & n14169 ) | ( n6506 & n14169 ) ;
  assign n14171 = n14170 ^ n9124 ^ 1'b0 ;
  assign n14172 = n14168 & ~n14171 ;
  assign n14173 = n9653 ^ n2476 ^ 1'b0 ;
  assign n14174 = n5546 ^ n3014 ^ 1'b0 ;
  assign n14175 = n14174 ^ n4264 ^ 1'b0 ;
  assign n14176 = ~n6039 & n13396 ;
  assign n14177 = ~n2471 & n14176 ;
  assign n14178 = n2059 | n14177 ;
  assign n14179 = n4315 | n7019 ;
  assign n14180 = ~n2429 & n12585 ;
  assign n14181 = n11052 & ~n14180 ;
  assign n14183 = ( ~n966 & n1485 ) | ( ~n966 & n1900 ) | ( n1485 & n1900 ) ;
  assign n14184 = n2433 & ~n14183 ;
  assign n14185 = n12990 & n14184 ;
  assign n14186 = n5404 & ~n7126 ;
  assign n14187 = n14185 & n14186 ;
  assign n14182 = ~n3762 & n8797 ;
  assign n14188 = n14187 ^ n14182 ^ 1'b0 ;
  assign n14189 = n14188 ^ n2816 ^ 1'b0 ;
  assign n14190 = n879 & ~n6273 ;
  assign n14191 = n14190 ^ n9620 ^ 1'b0 ;
  assign n14192 = n8830 & ~n14191 ;
  assign n14193 = n14192 ^ n1547 ^ 1'b0 ;
  assign n14194 = n6399 | n6941 ;
  assign n14195 = n6521 ^ n6091 ^ 1'b0 ;
  assign n14196 = n14194 | n14195 ;
  assign n14197 = n14196 ^ n10810 ^ 1'b0 ;
  assign n14198 = n14197 ^ n5420 ^ 1'b0 ;
  assign n14203 = n2544 ^ n2202 ^ 1'b0 ;
  assign n14204 = n3635 & ~n14203 ;
  assign n14205 = ~n3482 & n8904 ;
  assign n14206 = ~n14204 & n14205 ;
  assign n14207 = n14206 ^ n6120 ^ n1015 ;
  assign n14199 = n3840 ^ n2677 ^ 1'b0 ;
  assign n14200 = n3717 | n14199 ;
  assign n14201 = ~n10323 & n14200 ;
  assign n14202 = n14201 ^ n2553 ^ 1'b0 ;
  assign n14208 = n14207 ^ n14202 ^ n4743 ;
  assign n14209 = n1742 | n7873 ;
  assign n14210 = n7951 | n14209 ;
  assign n14211 = ( n2192 & ~n6095 ) | ( n2192 & n14210 ) | ( ~n6095 & n14210 ) ;
  assign n14212 = ( n9610 & n14135 ) | ( n9610 & n14211 ) | ( n14135 & n14211 ) ;
  assign n14213 = n1793 ^ x3 ^ 1'b0 ;
  assign n14214 = n14213 ^ n7804 ^ 1'b0 ;
  assign n14215 = n12321 ^ n3781 ^ 1'b0 ;
  assign n14216 = n11749 & ~n14215 ;
  assign n14217 = n3385 & ~n11795 ;
  assign n14218 = ~n11626 & n14217 ;
  assign n14219 = n3242 ^ n850 ^ 1'b0 ;
  assign n14220 = n14219 ^ n11272 ^ n5776 ;
  assign n14221 = n4465 & n7029 ;
  assign n14222 = n2840 & n14221 ;
  assign n14223 = n3684 & ~n14222 ;
  assign n14224 = n13927 & n14223 ;
  assign n14225 = n14224 ^ n3946 ^ 1'b0 ;
  assign n14226 = ~n8420 & n14225 ;
  assign n14227 = n1569 | n4659 ;
  assign n14228 = n1015 & n1147 ;
  assign n14229 = ( n3217 & ~n4400 ) | ( n3217 & n14228 ) | ( ~n4400 & n14228 ) ;
  assign n14230 = n5890 ^ n2818 ^ 1'b0 ;
  assign n14231 = n2021 & n14230 ;
  assign n14232 = n8725 ^ n4842 ^ 1'b0 ;
  assign n14233 = n14231 & ~n14232 ;
  assign n14234 = n14229 & n14233 ;
  assign n14235 = n14234 ^ n2162 ^ 1'b0 ;
  assign n14236 = n7970 & ~n14235 ;
  assign n14237 = n9829 ^ n2944 ^ 1'b0 ;
  assign n14238 = n10968 & ~n14237 ;
  assign n14239 = n14238 ^ n12638 ^ 1'b0 ;
  assign n14240 = n1815 | n9444 ;
  assign n14241 = ~n12028 & n14240 ;
  assign n14242 = n1672 & n3481 ;
  assign n14243 = n14242 ^ n6596 ^ 1'b0 ;
  assign n14244 = n1857 ^ n1153 ^ n919 ;
  assign n14245 = n931 & n4093 ;
  assign n14246 = n14244 & n14245 ;
  assign n14247 = n14246 ^ n1311 ^ 1'b0 ;
  assign n14248 = n3151 & n14247 ;
  assign n14249 = n14248 ^ n5261 ^ 1'b0 ;
  assign n14250 = ~n6027 & n12987 ;
  assign n14251 = n14250 ^ n10490 ^ 1'b0 ;
  assign n14252 = n4421 & n11495 ;
  assign n14253 = ~n5925 & n11062 ;
  assign n14254 = n14253 ^ n9117 ^ 1'b0 ;
  assign n14255 = n3384 | n5724 ;
  assign n14256 = n6004 ^ n3364 ^ n1033 ;
  assign n14257 = n14256 ^ n10664 ^ 1'b0 ;
  assign n14258 = n2515 ^ n1040 ^ n91 ;
  assign n14259 = n14258 ^ n4300 ^ 1'b0 ;
  assign n14260 = n9621 ^ n8119 ^ 1'b0 ;
  assign n14261 = n8061 | n14260 ;
  assign n14262 = ~n1937 & n12921 ;
  assign n14263 = n754 & n14262 ;
  assign n14264 = n6098 ^ n2393 ^ 1'b0 ;
  assign n14265 = n5828 ^ n3387 ^ 1'b0 ;
  assign n14266 = n6551 & n14265 ;
  assign n14268 = n130 & ~n3546 ;
  assign n14269 = n3546 & n14268 ;
  assign n14267 = ~n9426 & n12779 ;
  assign n14270 = n14269 ^ n14267 ^ 1'b0 ;
  assign n14271 = n6656 ^ n3313 ^ 1'b0 ;
  assign n14272 = n6477 & n14271 ;
  assign n14273 = n14272 ^ n3722 ^ 1'b0 ;
  assign n14274 = n13768 | n14273 ;
  assign n14275 = n10304 & ~n14274 ;
  assign n14276 = n9817 ^ n2496 ^ 1'b0 ;
  assign n14277 = ~n989 & n14276 ;
  assign n14278 = n8120 & ~n14277 ;
  assign n14279 = n3240 ^ n995 ^ 1'b0 ;
  assign n14280 = n14279 ^ n4375 ^ 1'b0 ;
  assign n14281 = n12969 | n14280 ;
  assign n14282 = n3106 ^ n42 ^ 1'b0 ;
  assign n14283 = n4560 ^ n2698 ^ 1'b0 ;
  assign n14284 = n14283 ^ n1231 ^ 1'b0 ;
  assign n14285 = n5478 | n14284 ;
  assign n14286 = ( n2728 & n14282 ) | ( n2728 & n14285 ) | ( n14282 & n14285 ) ;
  assign n14287 = n9519 & ~n14286 ;
  assign n14288 = n13988 ^ n1026 ^ 1'b0 ;
  assign n14289 = ( ~n4450 & n5684 ) | ( ~n4450 & n11642 ) | ( n5684 & n11642 ) ;
  assign n14290 = n14289 ^ n10816 ^ n2607 ;
  assign n14291 = ( ~n2074 & n5223 ) | ( ~n2074 & n12368 ) | ( n5223 & n12368 ) ;
  assign n14292 = ~n12259 & n14291 ;
  assign n14293 = ( n814 & n6093 ) | ( n814 & ~n14292 ) | ( n6093 & ~n14292 ) ;
  assign n14294 = n3851 | n4557 ;
  assign n14295 = n4911 ^ n3817 ^ 1'b0 ;
  assign n14296 = ( n11836 & n14294 ) | ( n11836 & n14295 ) | ( n14294 & n14295 ) ;
  assign n14297 = n10745 & n13206 ;
  assign n14298 = n6754 | n14297 ;
  assign n14299 = n2832 ^ n121 ^ 1'b0 ;
  assign n14300 = n14299 ^ n1924 ^ 1'b0 ;
  assign n14301 = n1786 & ~n14300 ;
  assign n14302 = n2818 ^ n696 ^ 1'b0 ;
  assign n14303 = n2176 & n14302 ;
  assign n14304 = ~n6947 & n7054 ;
  assign n14305 = ~n6098 & n14304 ;
  assign n14306 = n799 | n12801 ;
  assign n14307 = n14305 & ~n14306 ;
  assign n14308 = ( n2787 & n4567 ) | ( n2787 & n4584 ) | ( n4567 & n4584 ) ;
  assign n14309 = n3054 | n14308 ;
  assign n14310 = n14309 ^ n10123 ^ n8440 ;
  assign n14311 = n7116 & ~n9898 ;
  assign n14312 = n14311 ^ n7312 ^ 1'b0 ;
  assign n14313 = ( n1912 & n12481 ) | ( n1912 & n14312 ) | ( n12481 & n14312 ) ;
  assign n14314 = n10479 ^ n9912 ^ 1'b0 ;
  assign n14315 = n11460 | n14314 ;
  assign n14316 = n6789 & ~n14315 ;
  assign n14317 = n3235 | n4021 ;
  assign n14318 = n14317 ^ n9330 ^ 1'b0 ;
  assign n14319 = ~n3087 & n14318 ;
  assign n14320 = n14319 ^ n5329 ^ 1'b0 ;
  assign n14321 = n1170 & ~n14320 ;
  assign n14322 = n14321 ^ n13503 ^ 1'b0 ;
  assign n14323 = ~n115 & n14322 ;
  assign n14324 = n6958 & n13736 ;
  assign n14325 = n5341 | n6062 ;
  assign n14326 = n14325 ^ n13582 ^ 1'b0 ;
  assign n14328 = n13643 ^ n8754 ^ 1'b0 ;
  assign n14327 = n9798 & n12789 ;
  assign n14329 = n14328 ^ n14327 ^ 1'b0 ;
  assign n14332 = n2755 | n12569 ;
  assign n14330 = n2176 & ~n9497 ;
  assign n14331 = n14330 ^ n1463 ^ 1'b0 ;
  assign n14333 = n14332 ^ n14331 ^ 1'b0 ;
  assign n14334 = n6285 ^ n3145 ^ 1'b0 ;
  assign n14335 = n13470 & n14334 ;
  assign n14336 = n1516 | n8181 ;
  assign n14337 = n3211 & ~n14336 ;
  assign n14338 = n11267 ^ n91 ^ 1'b0 ;
  assign n14339 = n14338 ^ n2503 ^ 1'b0 ;
  assign n14340 = n11243 & ~n14339 ;
  assign n14341 = n1024 & n14340 ;
  assign n14342 = ~n14106 & n14341 ;
  assign n14343 = n4701 & n13180 ;
  assign n14344 = n12553 ^ n4686 ^ n494 ;
  assign n14347 = n3665 & n5092 ;
  assign n14345 = n4785 ^ n2666 ^ 1'b0 ;
  assign n14346 = n1628 & n14345 ;
  assign n14348 = n14347 ^ n14346 ^ 1'b0 ;
  assign n14349 = n6037 & n10871 ;
  assign n14350 = ~n6890 & n14349 ;
  assign n14351 = n5380 & ~n14350 ;
  assign n14352 = ( n879 & n2999 ) | ( n879 & ~n9775 ) | ( n2999 & ~n9775 ) ;
  assign n14353 = n14352 ^ n9781 ^ 1'b0 ;
  assign n14354 = ~n7315 & n14353 ;
  assign n14355 = ~n1399 & n14354 ;
  assign n14356 = n1426 & n14355 ;
  assign n14357 = n3858 ^ n3709 ^ 1'b0 ;
  assign n14358 = ~n1043 & n14357 ;
  assign n14359 = n6242 ^ n3818 ^ 1'b0 ;
  assign n14360 = n14358 & n14359 ;
  assign n14361 = n14360 ^ n4900 ^ 1'b0 ;
  assign n14362 = n2827 | n4915 ;
  assign n14363 = n14361 | n14362 ;
  assign n14364 = n7278 & n14363 ;
  assign n14365 = n11391 ^ n4599 ^ 1'b0 ;
  assign n14366 = n14365 ^ n5395 ^ 1'b0 ;
  assign n14367 = ~n1040 & n10054 ;
  assign n14368 = n1729 ^ n26 ^ 1'b0 ;
  assign n14369 = ~n5524 & n14368 ;
  assign n14370 = n14369 ^ n10200 ^ 1'b0 ;
  assign n14371 = ( n40 & n7721 ) | ( n40 & ~n14370 ) | ( n7721 & ~n14370 ) ;
  assign n14372 = n678 & n12548 ;
  assign n14373 = ~n3606 & n14372 ;
  assign n14374 = ( n4706 & ~n13462 ) | ( n4706 & n14373 ) | ( ~n13462 & n14373 ) ;
  assign n14375 = ~n2305 & n13099 ;
  assign n14376 = n8701 & n14375 ;
  assign n14377 = ~n922 & n14376 ;
  assign n14378 = n1135 | n10068 ;
  assign n14379 = n6083 ^ n4066 ^ 1'b0 ;
  assign n14380 = n16 | n14379 ;
  assign n14381 = n14380 ^ n1143 ^ n57 ;
  assign n14382 = n4738 & ~n5987 ;
  assign n14383 = n14382 ^ n8215 ^ 1'b0 ;
  assign n14384 = n115 & n1085 ;
  assign n14385 = ~n3590 & n14384 ;
  assign n14386 = n4324 ^ n3493 ^ n2667 ;
  assign n14387 = n2460 & n14386 ;
  assign n14388 = ~n2649 & n14387 ;
  assign n14389 = n5967 & ~n14388 ;
  assign n14390 = n1545 & ~n2646 ;
  assign n14391 = ~n14389 & n14390 ;
  assign n14392 = n10428 ^ n7358 ^ 1'b0 ;
  assign n14393 = ~n7496 & n14392 ;
  assign n14394 = n5164 ^ n1109 ^ 1'b0 ;
  assign n14395 = n14394 ^ n1783 ^ 1'b0 ;
  assign n14396 = n14395 ^ n12286 ^ 1'b0 ;
  assign n14397 = ~n4918 & n14396 ;
  assign n14398 = ~n5963 & n14397 ;
  assign n14399 = n14398 ^ n461 ^ 1'b0 ;
  assign n14400 = n1562 & ~n6457 ;
  assign n14401 = n14400 ^ n9165 ^ 1'b0 ;
  assign n14402 = n6583 & n14401 ;
  assign n14403 = ~n4570 & n14402 ;
  assign n14404 = n8303 & ~n14403 ;
  assign n14405 = n14404 ^ n8551 ^ 1'b0 ;
  assign n14406 = ~n5051 & n5285 ;
  assign n14407 = ( ~n4111 & n11662 ) | ( ~n4111 & n14406 ) | ( n11662 & n14406 ) ;
  assign n14408 = n3066 ^ n1022 ^ 1'b0 ;
  assign n14409 = n1064 | n14408 ;
  assign n14410 = n12682 ^ n299 ^ 1'b0 ;
  assign n14411 = n13165 | n14410 ;
  assign n14412 = n6131 & n12784 ;
  assign n14413 = n14412 ^ n7086 ^ 1'b0 ;
  assign n14414 = n14102 ^ n1437 ^ 1'b0 ;
  assign n14415 = ~n1339 & n14414 ;
  assign n14416 = ( n3127 & n5903 ) | ( n3127 & n6890 ) | ( n5903 & n6890 ) ;
  assign n14417 = n1212 & ~n14416 ;
  assign n14418 = ~n7292 & n14417 ;
  assign n14419 = ~n243 & n3784 ;
  assign n14420 = n14418 & ~n14419 ;
  assign n14421 = n1040 & n14420 ;
  assign n14422 = ( n6227 & ~n6743 ) | ( n6227 & n13151 ) | ( ~n6743 & n13151 ) ;
  assign n14425 = n1823 & n11149 ;
  assign n14426 = n2284 & ~n14425 ;
  assign n14423 = n289 & n4548 ;
  assign n14424 = n14423 ^ n4647 ^ 1'b0 ;
  assign n14427 = n14426 ^ n14424 ^ n12638 ;
  assign n14428 = n5140 & n9655 ;
  assign n14430 = n8763 ^ n3246 ^ 1'b0 ;
  assign n14431 = n2048 & n14430 ;
  assign n14429 = n8884 ^ n5496 ^ 1'b0 ;
  assign n14432 = n14431 ^ n14429 ^ 1'b0 ;
  assign n14433 = n7055 & n14432 ;
  assign n14434 = n2313 | n2725 ;
  assign n14436 = n611 & n1488 ;
  assign n14437 = ~n3789 & n14436 ;
  assign n14435 = ~n996 & n4252 ;
  assign n14438 = n14437 ^ n14435 ^ 1'b0 ;
  assign n14439 = n14438 ^ n6511 ^ n2497 ;
  assign n14440 = n91 & n1596 ;
  assign n14441 = n13262 ^ n1694 ^ 1'b0 ;
  assign n14442 = n3949 ^ n2176 ^ 1'b0 ;
  assign n14443 = n10623 ^ n7859 ^ 1'b0 ;
  assign n14444 = n5584 | n7218 ;
  assign n14445 = n1928 & ~n14444 ;
  assign n14446 = n14445 ^ n3710 ^ n2039 ;
  assign n14447 = ( n3187 & n14443 ) | ( n3187 & n14446 ) | ( n14443 & n14446 ) ;
  assign n14448 = n10180 ^ n5118 ^ n1439 ;
  assign n14449 = n14448 ^ n12548 ^ n4319 ;
  assign n14453 = ( ~n1807 & n5446 ) | ( ~n1807 & n5522 ) | ( n5446 & n5522 ) ;
  assign n14450 = ~n1660 & n3569 ;
  assign n14451 = n6576 & n13611 ;
  assign n14452 = n14450 & n14451 ;
  assign n14454 = n14453 ^ n14452 ^ 1'b0 ;
  assign n14455 = n421 | n1787 ;
  assign n14456 = n4521 | n14455 ;
  assign n14457 = n14456 ^ n7702 ^ 1'b0 ;
  assign n14458 = n12532 & ~n14457 ;
  assign n14459 = n7988 ^ n6590 ^ 1'b0 ;
  assign n14460 = n5470 & n9085 ;
  assign n14461 = n13739 & ~n14460 ;
  assign n14462 = n14461 ^ n11278 ^ 1'b0 ;
  assign n14463 = n4325 | n6845 ;
  assign n14464 = n14463 ^ n10433 ^ n1594 ;
  assign n14465 = n11700 ^ n5264 ^ 1'b0 ;
  assign n14469 = n6565 ^ n3130 ^ 1'b0 ;
  assign n14470 = n713 | n14469 ;
  assign n14468 = n8896 ^ n8894 ^ 1'b0 ;
  assign n14471 = n14470 ^ n14468 ^ 1'b0 ;
  assign n14466 = n355 & ~n4102 ;
  assign n14467 = n5725 & n14466 ;
  assign n14472 = n14471 ^ n14467 ^ 1'b0 ;
  assign n14473 = ( ~n1295 & n10315 ) | ( ~n1295 & n14472 ) | ( n10315 & n14472 ) ;
  assign n14475 = n1122 | n5565 ;
  assign n14474 = ~n3284 & n13676 ;
  assign n14476 = n14475 ^ n14474 ^ 1'b0 ;
  assign n14477 = n255 | n14476 ;
  assign n14478 = n9964 ^ n6324 ^ 1'b0 ;
  assign n14479 = n8390 ^ n431 ^ 1'b0 ;
  assign n14480 = n14479 ^ n12627 ^ 1'b0 ;
  assign n14481 = ( n6487 & ~n9148 ) | ( n6487 & n13839 ) | ( ~n9148 & n13839 ) ;
  assign n14482 = n5768 | n14481 ;
  assign n14483 = n8885 ^ n8676 ^ 1'b0 ;
  assign n14484 = n2986 ^ n2633 ^ 1'b0 ;
  assign n14485 = n14484 ^ n1245 ^ 1'b0 ;
  assign n14486 = n3819 & n5559 ;
  assign n14487 = n14486 ^ n4491 ^ 1'b0 ;
  assign n14488 = n12025 | n14487 ;
  assign n14489 = n1664 & ~n6689 ;
  assign n14490 = n14489 ^ n1439 ^ 1'b0 ;
  assign n14491 = n3700 | n14490 ;
  assign n14492 = n14491 ^ n4062 ^ 1'b0 ;
  assign n14493 = n10170 ^ n216 ^ 1'b0 ;
  assign n14494 = n3987 & n12664 ;
  assign n14495 = n14494 ^ n1202 ^ 1'b0 ;
  assign n14496 = n1896 | n14495 ;
  assign n14497 = n14493 & ~n14496 ;
  assign n14498 = ( n93 & n1577 ) | ( n93 & ~n14497 ) | ( n1577 & ~n14497 ) ;
  assign n14499 = n2440 | n4019 ;
  assign n14500 = n8407 ^ n7360 ^ 1'b0 ;
  assign n14501 = n14500 ^ n8051 ^ 1'b0 ;
  assign n14502 = n14083 & n14501 ;
  assign n14503 = n8880 & n14502 ;
  assign n14504 = n4699 & ~n10196 ;
  assign n14505 = n1182 & ~n9350 ;
  assign n14506 = n9839 | n14505 ;
  assign n14507 = n8532 ^ n3660 ^ n514 ;
  assign n14508 = n14507 ^ n10233 ^ 1'b0 ;
  assign n14509 = n684 ^ n202 ^ 1'b0 ;
  assign n14510 = n14509 ^ n2305 ^ 1'b0 ;
  assign n14511 = n14510 ^ n396 ^ 1'b0 ;
  assign n14512 = n14508 & n14511 ;
  assign n14513 = n6080 ^ n3406 ^ 1'b0 ;
  assign n14514 = n4743 & ~n14513 ;
  assign n14515 = n14514 ^ n12033 ^ 1'b0 ;
  assign n14516 = n14491 | n14515 ;
  assign n14517 = n14516 ^ n11762 ^ n2034 ;
  assign n14518 = n8058 ^ n668 ^ n313 ;
  assign n14519 = n13270 ^ n1875 ^ 1'b0 ;
  assign n14520 = n4271 | n14519 ;
  assign n14521 = n2566 & ~n14520 ;
  assign n14522 = n496 & n14521 ;
  assign n14526 = n13329 ^ n9490 ^ n969 ;
  assign n14523 = n6583 ^ n4426 ^ 1'b0 ;
  assign n14524 = n14523 ^ n1181 ^ 1'b0 ;
  assign n14525 = ~n10223 & n14524 ;
  assign n14527 = n14526 ^ n14525 ^ 1'b0 ;
  assign n14528 = n1083 & ~n7446 ;
  assign n14529 = n14528 ^ n1491 ^ 1'b0 ;
  assign n14530 = ( ~n111 & n749 ) | ( ~n111 & n7468 ) | ( n749 & n7468 ) ;
  assign n14531 = n7790 | n14530 ;
  assign n14532 = n757 & n2060 ;
  assign n14533 = n14532 ^ n8655 ^ n4147 ;
  assign n14534 = n9998 ^ n7448 ^ 1'b0 ;
  assign n14535 = n7014 ^ n3475 ^ n2650 ;
  assign n14536 = n6435 | n14535 ;
  assign n14537 = n14536 ^ n6745 ^ 1'b0 ;
  assign n14538 = ~n14534 & n14537 ;
  assign n14539 = ~n5099 & n14538 ;
  assign n14540 = n5387 | n10230 ;
  assign n14541 = n6872 & ~n14540 ;
  assign n14542 = n14541 ^ n1893 ^ 1'b0 ;
  assign n14543 = ( ~n9471 & n10108 ) | ( ~n9471 & n11748 ) | ( n10108 & n11748 ) ;
  assign n14544 = n11129 ^ n10535 ^ 1'b0 ;
  assign n14545 = n6287 ^ n3515 ^ 1'b0 ;
  assign n14546 = n3959 ^ n1838 ^ 1'b0 ;
  assign n14547 = ~n3575 & n14546 ;
  assign n14548 = n14547 ^ n5874 ^ n5708 ;
  assign n14549 = n944 & n1253 ;
  assign n14550 = ~n14548 & n14549 ;
  assign n14551 = ~n839 & n1406 ;
  assign n14552 = ~n4095 & n10260 ;
  assign n14553 = n10197 & n14552 ;
  assign n14554 = ( n2280 & n14551 ) | ( n2280 & n14553 ) | ( n14551 & n14553 ) ;
  assign n14555 = ~n1175 & n7130 ;
  assign n14556 = n14555 ^ n4052 ^ 1'b0 ;
  assign n14557 = n14530 & n14556 ;
  assign n14558 = n5552 ^ n2463 ^ 1'b0 ;
  assign n14559 = ~n5768 & n14558 ;
  assign n14560 = ( n823 & ~n14557 ) | ( n823 & n14559 ) | ( ~n14557 & n14559 ) ;
  assign n14563 = n8945 ^ n1586 ^ 1'b0 ;
  assign n14564 = n1280 & ~n14563 ;
  assign n14561 = n5016 ^ n4093 ^ 1'b0 ;
  assign n14562 = n4055 & n14561 ;
  assign n14565 = n14564 ^ n14562 ^ 1'b0 ;
  assign n14566 = n2570 | n13032 ;
  assign n14567 = ~n6353 & n8448 ;
  assign n14570 = n63 | n13155 ;
  assign n14568 = ~n483 & n8002 ;
  assign n14569 = ~n6620 & n14568 ;
  assign n14571 = n14570 ^ n14569 ^ 1'b0 ;
  assign n14572 = n8007 | n14571 ;
  assign n14573 = ( n57 & ~n4795 ) | ( n57 & n14572 ) | ( ~n4795 & n14572 ) ;
  assign n14574 = ~n6607 & n13980 ;
  assign n14575 = ~n14573 & n14574 ;
  assign n14576 = n8784 ^ n4100 ^ n3772 ;
  assign n14577 = n2088 | n13815 ;
  assign n14578 = n14577 ^ n5316 ^ 1'b0 ;
  assign n14579 = n14578 ^ n8291 ^ 1'b0 ;
  assign n14580 = ~n14576 & n14579 ;
  assign n14581 = ~n134 & n2935 ;
  assign n14582 = n14581 ^ n12855 ^ 1'b0 ;
  assign n14583 = n14580 & n14582 ;
  assign n14584 = ( n2994 & ~n3037 ) | ( n2994 & n12854 ) | ( ~n3037 & n12854 ) ;
  assign n14585 = ~n9344 & n10165 ;
  assign n14586 = n3568 ^ n1018 ^ 1'b0 ;
  assign n14587 = n14586 ^ n11149 ^ 1'b0 ;
  assign n14588 = n12963 ^ n10977 ^ 1'b0 ;
  assign n14589 = ~n14587 & n14588 ;
  assign n14590 = n2339 & ~n13072 ;
  assign n14591 = n13903 ^ n11884 ^ 1'b0 ;
  assign n14592 = n6245 & ~n14591 ;
  assign n14595 = n12569 ^ n68 ^ 1'b0 ;
  assign n14596 = n14595 ^ n5524 ^ 1'b0 ;
  assign n14597 = n750 & ~n14596 ;
  assign n14593 = ( n5464 & n8542 ) | ( n5464 & ~n13243 ) | ( n8542 & ~n13243 ) ;
  assign n14594 = n3508 & n14593 ;
  assign n14598 = n14597 ^ n14594 ^ 1'b0 ;
  assign n14599 = n14598 ^ n1431 ^ 1'b0 ;
  assign n14600 = n7514 & ~n14599 ;
  assign n14602 = n4925 & ~n9956 ;
  assign n14603 = n14602 ^ n6008 ^ 1'b0 ;
  assign n14601 = n954 | n10922 ;
  assign n14604 = n14603 ^ n14601 ^ 1'b0 ;
  assign n14605 = n14600 & ~n14604 ;
  assign n14614 = n5205 ^ n1446 ^ 1'b0 ;
  assign n14615 = n16 & ~n14614 ;
  assign n14616 = n14615 ^ n4872 ^ 1'b0 ;
  assign n14613 = n2422 | n5241 ;
  assign n14617 = n14616 ^ n14613 ^ 1'b0 ;
  assign n14606 = n3339 ^ n1558 ^ 1'b0 ;
  assign n14607 = n1489 & n14606 ;
  assign n14608 = ~n1311 & n14607 ;
  assign n14609 = ~n376 & n14608 ;
  assign n14610 = n6333 & n14609 ;
  assign n14611 = ~n4142 & n14610 ;
  assign n14612 = n14611 ^ n6951 ^ n4846 ;
  assign n14618 = n14617 ^ n14612 ^ 1'b0 ;
  assign n14619 = n609 & ~n14618 ;
  assign n14620 = n10023 ^ n5315 ^ n2583 ;
  assign n14628 = n3245 ^ n2044 ^ 1'b0 ;
  assign n14625 = ~n3001 & n4422 ;
  assign n14626 = n14625 ^ n11888 ^ 1'b0 ;
  assign n14627 = n8890 & n14626 ;
  assign n14629 = n14628 ^ n14627 ^ 1'b0 ;
  assign n14622 = n12290 ^ n7989 ^ n3382 ;
  assign n14623 = n14622 ^ n5735 ^ 1'b0 ;
  assign n14621 = n1800 | n6026 ;
  assign n14624 = n14623 ^ n14621 ^ 1'b0 ;
  assign n14630 = n14629 ^ n14624 ^ n2524 ;
  assign n14631 = n1247 | n1718 ;
  assign n14632 = n14631 ^ n6313 ^ 1'b0 ;
  assign n14633 = n14632 ^ n494 ^ 1'b0 ;
  assign n14634 = n14630 | n14633 ;
  assign n14635 = n14013 ^ n11255 ^ 1'b0 ;
  assign n14636 = n10328 ^ n8275 ^ 1'b0 ;
  assign n14637 = n914 & n4858 ;
  assign n14638 = n1818 & n14637 ;
  assign n14639 = ~n401 & n7869 ;
  assign n14640 = n14638 | n14639 ;
  assign n14641 = n8866 ^ n7765 ^ n6280 ;
  assign n14642 = n554 & n14641 ;
  assign n14643 = n6563 & ~n6727 ;
  assign n14644 = n14643 ^ n3778 ^ 1'b0 ;
  assign n14645 = n9588 & ~n14644 ;
  assign n14648 = n2021 & ~n9937 ;
  assign n14649 = n14648 ^ n4195 ^ 1'b0 ;
  assign n14646 = n1009 ^ n691 ^ 1'b0 ;
  assign n14647 = ~n9283 & n14646 ;
  assign n14650 = n14649 ^ n14647 ^ 1'b0 ;
  assign n14651 = n2228 | n8432 ;
  assign n14652 = n14651 ^ n7304 ^ 1'b0 ;
  assign n14653 = ~n10815 & n14652 ;
  assign n14654 = n4461 ^ n3387 ^ 1'b0 ;
  assign n14655 = ~n707 & n14654 ;
  assign n14656 = n14655 ^ n12397 ^ 1'b0 ;
  assign n14657 = n2535 & n6603 ;
  assign n14658 = n1509 ^ n983 ^ 1'b0 ;
  assign n14659 = ~n1531 & n4097 ;
  assign n14660 = n3883 & ~n8346 ;
  assign n14661 = ~n14659 & n14660 ;
  assign n14662 = n14661 ^ n12987 ^ 1'b0 ;
  assign n14663 = n1900 & n10197 ;
  assign n14664 = ~n7121 & n8903 ;
  assign n14665 = n7335 ^ n3790 ^ n3094 ;
  assign n14666 = n2542 & ~n14665 ;
  assign n14667 = ~n713 & n14666 ;
  assign n14668 = ~n443 & n14667 ;
  assign n14669 = n4055 & ~n14668 ;
  assign n14670 = n14669 ^ n3016 ^ 1'b0 ;
  assign n14671 = n12488 ^ n366 ^ 1'b0 ;
  assign n14678 = n9889 ^ n1542 ^ n1145 ;
  assign n14679 = n772 & n4998 ;
  assign n14680 = n14679 ^ n8585 ^ 1'b0 ;
  assign n14681 = n9443 & ~n14680 ;
  assign n14682 = n14681 ^ n7869 ^ 1'b0 ;
  assign n14683 = n14678 & n14682 ;
  assign n14672 = n2296 ^ n1105 ^ 1'b0 ;
  assign n14673 = n1715 | n11387 ;
  assign n14674 = n4591 & ~n14673 ;
  assign n14675 = n14672 | n14674 ;
  assign n14676 = ~n3384 & n12567 ;
  assign n14677 = n14675 & n14676 ;
  assign n14684 = n14683 ^ n14677 ^ 1'b0 ;
  assign n14685 = n7896 ^ n203 ^ 1'b0 ;
  assign n14686 = n11931 & ~n14685 ;
  assign n14687 = n11754 ^ n1869 ^ 1'b0 ;
  assign n14688 = n13 & ~n9946 ;
  assign n14689 = n5916 & ~n7726 ;
  assign n14690 = ~n14607 & n14689 ;
  assign n14691 = n14690 ^ n9876 ^ 1'b0 ;
  assign n14692 = n8575 & n14691 ;
  assign n14693 = n14692 ^ n7360 ^ 1'b0 ;
  assign n14694 = ~n8911 & n14693 ;
  assign n14695 = ( n2781 & n3066 ) | ( n2781 & n12002 ) | ( n3066 & n12002 ) ;
  assign n14696 = n3035 ^ n1105 ^ 1'b0 ;
  assign n14697 = ~n5748 & n9172 ;
  assign n14698 = n14697 ^ n4475 ^ 1'b0 ;
  assign n14700 = ( n2447 & n4338 ) | ( n2447 & n14373 ) | ( n4338 & n14373 ) ;
  assign n14699 = n8125 ^ n99 ^ 1'b0 ;
  assign n14701 = n14700 ^ n14699 ^ n5356 ;
  assign n14702 = n3079 & n6947 ;
  assign n14703 = n14702 ^ n9115 ^ 1'b0 ;
  assign n14708 = ~n5764 & n6555 ;
  assign n14709 = n14708 ^ n5534 ^ 1'b0 ;
  assign n14705 = n4620 ^ n3932 ^ 1'b0 ;
  assign n14706 = ~n12522 & n14705 ;
  assign n14704 = ~n1752 & n11437 ;
  assign n14707 = n14706 ^ n14704 ^ 1'b0 ;
  assign n14710 = n14709 ^ n14707 ^ 1'b0 ;
  assign n14711 = n6392 | n14051 ;
  assign n14712 = n3569 ^ n2004 ^ 1'b0 ;
  assign n14713 = ~n44 & n14712 ;
  assign n14714 = n14713 ^ n6289 ^ 1'b0 ;
  assign n14715 = n4251 | n10180 ;
  assign n14716 = n14715 ^ n8688 ^ n1566 ;
  assign n14717 = n14716 ^ n2067 ^ 1'b0 ;
  assign n14718 = n8671 & ~n14717 ;
  assign n14719 = ~n1561 & n2583 ;
  assign n14720 = n14719 ^ n1315 ^ 1'b0 ;
  assign n14721 = n3241 | n14720 ;
  assign n14722 = n14721 ^ n9137 ^ 1'b0 ;
  assign n14723 = n63 & n14722 ;
  assign n14724 = n10793 ^ n6227 ^ 1'b0 ;
  assign n14725 = n7554 | n14724 ;
  assign n14726 = n1693 ^ n1175 ^ 1'b0 ;
  assign n14727 = n2906 & ~n14726 ;
  assign n14728 = n11672 ^ n3092 ^ 1'b0 ;
  assign n14729 = n14727 & ~n14728 ;
  assign n14730 = n654 & n2964 ;
  assign n14731 = n14730 ^ n59 ^ 1'b0 ;
  assign n14732 = n14731 ^ n5935 ^ 1'b0 ;
  assign n14733 = n12469 ^ n6451 ^ 1'b0 ;
  assign n14734 = n14732 | n14733 ;
  assign n14735 = n852 & n974 ;
  assign n14736 = n14735 ^ n8234 ^ 1'b0 ;
  assign n14737 = n5323 & n14736 ;
  assign n14738 = ~n823 & n963 ;
  assign n14739 = n97 | n299 ;
  assign n14740 = n14738 | n14739 ;
  assign n14741 = ~n14737 & n14740 ;
  assign n14742 = n5898 ^ n1502 ^ 1'b0 ;
  assign n14743 = n10958 & ~n14742 ;
  assign n14747 = ~n2943 & n9230 ;
  assign n14748 = n14747 ^ n10550 ^ 1'b0 ;
  assign n14744 = n2942 ^ n1054 ^ 1'b0 ;
  assign n14745 = n9552 ^ n3660 ^ 1'b0 ;
  assign n14746 = n14744 & n14745 ;
  assign n14749 = n14748 ^ n14746 ^ 1'b0 ;
  assign n14750 = n12921 ^ n5882 ^ 1'b0 ;
  assign n14751 = ~n944 & n4331 ;
  assign n14752 = n14751 ^ n2217 ^ 1'b0 ;
  assign n14753 = n3016 & n14752 ;
  assign n14757 = n2846 | n6062 ;
  assign n14754 = n65 | n3144 ;
  assign n14755 = n14754 ^ n3496 ^ 1'b0 ;
  assign n14756 = n14755 ^ n5657 ^ 1'b0 ;
  assign n14758 = n14757 ^ n14756 ^ 1'b0 ;
  assign n14759 = n14755 ^ n4113 ^ 1'b0 ;
  assign n14760 = ~n2447 & n14759 ;
  assign n14761 = n558 & n4925 ;
  assign n14762 = n14760 & n14761 ;
  assign n14763 = n14762 ^ n8353 ^ 1'b0 ;
  assign n14764 = n6389 | n14763 ;
  assign n14765 = n3101 & ~n5568 ;
  assign n14766 = n8838 ^ n1838 ^ 1'b0 ;
  assign n14767 = ~n8326 & n14228 ;
  assign n14768 = ~n14766 & n14767 ;
  assign n14769 = n2877 | n11568 ;
  assign n14770 = n14769 ^ n13550 ^ 1'b0 ;
  assign n14771 = n12030 & n14770 ;
  assign n14772 = ~n741 & n1072 ;
  assign n14773 = n5503 | n11643 ;
  assign n14774 = n13209 | n14773 ;
  assign n14775 = n972 ^ n849 ^ 1'b0 ;
  assign n14776 = n14775 ^ n9014 ^ n4689 ;
  assign n14777 = n1666 | n14776 ;
  assign n14778 = n5533 ^ n2665 ^ 1'b0 ;
  assign n14779 = n14778 ^ n1122 ^ 1'b0 ;
  assign n14780 = n4460 ^ n886 ^ 1'b0 ;
  assign n14781 = n946 | n14780 ;
  assign n14782 = n4043 & ~n4066 ;
  assign n14783 = n6272 & n14782 ;
  assign n14784 = ( n5720 & n14781 ) | ( n5720 & n14783 ) | ( n14781 & n14783 ) ;
  assign n14785 = n2402 | n14784 ;
  assign n14786 = n14785 ^ n12847 ^ 1'b0 ;
  assign n14787 = n6021 ^ n4333 ^ 1'b0 ;
  assign n14788 = ~n6111 & n14787 ;
  assign n14789 = n13600 ^ n2883 ^ 1'b0 ;
  assign n14790 = n7391 | n14789 ;
  assign n14791 = ( n4872 & n10136 ) | ( n4872 & ~n10968 ) | ( n10136 & ~n10968 ) ;
  assign n14792 = ~n3107 & n11647 ;
  assign n14793 = ~n8741 & n14792 ;
  assign n14794 = ~n14791 & n14793 ;
  assign n14795 = n2110 & n4127 ;
  assign n14796 = n14795 ^ n1622 ^ 1'b0 ;
  assign n14797 = n14796 ^ n12985 ^ n8046 ;
  assign n14798 = n9996 ^ n1835 ^ 1'b0 ;
  assign n14799 = n571 & ~n4369 ;
  assign n14800 = n14784 ^ n3741 ^ 1'b0 ;
  assign n14801 = ~n7652 & n14800 ;
  assign n14802 = ~n1957 & n5694 ;
  assign n14803 = n14802 ^ n11091 ^ 1'b0 ;
  assign n14804 = n2428 & n5103 ;
  assign n14805 = n7523 & n14804 ;
  assign n14806 = n7617 ^ n661 ^ 1'b0 ;
  assign n14807 = ~n3779 & n14806 ;
  assign n14808 = ( ~n3918 & n14805 ) | ( ~n3918 & n14807 ) | ( n14805 & n14807 ) ;
  assign n14809 = ( ~n381 & n1079 ) | ( ~n381 & n14272 ) | ( n1079 & n14272 ) ;
  assign n14810 = ~n2108 & n14809 ;
  assign n14811 = n14808 & n14810 ;
  assign n14812 = ( ~n887 & n6956 ) | ( ~n887 & n14811 ) | ( n6956 & n14811 ) ;
  assign n14815 = n9012 ^ n4193 ^ 1'b0 ;
  assign n14816 = n14815 ^ n9193 ^ 1'b0 ;
  assign n14813 = ~n1167 & n7288 ;
  assign n14814 = ~n3305 & n14813 ;
  assign n14817 = n14816 ^ n14814 ^ 1'b0 ;
  assign n14818 = n2140 | n5286 ;
  assign n14837 = n11832 | n11994 ;
  assign n14838 = n4327 & ~n14837 ;
  assign n14839 = n14838 ^ n9858 ^ 1'b0 ;
  assign n14823 = n57 & ~n1296 ;
  assign n14824 = ~n154 & n14823 ;
  assign n14825 = ( ~n1470 & n4626 ) | ( ~n1470 & n14824 ) | ( n4626 & n14824 ) ;
  assign n14819 = n6775 ^ n2233 ^ 1'b0 ;
  assign n14820 = ~n3001 & n14819 ;
  assign n14821 = n6144 | n14820 ;
  assign n14822 = n10288 & n14821 ;
  assign n14826 = n14825 ^ n14822 ^ 1'b0 ;
  assign n14827 = n13257 ^ n8469 ^ n5178 ;
  assign n14828 = n3429 ^ n1523 ^ 1'b0 ;
  assign n14829 = n13561 & ~n14828 ;
  assign n14830 = n14829 ^ n3398 ^ 1'b0 ;
  assign n14831 = ~n3774 & n14830 ;
  assign n14832 = n14827 | n14831 ;
  assign n14833 = n9414 ^ n6929 ^ 1'b0 ;
  assign n14834 = n14833 ^ n3564 ^ 1'b0 ;
  assign n14835 = ~n14832 & n14834 ;
  assign n14836 = n14826 & n14835 ;
  assign n14840 = n14839 ^ n14836 ^ 1'b0 ;
  assign n14841 = ( n5036 & ~n9113 ) | ( n5036 & n11268 ) | ( ~n9113 & n11268 ) ;
  assign n14842 = ~n2474 & n6431 ;
  assign n14843 = n2918 & n5393 ;
  assign n14844 = n8680 & n9191 ;
  assign n14845 = n14844 ^ n2885 ^ 1'b0 ;
  assign n14846 = n14845 ^ n9251 ^ 1'b0 ;
  assign n14847 = n3840 & ~n8212 ;
  assign n14848 = n5554 | n14332 ;
  assign n14849 = n14848 ^ n3579 ^ n1462 ;
  assign n14850 = n10668 ^ n6278 ^ 1'b0 ;
  assign n14851 = n14850 ^ n14029 ^ 1'b0 ;
  assign n14852 = n690 & ~n3393 ;
  assign n14853 = ~n2447 & n14852 ;
  assign n14854 = n6597 & n14853 ;
  assign n14855 = n14854 ^ n13453 ^ n13097 ;
  assign n14856 = ~n11778 & n13186 ;
  assign n14857 = ( n8079 & ~n10129 ) | ( n8079 & n12056 ) | ( ~n10129 & n12056 ) ;
  assign n14858 = n14097 & ~n14857 ;
  assign n14859 = n6660 ^ n6384 ^ 1'b0 ;
  assign n14860 = n14858 | n14859 ;
  assign n14861 = n9487 & ~n14860 ;
  assign n14862 = n14861 ^ n9072 ^ 1'b0 ;
  assign n14863 = n7661 ^ n3564 ^ 1'b0 ;
  assign n14864 = ~n68 & n14863 ;
  assign n14865 = ~n8267 & n14864 ;
  assign n14866 = n14865 ^ n4720 ^ 1'b0 ;
  assign n14867 = ( n2526 & n11774 ) | ( n2526 & ~n14866 ) | ( n11774 & ~n14866 ) ;
  assign n14868 = n4488 | n12066 ;
  assign n14869 = n648 & ~n14868 ;
  assign n14870 = n14869 ^ n13469 ^ 1'b0 ;
  assign n14871 = n10865 ^ n7479 ^ 1'b0 ;
  assign n14872 = n4696 ^ n3109 ^ 1'b0 ;
  assign n14873 = n4264 ^ n3776 ^ 1'b0 ;
  assign n14874 = n8973 & ~n11685 ;
  assign n14875 = n1391 & n14874 ;
  assign n14876 = ( n10479 & n14873 ) | ( n10479 & ~n14875 ) | ( n14873 & ~n14875 ) ;
  assign n14877 = n14872 & n14876 ;
  assign n14878 = n4914 & n14877 ;
  assign n14879 = n14878 ^ n7668 ^ n517 ;
  assign n14881 = ~n36 & n4067 ;
  assign n14882 = n8678 & ~n14881 ;
  assign n14880 = n6302 ^ n1260 ^ 1'b0 ;
  assign n14883 = n14882 ^ n14880 ^ n9839 ;
  assign n14884 = ~n57 & n4882 ;
  assign n14885 = n14884 ^ n2860 ^ 1'b0 ;
  assign n14886 = ~n13400 & n14885 ;
  assign n14887 = n14886 ^ n13632 ^ n10106 ;
  assign n14888 = n6979 ^ n5047 ^ 1'b0 ;
  assign n14889 = n20 | n14888 ;
  assign n14890 = n4416 | n14889 ;
  assign n14891 = n14890 ^ n14119 ^ 1'b0 ;
  assign n14892 = n14891 ^ n940 ^ 1'b0 ;
  assign n14893 = n7763 ^ n2835 ^ 1'b0 ;
  assign n14894 = n14893 ^ n6453 ^ 1'b0 ;
  assign n14895 = n1694 & n14894 ;
  assign n14896 = ~n9548 & n10031 ;
  assign n14897 = n9879 & n14896 ;
  assign n14898 = n5961 & n9372 ;
  assign n14899 = n368 & ~n14057 ;
  assign n14900 = n14898 & n14899 ;
  assign n14901 = n13560 | n14900 ;
  assign n14902 = n8938 | n14901 ;
  assign n14903 = ~n1407 & n6406 ;
  assign n14904 = n14903 ^ n4661 ^ 1'b0 ;
  assign n14905 = n159 | n14904 ;
  assign n14906 = ~n2084 & n5441 ;
  assign n14907 = ( ~n7208 & n7280 ) | ( ~n7208 & n12931 ) | ( n7280 & n12931 ) ;
  assign n14908 = n14907 ^ n13865 ^ 1'b0 ;
  assign n14909 = n11120 & ~n14908 ;
  assign n14910 = n10264 ^ n2184 ^ 1'b0 ;
  assign n14911 = n3351 ^ n1547 ^ 1'b0 ;
  assign n14912 = n14910 & n14911 ;
  assign n14913 = n14912 ^ n3770 ^ 1'b0 ;
  assign n14914 = n4286 | n8139 ;
  assign n14915 = n14914 ^ n6213 ^ n251 ;
  assign n14916 = n11841 | n14915 ;
  assign n14917 = n12180 ^ n6761 ^ 1'b0 ;
  assign n14918 = n9601 ^ n4099 ^ 1'b0 ;
  assign n14919 = ~n3765 & n6791 ;
  assign n14920 = n14918 | n14919 ;
  assign n14921 = n14917 & n14920 ;
  assign n14922 = ~n14916 & n14921 ;
  assign n14923 = n1339 | n2108 ;
  assign n14924 = n14923 ^ n13196 ^ 1'b0 ;
  assign n14925 = n6328 & n14924 ;
  assign n14926 = n1424 & n4228 ;
  assign n14927 = n7867 ^ n4894 ^ 1'b0 ;
  assign n14928 = ~n1172 & n14927 ;
  assign n14929 = n14926 | n14928 ;
  assign n14930 = ~n5961 & n14824 ;
  assign n14931 = n2760 & n12543 ;
  assign n14932 = n10449 | n12914 ;
  assign n14933 = n3119 ^ n37 ^ 1'b0 ;
  assign n14934 = n1495 & n14933 ;
  assign n14935 = n3007 ^ n1811 ^ 1'b0 ;
  assign n14936 = n5175 | n14935 ;
  assign n14937 = ( ~n3939 & n8662 ) | ( ~n3939 & n14936 ) | ( n8662 & n14936 ) ;
  assign n14938 = n2890 & ~n14937 ;
  assign n14939 = n7338 | n14764 ;
  assign n14940 = n4294 & ~n4689 ;
  assign n14941 = n883 & n14940 ;
  assign n14942 = n3984 | n7234 ;
  assign n14943 = n14942 ^ n13504 ^ 1'b0 ;
  assign n14944 = ~n8750 & n13157 ;
  assign n14945 = n14944 ^ n13992 ^ 1'b0 ;
  assign n14946 = ~n9192 & n14945 ;
  assign n14947 = ~n1426 & n14946 ;
  assign n14948 = ~n150 & n14299 ;
  assign n14949 = ~n7571 & n14948 ;
  assign n14950 = ~n14947 & n14949 ;
  assign n14951 = n2447 | n6420 ;
  assign n14953 = n12082 ^ n2354 ^ 1'b0 ;
  assign n14952 = n1024 & ~n14616 ;
  assign n14954 = n14953 ^ n14952 ^ 1'b0 ;
  assign n14955 = n5055 & ~n14825 ;
  assign n14956 = n14955 ^ n9224 ^ 1'b0 ;
  assign n14957 = n6021 & n6049 ;
  assign n14958 = n14957 ^ n9146 ^ 1'b0 ;
  assign n14959 = n3348 & ~n6430 ;
  assign n14960 = n13283 & n14959 ;
  assign n14961 = n5683 ^ n2124 ^ 1'b0 ;
  assign n14962 = ( n10215 & n11400 ) | ( n10215 & ~n14961 ) | ( n11400 & ~n14961 ) ;
  assign n14963 = n7203 & ~n14962 ;
  assign n14964 = n2696 & n14963 ;
  assign n14965 = n14964 ^ n8485 ^ 1'b0 ;
  assign n14966 = n2142 | n14965 ;
  assign n14967 = n935 | n14966 ;
  assign n14968 = n14967 ^ n6302 ^ n1173 ;
  assign n14969 = n14968 ^ n7752 ^ 1'b0 ;
  assign n14970 = n14238 ^ n3685 ^ 1'b0 ;
  assign n14971 = n678 & ~n3861 ;
  assign n14972 = ~n1729 & n14971 ;
  assign n14973 = n1367 & n14972 ;
  assign n14974 = ( n3370 & ~n8911 ) | ( n3370 & n14973 ) | ( ~n8911 & n14973 ) ;
  assign n14975 = n434 | n4520 ;
  assign n14976 = n4637 & n14975 ;
  assign n14977 = n14976 ^ n5707 ^ 1'b0 ;
  assign n14978 = ~n2403 & n4823 ;
  assign n14979 = n14978 ^ n1328 ^ 1'b0 ;
  assign n14980 = n654 & ~n7872 ;
  assign n14981 = n13992 ^ n469 ^ 1'b0 ;
  assign n14982 = n14981 ^ n6766 ^ 1'b0 ;
  assign n14983 = n14980 & ~n14982 ;
  assign n14984 = ~n4071 & n14983 ;
  assign n14985 = ~n14979 & n14984 ;
  assign n14986 = n8129 & ~n14985 ;
  assign n14987 = n14977 & n14986 ;
  assign n14988 = n6821 ^ n3254 ^ 1'b0 ;
  assign n14989 = n152 & n14988 ;
  assign n14990 = n14989 ^ n11853 ^ 1'b0 ;
  assign n14991 = n10795 ^ n2239 ^ n505 ;
  assign n14992 = n4338 ^ n959 ^ 1'b0 ;
  assign n14993 = ~n1423 & n14992 ;
  assign n14994 = ( n3615 & n4365 ) | ( n3615 & ~n14993 ) | ( n4365 & ~n14993 ) ;
  assign n14995 = n647 | n14994 ;
  assign n14996 = n14995 ^ n7455 ^ n3866 ;
  assign n14997 = n8301 ^ n373 ^ 1'b0 ;
  assign n15017 = n4311 | n13188 ;
  assign n15014 = n878 ^ n706 ^ 1'b0 ;
  assign n15015 = n3466 & n5280 ;
  assign n15016 = ~n15014 & n15015 ;
  assign n15018 = n15017 ^ n15016 ^ n8521 ;
  assign n14998 = n6561 ^ n3465 ^ 1'b0 ;
  assign n14999 = ~n5987 & n14998 ;
  assign n15000 = n7269 & n14999 ;
  assign n15001 = n11982 & n15000 ;
  assign n15002 = n340 & n7367 ;
  assign n15003 = n1956 & n15002 ;
  assign n15004 = n1249 & ~n15003 ;
  assign n15005 = ~n4699 & n15004 ;
  assign n15006 = ( n91 & ~n15001 ) | ( n91 & n15005 ) | ( ~n15001 & n15005 ) ;
  assign n15007 = ~n396 & n2695 ;
  assign n15008 = n5414 | n15007 ;
  assign n15009 = n4856 | n15008 ;
  assign n15010 = ~n15006 & n15009 ;
  assign n15011 = n1183 & n15010 ;
  assign n15012 = n2604 & ~n15011 ;
  assign n15013 = n13344 & n15012 ;
  assign n15019 = n15018 ^ n15013 ^ 1'b0 ;
  assign n15020 = n14997 & ~n15019 ;
  assign n15021 = n13408 ^ n12567 ^ 1'b0 ;
  assign n15022 = n9592 ^ n1856 ^ 1'b0 ;
  assign n15023 = n7280 ^ n1744 ^ 1'b0 ;
  assign n15024 = ~n12704 & n15023 ;
  assign n15025 = n9184 & n15024 ;
  assign n15026 = n4646 ^ n2418 ^ 1'b0 ;
  assign n15027 = n3982 | n15026 ;
  assign n15028 = n10441 ^ n9386 ^ 1'b0 ;
  assign n15029 = n2878 & n8292 ;
  assign n15030 = n12698 & n15029 ;
  assign n15031 = ( ~n736 & n3254 ) | ( ~n736 & n10124 ) | ( n3254 & n10124 ) ;
  assign n15032 = n14664 ^ n250 ^ 1'b0 ;
  assign n15033 = ~n374 & n14106 ;
  assign n15034 = n15033 ^ n10217 ^ 1'b0 ;
  assign n15035 = n10219 ^ n8884 ^ 1'b0 ;
  assign n15036 = ~n7272 & n15035 ;
  assign n15037 = n7020 | n13690 ;
  assign n15039 = ~n14294 & n14831 ;
  assign n15040 = n1619 & n15039 ;
  assign n15038 = n4607 | n10139 ;
  assign n15041 = n15040 ^ n15038 ^ 1'b0 ;
  assign n15042 = ( n13131 & ~n14634 ) | ( n13131 & n15041 ) | ( ~n14634 & n15041 ) ;
  assign n15043 = ( n2650 & n4801 ) | ( n2650 & n6725 ) | ( n4801 & n6725 ) ;
  assign n15044 = ( ~n15037 & n15042 ) | ( ~n15037 & n15043 ) | ( n15042 & n15043 ) ;
  assign n15045 = n13490 ^ n5418 ^ 1'b0 ;
  assign n15046 = ~n879 & n15045 ;
  assign n15047 = n12765 ^ n7011 ^ n1171 ;
  assign n15048 = ( ~n6412 & n8683 ) | ( ~n6412 & n15047 ) | ( n8683 & n15047 ) ;
  assign n15049 = n10397 & ~n14523 ;
  assign n15050 = n10111 ^ n5313 ^ 1'b0 ;
  assign n15051 = n6542 ^ n57 ^ 1'b0 ;
  assign n15052 = n9904 & ~n13155 ;
  assign n15053 = ~n6073 & n15052 ;
  assign n15054 = n3524 & ~n15053 ;
  assign n15055 = ~n15051 & n15054 ;
  assign n15056 = n7707 ^ n7400 ^ 1'b0 ;
  assign n15057 = n6781 & n15056 ;
  assign n15058 = n15057 ^ n6510 ^ 1'b0 ;
  assign n15059 = n14289 & ~n15058 ;
  assign n15060 = n15059 ^ n63 ^ 1'b0 ;
  assign n15061 = n11806 ^ n3754 ^ 1'b0 ;
  assign n15062 = ~n877 & n5173 ;
  assign n15063 = ~n15061 & n15062 ;
  assign n15064 = ( ~n909 & n1442 ) | ( ~n909 & n12339 ) | ( n1442 & n12339 ) ;
  assign n15065 = ~n12307 & n12470 ;
  assign n15066 = n696 | n10091 ;
  assign n15067 = ~n9759 & n15066 ;
  assign n15068 = n15065 & n15067 ;
  assign n15070 = n8555 ^ n1196 ^ n141 ;
  assign n15069 = n2074 & n8482 ;
  assign n15071 = n15070 ^ n15069 ^ 1'b0 ;
  assign n15072 = ( ~n1079 & n2826 ) | ( ~n1079 & n9160 ) | ( n2826 & n9160 ) ;
  assign n15073 = ~n4574 & n10865 ;
  assign n15074 = ~n9577 & n15073 ;
  assign n15075 = ( n9437 & ~n15072 ) | ( n9437 & n15074 ) | ( ~n15072 & n15074 ) ;
  assign n15076 = ~n360 & n6628 ;
  assign n15077 = n15076 ^ n7328 ^ n5541 ;
  assign n15078 = n8351 ^ n3179 ^ 1'b0 ;
  assign n15079 = n15077 | n15078 ;
  assign n15083 = n4584 ^ n4469 ^ 1'b0 ;
  assign n15084 = ~n12079 & n15083 ;
  assign n15080 = ( n1470 & n5816 ) | ( n1470 & n11241 ) | ( n5816 & n11241 ) ;
  assign n15081 = n15080 ^ n4506 ^ 1'b0 ;
  assign n15082 = n121 & ~n15081 ;
  assign n15085 = n15084 ^ n15082 ^ 1'b0 ;
  assign n15094 = n1023 | n12879 ;
  assign n15087 = n813 & n6241 ;
  assign n15088 = n5099 ^ n2993 ^ 1'b0 ;
  assign n15089 = n2072 | n15088 ;
  assign n15090 = n2084 | n15089 ;
  assign n15091 = n15090 ^ n9397 ^ 1'b0 ;
  assign n15092 = ( n575 & ~n15087 ) | ( n575 & n15091 ) | ( ~n15087 & n15091 ) ;
  assign n15093 = n9228 & n15092 ;
  assign n15095 = n15094 ^ n15093 ^ 1'b0 ;
  assign n15086 = ~n884 & n1314 ;
  assign n15096 = n15095 ^ n15086 ^ 1'b0 ;
  assign n15097 = n452 & n3637 ;
  assign n15098 = n15097 ^ n6761 ^ 1'b0 ;
  assign n15099 = n776 | n15098 ;
  assign n15100 = n1311 & ~n15099 ;
  assign n15101 = n8508 ^ n5982 ^ n156 ;
  assign n15102 = n3510 ^ n352 ^ 1'b0 ;
  assign n15103 = x0 & n7118 ;
  assign n15104 = n14073 & ~n15103 ;
  assign n15105 = n15104 ^ n2528 ^ 1'b0 ;
  assign n15106 = n15105 ^ n5370 ^ 1'b0 ;
  assign n15107 = n12515 ^ n4809 ^ 1'b0 ;
  assign n15108 = n947 | n4761 ;
  assign n15109 = ( ~n112 & n2044 ) | ( ~n112 & n15108 ) | ( n2044 & n15108 ) ;
  assign n15110 = n9457 & ~n15109 ;
  assign n15111 = n15110 ^ n9091 ^ 1'b0 ;
  assign n15112 = ( n461 & n982 ) | ( n461 & n3045 ) | ( n982 & n3045 ) ;
  assign n15113 = n4686 & ~n15112 ;
  assign n15114 = ~n10123 & n15113 ;
  assign n15115 = n15114 ^ n2995 ^ 1'b0 ;
  assign n15116 = ~n5616 & n13050 ;
  assign n15117 = n6690 & n15116 ;
  assign n15118 = n12028 | n15117 ;
  assign n15119 = n1357 ^ n1319 ^ n346 ;
  assign n15120 = ( ~n1737 & n3981 ) | ( ~n1737 & n7482 ) | ( n3981 & n7482 ) ;
  assign n15121 = n1545 | n15120 ;
  assign n15122 = n5845 | n15121 ;
  assign n15123 = ( n13766 & n15119 ) | ( n13766 & ~n15122 ) | ( n15119 & ~n15122 ) ;
  assign n15124 = n15123 ^ n14664 ^ n11952 ;
  assign n15127 = n3878 | n13778 ;
  assign n15125 = n1309 ^ n609 ^ 1'b0 ;
  assign n15126 = ~n4641 & n15125 ;
  assign n15128 = n15127 ^ n15126 ^ 1'b0 ;
  assign n15129 = n7862 & ~n15128 ;
  assign n15130 = n2453 | n11526 ;
  assign n15131 = ( n5651 & n8060 ) | ( n5651 & n15130 ) | ( n8060 & n15130 ) ;
  assign n15132 = n10919 | n15131 ;
  assign n15133 = n15132 ^ n6381 ^ 1'b0 ;
  assign n15134 = n2618 & ~n9743 ;
  assign n15135 = ~n890 & n7749 ;
  assign n15136 = n15135 ^ n5272 ^ 1'b0 ;
  assign n15137 = n15134 | n15136 ;
  assign n15138 = n15137 ^ n6369 ^ 1'b0 ;
  assign n15139 = n15138 ^ n14101 ^ 1'b0 ;
  assign n15140 = ~n14421 & n15139 ;
  assign n15141 = n12320 ^ n2687 ^ 1'b0 ;
  assign n15142 = n14937 & ~n15141 ;
  assign n15144 = n3749 ^ n2140 ^ 1'b0 ;
  assign n15143 = ~n5234 & n7058 ;
  assign n15145 = n15144 ^ n15143 ^ 1'b0 ;
  assign n15146 = n26 & n4626 ;
  assign n15151 = n1055 & ~n1895 ;
  assign n15152 = n14073 & n15151 ;
  assign n15147 = n12119 & n12285 ;
  assign n15148 = n15147 ^ n70 ^ 1'b0 ;
  assign n15149 = n13717 & ~n15148 ;
  assign n15150 = ~n10816 & n15149 ;
  assign n15153 = n15152 ^ n15150 ^ 1'b0 ;
  assign n15154 = n5803 & n6809 ;
  assign n15155 = n4233 & ~n14866 ;
  assign n15156 = ~n15154 & n15155 ;
  assign n15157 = n1177 | n15156 ;
  assign n15158 = n41 & n2529 ;
  assign n15159 = n15158 ^ n10804 ^ 1'b0 ;
  assign n15160 = ~n11729 & n15159 ;
  assign n15161 = n439 & ~n11815 ;
  assign n15162 = n10849 ^ n4574 ^ 1'b0 ;
  assign n15163 = n15161 | n15162 ;
  assign n15164 = n9494 | n15163 ;
  assign n15165 = n15164 ^ n10136 ^ n5563 ;
  assign n15166 = n6969 | n11915 ;
  assign n15167 = n289 | n1463 ;
  assign n15168 = n15167 ^ n7298 ^ n2944 ;
  assign n15169 = n4024 & n10835 ;
  assign n15170 = n15168 & n15169 ;
  assign n15171 = n7649 ^ n1436 ^ 1'b0 ;
  assign n15172 = n3355 & n15171 ;
  assign n15173 = n2479 & ~n15172 ;
  assign n15174 = n10220 ^ n8826 ^ 1'b0 ;
  assign n15175 = n15173 | n15174 ;
  assign n15176 = n13217 ^ n2885 ^ 1'b0 ;
  assign n15177 = n6166 ^ n1094 ^ 1'b0 ;
  assign n15178 = n6827 ^ n267 ^ 1'b0 ;
  assign n15179 = n3577 & ~n15178 ;
  assign n15180 = ( n5881 & n12089 ) | ( n5881 & ~n15179 ) | ( n12089 & ~n15179 ) ;
  assign n15181 = n2902 ^ n2147 ^ 1'b0 ;
  assign n15182 = n10267 ^ n3968 ^ 1'b0 ;
  assign n15183 = n10342 & ~n15182 ;
  assign n15184 = n5185 | n11708 ;
  assign n15185 = n15184 ^ n8491 ^ 1'b0 ;
  assign n15186 = n10656 & n15185 ;
  assign n15187 = ( ~n5859 & n12619 ) | ( ~n5859 & n15186 ) | ( n12619 & n15186 ) ;
  assign n15189 = n4696 ^ n2885 ^ 1'b0 ;
  assign n15188 = ~n2645 & n6551 ;
  assign n15190 = n15189 ^ n15188 ^ 1'b0 ;
  assign n15191 = ( ~n101 & n1367 ) | ( ~n101 & n7788 ) | ( n1367 & n7788 ) ;
  assign n15192 = ( n859 & n2184 ) | ( n859 & n3422 ) | ( n2184 & n3422 ) ;
  assign n15193 = ( n15190 & n15191 ) | ( n15190 & ~n15192 ) | ( n15191 & ~n15192 ) ;
  assign n15194 = ~n553 & n7465 ;
  assign n15195 = ~n2859 & n14107 ;
  assign n15196 = n8986 & ~n10830 ;
  assign n15197 = ~n14480 & n15196 ;
  assign n15198 = n9200 ^ n4052 ^ 1'b0 ;
  assign n15199 = ~n176 & n11076 ;
  assign n15200 = ( n10337 & n15198 ) | ( n10337 & n15199 ) | ( n15198 & n15199 ) ;
  assign n15201 = n637 & n5149 ;
  assign n15202 = n765 | n3370 ;
  assign n15203 = n766 | n15202 ;
  assign n15204 = n13343 & n15203 ;
  assign n15205 = n15204 ^ n2764 ^ 1'b0 ;
  assign n15206 = n11250 ^ n5202 ^ 1'b0 ;
  assign n15207 = n3519 | n10915 ;
  assign n15208 = n11908 & n15207 ;
  assign n15209 = ~n3658 & n3946 ;
  assign n15210 = n5985 & n14115 ;
  assign n15211 = n10428 & n14509 ;
  assign n15212 = ~n3888 & n15211 ;
  assign n15213 = n6535 ^ n3253 ^ 1'b0 ;
  assign n15216 = n762 & n3377 ;
  assign n15217 = n672 & n15216 ;
  assign n15214 = n3049 ^ n962 ^ 1'b0 ;
  assign n15215 = n2271 & ~n15214 ;
  assign n15218 = n15217 ^ n15215 ^ 1'b0 ;
  assign n15219 = ~n4518 & n15218 ;
  assign n15220 = n15219 ^ n2257 ^ 1'b0 ;
  assign n15221 = n7534 ^ n1011 ^ 1'b0 ;
  assign n15222 = n15220 | n15221 ;
  assign n15223 = n15213 & ~n15222 ;
  assign n15224 = n15212 & n15223 ;
  assign n15225 = n6795 ^ n6164 ^ 1'b0 ;
  assign n15226 = n6667 ^ n5665 ^ 1'b0 ;
  assign n15227 = n2751 & n15226 ;
  assign n15228 = ~n1630 & n7471 ;
  assign n15229 = ~n4275 & n7096 ;
  assign n15230 = ( n4047 & n9974 ) | ( n4047 & ~n11060 ) | ( n9974 & ~n11060 ) ;
  assign n15231 = n8818 ^ n7876 ^ 1'b0 ;
  assign n15232 = ~n15046 & n15231 ;
  assign n15233 = n12219 ^ n3305 ^ 1'b0 ;
  assign n15234 = n9740 ^ n73 ^ 1'b0 ;
  assign n15235 = ( n1186 & ~n7227 ) | ( n1186 & n15234 ) | ( ~n7227 & n15234 ) ;
  assign n15236 = ~n7471 & n15235 ;
  assign n15237 = ~n10781 & n15236 ;
  assign n15238 = n9213 ^ n3564 ^ 1'b0 ;
  assign n15239 = n1088 & ~n15238 ;
  assign n15240 = n15239 ^ n1147 ^ 1'b0 ;
  assign n15241 = ~n2143 & n6222 ;
  assign n15242 = n7763 & ~n13090 ;
  assign n15243 = n15242 ^ n4275 ^ 1'b0 ;
  assign n15244 = ( n3810 & n7742 ) | ( n3810 & ~n9296 ) | ( n7742 & ~n9296 ) ;
  assign n15245 = n687 & ~n6646 ;
  assign n15246 = ~n1666 & n15245 ;
  assign n15247 = n4427 | n6814 ;
  assign n15248 = n15246 & ~n15247 ;
  assign n15249 = ( ~n2011 & n4066 ) | ( ~n2011 & n15248 ) | ( n4066 & n15248 ) ;
  assign n15250 = n15244 & n15249 ;
  assign n15251 = n13438 & ~n15250 ;
  assign n15252 = ~n4648 & n13342 ;
  assign n15253 = n1135 | n3647 ;
  assign n15254 = n15253 ^ n1959 ^ 1'b0 ;
  assign n15255 = n15254 ^ n2993 ^ 1'b0 ;
  assign n15256 = n9933 & n15255 ;
  assign n15257 = ~n7773 & n15256 ;
  assign n15258 = n10352 ^ n8996 ^ 1'b0 ;
  assign n15259 = n2231 & n15097 ;
  assign n15260 = n9162 & n15259 ;
  assign n15261 = n15260 ^ n12388 ^ 1'b0 ;
  assign n15262 = n406 & ~n15261 ;
  assign n15263 = ~n8812 & n9358 ;
  assign n15264 = n15263 ^ n14915 ^ n7318 ;
  assign n15267 = n214 | n2731 ;
  assign n15265 = n11626 ^ n361 ^ 1'b0 ;
  assign n15266 = n4055 & n15265 ;
  assign n15268 = n15267 ^ n15266 ^ 1'b0 ;
  assign n15269 = ~n6236 & n15268 ;
  assign n15270 = n5236 ^ n3061 ^ 1'b0 ;
  assign n15271 = n5707 & ~n15270 ;
  assign n15272 = ( n349 & n12017 ) | ( n349 & n15271 ) | ( n12017 & n15271 ) ;
  assign n15273 = n8298 & ~n15272 ;
  assign n15274 = n15273 ^ n6153 ^ 1'b0 ;
  assign n15277 = n15 & n1647 ;
  assign n15275 = n2541 & n6767 ;
  assign n15276 = n713 & n15275 ;
  assign n15278 = n15277 ^ n15276 ^ 1'b0 ;
  assign n15279 = ~n9326 & n15278 ;
  assign n15280 = n15279 ^ n13569 ^ n8557 ;
  assign n15281 = n4388 & ~n11169 ;
  assign n15282 = n15281 ^ n1031 ^ 1'b0 ;
  assign n15283 = n10942 ^ n8856 ^ 1'b0 ;
  assign n15284 = n8421 ^ n2538 ^ 1'b0 ;
  assign n15285 = ~n9724 & n15284 ;
  assign n15286 = ~n12818 & n15285 ;
  assign n15287 = ~n15283 & n15286 ;
  assign n15288 = n6004 ^ n863 ^ 1'b0 ;
  assign n15289 = n1386 & n15288 ;
  assign n15290 = n15289 ^ n621 ^ 1'b0 ;
  assign n15291 = ~n3966 & n12545 ;
  assign n15292 = n7384 | n7812 ;
  assign n15293 = ~n1751 & n3720 ;
  assign n15294 = ~n7921 & n15293 ;
  assign n15295 = n13335 | n15294 ;
  assign n15296 = n15295 ^ n11258 ^ 1'b0 ;
  assign n15297 = ( n1930 & n5766 ) | ( n1930 & ~n11610 ) | ( n5766 & ~n11610 ) ;
  assign n15298 = n9519 | n15297 ;
  assign n15299 = n4192 & ~n15298 ;
  assign n15300 = n4785 ^ n503 ^ 1'b0 ;
  assign n15301 = n7192 | n15300 ;
  assign n15302 = n12051 ^ n8633 ^ 1'b0 ;
  assign n15303 = ~n15301 & n15302 ;
  assign n15304 = ~n3883 & n15303 ;
  assign n15306 = n2129 | n14112 ;
  assign n15307 = n15306 ^ n11718 ^ 1'b0 ;
  assign n15308 = n8748 & ~n15307 ;
  assign n15305 = n5533 & n10239 ;
  assign n15309 = n15308 ^ n15305 ^ 1'b0 ;
  assign n15310 = n11155 ^ n11128 ^ 1'b0 ;
  assign n15311 = n2305 & ~n15310 ;
  assign n15312 = n1804 & ~n8390 ;
  assign n15313 = n15312 ^ n82 ^ 1'b0 ;
  assign n15314 = n10631 ^ n8936 ^ 1'b0 ;
  assign n15317 = n11815 ^ n3235 ^ 1'b0 ;
  assign n15315 = n902 ^ n526 ^ 1'b0 ;
  assign n15316 = ( n2693 & n4350 ) | ( n2693 & n15315 ) | ( n4350 & n15315 ) ;
  assign n15318 = n15317 ^ n15316 ^ n3867 ;
  assign n15319 = ( n6510 & n10568 ) | ( n6510 & ~n15318 ) | ( n10568 & ~n15318 ) ;
  assign n15320 = n8911 ^ n8792 ^ n2421 ;
  assign n15321 = n15320 ^ n15066 ^ n3290 ;
  assign n15322 = n13975 ^ n3027 ^ 1'b0 ;
  assign n15323 = n15321 | n15322 ;
  assign n15324 = ( ~n2413 & n5206 ) | ( ~n2413 & n10523 ) | ( n5206 & n10523 ) ;
  assign n15325 = n1548 ^ n523 ^ 1'b0 ;
  assign n15326 = ( n9450 & ~n15324 ) | ( n9450 & n15325 ) | ( ~n15324 & n15325 ) ;
  assign n15327 = ( n2159 & ~n6101 ) | ( n2159 & n13754 ) | ( ~n6101 & n13754 ) ;
  assign n15328 = n2412 & ~n6345 ;
  assign n15329 = n1472 & ~n3828 ;
  assign n15330 = n15329 ^ n5064 ^ 1'b0 ;
  assign n15331 = n15330 ^ n13101 ^ 1'b0 ;
  assign n15332 = n601 & n7288 ;
  assign n15333 = ~n3901 & n15332 ;
  assign n15334 = ~n2334 & n12290 ;
  assign n15335 = ~n9072 & n15334 ;
  assign n15336 = n1188 & n3570 ;
  assign n15337 = n15336 ^ n14879 ^ 1'b0 ;
  assign n15338 = n1296 & n13550 ;
  assign n15339 = n14456 ^ n6302 ^ 1'b0 ;
  assign n15340 = n15338 & n15339 ;
  assign n15341 = n15340 ^ n1623 ^ 1'b0 ;
  assign n15342 = n5673 | n15341 ;
  assign n15343 = n15342 ^ n2568 ^ 1'b0 ;
  assign n15344 = n10451 ^ n4043 ^ n3883 ;
  assign n15345 = n7598 & n15344 ;
  assign n15346 = n2028 | n5748 ;
  assign n15347 = n1482 & n5202 ;
  assign n15348 = n15347 ^ n8229 ^ 1'b0 ;
  assign n15349 = ( ~n9444 & n15346 ) | ( ~n9444 & n15348 ) | ( n15346 & n15348 ) ;
  assign n15350 = n1135 | n15349 ;
  assign n15351 = n15350 ^ n13882 ^ 1'b0 ;
  assign n15352 = n15351 ^ n366 ^ 1'b0 ;
  assign n15353 = n15345 & ~n15352 ;
  assign n15354 = n678 & n7293 ;
  assign n15355 = n4657 & n15354 ;
  assign n15358 = n5001 ^ n855 ^ 1'b0 ;
  assign n15359 = ~n6460 & n15358 ;
  assign n15356 = n5924 ^ n3125 ^ 1'b0 ;
  assign n15357 = n4648 | n15356 ;
  assign n15360 = n15359 ^ n15357 ^ 1'b0 ;
  assign n15361 = n3866 | n12289 ;
  assign n15362 = n3912 | n15361 ;
  assign n15363 = ~n2664 & n15362 ;
  assign n15364 = n15363 ^ n7716 ^ 1'b0 ;
  assign n15365 = ~n5051 & n15235 ;
  assign n15366 = n12657 & n15365 ;
  assign n15369 = ~n996 & n7762 ;
  assign n15370 = ~n41 & n15369 ;
  assign n15371 = n7854 & ~n15370 ;
  assign n15372 = ( n1084 & n8491 ) | ( n1084 & ~n15371 ) | ( n8491 & ~n15371 ) ;
  assign n15367 = n14491 ^ n3959 ^ n97 ;
  assign n15368 = n3660 & n15367 ;
  assign n15373 = n15372 ^ n15368 ^ 1'b0 ;
  assign n15374 = n2995 | n6443 ;
  assign n15375 = n15373 & ~n15374 ;
  assign n15376 = n13643 ^ n4703 ^ 1'b0 ;
  assign n15377 = n15376 ^ n13131 ^ 1'b0 ;
  assign n15378 = n1826 & n15377 ;
  assign n15379 = n15378 ^ n11680 ^ 1'b0 ;
  assign n15380 = n5128 ^ n4077 ^ 1'b0 ;
  assign n15381 = n15380 ^ n2427 ^ 1'b0 ;
  assign n15382 = n4102 ^ n3397 ^ 1'b0 ;
  assign n15383 = ( ~n6639 & n9107 ) | ( ~n6639 & n15382 ) | ( n9107 & n15382 ) ;
  assign n15384 = n9496 | n13766 ;
  assign n15385 = n9829 & ~n15384 ;
  assign n15386 = n3608 | n11782 ;
  assign n15387 = ~n10685 & n15386 ;
  assign n15388 = n15385 & n15387 ;
  assign n15389 = n2679 & n5817 ;
  assign n15390 = n4259 & n15389 ;
  assign n15391 = ~n2541 & n15390 ;
  assign n15392 = ( n1122 & n6243 ) | ( n1122 & ~n15391 ) | ( n6243 & ~n15391 ) ;
  assign n15393 = n15392 ^ n2475 ^ 1'b0 ;
  assign n15394 = n15388 | n15393 ;
  assign n15395 = ~n2277 & n9437 ;
  assign n15396 = n10867 ^ n2259 ^ 1'b0 ;
  assign n15397 = n15396 ^ n1166 ^ 1'b0 ;
  assign n15398 = n15395 & ~n15397 ;
  assign n15399 = ~n4967 & n15398 ;
  assign n15400 = n697 & ~n10935 ;
  assign n15401 = n15400 ^ n3163 ^ 1'b0 ;
  assign n15402 = n4273 & n5712 ;
  assign n15403 = n750 | n8950 ;
  assign n15404 = n15402 & n15403 ;
  assign n15405 = ~n1700 & n14440 ;
  assign n15406 = n2123 & ~n9118 ;
  assign n15407 = ( x11 & ~n3473 ) | ( x11 & n8848 ) | ( ~n3473 & n8848 ) ;
  assign n15408 = n13547 ^ n9872 ^ 1'b0 ;
  assign n15409 = n12282 & ~n15408 ;
  assign n15410 = n15409 ^ n8182 ^ 1'b0 ;
  assign n15413 = n2070 | n4648 ;
  assign n15414 = n15413 ^ n7130 ^ 1'b0 ;
  assign n15411 = n6664 ^ n801 ^ n750 ;
  assign n15412 = n2296 & n15411 ;
  assign n15415 = n15414 ^ n15412 ^ 1'b0 ;
  assign n15416 = n6383 | n15415 ;
  assign n15417 = n3840 & n5660 ;
  assign n15418 = n12241 & n15417 ;
  assign n15419 = n13854 ^ n11984 ^ 1'b0 ;
  assign n15420 = n5854 & ~n15419 ;
  assign n15421 = n5309 ^ n4411 ^ 1'b0 ;
  assign n15422 = n15421 ^ n7236 ^ 1'b0 ;
  assign n15423 = ~n14452 & n15422 ;
  assign n15424 = ( ~n44 & n1638 ) | ( ~n44 & n8254 ) | ( n1638 & n8254 ) ;
  assign n15425 = ~n4516 & n10679 ;
  assign n15426 = n15425 ^ n8672 ^ 1'b0 ;
  assign n15427 = n15426 ^ n11018 ^ 1'b0 ;
  assign n15428 = n15424 | n15427 ;
  assign n15429 = n6656 & ~n10423 ;
  assign n15430 = ~n11652 & n15429 ;
  assign n15431 = n15430 ^ n2143 ^ 1'b0 ;
  assign n15435 = ~n7126 & n8747 ;
  assign n15432 = n7565 ^ n442 ^ 1'b0 ;
  assign n15433 = n15432 ^ n1638 ^ 1'b0 ;
  assign n15434 = n860 & ~n15433 ;
  assign n15436 = n15435 ^ n15434 ^ 1'b0 ;
  assign n15437 = n1207 ^ n134 ^ 1'b0 ;
  assign n15438 = n732 & ~n4799 ;
  assign n15439 = n15438 ^ n8647 ^ 1'b0 ;
  assign n15440 = n15439 ^ n9432 ^ 1'b0 ;
  assign n15441 = n15437 | n15440 ;
  assign n15442 = n3501 ^ n2934 ^ 1'b0 ;
  assign n15443 = n15442 ^ n4260 ^ 1'b0 ;
  assign n15444 = n15443 ^ n4161 ^ 1'b0 ;
  assign n15445 = n15444 ^ n4875 ^ 1'b0 ;
  assign n15446 = n7438 & n15445 ;
  assign n15447 = n2460 ^ n1180 ^ 1'b0 ;
  assign n15448 = n4515 | n15447 ;
  assign n15449 = n3271 & ~n15448 ;
  assign n15450 = ~n12382 & n15449 ;
  assign n15452 = n9683 ^ n2944 ^ n698 ;
  assign n15453 = ~n686 & n15452 ;
  assign n15454 = n1465 & n15453 ;
  assign n15451 = n1945 | n2760 ;
  assign n15455 = n15454 ^ n15451 ^ 1'b0 ;
  assign n15456 = n10356 ^ n5888 ^ n5706 ;
  assign n15457 = n15326 ^ n1875 ^ 1'b0 ;
  assign n15461 = n8801 ^ n7418 ^ n91 ;
  assign n15458 = ~n2692 & n7245 ;
  assign n15459 = n15458 ^ n4887 ^ 1'b0 ;
  assign n15460 = n11798 & ~n15459 ;
  assign n15462 = n15461 ^ n15460 ^ 1'b0 ;
  assign n15463 = ~n2787 & n7804 ;
  assign n15464 = n15463 ^ n11724 ^ 1'b0 ;
  assign n15465 = n13031 ^ n2113 ^ 1'b0 ;
  assign n15466 = n11830 & n15465 ;
  assign n15467 = n3252 | n4465 ;
  assign n15468 = n3202 & n15467 ;
  assign n15471 = n6474 ^ n6003 ^ 1'b0 ;
  assign n15472 = n2649 & n15471 ;
  assign n15469 = n1891 | n8885 ;
  assign n15470 = n13265 | n15469 ;
  assign n15473 = n15472 ^ n15470 ^ 1'b0 ;
  assign n15474 = ~n4308 & n14238 ;
  assign n15475 = n15474 ^ n4830 ^ 1'b0 ;
  assign n15476 = n451 | n2101 ;
  assign n15477 = ~n9857 & n15476 ;
  assign n15478 = ~n1348 & n14170 ;
  assign n15479 = ( ~n2993 & n5517 ) | ( ~n2993 & n13881 ) | ( n5517 & n13881 ) ;
  assign n15480 = ~n3292 & n8920 ;
  assign n15481 = n10722 & n15480 ;
  assign n15482 = n1425 | n2614 ;
  assign n15483 = n1794 | n15482 ;
  assign n15484 = n6082 | n6608 ;
  assign n15485 = n13620 & ~n15484 ;
  assign n15486 = n15483 | n15485 ;
  assign n15487 = n15486 ^ n2032 ^ n697 ;
  assign n15488 = ~n195 & n6376 ;
  assign n15489 = n15488 ^ n12495 ^ n3647 ;
  assign n15490 = n7242 ^ n208 ^ 1'b0 ;
  assign n15491 = ~n3787 & n15490 ;
  assign n15492 = ~n11762 & n15491 ;
  assign n15493 = n9959 ^ n411 ^ 1'b0 ;
  assign n15494 = n4322 & n15493 ;
  assign n15495 = n3753 & n15494 ;
  assign n15496 = n2284 & n8989 ;
  assign n15497 = n15496 ^ n9600 ^ n3170 ;
  assign n15498 = n14427 ^ n3592 ^ 1'b0 ;
  assign n15499 = n9557 ^ n4404 ^ 1'b0 ;
  assign n15500 = n2040 | n15499 ;
  assign n15501 = n15500 ^ n12878 ^ 1'b0 ;
  assign n15502 = n6133 | n6516 ;
  assign n15503 = n15502 ^ n11074 ^ 1'b0 ;
  assign n15504 = n7633 ^ n7419 ^ 1'b0 ;
  assign n15505 = ~n8449 & n15504 ;
  assign n15506 = n839 & ~n3229 ;
  assign n15507 = n15506 ^ n14902 ^ 1'b0 ;
  assign n15510 = n6978 ^ n3276 ^ 1'b0 ;
  assign n15511 = n2859 & n15510 ;
  assign n15512 = n15511 ^ n6201 ^ 1'b0 ;
  assign n15509 = n3407 ^ n2449 ^ 1'b0 ;
  assign n15508 = ~n6433 & n14418 ;
  assign n15513 = n15512 ^ n15509 ^ n15508 ;
  assign n15515 = n10851 ^ n4962 ^ 1'b0 ;
  assign n15516 = n15461 | n15515 ;
  assign n15514 = ~n296 & n9507 ;
  assign n15517 = n15516 ^ n15514 ^ 1'b0 ;
  assign n15518 = ( ~n145 & n9110 ) | ( ~n145 & n15517 ) | ( n9110 & n15517 ) ;
  assign n15519 = n10857 ^ n6431 ^ 1'b0 ;
  assign n15520 = n6607 | n15519 ;
  assign n15521 = n4622 & n8998 ;
  assign n15522 = n514 & n15521 ;
  assign n15523 = n10898 ^ n8017 ^ n352 ;
  assign n15524 = n13103 & n13136 ;
  assign n15525 = n10744 & n15524 ;
  assign n15526 = n2471 & n14365 ;
  assign n15527 = n15526 ^ n1546 ^ 1'b0 ;
  assign n15528 = n10807 ^ n5157 ^ 1'b0 ;
  assign n15529 = n3564 ^ n2619 ^ n41 ;
  assign n15530 = n471 | n8952 ;
  assign n15531 = n3787 & ~n15530 ;
  assign n15532 = n13404 ^ n4944 ^ 1'b0 ;
  assign n15533 = ~n15531 & n15532 ;
  assign n15534 = n11450 ^ n2334 ^ 1'b0 ;
  assign n15535 = n6973 & ~n8826 ;
  assign n15536 = n10700 ^ n5301 ^ 1'b0 ;
  assign n15537 = n15535 & n15536 ;
  assign n15538 = n631 | n756 ;
  assign n15539 = n631 & ~n15538 ;
  assign n15540 = n4120 & ~n15539 ;
  assign n15541 = n15539 & n15540 ;
  assign n15542 = ( n2923 & ~n3307 ) | ( n2923 & n14772 ) | ( ~n3307 & n14772 ) ;
  assign n15543 = n3312 & n15542 ;
  assign n15544 = n15543 ^ n2618 ^ 1'b0 ;
  assign n15545 = n15544 ^ n7659 ^ 1'b0 ;
  assign n15546 = ~n15541 & n15545 ;
  assign n15547 = n2569 & ~n2923 ;
  assign n15548 = ~n5969 & n15547 ;
  assign n15549 = n1591 | n15548 ;
  assign n15550 = n11227 & ~n15549 ;
  assign n15551 = ~n2466 & n3888 ;
  assign n15552 = n15551 ^ n2104 ^ 1'b0 ;
  assign n15553 = n12509 ^ n3343 ^ 1'b0 ;
  assign n15554 = n15552 & ~n15553 ;
  assign n15555 = n9929 & n12854 ;
  assign n15556 = n15555 ^ n4562 ^ 1'b0 ;
  assign n15557 = n6949 | n15556 ;
  assign n15558 = n15454 ^ n14504 ^ n2831 ;
  assign n15559 = n9452 ^ n9220 ^ 1'b0 ;
  assign n15560 = n5543 & ~n15559 ;
  assign n15561 = n8863 ^ n1089 ^ 1'b0 ;
  assign n15562 = n1414 | n15561 ;
  assign n15563 = ( n2601 & n2678 ) | ( n2601 & n3202 ) | ( n2678 & n3202 ) ;
  assign n15564 = n786 & n15563 ;
  assign n15565 = n15562 | n15564 ;
  assign n15566 = n2677 & n5645 ;
  assign n15567 = n6098 ^ n2989 ^ 1'b0 ;
  assign n15568 = n627 | n15567 ;
  assign n15569 = n10094 & n15568 ;
  assign n15570 = n2686 & ~n15569 ;
  assign n15571 = ~n13084 & n15570 ;
  assign n15572 = n5745 | n8881 ;
  assign n15573 = n5854 & ~n15572 ;
  assign n15574 = ( n4544 & n11701 ) | ( n4544 & n14097 ) | ( n11701 & n14097 ) ;
  assign n15575 = n4640 & ~n9281 ;
  assign n15576 = n8130 & n15575 ;
  assign n15577 = n1616 | n15576 ;
  assign n15578 = n1658 | n2304 ;
  assign n15579 = ( x3 & n15577 ) | ( x3 & ~n15578 ) | ( n15577 & ~n15578 ) ;
  assign n15580 = ( n4220 & n7089 ) | ( n4220 & n12269 ) | ( n7089 & n12269 ) ;
  assign n15581 = n6221 | n15580 ;
  assign n15582 = n6034 ^ n452 ^ 1'b0 ;
  assign n15583 = n839 ^ n645 ^ 1'b0 ;
  assign n15584 = n2731 & n15583 ;
  assign n15585 = n15584 ^ n14343 ^ n14035 ;
  assign n15586 = n6466 ^ n1591 ^ 1'b0 ;
  assign n15587 = ~n3295 & n15586 ;
  assign n15588 = n1000 & n15587 ;
  assign n15589 = n9750 & n15588 ;
  assign n15590 = n995 & n2258 ;
  assign n15591 = ( n6787 & n10824 ) | ( n6787 & ~n11757 ) | ( n10824 & ~n11757 ) ;
  assign n15592 = n15591 ^ n11798 ^ 1'b0 ;
  assign n15599 = n1250 | n6350 ;
  assign n15600 = n15599 ^ n13509 ^ 1'b0 ;
  assign n15593 = n1463 | n6991 ;
  assign n15594 = n596 | n15593 ;
  assign n15595 = n12097 | n15594 ;
  assign n15596 = n1791 & n15595 ;
  assign n15597 = n5048 & n15596 ;
  assign n15598 = n3864 & ~n15597 ;
  assign n15601 = n15600 ^ n15598 ^ 1'b0 ;
  assign n15602 = n7495 ^ n2986 ^ 1'b0 ;
  assign n15603 = n15602 ^ n3635 ^ 1'b0 ;
  assign n15604 = n15601 | n15603 ;
  assign n15605 = n8077 ^ n6336 ^ 1'b0 ;
  assign n15606 = n4197 ^ n3245 ^ 1'b0 ;
  assign n15607 = ~n2075 & n15606 ;
  assign n15608 = n15605 & n15607 ;
  assign n15610 = n1444 & ~n1815 ;
  assign n15611 = ( n3619 & n8727 ) | ( n3619 & ~n8902 ) | ( n8727 & ~n8902 ) ;
  assign n15612 = n15610 & ~n15611 ;
  assign n15609 = n7292 | n13426 ;
  assign n15613 = n15612 ^ n15609 ^ 1'b0 ;
  assign n15614 = ( n408 & n2214 ) | ( n408 & n11763 ) | ( n2214 & n11763 ) ;
  assign n15615 = n15614 ^ n12730 ^ n418 ;
  assign n15616 = n10758 ^ n78 ^ 1'b0 ;
  assign n15617 = n2544 & n15616 ;
  assign n15618 = ( n5233 & ~n8126 ) | ( n5233 & n15617 ) | ( ~n8126 & n15617 ) ;
  assign n15619 = n9113 & n15618 ;
  assign n15620 = n15619 ^ n13009 ^ 1'b0 ;
  assign n15621 = ( n9485 & ~n15615 ) | ( n9485 & n15620 ) | ( ~n15615 & n15620 ) ;
  assign n15622 = n12180 ^ n5175 ^ 1'b0 ;
  assign n15623 = n2428 & ~n15622 ;
  assign n15624 = n15623 ^ n11718 ^ 1'b0 ;
  assign n15625 = n4971 ^ n3510 ^ 1'b0 ;
  assign n15626 = ~n448 & n15625 ;
  assign n15627 = n15626 ^ n4605 ^ 1'b0 ;
  assign n15628 = n15627 ^ n13697 ^ 1'b0 ;
  assign n15629 = n11905 ^ n6050 ^ 1'b0 ;
  assign n15630 = n6827 | n15629 ;
  assign n15631 = n8976 ^ n1263 ^ 1'b0 ;
  assign n15632 = n5323 & ~n11779 ;
  assign n15633 = n398 | n6509 ;
  assign n15634 = n15632 & ~n15633 ;
  assign n15635 = n15631 | n15634 ;
  assign n15636 = n6036 & ~n15635 ;
  assign n15637 = n15630 & ~n15636 ;
  assign n15638 = n5781 & n13218 ;
  assign n15639 = n4477 | n15638 ;
  assign n15640 = n4041 | n15639 ;
  assign n15641 = ( n3027 & ~n3114 ) | ( n3027 & n3923 ) | ( ~n3114 & n3923 ) ;
  assign n15642 = n4650 & ~n15641 ;
  assign n15643 = ~n3976 & n15642 ;
  assign n15644 = n6071 ^ n1181 ^ 1'b0 ;
  assign n15645 = ~n672 & n15644 ;
  assign n15646 = n15391 | n15645 ;
  assign n15647 = ( ~n13263 & n15643 ) | ( ~n13263 & n15646 ) | ( n15643 & n15646 ) ;
  assign n15648 = n2597 & n15198 ;
  assign n15649 = n15648 ^ n7639 ^ 1'b0 ;
  assign n15650 = n13019 & n15649 ;
  assign n15651 = n10467 ^ n3832 ^ 1'b0 ;
  assign n15652 = n10835 ^ n7492 ^ n7388 ;
  assign n15653 = ( ~n6846 & n8260 ) | ( ~n6846 & n11894 ) | ( n8260 & n11894 ) ;
  assign n15656 = ~n2264 & n2665 ;
  assign n15657 = n1545 & n15656 ;
  assign n15658 = n8164 | n15657 ;
  assign n15659 = n4920 & ~n15658 ;
  assign n15654 = n11769 ^ n8976 ^ n3437 ;
  assign n15655 = n14272 & ~n15654 ;
  assign n15660 = n15659 ^ n15655 ^ 1'b0 ;
  assign n15661 = n10459 & n11781 ;
  assign n15662 = n9097 & n15661 ;
  assign n15663 = n4345 & n15662 ;
  assign n15664 = n14144 ^ n2591 ^ 1'b0 ;
  assign n15665 = n7493 | n15664 ;
  assign n15666 = n15665 ^ n5607 ^ n157 ;
  assign n15667 = ( n4577 & n7198 ) | ( n4577 & ~n13899 ) | ( n7198 & ~n13899 ) ;
  assign n15668 = n6770 ^ n75 ^ 1'b0 ;
  assign n15669 = ~n15667 & n15668 ;
  assign n15670 = n8607 ^ n1436 ^ 1'b0 ;
  assign n15671 = n15670 ^ n13184 ^ 1'b0 ;
  assign n15672 = n9143 ^ n7584 ^ 1'b0 ;
  assign n15675 = n4977 ^ n2705 ^ 1'b0 ;
  assign n15676 = n3923 & ~n15675 ;
  assign n15677 = n15676 ^ n9042 ^ 1'b0 ;
  assign n15673 = n1218 & ~n2248 ;
  assign n15674 = n9528 & n15673 ;
  assign n15678 = n15677 ^ n15674 ^ 1'b0 ;
  assign n15679 = n4590 | n12800 ;
  assign n15680 = n3713 ^ n67 ^ 1'b0 ;
  assign n15681 = n12084 ^ n991 ^ 1'b0 ;
  assign n15682 = n4144 & n15681 ;
  assign n15683 = n14665 | n15682 ;
  assign n15684 = ( n208 & n2944 ) | ( n208 & ~n3043 ) | ( n2944 & ~n3043 ) ;
  assign n15685 = n13932 ^ n12717 ^ n5085 ;
  assign n15686 = n3336 ^ n541 ^ 1'b0 ;
  assign n15687 = ~n5885 & n15686 ;
  assign n15688 = n2067 ^ n465 ^ 1'b0 ;
  assign n15689 = n15688 ^ n1764 ^ 1'b0 ;
  assign n15690 = n15687 & ~n15689 ;
  assign n15691 = n15690 ^ n5017 ^ 1'b0 ;
  assign n15692 = n3812 & ~n15691 ;
  assign n15693 = n5745 | n6440 ;
  assign n15694 = n11562 & ~n15693 ;
  assign n15695 = n15694 ^ n3056 ^ 1'b0 ;
  assign n15696 = n12024 ^ n4607 ^ 1'b0 ;
  assign n15697 = n1959 ^ n306 ^ 1'b0 ;
  assign n15699 = n324 & n2431 ;
  assign n15700 = n1201 & n15699 ;
  assign n15701 = n15700 ^ n649 ^ 1'b0 ;
  assign n15698 = n1596 & ~n6727 ;
  assign n15702 = n15701 ^ n15698 ^ 1'b0 ;
  assign n15703 = n15697 | n15702 ;
  assign n15704 = n15703 ^ n5113 ^ 1'b0 ;
  assign n15713 = n955 | n7325 ;
  assign n15714 = n797 & ~n15713 ;
  assign n15711 = n1943 & ~n5156 ;
  assign n15712 = n15711 ^ n8409 ^ 1'b0 ;
  assign n15715 = n15714 ^ n15712 ^ n12728 ;
  assign n15708 = n3174 ^ n2372 ^ 1'b0 ;
  assign n15705 = n4791 | n9362 ;
  assign n15706 = n12635 ^ n3085 ^ 1'b0 ;
  assign n15707 = n15705 | n15706 ;
  assign n15709 = n15708 ^ n15707 ^ 1'b0 ;
  assign n15710 = ~n11833 & n15709 ;
  assign n15716 = n15715 ^ n15710 ^ 1'b0 ;
  assign n15721 = n592 & n4167 ;
  assign n15722 = ~n592 & n15721 ;
  assign n15717 = n542 | n8210 ;
  assign n15718 = n15717 ^ n5014 ^ 1'b0 ;
  assign n15719 = n15718 ^ n1912 ^ 1'b0 ;
  assign n15720 = ~n13726 & n15719 ;
  assign n15723 = n15722 ^ n15720 ^ 1'b0 ;
  assign n15724 = n7927 & ~n15723 ;
  assign n15725 = n1395 | n9583 ;
  assign n15726 = n15725 ^ n1457 ^ 1'b0 ;
  assign n15727 = n13528 ^ n6551 ^ 1'b0 ;
  assign n15728 = n15726 & n15727 ;
  assign n15729 = n3332 ^ n2102 ^ n1206 ;
  assign n15730 = ( ~n208 & n9973 ) | ( ~n208 & n15729 ) | ( n9973 & n15729 ) ;
  assign n15731 = ~n72 & n11571 ;
  assign n15732 = n15731 ^ n6743 ^ 1'b0 ;
  assign n15733 = n15732 ^ n3987 ^ 1'b0 ;
  assign n15734 = ( ~n2005 & n2186 ) | ( ~n2005 & n4399 ) | ( n2186 & n4399 ) ;
  assign n15735 = ( ~n8861 & n8970 ) | ( ~n8861 & n15734 ) | ( n8970 & n15734 ) ;
  assign n15736 = n1586 & n3435 ;
  assign n15737 = ( n1023 & n11701 ) | ( n1023 & ~n15736 ) | ( n11701 & ~n15736 ) ;
  assign n15738 = n15737 ^ n11288 ^ 1'b0 ;
  assign n15739 = n15735 | n15738 ;
  assign n15740 = ~n14409 & n15715 ;
  assign n15741 = n15740 ^ n9827 ^ 1'b0 ;
  assign n15742 = ~n3373 & n10452 ;
  assign n15743 = ~n1461 & n8622 ;
  assign n15744 = ~n5693 & n15743 ;
  assign n15745 = n2377 & ~n12936 ;
  assign n15746 = n15745 ^ n12954 ^ 1'b0 ;
  assign n15747 = n15744 | n15746 ;
  assign n15748 = n14548 & ~n15747 ;
  assign n15749 = n5225 | n13545 ;
  assign n15750 = n7386 | n12347 ;
  assign n15751 = n6107 | n15750 ;
  assign n15752 = n8110 & ~n15751 ;
  assign n15753 = n251 | n5545 ;
  assign n15754 = n2130 & n15753 ;
  assign n15755 = n3127 ^ n270 ^ 1'b0 ;
  assign n15756 = n5465 & n15755 ;
  assign n15757 = n7550 ^ n2678 ^ 1'b0 ;
  assign n15758 = ~n4230 & n15757 ;
  assign n15759 = ~n15756 & n15758 ;
  assign n15760 = n5159 & ~n6711 ;
  assign n15761 = n15760 ^ n1967 ^ 1'b0 ;
  assign n15762 = n5377 | n15761 ;
  assign n15763 = n15762 ^ n1959 ^ 1'b0 ;
  assign n15764 = n10037 ^ n1255 ^ 1'b0 ;
  assign n15765 = n15763 & ~n15764 ;
  assign n15766 = n6134 | n13107 ;
  assign n15767 = n15766 ^ n7676 ^ 1'b0 ;
  assign n15768 = n1784 & ~n15767 ;
  assign n15769 = n15768 ^ n481 ^ 1'b0 ;
  assign n15770 = n15769 ^ n15231 ^ 1'b0 ;
  assign n15771 = n11632 ^ n2338 ^ 1'b0 ;
  assign n15772 = n3216 | n15771 ;
  assign n15773 = n2979 & n5603 ;
  assign n15774 = n15772 & n15773 ;
  assign n15775 = ( n12548 & ~n12787 ) | ( n12548 & n15774 ) | ( ~n12787 & n15774 ) ;
  assign n15776 = n1572 ^ n501 ^ 1'b0 ;
  assign n15777 = n156 | n15776 ;
  assign n15778 = n4104 & n9955 ;
  assign n15779 = ~n415 & n15778 ;
  assign n15780 = n15779 ^ n2832 ^ 1'b0 ;
  assign n15781 = n656 & ~n6424 ;
  assign n15782 = ~n14219 & n15781 ;
  assign n15783 = n15780 & n15782 ;
  assign n15784 = n15783 ^ n11387 ^ 1'b0 ;
  assign n15785 = n2939 ^ n611 ^ 1'b0 ;
  assign n15786 = n8920 ^ n5504 ^ 1'b0 ;
  assign n15787 = ~n5488 & n15786 ;
  assign n15788 = n372 | n7876 ;
  assign n15789 = ( ~n3575 & n15787 ) | ( ~n3575 & n15788 ) | ( n15787 & n15788 ) ;
  assign n15790 = n276 | n3523 ;
  assign n15791 = n1988 & ~n15790 ;
  assign n15792 = n15791 ^ n4720 ^ 1'b0 ;
  assign n15793 = n11688 & ~n12187 ;
  assign n15794 = n15793 ^ n14484 ^ 1'b0 ;
  assign n15795 = n8099 & ~n15794 ;
  assign n15796 = ~n326 & n15795 ;
  assign n15797 = n8612 ^ n6369 ^ 1'b0 ;
  assign n15800 = n3776 & ~n6024 ;
  assign n15801 = n12375 & ~n15800 ;
  assign n15802 = ( n954 & ~n10129 ) | ( n954 & n15801 ) | ( ~n10129 & n15801 ) ;
  assign n15798 = ~n220 & n4281 ;
  assign n15799 = ~n13279 & n15798 ;
  assign n15803 = n15802 ^ n15799 ^ 1'b0 ;
  assign n15804 = n10145 ^ n1336 ^ 1'b0 ;
  assign n15805 = n12166 ^ n4394 ^ n844 ;
  assign n15806 = n15805 ^ n9526 ^ 1'b0 ;
  assign n15807 = ~n15804 & n15806 ;
  assign n15808 = ~x3 & n8595 ;
  assign n15809 = n12038 & n15808 ;
  assign n15810 = ~n736 & n8662 ;
  assign n15811 = n15810 ^ n4369 ^ 1'b0 ;
  assign n15812 = ~n6816 & n10780 ;
  assign n15813 = n15811 & n15812 ;
  assign n15814 = n7798 ^ n4830 ^ 1'b0 ;
  assign n15815 = n108 & ~n15814 ;
  assign n15816 = n4280 ^ n3995 ^ n57 ;
  assign n15817 = n5380 ^ n191 ^ 1'b0 ;
  assign n15818 = n2211 & ~n5045 ;
  assign n15819 = ~n2176 & n15818 ;
  assign n15820 = ( n2825 & ~n15568 ) | ( n2825 & n15819 ) | ( ~n15568 & n15819 ) ;
  assign n15824 = n4158 ^ n947 ^ 1'b0 ;
  assign n15825 = n7752 & n15824 ;
  assign n15826 = n15825 ^ n5350 ^ 1'b0 ;
  assign n15827 = ( ~n82 & n9175 ) | ( ~n82 & n15826 ) | ( n9175 & n15826 ) ;
  assign n15828 = n1122 | n10509 ;
  assign n15829 = n3661 & ~n15828 ;
  assign n15830 = ( n149 & n7130 ) | ( n149 & n15829 ) | ( n7130 & n15829 ) ;
  assign n15831 = n2986 | n15830 ;
  assign n15832 = ( n5098 & n15827 ) | ( n5098 & n15831 ) | ( n15827 & n15831 ) ;
  assign n15821 = n7931 ^ n5591 ^ n3517 ;
  assign n15822 = n13594 & n15821 ;
  assign n15823 = ~n2644 & n15822 ;
  assign n15833 = n15832 ^ n15823 ^ 1'b0 ;
  assign n15834 = n12717 ^ n11137 ^ 1'b0 ;
  assign n15835 = n4024 | n15834 ;
  assign n15836 = ( ~n6341 & n11798 ) | ( ~n6341 & n12162 ) | ( n11798 & n12162 ) ;
  assign n15837 = n5841 ^ n1760 ^ n376 ;
  assign n15838 = ( ~n7653 & n12853 ) | ( ~n7653 & n15837 ) | ( n12853 & n15837 ) ;
  assign n15839 = n15838 ^ n287 ^ 1'b0 ;
  assign n15840 = n5934 | n8356 ;
  assign n15841 = n8919 & ~n15840 ;
  assign n15842 = n1453 & ~n15841 ;
  assign n15843 = n15842 ^ n12657 ^ 1'b0 ;
  assign n15844 = n13280 & ~n15388 ;
  assign n15845 = n15844 ^ n62 ^ 1'b0 ;
  assign n15846 = n4551 | n10533 ;
  assign n15848 = n3345 | n6833 ;
  assign n15849 = n15848 ^ n1752 ^ 1'b0 ;
  assign n15847 = n523 & ~n3303 ;
  assign n15850 = n15849 ^ n15847 ^ 1'b0 ;
  assign n15851 = n15850 ^ n4880 ^ n1118 ;
  assign n15852 = n80 & n15851 ;
  assign n15853 = n8479 ^ n4982 ^ 1'b0 ;
  assign n15854 = n14002 | n15853 ;
  assign n15855 = n100 & n4970 ;
  assign n15856 = n15855 ^ n6221 ^ 1'b0 ;
  assign n15857 = ~n15854 & n15856 ;
  assign n15858 = n676 & ~n12515 ;
  assign n15859 = n104 & n15858 ;
  assign n15860 = n15859 ^ n10721 ^ 1'b0 ;
  assign n15861 = n3022 & n15860 ;
  assign n15862 = n1483 & ~n4797 ;
  assign n15863 = ~n11698 & n15862 ;
  assign n15864 = n1900 ^ n961 ^ 1'b0 ;
  assign n15867 = n9020 ^ n6895 ^ 1'b0 ;
  assign n15868 = n1658 ^ n1048 ^ 1'b0 ;
  assign n15869 = ~n13721 & n15868 ;
  assign n15870 = n15867 & n15869 ;
  assign n15865 = n2067 & ~n2859 ;
  assign n15866 = ~n1596 & n15865 ;
  assign n15871 = n15870 ^ n15866 ^ n5178 ;
  assign n15872 = n2919 | n10737 ;
  assign n15873 = n7921 & ~n15872 ;
  assign n15874 = ~n13537 & n15873 ;
  assign n15875 = n2228 & ~n8442 ;
  assign n15876 = n15874 & n15875 ;
  assign n15877 = n15490 ^ n8298 ^ 1'b0 ;
  assign n15878 = n12321 & n15877 ;
  assign n15879 = n15878 ^ n9743 ^ 1'b0 ;
  assign n15880 = n12006 | n13703 ;
  assign n15881 = n6554 & n8587 ;
  assign n15882 = n15881 ^ n11612 ^ 1'b0 ;
  assign n15883 = ~n9450 & n13239 ;
  assign n15884 = n5965 & n15883 ;
  assign n15885 = n7778 ^ n4612 ^ n3792 ;
  assign n15886 = n525 & n15885 ;
  assign n15888 = n1245 & ~n5017 ;
  assign n15889 = n15888 ^ n7678 ^ 1'b0 ;
  assign n15887 = n8590 & ~n13567 ;
  assign n15890 = n15889 ^ n15887 ^ 1'b0 ;
  assign n15893 = ~n3459 & n13968 ;
  assign n15894 = ~n14918 & n15893 ;
  assign n15891 = n6196 & n13198 ;
  assign n15892 = n15891 ^ n8622 ^ 1'b0 ;
  assign n15895 = n15894 ^ n15892 ^ 1'b0 ;
  assign n15896 = n1432 & ~n2858 ;
  assign n15897 = n15896 ^ n14102 ^ 1'b0 ;
  assign n15898 = ( ~n2187 & n2648 ) | ( ~n2187 & n3343 ) | ( n2648 & n3343 ) ;
  assign n15902 = ~n1461 & n12304 ;
  assign n15903 = n15902 ^ n1809 ^ 1'b0 ;
  assign n15899 = n2695 | n11892 ;
  assign n15900 = n15899 ^ n3241 ^ 1'b0 ;
  assign n15901 = n15272 | n15900 ;
  assign n15904 = n15903 ^ n15901 ^ 1'b0 ;
  assign n15905 = n15904 ^ n4450 ^ 1'b0 ;
  assign n15906 = ~n5339 & n15905 ;
  assign n15907 = ~n11363 & n15906 ;
  assign n15908 = n6340 & ~n15907 ;
  assign n15909 = ~n15898 & n15908 ;
  assign n15910 = n15909 ^ n13760 ^ 1'b0 ;
  assign n15911 = n2330 & n7902 ;
  assign n15912 = n2457 & n11283 ;
  assign n15913 = ~n2645 & n8342 ;
  assign n15914 = n13567 & n15913 ;
  assign n15915 = n4088 & ~n15914 ;
  assign n15916 = ( n3693 & ~n8041 ) | ( n3693 & n15915 ) | ( ~n8041 & n15915 ) ;
  assign n15917 = ~n545 & n5249 ;
  assign n15918 = n15917 ^ n9401 ^ 1'b0 ;
  assign n15919 = n13580 ^ n1779 ^ 1'b0 ;
  assign n15920 = n7203 ^ n4086 ^ 1'b0 ;
  assign n15921 = n563 | n15920 ;
  assign n15922 = n8031 & n13503 ;
  assign n15923 = n15922 ^ n10217 ^ 1'b0 ;
  assign n15924 = n13504 | n15923 ;
  assign n15925 = n1818 & ~n15924 ;
  assign n15926 = ~n6221 & n12932 ;
  assign n15927 = n63 & n7225 ;
  assign n15928 = n15927 ^ n2878 ^ 1'b0 ;
  assign n15929 = n7150 & ~n15928 ;
  assign n15930 = n15929 ^ n7689 ^ 1'b0 ;
  assign n15931 = ~n3725 & n6208 ;
  assign n15932 = n6380 ^ n6091 ^ 1'b0 ;
  assign n15933 = n4085 & n15932 ;
  assign n15934 = n11169 | n15933 ;
  assign n15935 = ~n6584 & n15934 ;
  assign n15936 = ~n7427 & n15935 ;
  assign n15937 = n8655 ^ n3134 ^ n892 ;
  assign n15938 = n346 & ~n4490 ;
  assign n15939 = n11782 & n15938 ;
  assign n15940 = n15939 ^ n10053 ^ 1'b0 ;
  assign n15941 = n15940 ^ n2920 ^ 1'b0 ;
  assign n15942 = n3093 | n15941 ;
  assign n15943 = n13121 & n15942 ;
  assign n15944 = n3817 ^ n126 ^ 1'b0 ;
  assign n15945 = n3127 ^ n2989 ^ 1'b0 ;
  assign n15946 = n15944 & ~n15945 ;
  assign n15947 = n15946 ^ n2139 ^ 1'b0 ;
  assign n15948 = n11609 & ~n15947 ;
  assign n15949 = ~n1709 & n15948 ;
  assign n15950 = n10998 ^ n915 ^ n287 ;
  assign n15951 = n15950 ^ n9595 ^ n2169 ;
  assign n15952 = n15951 ^ n8188 ^ n5311 ;
  assign n15953 = n11897 ^ n1751 ^ n533 ;
  assign n15954 = n2223 | n15953 ;
  assign n15955 = n9659 | n15954 ;
  assign n15956 = ~n3455 & n8885 ;
  assign n15957 = n854 & n15956 ;
  assign n15958 = n15957 ^ n4454 ^ 1'b0 ;
  assign n15959 = ( n1503 & n13493 ) | ( n1503 & n15958 ) | ( n13493 & n15958 ) ;
  assign n15960 = n8138 ^ n7943 ^ 1'b0 ;
  assign n15961 = n13228 ^ n1276 ^ 1'b0 ;
  assign n15962 = n4823 & n15961 ;
  assign n15963 = ~n7051 & n8676 ;
  assign n15964 = ~n7598 & n11608 ;
  assign n15965 = ~n15042 & n15964 ;
  assign n15966 = ( n5003 & ~n15963 ) | ( n5003 & n15965 ) | ( ~n15963 & n15965 ) ;
  assign n15967 = n7053 & n14052 ;
  assign n15969 = n6159 ^ n2713 ^ 1'b0 ;
  assign n15968 = ~n216 & n10529 ;
  assign n15970 = n15969 ^ n15968 ^ 1'b0 ;
  assign n15971 = n4239 & ~n15970 ;
  assign n15972 = n11954 ^ n11608 ^ 1'b0 ;
  assign n15973 = n2182 ^ n823 ^ n414 ;
  assign n15974 = n294 | n3293 ;
  assign n15975 = n4351 & ~n15974 ;
  assign n15976 = n9713 | n15975 ;
  assign n15977 = n8621 ^ n2756 ^ 1'b0 ;
  assign n15978 = n1448 | n2276 ;
  assign n15979 = n15978 ^ n962 ^ 1'b0 ;
  assign n15980 = ~n6262 & n15979 ;
  assign n15981 = n15980 ^ n15385 ^ 1'b0 ;
  assign n15982 = ( n1234 & n1781 ) | ( n1234 & n5699 ) | ( n1781 & n5699 ) ;
  assign n15983 = n8474 & n15982 ;
  assign n15984 = n8275 & n15983 ;
  assign n15986 = n204 ^ n192 ^ 1'b0 ;
  assign n15987 = n15986 ^ n4010 ^ n2118 ;
  assign n15985 = ~n4754 & n13754 ;
  assign n15988 = n15987 ^ n15985 ^ 1'b0 ;
  assign n15989 = n15574 ^ n6485 ^ 1'b0 ;
  assign n15990 = n6614 ^ n26 ^ 1'b0 ;
  assign n15991 = n14125 ^ n1228 ^ n670 ;
  assign n15992 = n2374 & ~n10017 ;
  assign n15993 = n859 & n15992 ;
  assign n15994 = n1436 & n15993 ;
  assign n15995 = n11924 ^ n5240 ^ 1'b0 ;
  assign n15996 = n361 | n4341 ;
  assign n15997 = n2651 & n15359 ;
  assign n15998 = n2114 & n10267 ;
  assign n15999 = n15998 ^ n1666 ^ 1'b0 ;
  assign n16000 = n15999 ^ n14462 ^ n2560 ;
  assign n16001 = n4165 ^ n661 ^ 1'b0 ;
  assign n16002 = n16001 ^ n10701 ^ 1'b0 ;
  assign n16003 = n7545 & n16002 ;
  assign n16004 = ( n3016 & n5774 ) | ( n3016 & ~n16003 ) | ( n5774 & ~n16003 ) ;
  assign n16005 = n1926 | n9164 ;
  assign n16006 = n13542 ^ n12622 ^ 1'b0 ;
  assign n16007 = n14824 ^ n1647 ^ 1'b0 ;
  assign n16008 = ( n711 & n2994 ) | ( n711 & ~n16007 ) | ( n2994 & ~n16007 ) ;
  assign n16010 = n12935 ^ n6522 ^ 1'b0 ;
  assign n16009 = n6766 & n14514 ;
  assign n16011 = n16010 ^ n16009 ^ 1'b0 ;
  assign n16012 = n9027 & n10212 ;
  assign n16013 = n502 | n15602 ;
  assign n16014 = n16012 | n16013 ;
  assign n16015 = n906 | n11690 ;
  assign n16016 = n16015 ^ n8379 ^ 1'b0 ;
  assign n16017 = n797 & ~n2561 ;
  assign n16018 = ~n16016 & n16017 ;
  assign n16019 = n16018 ^ n2447 ^ 1'b0 ;
  assign n16020 = n7858 ^ n583 ^ 1'b0 ;
  assign n16021 = n1706 & ~n16020 ;
  assign n16022 = n5508 | n6205 ;
  assign n16023 = n16021 | n16022 ;
  assign n16024 = n13210 ^ n159 ^ 1'b0 ;
  assign n16025 = n10527 | n14597 ;
  assign n16026 = n4485 & n16025 ;
  assign n16027 = n16026 ^ n10751 ^ 1'b0 ;
  assign n16028 = n15493 ^ n6296 ^ 1'b0 ;
  assign n16029 = n2503 | n16028 ;
  assign n16030 = n1039 & ~n16029 ;
  assign n16031 = n15074 ^ n4387 ^ 1'b0 ;
  assign n16032 = n9433 & ~n16031 ;
  assign n16033 = n12415 ^ n11538 ^ 1'b0 ;
  assign n16034 = n1167 & n13257 ;
  assign n16035 = n16034 ^ n10254 ^ 1'b0 ;
  assign n16036 = n12693 | n13124 ;
  assign n16037 = n10839 ^ n6732 ^ 1'b0 ;
  assign n16038 = n6435 | n16037 ;
  assign n16039 = n16038 ^ n3261 ^ 1'b0 ;
  assign n16040 = n14531 & ~n16039 ;
  assign n16041 = ~n7790 & n16040 ;
  assign n16042 = n3264 & n8542 ;
  assign n16043 = n2766 & n4633 ;
  assign n16044 = n3812 & n16043 ;
  assign n16045 = n16044 ^ n11130 ^ 1'b0 ;
  assign n16046 = n16042 | n16045 ;
  assign n16048 = n3071 & ~n5520 ;
  assign n16049 = n16048 ^ n8033 ^ 1'b0 ;
  assign n16047 = n6285 & n15080 ;
  assign n16050 = n16049 ^ n16047 ^ n5631 ;
  assign n16051 = n5266 ^ n4799 ^ 1'b0 ;
  assign n16052 = n16051 ^ n605 ^ 1'b0 ;
  assign n16053 = n11852 & n16052 ;
  assign n16054 = ( n3699 & ~n4082 ) | ( n3699 & n5209 ) | ( ~n4082 & n5209 ) ;
  assign n16055 = n8314 | n16054 ;
  assign n16056 = n16055 ^ n3790 ^ 1'b0 ;
  assign n16057 = n16056 ^ n4461 ^ 1'b0 ;
  assign n16058 = ~n8655 & n16057 ;
  assign n16059 = ( n77 & n2181 ) | ( n77 & ~n13441 ) | ( n2181 & ~n13441 ) ;
  assign n16060 = n14953 ^ n2953 ^ 1'b0 ;
  assign n16061 = n4563 & ~n8715 ;
  assign n16062 = ~n1311 & n16061 ;
  assign n16063 = n16062 ^ n1815 ^ 1'b0 ;
  assign n16064 = n6125 ^ n1465 ^ 1'b0 ;
  assign n16065 = n16064 ^ n13698 ^ 1'b0 ;
  assign n16066 = n2670 & ~n3916 ;
  assign n16067 = n7019 & ~n8016 ;
  assign n16068 = ( ~n61 & n2864 ) | ( ~n61 & n6262 ) | ( n2864 & n6262 ) ;
  assign n16069 = n1822 & n16068 ;
  assign n16070 = n16069 ^ n1276 ^ 1'b0 ;
  assign n16071 = n1037 & ~n16070 ;
  assign n16072 = n2573 ^ n2356 ^ 1'b0 ;
  assign n16073 = n7400 | n16072 ;
  assign n16074 = n3141 & n5673 ;
  assign n16075 = ( ~n11249 & n16073 ) | ( ~n11249 & n16074 ) | ( n16073 & n16074 ) ;
  assign n16076 = n9241 ^ n1387 ^ 1'b0 ;
  assign n16077 = n953 & n16076 ;
  assign n16078 = n176 & n840 ;
  assign n16079 = n16078 ^ n1314 ^ 1'b0 ;
  assign n16080 = n16079 ^ n10894 ^ 1'b0 ;
  assign n16081 = n1766 | n16080 ;
  assign n16082 = n2734 ^ n91 ^ 1'b0 ;
  assign n16083 = n9718 ^ n3011 ^ 1'b0 ;
  assign n16084 = ( n8494 & n16082 ) | ( n8494 & n16083 ) | ( n16082 & n16083 ) ;
  assign n16085 = ~n11646 & n16084 ;
  assign n16086 = n16085 ^ n732 ^ 1'b0 ;
  assign n16087 = n12384 & ~n16086 ;
  assign n16089 = n1046 & ~n9594 ;
  assign n16088 = ~n2873 & n13821 ;
  assign n16090 = n16089 ^ n16088 ^ 1'b0 ;
  assign n16091 = n16090 ^ n9858 ^ 1'b0 ;
  assign n16092 = n2584 & n3079 ;
  assign n16093 = n16092 ^ n5263 ^ 1'b0 ;
  assign n16094 = n11140 ^ n3481 ^ 1'b0 ;
  assign n16095 = ~n2095 & n16094 ;
  assign n16096 = n3811 & n16095 ;
  assign n16097 = n14167 & n14231 ;
  assign n16098 = n5791 & n8171 ;
  assign n16099 = n580 & ~n6576 ;
  assign n16100 = n16099 ^ n4147 ^ 1'b0 ;
  assign n16101 = n10123 & n16100 ;
  assign n16102 = n16101 ^ n14019 ^ 1'b0 ;
  assign n16103 = n848 & ~n7013 ;
  assign n16104 = n16103 ^ n1902 ^ 1'b0 ;
  assign n16105 = ~n593 & n5596 ;
  assign n16106 = n13747 & n16105 ;
  assign n16107 = n933 ^ n294 ^ 1'b0 ;
  assign n16108 = n3100 & n16107 ;
  assign n16109 = ~n1206 & n1621 ;
  assign n16110 = n16109 ^ n6787 ^ 1'b0 ;
  assign n16112 = n10415 ^ n3635 ^ 1'b0 ;
  assign n16111 = ~n3455 & n8074 ;
  assign n16113 = n16112 ^ n16111 ^ 1'b0 ;
  assign n16114 = n5625 & n16113 ;
  assign n16115 = ~n16110 & n16114 ;
  assign n16116 = ( n11782 & n16108 ) | ( n11782 & ~n16115 ) | ( n16108 & ~n16115 ) ;
  assign n16117 = ~n10682 & n16116 ;
  assign n16118 = n6074 ^ n3919 ^ 1'b0 ;
  assign n16119 = n12684 & n16118 ;
  assign n16120 = n16119 ^ n8953 ^ 1'b0 ;
  assign n16121 = n16120 ^ n113 ^ 1'b0 ;
  assign n16122 = n9615 | n16121 ;
  assign n16123 = n13739 ^ n10478 ^ n5393 ;
  assign n16124 = ~n772 & n11904 ;
  assign n16125 = n8265 & n16124 ;
  assign n16126 = ~n12214 & n16125 ;
  assign n16127 = n3732 ^ n2463 ^ 1'b0 ;
  assign n16128 = n4531 | n10830 ;
  assign n16129 = n464 | n16128 ;
  assign n16130 = n8306 | n16129 ;
  assign n16132 = n3190 ^ n2992 ^ 1'b0 ;
  assign n16131 = n11451 ^ n3383 ^ n1000 ;
  assign n16133 = n16132 ^ n16131 ^ n4054 ;
  assign n16138 = n8911 ^ n3467 ^ 1'b0 ;
  assign n16139 = n645 & n16138 ;
  assign n16134 = ~n5085 & n8539 ;
  assign n16135 = n8952 ^ n98 ^ 1'b0 ;
  assign n16136 = n16134 & n16135 ;
  assign n16137 = n9799 & n16136 ;
  assign n16140 = n16139 ^ n16137 ^ 1'b0 ;
  assign n16141 = ~n374 & n10279 ;
  assign n16142 = n16141 ^ n9208 ^ 1'b0 ;
  assign n16143 = n41 | n16142 ;
  assign n16144 = n13943 ^ n4765 ^ 1'b0 ;
  assign n16145 = ~n16143 & n16144 ;
  assign n16146 = n16145 ^ n10647 ^ n1527 ;
  assign n16149 = n7872 ^ n5028 ^ 1'b0 ;
  assign n16148 = ~n5815 & n7707 ;
  assign n16150 = n16149 ^ n16148 ^ 1'b0 ;
  assign n16147 = n7398 & n11764 ;
  assign n16151 = n16150 ^ n16147 ^ 1'b0 ;
  assign n16152 = n3539 ^ n1350 ^ 1'b0 ;
  assign n16153 = ~n16151 & n16152 ;
  assign n16154 = n16153 ^ n9351 ^ n7190 ;
  assign n16155 = n3137 | n7443 ;
  assign n16156 = n4489 ^ n1540 ^ 1'b0 ;
  assign n16157 = n16155 & n16156 ;
  assign n16158 = n2615 & ~n3557 ;
  assign n16159 = ~n5256 & n16158 ;
  assign n16160 = ( n547 & ~n3798 ) | ( n547 & n13627 ) | ( ~n3798 & n13627 ) ;
  assign n16161 = n1064 | n16160 ;
  assign n16162 = n2869 & ~n16161 ;
  assign n16163 = ~n7393 & n10356 ;
  assign n16164 = n16162 & n16163 ;
  assign n16165 = n16159 | n16164 ;
  assign n16166 = n16165 ^ n6662 ^ 1'b0 ;
  assign n16167 = n3769 ^ n3531 ^ 1'b0 ;
  assign n16168 = n6386 | n16167 ;
  assign n16169 = n16168 ^ n6698 ^ n350 ;
  assign n16170 = ( n4674 & ~n9002 ) | ( n4674 & n16169 ) | ( ~n9002 & n16169 ) ;
  assign n16171 = ~n3229 & n11587 ;
  assign n16172 = n7300 ^ n4914 ^ 1'b0 ;
  assign n16173 = ~n10199 & n16172 ;
  assign n16174 = n16173 ^ n9680 ^ 1'b0 ;
  assign n16175 = ~n10722 & n16174 ;
  assign n16176 = ( ~n2484 & n4043 ) | ( ~n2484 & n5103 ) | ( n4043 & n5103 ) ;
  assign n16177 = ~n8154 & n16176 ;
  assign n16178 = n6609 & ~n16177 ;
  assign n16179 = n8323 & n16178 ;
  assign n16180 = n16175 & ~n16179 ;
  assign n16181 = n16180 ^ n1661 ^ 1'b0 ;
  assign n16182 = n4183 ^ n3201 ^ n2705 ;
  assign n16184 = n5142 ^ n3526 ^ 1'b0 ;
  assign n16185 = n1303 & n16184 ;
  assign n16183 = n3407 & ~n11066 ;
  assign n16186 = n16185 ^ n16183 ^ 1'b0 ;
  assign n16192 = n9263 ^ n8467 ^ 1'b0 ;
  assign n16187 = ~n3218 & n11555 ;
  assign n16188 = n695 & ~n6236 ;
  assign n16189 = ~n1350 & n16188 ;
  assign n16190 = n5948 | n16189 ;
  assign n16191 = n16187 & ~n16190 ;
  assign n16193 = n16192 ^ n16191 ^ 1'b0 ;
  assign n16194 = n15271 & ~n16193 ;
  assign n16195 = n1686 & n12588 ;
  assign n16196 = n2895 & ~n9866 ;
  assign n16197 = n11959 & ~n14721 ;
  assign n16198 = n1269 | n16197 ;
  assign n16199 = n4335 ^ n494 ^ n434 ;
  assign n16200 = n2828 & n14509 ;
  assign n16201 = n16200 ^ n15364 ^ 1'b0 ;
  assign n16202 = n9789 ^ n197 ^ 1'b0 ;
  assign n16203 = n16112 | n16202 ;
  assign n16204 = ~n1003 & n7397 ;
  assign n16205 = n5169 & ~n16204 ;
  assign n16206 = n379 | n4334 ;
  assign n16207 = n16206 ^ n2686 ^ 1'b0 ;
  assign n16208 = n523 | n16207 ;
  assign n16209 = n4966 & n8486 ;
  assign n16210 = n16209 ^ n2174 ^ 1'b0 ;
  assign n16211 = n2720 ^ n2544 ^ 1'b0 ;
  assign n16212 = n2980 & ~n16211 ;
  assign n16213 = n7158 | n16212 ;
  assign n16214 = n11117 & ~n16213 ;
  assign n16215 = n5921 ^ n5711 ^ n4543 ;
  assign n16216 = n16215 ^ n10817 ^ 1'b0 ;
  assign n16217 = ~n16214 & n16216 ;
  assign n16218 = ( n1155 & n2045 ) | ( n1155 & n16217 ) | ( n2045 & n16217 ) ;
  assign n16219 = n11894 ^ n5107 ^ 1'b0 ;
  assign n16220 = n320 & n1200 ;
  assign n16221 = n101 & n2773 ;
  assign n16222 = n16221 ^ n15737 ^ 1'b0 ;
  assign n16223 = n2791 & n16222 ;
  assign n16224 = ( n9717 & ~n11734 ) | ( n9717 & n16223 ) | ( ~n11734 & n16223 ) ;
  assign n16225 = ( ~n2168 & n16220 ) | ( ~n2168 & n16224 ) | ( n16220 & n16224 ) ;
  assign n16226 = n2594 ^ n1305 ^ 1'b0 ;
  assign n16227 = n9373 ^ n5062 ^ 1'b0 ;
  assign n16228 = n5965 | n16227 ;
  assign n16229 = n5648 | n16228 ;
  assign n16230 = n231 & ~n16229 ;
  assign n16231 = ~n1522 & n13766 ;
  assign n16232 = n200 | n1606 ;
  assign n16233 = ( n4715 & n7441 ) | ( n4715 & n15344 ) | ( n7441 & n15344 ) ;
  assign n16234 = n8231 & n16233 ;
  assign n16235 = n16234 ^ n6674 ^ 1'b0 ;
  assign n16236 = n7092 ^ n3779 ^ 1'b0 ;
  assign n16237 = n10768 | n16236 ;
  assign n16238 = n16237 ^ n3853 ^ 1'b0 ;
  assign n16239 = n9120 ^ n6866 ^ 1'b0 ;
  assign n16240 = n6520 & n16239 ;
  assign n16241 = n13970 ^ n13850 ^ 1'b0 ;
  assign n16242 = ~n8085 & n16241 ;
  assign n16243 = ~n14125 & n16242 ;
  assign n16244 = n16243 ^ n717 ^ 1'b0 ;
  assign n16245 = n379 & ~n4750 ;
  assign n16246 = n2864 ^ n122 ^ 1'b0 ;
  assign n16247 = ( n1125 & ~n3442 ) | ( n1125 & n16246 ) | ( ~n3442 & n16246 ) ;
  assign n16248 = n394 & ~n16247 ;
  assign n16249 = n12161 & ~n16248 ;
  assign n16250 = n16245 & n16249 ;
  assign n16251 = ~n9134 & n14148 ;
  assign n16252 = n16251 ^ n594 ^ 1'b0 ;
  assign n16253 = ~n10229 & n10263 ;
  assign n16254 = n16252 & n16253 ;
  assign n16255 = n4495 & ~n16254 ;
  assign n16256 = n14605 ^ n3330 ^ 1'b0 ;
  assign n16257 = n2986 ^ n2058 ^ 1'b0 ;
  assign n16258 = n5107 & n16257 ;
  assign n16259 = ( ~n11615 & n15148 ) | ( ~n11615 & n16258 ) | ( n15148 & n16258 ) ;
  assign n16260 = n3066 | n9453 ;
  assign n16261 = n922 & ~n15693 ;
  assign n16262 = ( n332 & ~n1448 ) | ( n332 & n16261 ) | ( ~n1448 & n16261 ) ;
  assign n16263 = n844 & n12097 ;
  assign n16264 = n16263 ^ n4002 ^ n505 ;
  assign n16265 = n7061 & n9261 ;
  assign n16266 = n9428 ^ n3274 ^ 1'b0 ;
  assign n16267 = n6911 & ~n16266 ;
  assign n16268 = n7848 ^ n1535 ^ n57 ;
  assign n16269 = ( n5562 & ~n16267 ) | ( n5562 & n16268 ) | ( ~n16267 & n16268 ) ;
  assign n16270 = n3361 ^ n2483 ^ 1'b0 ;
  assign n16271 = n16269 & n16270 ;
  assign n16272 = n12938 & n16271 ;
  assign n16273 = n16265 & n16272 ;
  assign n16274 = ~n7455 & n13380 ;
  assign n16275 = n257 | n10815 ;
  assign n16276 = n12348 & ~n15102 ;
  assign n16277 = n16275 & n16276 ;
  assign n16278 = n10957 & ~n13891 ;
  assign n16279 = n3170 | n9864 ;
  assign n16280 = ~n5444 & n12451 ;
  assign n16281 = n8232 ^ n4848 ^ 1'b0 ;
  assign n16282 = ~n14964 & n16281 ;
  assign n16283 = ~n2113 & n4014 ;
  assign n16284 = n16283 ^ n11874 ^ 1'b0 ;
  assign n16285 = n16284 ^ n5234 ^ 1'b0 ;
  assign n16286 = n16282 & ~n16285 ;
  assign n16287 = n2984 | n7240 ;
  assign n16288 = n6676 & ~n16287 ;
  assign n16289 = n1233 | n16288 ;
  assign n16290 = n11792 & ~n16289 ;
  assign n16291 = n7998 ^ n5853 ^ n3973 ;
  assign n16292 = n646 & ~n5996 ;
  assign n16293 = ~n4757 & n16292 ;
  assign n16294 = n5399 | n6428 ;
  assign n16295 = n16294 ^ n9981 ^ n7445 ;
  assign n16296 = n16295 ^ n9755 ^ n8344 ;
  assign n16298 = n8624 ^ n8103 ^ n6122 ;
  assign n16297 = n4204 & n11955 ;
  assign n16299 = n16298 ^ n16297 ^ 1'b0 ;
  assign n16300 = n3408 & n4608 ;
  assign n16301 = n1283 & n16300 ;
  assign n16302 = n603 & ~n16301 ;
  assign n16303 = ( ~n3624 & n7454 ) | ( ~n3624 & n13330 ) | ( n7454 & n13330 ) ;
  assign n16304 = n2411 & ~n16303 ;
  assign n16305 = n1775 & n6546 ;
  assign n16306 = n1110 & n16305 ;
  assign n16307 = ~n4512 & n16306 ;
  assign n16308 = n16307 ^ n13346 ^ 1'b0 ;
  assign n16309 = n8887 & n16308 ;
  assign n16310 = n7308 & n9896 ;
  assign n16311 = n16309 & ~n16310 ;
  assign n16312 = n2050 & ~n2139 ;
  assign n16313 = ~n2435 & n16312 ;
  assign n16314 = n8047 & ~n16313 ;
  assign n16315 = ~n5727 & n7770 ;
  assign n16316 = n16315 ^ n4009 ^ 1'b0 ;
  assign n16317 = n2150 & ~n16316 ;
  assign n16318 = n15509 ^ n12936 ^ n5169 ;
  assign n16325 = n6576 ^ n2072 ^ 1'b0 ;
  assign n16326 = ~n1856 & n16325 ;
  assign n16319 = n1842 & ~n3928 ;
  assign n16320 = n3926 & n16319 ;
  assign n16321 = ~n5724 & n16320 ;
  assign n16322 = n13205 | n16321 ;
  assign n16323 = n4673 & ~n16322 ;
  assign n16324 = ( n245 & n10307 ) | ( n245 & n16323 ) | ( n10307 & n16323 ) ;
  assign n16327 = n16326 ^ n16324 ^ 1'b0 ;
  assign n16328 = n13738 ^ n4736 ^ 1'b0 ;
  assign n16329 = ~n2433 & n4584 ;
  assign n16330 = ( n187 & n15389 ) | ( n187 & ~n16329 ) | ( n15389 & ~n16329 ) ;
  assign n16331 = n283 & ~n14437 ;
  assign n16332 = n436 & n16331 ;
  assign n16333 = n601 & n1353 ;
  assign n16334 = n16333 ^ n1031 ^ 1'b0 ;
  assign n16335 = n8555 ^ n8438 ^ 1'b0 ;
  assign n16336 = ~n16334 & n16335 ;
  assign n16337 = n3467 ^ n299 ^ 1'b0 ;
  assign n16338 = n4185 & ~n5580 ;
  assign n16339 = n16338 ^ n9451 ^ 1'b0 ;
  assign n16340 = n16339 ^ n9003 ^ 1'b0 ;
  assign n16341 = ( n9862 & ~n16337 ) | ( n9862 & n16340 ) | ( ~n16337 & n16340 ) ;
  assign n16342 = n9052 ^ n107 ^ 1'b0 ;
  assign n16343 = n12143 & ~n14671 ;
  assign n16344 = n678 & ~n1137 ;
  assign n16345 = n16344 ^ n6221 ^ 1'b0 ;
  assign n16346 = n9339 ^ n7242 ^ n1818 ;
  assign n16347 = n7971 | n9667 ;
  assign n16348 = n16346 & n16347 ;
  assign n16349 = n16348 ^ n12517 ^ 1'b0 ;
  assign n16350 = n16345 & ~n16349 ;
  assign n16351 = n11253 ^ n8282 ^ 1'b0 ;
  assign n16352 = n16351 ^ n6107 ^ 1'b0 ;
  assign n16353 = n12452 & n16352 ;
  assign n16355 = n2884 & ~n7535 ;
  assign n16354 = n6466 & ~n9065 ;
  assign n16356 = n16355 ^ n16354 ^ 1'b0 ;
  assign n16357 = n16356 ^ n15420 ^ n13428 ;
  assign n16358 = n14187 ^ n10775 ^ 1'b0 ;
  assign n16359 = n8678 | n16358 ;
  assign n16360 = ( n3890 & ~n12844 ) | ( n3890 & n16359 ) | ( ~n12844 & n16359 ) ;
  assign n16361 = ~n3404 & n9424 ;
  assign n16362 = ~n6337 & n16361 ;
  assign n16363 = n5302 | n9141 ;
  assign n16364 = ~n11307 & n16363 ;
  assign n16365 = ~n8292 & n16364 ;
  assign n16366 = ( n2350 & n11976 ) | ( n2350 & n16309 ) | ( n11976 & n16309 ) ;
  assign n16367 = n13997 ^ n2354 ^ 1'b0 ;
  assign n16368 = n5872 ^ n2097 ^ 1'b0 ;
  assign n16371 = n453 & n2493 ;
  assign n16369 = n1690 & ~n5673 ;
  assign n16370 = n16369 ^ n9517 ^ 1'b0 ;
  assign n16372 = n16371 ^ n16370 ^ n2648 ;
  assign n16373 = n16368 & ~n16372 ;
  assign n16374 = n12004 ^ n9079 ^ n8466 ;
  assign n16375 = ~n2591 & n6561 ;
  assign n16376 = n16375 ^ n10982 ^ 1'b0 ;
  assign n16377 = ~n719 & n11341 ;
  assign n16378 = n9344 & n16377 ;
  assign n16379 = n8074 ^ n2368 ^ 1'b0 ;
  assign n16380 = n16379 ^ n6630 ^ 1'b0 ;
  assign n16381 = n16378 | n16380 ;
  assign n16382 = n4638 & n14066 ;
  assign n16383 = n16382 ^ n9416 ^ 1'b0 ;
  assign n16384 = n9045 ^ n5092 ^ 1'b0 ;
  assign n16385 = ~n1134 & n16384 ;
  assign n16386 = ~n2980 & n4684 ;
  assign n16387 = n16386 ^ n2728 ^ 1'b0 ;
  assign n16388 = ~n10023 & n16387 ;
  assign n16389 = n16388 ^ n16045 ^ 1'b0 ;
  assign n16390 = n4142 | n16389 ;
  assign n16391 = n1744 & n16390 ;
  assign n16392 = n3991 ^ n3071 ^ 1'b0 ;
  assign n16393 = n12089 & ~n16392 ;
  assign n16394 = n13215 | n16101 ;
  assign n16395 = n13073 ^ n2682 ^ 1'b0 ;
  assign n16396 = ~n4896 & n16395 ;
  assign n16397 = n7633 ^ n3073 ^ 1'b0 ;
  assign n16398 = n3446 | n16397 ;
  assign n16399 = n4618 & n6475 ;
  assign n16400 = n16014 ^ n8383 ^ n5218 ;
  assign n16401 = x1 & n14755 ;
  assign n16402 = n16401 ^ n2597 ^ 1'b0 ;
  assign n16403 = n16402 ^ n10029 ^ 1'b0 ;
  assign n16404 = n1334 & ~n16403 ;
  assign n16405 = n2880 & n9852 ;
  assign n16406 = n9224 | n16405 ;
  assign n16407 = ( ~n1775 & n13605 ) | ( ~n1775 & n13876 ) | ( n13605 & n13876 ) ;
  assign n16408 = n3045 | n6412 ;
  assign n16409 = n16408 ^ n374 ^ 1'b0 ;
  assign n16410 = n14578 | n16409 ;
  assign n16411 = n16407 & ~n16410 ;
  assign n16412 = ~n4181 & n5491 ;
  assign n16413 = ( n1937 & ~n16411 ) | ( n1937 & n16412 ) | ( ~n16411 & n16412 ) ;
  assign n16415 = n13034 ^ n9397 ^ n8129 ;
  assign n16414 = n8033 & ~n11447 ;
  assign n16416 = n16415 ^ n16414 ^ 1'b0 ;
  assign n16417 = n9997 | n16416 ;
  assign n16418 = n1214 | n7335 ;
  assign n16419 = n16418 ^ n10425 ^ 1'b0 ;
  assign n16420 = n16419 ^ n2137 ^ n1980 ;
  assign n16421 = n12734 ^ n10569 ^ 1'b0 ;
  assign n16423 = n11195 ^ n9195 ^ 1'b0 ;
  assign n16424 = n8245 & ~n16423 ;
  assign n16422 = ~n1026 & n15407 ;
  assign n16425 = n16424 ^ n16422 ^ 1'b0 ;
  assign n16426 = n10975 ^ n3989 ^ n2123 ;
  assign n16427 = n11220 & n16426 ;
  assign n16428 = n16427 ^ n3656 ^ 1'b0 ;
  assign n16429 = n14845 ^ n63 ^ 1'b0 ;
  assign n16430 = n7615 & n16429 ;
  assign n16435 = n1053 & n1241 ;
  assign n16436 = ~n1241 & n16435 ;
  assign n16433 = n141 & ~n8692 ;
  assign n16434 = ~n141 & n16433 ;
  assign n16437 = n16436 ^ n16434 ^ 1'b0 ;
  assign n16431 = n230 & ~n2469 ;
  assign n16432 = n2469 & n16431 ;
  assign n16438 = n16437 ^ n16432 ^ 1'b0 ;
  assign n16439 = n13676 & ~n16438 ;
  assign n16442 = n1932 & ~n3624 ;
  assign n16443 = ~n13101 & n16442 ;
  assign n16440 = n9227 ^ n2827 ^ n63 ;
  assign n16441 = n16440 ^ n1487 ^ n23 ;
  assign n16444 = n16443 ^ n16441 ^ 1'b0 ;
  assign n16445 = n3684 ^ n1645 ^ 1'b0 ;
  assign n16446 = n14962 ^ n7817 ^ 1'b0 ;
  assign n16447 = n16445 & ~n16446 ;
  assign n16448 = n3838 & ~n8560 ;
  assign n16449 = ~n3016 & n16448 ;
  assign n16450 = n16449 ^ n6622 ^ n6574 ;
  assign n16451 = n16450 ^ n14487 ^ n11415 ;
  assign n16452 = ~n4442 & n6614 ;
  assign n16453 = ( ~n134 & n3326 ) | ( ~n134 & n3868 ) | ( n3326 & n3868 ) ;
  assign n16454 = n5732 | n16453 ;
  assign n16455 = ~n9151 & n11707 ;
  assign n16456 = ~n2563 & n16455 ;
  assign n16457 = n16454 | n16456 ;
  assign n16458 = n889 & n9686 ;
  assign n16459 = n16458 ^ n1754 ^ 1'b0 ;
  assign n16460 = n3916 & ~n8565 ;
  assign n16461 = ( ~n1289 & n7914 ) | ( ~n1289 & n16460 ) | ( n7914 & n16460 ) ;
  assign n16462 = ~n6842 & n10239 ;
  assign n16463 = n16462 ^ n13257 ^ 1'b0 ;
  assign n16464 = ~n10846 & n16463 ;
  assign n16465 = ( ~n4084 & n13137 ) | ( ~n4084 & n16464 ) | ( n13137 & n16464 ) ;
  assign n16466 = n640 | n3855 ;
  assign n16467 = n16466 ^ n12369 ^ 1'b0 ;
  assign n16468 = n16467 ^ n844 ^ 1'b0 ;
  assign n16469 = n5568 & n13177 ;
  assign n16470 = n16469 ^ n7003 ^ 1'b0 ;
  assign n16475 = n2475 ^ n1613 ^ 1'b0 ;
  assign n16474 = n14975 ^ n6181 ^ 1'b0 ;
  assign n16473 = n5836 ^ n3310 ^ 1'b0 ;
  assign n16476 = n16475 ^ n16474 ^ n16473 ;
  assign n16471 = n569 & n5806 ;
  assign n16472 = n6125 & ~n16471 ;
  assign n16477 = n16476 ^ n16472 ^ 1'b0 ;
  assign n16479 = n9295 ^ n3780 ^ 1'b0 ;
  assign n16480 = n12032 & ~n16479 ;
  assign n16481 = ( ~n436 & n14258 ) | ( ~n436 & n16480 ) | ( n14258 & n16480 ) ;
  assign n16478 = n1384 & ~n1791 ;
  assign n16482 = n16481 ^ n16478 ^ n6317 ;
  assign n16483 = n16482 ^ n2913 ^ 1'b0 ;
  assign n16484 = n13700 ^ n9800 ^ 1'b0 ;
  assign n16485 = n3560 | n4846 ;
  assign n16486 = ~n13462 & n16485 ;
  assign n16487 = n49 & n16486 ;
  assign n16488 = n1415 & n4615 ;
  assign n16489 = n16488 ^ n12662 ^ 1'b0 ;
  assign n16490 = n10660 ^ n4457 ^ 1'b0 ;
  assign n16491 = n1170 & ~n16490 ;
  assign n16492 = n3134 | n16491 ;
  assign n16493 = n918 & n10083 ;
  assign n16494 = n1196 | n16493 ;
  assign n16495 = n5329 & ~n16494 ;
  assign n16496 = ( n16489 & n16492 ) | ( n16489 & ~n16495 ) | ( n16492 & ~n16495 ) ;
  assign n16497 = n12050 ^ n2408 ^ 1'b0 ;
  assign n16498 = n4440 ^ n926 ^ 1'b0 ;
  assign n16499 = n4591 | n16498 ;
  assign n16500 = ( n1350 & n8978 ) | ( n1350 & ~n16499 ) | ( n8978 & ~n16499 ) ;
  assign n16501 = n10895 ^ n4689 ^ 1'b0 ;
  assign n16502 = n16500 | n16501 ;
  assign n16503 = n14057 ^ n41 ^ 1'b0 ;
  assign n16504 = n242 | n16503 ;
  assign n16505 = ( ~n4982 & n7760 ) | ( ~n4982 & n16504 ) | ( n7760 & n16504 ) ;
  assign n16508 = n11628 ^ n38 ^ 1'b0 ;
  assign n16509 = ~n2841 & n16508 ;
  assign n16506 = ( ~n1805 & n3894 ) | ( ~n1805 & n12527 ) | ( n3894 & n12527 ) ;
  assign n16507 = n14039 & ~n16506 ;
  assign n16510 = n16509 ^ n16507 ^ 1'b0 ;
  assign n16511 = n13096 ^ n8327 ^ n250 ;
  assign n16512 = n14851 ^ n6970 ^ 1'b0 ;
  assign n16513 = n9707 | n16512 ;
  assign n16514 = n2939 & ~n12914 ;
  assign n16515 = n14651 & n16514 ;
  assign n16516 = n16454 & n16515 ;
  assign n16517 = n12551 ^ n6076 ^ 1'b0 ;
  assign n16518 = ~n5468 & n5724 ;
  assign n16519 = n16518 ^ n11182 ^ 1'b0 ;
  assign n16520 = n16519 ^ n12375 ^ 1'b0 ;
  assign n16521 = n5883 | n16520 ;
  assign n16522 = n605 & ~n7038 ;
  assign n16523 = n16521 | n16522 ;
  assign n16525 = ( n3196 & n7103 ) | ( n3196 & ~n7211 ) | ( n7103 & ~n7211 ) ;
  assign n16524 = ~n2568 & n4134 ;
  assign n16526 = n16525 ^ n16524 ^ 1'b0 ;
  assign n16527 = n4835 ^ n3020 ^ 1'b0 ;
  assign n16528 = n16527 ^ n2932 ^ 1'b0 ;
  assign n16529 = n3439 | n16528 ;
  assign n16530 = n16529 ^ n16421 ^ 1'b0 ;
  assign n16531 = n5225 & ~n16530 ;
  assign n16532 = n4159 | n9538 ;
  assign n16533 = ~n135 & n4126 ;
  assign n16534 = ~n16532 & n16533 ;
  assign n16535 = n2922 & ~n16534 ;
  assign n16536 = n2528 & n16535 ;
  assign n16537 = n887 & n3481 ;
  assign n16538 = n16536 & n16537 ;
  assign n16539 = n10528 & n14603 ;
  assign n16540 = n5266 & ~n10850 ;
  assign n16541 = n11091 ^ n933 ^ 1'b0 ;
  assign n16542 = n16540 & ~n16541 ;
  assign n16543 = n9643 ^ n1148 ^ 1'b0 ;
  assign n16544 = n153 & n16543 ;
  assign n16545 = n6356 ^ n6188 ^ 1'b0 ;
  assign n16546 = n16545 ^ n16488 ^ 1'b0 ;
  assign n16547 = n392 | n16546 ;
  assign n16548 = n12000 | n16547 ;
  assign n16549 = n11209 ^ n2330 ^ 1'b0 ;
  assign n16550 = n3098 ^ n1983 ^ 1'b0 ;
  assign n16551 = ( n4272 & n4889 ) | ( n4272 & ~n16550 ) | ( n4889 & ~n16550 ) ;
  assign n16552 = n16551 ^ n3936 ^ 1'b0 ;
  assign n16553 = n11860 ^ n5796 ^ 1'b0 ;
  assign n16554 = n7590 & ~n16553 ;
  assign n16556 = ( ~n1249 & n3248 ) | ( ~n1249 & n5321 ) | ( n3248 & n5321 ) ;
  assign n16555 = ~n2832 & n7766 ;
  assign n16557 = n16556 ^ n16555 ^ 1'b0 ;
  assign n16558 = n16557 ^ n6491 ^ 1'b0 ;
  assign n16559 = n16554 & n16558 ;
  assign n16560 = n2051 & n16559 ;
  assign n16561 = n2745 ^ n2014 ^ 1'b0 ;
  assign n16562 = n16561 ^ n10973 ^ 1'b0 ;
  assign n16563 = n6490 & ~n16562 ;
  assign n16564 = n8338 & n13676 ;
  assign n16565 = ~n4215 & n16564 ;
  assign n16566 = n608 | n16565 ;
  assign n16567 = n11485 | n16566 ;
  assign n16568 = n16567 ^ n11374 ^ 1'b0 ;
  assign n16569 = n6128 ^ n4497 ^ 1'b0 ;
  assign n16570 = n2124 & n16569 ;
  assign n16571 = n2808 & n16570 ;
  assign n16572 = n1091 & ~n1373 ;
  assign n16573 = n1400 & n15190 ;
  assign n16574 = n4009 ^ n3557 ^ 1'b0 ;
  assign n16575 = ( ~n2025 & n7807 ) | ( ~n2025 & n13050 ) | ( n7807 & n13050 ) ;
  assign n16576 = n12583 ^ n1717 ^ 1'b0 ;
  assign n16577 = n8341 & ~n16576 ;
  assign n16578 = n8148 & n16577 ;
  assign n16579 = n2369 & ~n13727 ;
  assign n16580 = n16579 ^ n12028 ^ 1'b0 ;
  assign n16581 = n13771 ^ n11076 ^ n2525 ;
  assign n16582 = n10596 & ~n16581 ;
  assign n16583 = n7864 & n8157 ;
  assign n16584 = n16582 & n16583 ;
  assign n16585 = ~n2773 & n16584 ;
  assign n16586 = n1793 & ~n5314 ;
  assign n16587 = n1250 & n16586 ;
  assign n16588 = ~n2918 & n5570 ;
  assign n16589 = n16588 ^ n15557 ^ 1'b0 ;
  assign n16597 = n12272 ^ n7320 ^ n1346 ;
  assign n16598 = n16597 ^ n7963 ^ n6960 ;
  assign n16591 = n3365 ^ n3277 ^ 1'b0 ;
  assign n16590 = n1783 & n10038 ;
  assign n16592 = n16591 ^ n16590 ^ 1'b0 ;
  assign n16593 = n11927 | n16592 ;
  assign n16594 = n16593 ^ n7395 ^ 1'b0 ;
  assign n16595 = ~n3341 & n16594 ;
  assign n16596 = n2497 & n16595 ;
  assign n16599 = n16598 ^ n16596 ^ n5910 ;
  assign n16600 = ~n1777 & n6102 ;
  assign n16601 = n16600 ^ n13923 ^ 1'b0 ;
  assign n16602 = ~n6178 & n7603 ;
  assign n16603 = n16601 | n16602 ;
  assign n16608 = n2461 & ~n10140 ;
  assign n16609 = ~n13498 & n16608 ;
  assign n16604 = n1282 ^ n601 ^ 1'b0 ;
  assign n16605 = n786 | n16604 ;
  assign n16606 = n16605 ^ n11638 ^ n11485 ;
  assign n16607 = n8899 & ~n16606 ;
  assign n16610 = n16609 ^ n16607 ^ 1'b0 ;
  assign n16611 = n8695 ^ n2861 ^ 1'b0 ;
  assign n16612 = n10548 ^ n4088 ^ 1'b0 ;
  assign n16613 = n15590 ^ n15017 ^ 1'b0 ;
  assign n16614 = n8176 & n16613 ;
  assign n16615 = n2818 | n7908 ;
  assign n16616 = n9180 & n16615 ;
  assign n16617 = ~n12530 & n16616 ;
  assign n16618 = ~n3518 & n16617 ;
  assign n16619 = n4085 & n6426 ;
  assign n16620 = n16619 ^ n7108 ^ 1'b0 ;
  assign n16621 = n16620 ^ n4260 ^ 1'b0 ;
  assign n16622 = ~n7958 & n16621 ;
  assign n16623 = n15958 & ~n16622 ;
  assign n16624 = ( n2507 & n2702 ) | ( n2507 & n10703 ) | ( n2702 & n10703 ) ;
  assign n16625 = n14701 ^ n9232 ^ n4751 ;
  assign n16626 = n2186 & n8260 ;
  assign n16627 = n265 & n16626 ;
  assign n16628 = ~n4987 & n14445 ;
  assign n16629 = n16185 & ~n16628 ;
  assign n16630 = n13103 ^ n3317 ^ 1'b0 ;
  assign n16631 = n5316 | n16630 ;
  assign n16632 = n9866 & ~n16631 ;
  assign n16633 = ( n5771 & ~n7600 ) | ( n5771 & n9286 ) | ( ~n7600 & n9286 ) ;
  assign n16634 = ~n4246 & n16633 ;
  assign n16635 = ~n5160 & n16634 ;
  assign n16636 = n12749 ^ n10632 ^ n2880 ;
  assign n16637 = n5414 ^ n2992 ^ n830 ;
  assign n16638 = n14848 ^ n6018 ^ 1'b0 ;
  assign n16639 = n4340 | n16638 ;
  assign n16640 = n16637 & n16639 ;
  assign n16641 = n2370 & ~n6119 ;
  assign n16642 = n16641 ^ n10674 ^ n4864 ;
  assign n16650 = n11533 ^ n749 ^ 1'b0 ;
  assign n16646 = n166 & n3981 ;
  assign n16647 = n16646 ^ n405 ^ 1'b0 ;
  assign n16643 = n6091 ^ n1186 ^ 1'b0 ;
  assign n16644 = n1888 | n16643 ;
  assign n16645 = n4599 & ~n16644 ;
  assign n16648 = n16647 ^ n16645 ^ 1'b0 ;
  assign n16649 = n11902 & n16648 ;
  assign n16651 = n16650 ^ n16649 ^ 1'b0 ;
  assign n16652 = n1827 ^ n30 ^ 1'b0 ;
  assign n16653 = n16652 ^ n16130 ^ n10827 ;
  assign n16656 = n3732 ^ n1160 ^ 1'b0 ;
  assign n16657 = n15837 & n16656 ;
  assign n16654 = n8980 ^ n784 ^ 1'b0 ;
  assign n16655 = n2645 | n16654 ;
  assign n16658 = n16657 ^ n16655 ^ 1'b0 ;
  assign n16659 = ~n6457 & n8083 ;
  assign n16660 = ~n7750 & n16659 ;
  assign n16661 = n6899 ^ n2939 ^ n1622 ;
  assign n16662 = n5635 & ~n16661 ;
  assign n16663 = n16660 & n16662 ;
  assign n16664 = n9468 ^ n2620 ^ 1'b0 ;
  assign n16665 = n9555 ^ n1636 ^ 1'b0 ;
  assign n16666 = n16664 & ~n16665 ;
  assign n16667 = ~n10669 & n13262 ;
  assign n16668 = ~n12810 & n16667 ;
  assign n16669 = n11078 ^ n6123 ^ 1'b0 ;
  assign n16670 = n7870 ^ n5626 ^ n5001 ;
  assign n16671 = n63 & n4602 ;
  assign n16672 = ( n16449 & n16670 ) | ( n16449 & n16671 ) | ( n16670 & n16671 ) ;
  assign n16674 = n42 & n1629 ;
  assign n16675 = n7291 & ~n16674 ;
  assign n16676 = n6238 & ~n16675 ;
  assign n16677 = n1537 & n16676 ;
  assign n16673 = n628 | n8382 ;
  assign n16678 = n16677 ^ n16673 ^ 1'b0 ;
  assign n16679 = n16678 ^ n200 ^ 1'b0 ;
  assign n16680 = n16679 ^ n5717 ^ 1'b0 ;
  assign n16683 = n998 & n8344 ;
  assign n16684 = n16683 ^ n7513 ^ 1'b0 ;
  assign n16685 = n16684 ^ n6979 ^ 1'b0 ;
  assign n16681 = n9047 ^ n3019 ^ 1'b0 ;
  assign n16682 = n8497 & ~n16681 ;
  assign n16686 = n16685 ^ n16682 ^ 1'b0 ;
  assign n16687 = ( ~n16672 & n16680 ) | ( ~n16672 & n16686 ) | ( n16680 & n16686 ) ;
  assign n16688 = ~n2385 & n14303 ;
  assign n16689 = n14690 & n16688 ;
  assign n16703 = n13250 ^ n12668 ^ n5783 ;
  assign n16690 = ~n6316 & n6579 ;
  assign n16691 = n16690 ^ n9425 ^ 1'b0 ;
  assign n16696 = n13940 ^ n3789 ^ 1'b0 ;
  assign n16697 = ~n3788 & n16696 ;
  assign n16692 = n1274 & ~n2905 ;
  assign n16693 = n16692 ^ n1290 ^ 1'b0 ;
  assign n16694 = n6322 & ~n16693 ;
  assign n16695 = n16694 ^ n9393 ^ n1811 ;
  assign n16698 = n16697 ^ n16695 ^ n633 ;
  assign n16699 = n16698 ^ n1290 ^ 1'b0 ;
  assign n16700 = n16691 & ~n16699 ;
  assign n16701 = n16700 ^ n9232 ^ n6100 ;
  assign n16702 = n4197 & n16701 ;
  assign n16704 = n16703 ^ n16702 ^ 1'b0 ;
  assign n16705 = ( ~n3993 & n11196 ) | ( ~n3993 & n12475 ) | ( n11196 & n12475 ) ;
  assign n16706 = n8597 & ~n16705 ;
  assign n16707 = n11369 ^ n4809 ^ 1'b0 ;
  assign n16708 = n926 | n10079 ;
  assign n16709 = n16708 ^ n3561 ^ 1'b0 ;
  assign n16710 = n10345 | n12337 ;
  assign n16711 = n16710 ^ n6447 ^ 1'b0 ;
  assign n16712 = ~n4443 & n9360 ;
  assign n16713 = n16712 ^ n5617 ^ 1'b0 ;
  assign n16714 = n15378 & n16713 ;
  assign n16715 = n8910 | n12945 ;
  assign n16716 = n16714 & ~n16715 ;
  assign n16717 = n16716 ^ n14329 ^ 1'b0 ;
  assign n16718 = ~n1654 & n6326 ;
  assign n16719 = n102 & n16718 ;
  assign n16720 = n16719 ^ n14294 ^ n2873 ;
  assign n16721 = n10200 ^ n9358 ^ 1'b0 ;
  assign n16722 = n2190 & n16721 ;
  assign n16723 = n16722 ^ n8942 ^ n406 ;
  assign n16724 = n11691 ^ n3207 ^ 1'b0 ;
  assign n16725 = n16724 ^ n14112 ^ 1'b0 ;
  assign n16726 = n2303 | n16725 ;
  assign n16727 = n16407 ^ n6458 ^ n3216 ;
  assign n16728 = n8917 ^ n4243 ^ 1'b0 ;
  assign n16729 = n16124 & n16728 ;
  assign n16730 = n16727 & n16729 ;
  assign n16731 = n4112 | n11912 ;
  assign n16732 = n16546 ^ n4920 ^ 1'b0 ;
  assign n16733 = n14672 | n16732 ;
  assign n16734 = n16731 & ~n16733 ;
  assign n16735 = n16734 ^ n1495 ^ 1'b0 ;
  assign n16736 = n16735 ^ n16160 ^ n6714 ;
  assign n16737 = n687 & ~n1849 ;
  assign n16738 = n481 & n16737 ;
  assign n16739 = n16738 ^ n2890 ^ 1'b0 ;
  assign n16740 = ~n11825 & n16739 ;
  assign n16741 = n16740 ^ n4911 ^ 1'b0 ;
  assign n16742 = ~n332 & n586 ;
  assign n16743 = n16742 ^ n2556 ^ 1'b0 ;
  assign n16744 = n16743 ^ n6524 ^ 1'b0 ;
  assign n16745 = n16113 & ~n16744 ;
  assign n16746 = n16741 & n16745 ;
  assign n16747 = n8881 | n16746 ;
  assign n16748 = n16747 ^ n8375 ^ 1'b0 ;
  assign n16749 = n15706 ^ n7807 ^ 1'b0 ;
  assign n16750 = n8355 & ~n10023 ;
  assign n16751 = n3966 & ~n16750 ;
  assign n16752 = n2723 & n9664 ;
  assign n16753 = n3232 & n16752 ;
  assign n16754 = n1668 & n6941 ;
  assign n16755 = ~n6053 & n16754 ;
  assign n16756 = n16755 ^ n8306 ^ n597 ;
  assign n16757 = n6671 & n14178 ;
  assign n16758 = n16757 ^ n14533 ^ 1'b0 ;
  assign n16759 = n16756 | n16758 ;
  assign n16760 = n1589 | n8248 ;
  assign n16761 = n8024 | n16760 ;
  assign n16762 = n16761 ^ n5511 ^ 1'b0 ;
  assign n16763 = n3303 | n15027 ;
  assign n16764 = n6277 ^ n2937 ^ 1'b0 ;
  assign n16765 = ~n3176 & n16764 ;
  assign n16766 = n16765 ^ n3624 ^ 1'b0 ;
  assign n16767 = ( n7185 & n9134 ) | ( n7185 & n16766 ) | ( n9134 & n16766 ) ;
  assign n16768 = n16767 ^ n12162 ^ n11386 ;
  assign n16769 = ~n1640 & n7031 ;
  assign n16770 = n16769 ^ n4185 ^ 1'b0 ;
  assign n16771 = ( n1197 & n14397 ) | ( n1197 & n16770 ) | ( n14397 & n16770 ) ;
  assign n16772 = n6598 | n16771 ;
  assign n16773 = n998 & ~n15811 ;
  assign n16774 = n16773 ^ n5800 ^ 1'b0 ;
  assign n16776 = n2165 & n16345 ;
  assign n16777 = ( n4845 & n10412 ) | ( n4845 & n16776 ) | ( n10412 & n16776 ) ;
  assign n16775 = ~n4246 & n11239 ;
  assign n16778 = n16777 ^ n16775 ^ 1'b0 ;
  assign n16779 = ~n6269 & n15824 ;
  assign n16780 = ~n241 & n16779 ;
  assign n16781 = n1606 ^ n316 ^ 1'b0 ;
  assign n16782 = n8000 ^ n3334 ^ n1796 ;
  assign n16783 = ~n398 & n2490 ;
  assign n16784 = ~n16782 & n16783 ;
  assign n16785 = n16784 ^ n10488 ^ 1'b0 ;
  assign n16786 = ~n16781 & n16785 ;
  assign n16787 = n14101 ^ n7665 ^ 1'b0 ;
  assign n16788 = n5264 & ~n16787 ;
  assign n16789 = ~n9982 & n16788 ;
  assign n16790 = n3853 | n4417 ;
  assign n16791 = n16790 ^ n2954 ^ n1825 ;
  assign n16792 = n14049 ^ n4269 ^ 1'b0 ;
  assign n16793 = ( n1823 & n16791 ) | ( n1823 & ~n16792 ) | ( n16791 & ~n16792 ) ;
  assign n16794 = n5182 & ~n16793 ;
  assign n16795 = n5599 & n16794 ;
  assign n16796 = n9838 & n16795 ;
  assign n16797 = n16796 ^ n11288 ^ n6497 ;
  assign n16798 = n1017 & n1761 ;
  assign n16799 = ~n108 & n7249 ;
  assign n16800 = n7363 ^ n6306 ^ 1'b0 ;
  assign n16801 = n16799 | n16800 ;
  assign n16802 = ~n324 & n630 ;
  assign n16803 = n6662 & ~n16802 ;
  assign n16804 = ~n1482 & n16803 ;
  assign n16805 = ( n166 & n16801 ) | ( n166 & ~n16804 ) | ( n16801 & ~n16804 ) ;
  assign n16808 = n15246 ^ n9790 ^ 1'b0 ;
  assign n16809 = n14141 & n16808 ;
  assign n16806 = n11021 & n11769 ;
  assign n16807 = n1679 & ~n16806 ;
  assign n16810 = n16809 ^ n16807 ^ 1'b0 ;
  assign n16811 = ( n5488 & ~n9226 ) | ( n5488 & n12221 ) | ( ~n9226 & n12221 ) ;
  assign n16812 = n11908 ^ n4719 ^ 1'b0 ;
  assign n16813 = ~n503 & n16750 ;
  assign n16814 = n525 & n5908 ;
  assign n16815 = n9984 ^ n8712 ^ 1'b0 ;
  assign n16816 = n8849 & n16815 ;
  assign n16817 = ~n1492 & n7304 ;
  assign n16818 = ~n16816 & n16817 ;
  assign n16819 = ~n5311 & n11786 ;
  assign n16820 = n650 | n2080 ;
  assign n16821 = ~n6569 & n16820 ;
  assign n16822 = ( n141 & n3738 ) | ( n141 & n11754 ) | ( n3738 & n11754 ) ;
  assign n16823 = n4226 ^ n3173 ^ n1851 ;
  assign n16824 = ( n5508 & ~n16822 ) | ( n5508 & n16823 ) | ( ~n16822 & n16823 ) ;
  assign n16825 = n4620 & n16824 ;
  assign n16826 = n9206 ^ n5391 ^ 1'b0 ;
  assign n16827 = ( ~n2612 & n14261 ) | ( ~n2612 & n16826 ) | ( n14261 & n16826 ) ;
  assign n16828 = n6155 ^ n3663 ^ 1'b0 ;
  assign n16829 = n10018 & n16828 ;
  assign n16832 = ~n893 & n2011 ;
  assign n16830 = ( n130 & n13479 ) | ( n130 & ~n15950 ) | ( n13479 & ~n15950 ) ;
  assign n16831 = ~n734 & n16830 ;
  assign n16833 = n16832 ^ n16831 ^ 1'b0 ;
  assign n16834 = ~n2857 & n4019 ;
  assign n16835 = ~n16833 & n16834 ;
  assign n16836 = n8458 & n9257 ;
  assign n16837 = n13064 ^ n3313 ^ 1'b0 ;
  assign n16838 = n16837 ^ n16672 ^ n15153 ;
  assign n16839 = n9105 & ~n13881 ;
  assign n16840 = ~n13774 & n16839 ;
  assign n16842 = ~n4543 & n8780 ;
  assign n16843 = n16842 ^ n1858 ^ 1'b0 ;
  assign n16841 = n3367 ^ n1317 ^ 1'b0 ;
  assign n16844 = n16843 ^ n16841 ^ n11069 ;
  assign n16845 = n16517 & ~n16844 ;
  assign n16846 = n10049 & n16845 ;
  assign n16853 = n13315 ^ n5552 ^ 1'b0 ;
  assign n16849 = n5029 ^ n3920 ^ 1'b0 ;
  assign n16850 = n9967 & n16849 ;
  assign n16851 = n16850 ^ n16016 ^ 1'b0 ;
  assign n16847 = n67 & ~n2327 ;
  assign n16848 = n7273 | n16847 ;
  assign n16852 = n16851 ^ n16848 ^ 1'b0 ;
  assign n16854 = n16853 ^ n16852 ^ 1'b0 ;
  assign n16855 = n8239 ^ n2665 ^ n2403 ;
  assign n16856 = n16443 ^ n10695 ^ 1'b0 ;
  assign n16857 = ~n9770 & n16856 ;
  assign n16858 = n3229 & ~n16857 ;
  assign n16859 = n16858 ^ n12668 ^ n4737 ;
  assign n16860 = n2992 & ~n10115 ;
  assign n16861 = n16860 ^ n7166 ^ 1'b0 ;
  assign n16862 = n16861 ^ n4490 ^ 1'b0 ;
  assign n16863 = n1433 & ~n16862 ;
  assign n16864 = n3037 & ~n15920 ;
  assign n16865 = ( ~n4927 & n6641 ) | ( ~n4927 & n7529 ) | ( n6641 & n7529 ) ;
  assign n16866 = n16865 ^ n5800 ^ 1'b0 ;
  assign n16867 = ~n6116 & n16866 ;
  assign n16868 = ( n1109 & ~n3564 ) | ( n1109 & n12703 ) | ( ~n3564 & n12703 ) ;
  assign n16869 = n1956 | n3911 ;
  assign n16870 = n4077 & ~n16869 ;
  assign n16871 = n14211 ^ n13987 ^ 1'b0 ;
  assign n16872 = ~n16870 & n16871 ;
  assign n16873 = n16232 & n16872 ;
  assign n16874 = n8496 ^ n2070 ^ 1'b0 ;
  assign n16875 = ~n523 & n16874 ;
  assign n16876 = n16875 ^ n1195 ^ 1'b0 ;
  assign n16877 = n16876 ^ n12116 ^ 1'b0 ;
  assign n16878 = n6067 ^ n1506 ^ n310 ;
  assign n16879 = ~n15982 & n16091 ;
  assign n16880 = n2689 & ~n9683 ;
  assign n16881 = ~n1964 & n16880 ;
  assign n16882 = n13918 ^ n5051 ^ 1'b0 ;
  assign n16883 = n9783 ^ n9011 ^ n4313 ;
  assign n16884 = n15617 ^ n40 ^ 1'b0 ;
  assign n16885 = ~n16883 & n16884 ;
  assign n16886 = n1808 & n2190 ;
  assign n16887 = n6835 & n16886 ;
  assign n16888 = n10998 & ~n16887 ;
  assign n16889 = n1783 & n7740 ;
  assign n16890 = ( ~n4632 & n12115 ) | ( ~n4632 & n16889 ) | ( n12115 & n16889 ) ;
  assign n16891 = n6251 & n11671 ;
  assign n16892 = n8920 & ~n13548 ;
  assign n16893 = n13548 & n16892 ;
  assign n16894 = n10488 ^ n2471 ^ 1'b0 ;
  assign n16895 = n3938 ^ n2485 ^ 1'b0 ;
  assign n16896 = n4132 | n16895 ;
  assign n16897 = n2638 & ~n16896 ;
  assign n16898 = n16897 ^ n9279 ^ 1'b0 ;
  assign n16899 = n4192 | n11371 ;
  assign n16900 = ~n8435 & n16899 ;
  assign n16901 = n1845 & n16900 ;
  assign n16902 = n710 & ~n16901 ;
  assign n16903 = n16902 ^ n1348 ^ 1'b0 ;
  assign n16904 = ~n1339 & n15765 ;
  assign n16905 = n13747 ^ n3727 ^ 1'b0 ;
  assign n16906 = n8125 & n16905 ;
  assign n16907 = n12020 & ~n14526 ;
  assign n16910 = ~n3522 & n8342 ;
  assign n16908 = n590 & ~n14066 ;
  assign n16909 = n2960 & n16908 ;
  assign n16911 = n16910 ^ n16909 ^ 1'b0 ;
  assign n16912 = n3871 ^ n2858 ^ 1'b0 ;
  assign n16913 = ( n8917 & n10348 ) | ( n8917 & ~n16912 ) | ( n10348 & ~n16912 ) ;
  assign n16914 = ~n5573 & n8209 ;
  assign n16915 = n4260 | n16914 ;
  assign n16916 = n1600 & n12685 ;
  assign n16917 = ~n16915 & n16916 ;
  assign n16918 = n5237 & n16917 ;
  assign n16919 = n9120 ^ n6808 ^ 1'b0 ;
  assign n16920 = ~n16504 & n16919 ;
  assign n16921 = ~n670 & n4568 ;
  assign n16922 = n16921 ^ n1177 ^ 1'b0 ;
  assign n16923 = n1781 ^ n971 ^ 1'b0 ;
  assign n16924 = n3252 | n6315 ;
  assign n16925 = n16923 | n16924 ;
  assign n16926 = ~n16922 & n16925 ;
  assign n16927 = n16926 ^ n5312 ^ 1'b0 ;
  assign n16929 = n2607 | n3488 ;
  assign n16930 = n1125 | n16929 ;
  assign n16928 = n4422 & ~n15399 ;
  assign n16931 = n16930 ^ n16928 ^ 1'b0 ;
  assign n16932 = n9565 ^ n1182 ^ 1'b0 ;
  assign n16933 = n11139 | n16932 ;
  assign n16934 = n16933 ^ n12641 ^ 1'b0 ;
  assign n16935 = n187 & ~n16934 ;
  assign n16936 = n14192 & ~n16935 ;
  assign n16937 = n16126 ^ n9824 ^ 1'b0 ;
  assign n16938 = n838 | n16937 ;
  assign n16939 = n16331 ^ n14674 ^ n5115 ;
  assign n16940 = n1004 & n1960 ;
  assign n16941 = n2076 & ~n16940 ;
  assign n16942 = n16939 & n16941 ;
  assign n16943 = n10274 ^ n1493 ^ 1'b0 ;
  assign n16944 = n15589 & ~n16943 ;
  assign n16945 = ~n7234 & n16944 ;
  assign n16946 = n11715 & n16945 ;
  assign n16947 = ( n6635 & n11563 ) | ( n6635 & n14475 ) | ( n11563 & n14475 ) ;
  assign n16948 = n10309 ^ n4208 ^ n1700 ;
  assign n16949 = n11247 | n16948 ;
  assign n16950 = n16947 | n16949 ;
  assign n16951 = n14282 ^ n4769 ^ 1'b0 ;
  assign n16952 = n8355 ^ n804 ^ 1'b0 ;
  assign n16953 = n8145 & ~n16952 ;
  assign n16954 = ( n830 & n7270 ) | ( n830 & ~n9213 ) | ( n7270 & ~n9213 ) ;
  assign n16955 = ( n12119 & n14063 ) | ( n12119 & n16954 ) | ( n14063 & n16954 ) ;
  assign n16956 = ~n7930 & n8242 ;
  assign n16957 = n8582 & n16956 ;
  assign n16958 = n1875 | n16957 ;
  assign n16959 = n3041 & ~n16958 ;
  assign n16960 = n16279 ^ n14653 ^ 1'b0 ;
  assign n16961 = n14009 & ~n16960 ;
  assign n16962 = n1290 & n11300 ;
  assign n16963 = n466 & n16962 ;
  assign n16964 = n11164 ^ n2333 ^ 1'b0 ;
  assign n16965 = n4638 & ~n16964 ;
  assign n16966 = n2542 ^ x11 ^ 1'b0 ;
  assign n16967 = n16966 ^ n15061 ^ n2483 ;
  assign n16968 = ~n3603 & n4495 ;
  assign n16969 = ~n6119 & n16968 ;
  assign n16970 = n11543 | n16969 ;
  assign n16971 = n3966 | n16970 ;
  assign n16972 = n3868 | n7151 ;
  assign n16973 = n15701 | n16972 ;
  assign n16974 = n16973 ^ n4652 ^ n3803 ;
  assign n16975 = n7851 & n16974 ;
  assign n16976 = n16975 ^ n6201 ^ 1'b0 ;
  assign n16977 = ( n1029 & n5490 ) | ( n1029 & ~n13175 ) | ( n5490 & ~n13175 ) ;
  assign n16979 = ( ~n5175 & n8625 ) | ( ~n5175 & n11682 ) | ( n8625 & n11682 ) ;
  assign n16978 = n15488 | n16847 ;
  assign n16980 = n16979 ^ n16978 ^ 1'b0 ;
  assign n16981 = n16977 & n16980 ;
  assign n16982 = n16981 ^ n3712 ^ 1'b0 ;
  assign n16983 = n5111 | n16068 ;
  assign n16984 = n11426 ^ n9907 ^ 1'b0 ;
  assign n16985 = n15892 | n16984 ;
  assign n16986 = n16985 ^ n15581 ^ 1'b0 ;
  assign n16987 = n3824 ^ n383 ^ 1'b0 ;
  assign n16988 = n16986 & n16987 ;
  assign n16989 = n2992 | n3195 ;
  assign n16990 = n16989 ^ n1374 ^ 1'b0 ;
  assign n16991 = ( n8895 & ~n15347 ) | ( n8895 & n16990 ) | ( ~n15347 & n16990 ) ;
  assign n16992 = n6169 & ~n16991 ;
  assign n16993 = n11722 & n16992 ;
  assign n16995 = n12420 ^ n4700 ^ 1'b0 ;
  assign n16996 = ~n102 & n16995 ;
  assign n16994 = n1824 & ~n7440 ;
  assign n16997 = n16996 ^ n16994 ^ 1'b0 ;
  assign n16998 = n141 & ~n3976 ;
  assign n16999 = n10072 & ~n16998 ;
  assign n17000 = n6707 & n16999 ;
  assign n17001 = n4432 | n9939 ;
  assign n17002 = n16596 ^ n9168 ^ 1'b0 ;
  assign n17003 = n17001 | n17002 ;
  assign n17004 = n2899 & n8843 ;
  assign n17005 = n13772 & n17004 ;
  assign n17006 = n14781 ^ n9127 ^ 1'b0 ;
  assign n17007 = n6199 & ~n17006 ;
  assign n17008 = ~n1312 & n17007 ;
  assign n17009 = n17005 | n17008 ;
  assign n17010 = n15282 & ~n17009 ;
  assign n17011 = n6821 ^ n486 ^ 1'b0 ;
  assign n17012 = ~n434 & n17011 ;
  assign n17013 = n3979 ^ n3112 ^ 1'b0 ;
  assign n17014 = n17013 ^ n9224 ^ n183 ;
  assign n17015 = n469 & n6352 ;
  assign n17016 = n14462 ^ n4925 ^ 1'b0 ;
  assign n17023 = n560 ^ n125 ^ 1'b0 ;
  assign n17024 = n17023 ^ n7780 ^ n4272 ;
  assign n17025 = n17024 ^ n4059 ^ 1'b0 ;
  assign n17026 = ~n10897 & n17025 ;
  assign n17017 = n929 & n6099 ;
  assign n17018 = n17017 ^ n7004 ^ 1'b0 ;
  assign n17019 = n16068 & n17018 ;
  assign n17020 = ( ~n3016 & n5047 ) | ( ~n3016 & n15791 ) | ( n5047 & n15791 ) ;
  assign n17021 = ( n1904 & ~n12851 ) | ( n1904 & n17020 ) | ( ~n12851 & n17020 ) ;
  assign n17022 = ~n17019 & n17021 ;
  assign n17027 = n17026 ^ n17022 ^ 1'b0 ;
  assign n17028 = n4657 ^ n4192 ^ 1'b0 ;
  assign n17029 = ~n13965 & n17028 ;
  assign n17030 = n11269 ^ n8868 ^ 1'b0 ;
  assign n17031 = n17030 ^ n1658 ^ 1'b0 ;
  assign n17032 = n10267 ^ n6722 ^ 1'b0 ;
  assign n17033 = n13397 & ~n17032 ;
  assign n17037 = n3864 ^ n1481 ^ n1318 ;
  assign n17034 = n688 ^ n139 ^ 1'b0 ;
  assign n17035 = n3104 | n17034 ;
  assign n17036 = n17035 ^ n11196 ^ 1'b0 ;
  assign n17038 = n17037 ^ n17036 ^ n1168 ;
  assign n17039 = n17038 ^ n1511 ^ 1'b0 ;
  assign n17040 = n17033 & ~n17039 ;
  assign n17041 = n17040 ^ n15066 ^ 1'b0 ;
  assign n17042 = n7275 ^ n3288 ^ 1'b0 ;
  assign n17043 = n13688 & ~n13735 ;
  assign n17044 = n1800 & n17043 ;
  assign n17045 = n17044 ^ n2514 ^ 1'b0 ;
  assign n17048 = n10841 ^ n6251 ^ 1'b0 ;
  assign n17049 = n8239 & ~n17048 ;
  assign n17046 = ( n1374 & ~n1521 ) | ( n1374 & n13062 ) | ( ~n1521 & n13062 ) ;
  assign n17047 = n9072 & n17046 ;
  assign n17050 = n17049 ^ n17047 ^ 1'b0 ;
  assign n17051 = n9847 & ~n17050 ;
  assign n17052 = n4825 | n7988 ;
  assign n17053 = n8333 | n17052 ;
  assign n17054 = n2475 ^ n1232 ^ 1'b0 ;
  assign n17055 = n17054 ^ n11757 ^ 1'b0 ;
  assign n17056 = n3350 & ~n17055 ;
  assign n17057 = ~n5797 & n17056 ;
  assign n17058 = n11177 ^ n1929 ^ 1'b0 ;
  assign n17059 = n4057 | n13437 ;
  assign n17060 = ( n400 & n3443 ) | ( n400 & n17059 ) | ( n3443 & n17059 ) ;
  assign n17061 = n3000 & n8407 ;
  assign n17062 = ~n1932 & n17061 ;
  assign n17063 = n4827 | n17062 ;
  assign n17064 = n7307 | n17063 ;
  assign n17065 = ~n3530 & n17064 ;
  assign n17067 = n4647 ^ n3085 ^ 1'b0 ;
  assign n17068 = n3902 | n17067 ;
  assign n17069 = n3079 | n17068 ;
  assign n17066 = n4819 & ~n7040 ;
  assign n17070 = n17069 ^ n17066 ^ 1'b0 ;
  assign n17076 = n5051 & ~n10178 ;
  assign n17077 = n5538 & n17076 ;
  assign n17071 = n3637 & n7804 ;
  assign n17072 = ~n3637 & n17071 ;
  assign n17073 = n4796 | n17072 ;
  assign n17074 = n4796 & ~n17073 ;
  assign n17075 = ( n6415 & ~n11796 ) | ( n6415 & n17074 ) | ( ~n11796 & n17074 ) ;
  assign n17078 = n17077 ^ n17075 ^ 1'b0 ;
  assign n17079 = n1244 & ~n17078 ;
  assign n17080 = n11693 ^ n922 ^ 1'b0 ;
  assign n17081 = n17079 & ~n17080 ;
  assign n17082 = n16550 ^ n771 ^ 1'b0 ;
  assign n17083 = n1869 & ~n17082 ;
  assign n17084 = n2986 ^ n1590 ^ n101 ;
  assign n17085 = n17084 ^ n7393 ^ n6882 ;
  assign n17086 = ~n6024 & n6718 ;
  assign n17087 = n378 | n17086 ;
  assign n17088 = n17087 ^ n5163 ^ 1'b0 ;
  assign n17089 = ~n6067 & n9094 ;
  assign n17090 = n960 & ~n2385 ;
  assign n17091 = ~n2930 & n17090 ;
  assign n17092 = ~n17089 & n17091 ;
  assign n17093 = ~n2067 & n6128 ;
  assign n17094 = n17093 ^ n3275 ^ 1'b0 ;
  assign n17095 = n14032 ^ n13265 ^ 1'b0 ;
  assign n17096 = n13362 ^ n11500 ^ 1'b0 ;
  assign n17097 = n17096 ^ n9601 ^ 1'b0 ;
  assign n17099 = n5596 ^ n3997 ^ n1017 ;
  assign n17098 = n6369 & n7886 ;
  assign n17100 = n17099 ^ n17098 ^ 1'b0 ;
  assign n17101 = n1775 & n7860 ;
  assign n17102 = ~n13222 & n17101 ;
  assign n17103 = n6673 ^ n5428 ^ 1'b0 ;
  assign n17104 = ~n14881 & n17103 ;
  assign n17105 = n824 | n1553 ;
  assign n17106 = n122 | n17105 ;
  assign n17107 = n8988 | n17106 ;
  assign n17108 = ( n5269 & ~n17104 ) | ( n5269 & n17107 ) | ( ~n17104 & n17107 ) ;
  assign n17109 = ~n2581 & n6146 ;
  assign n17110 = n554 & ~n3270 ;
  assign n17111 = ~n3363 & n17110 ;
  assign n17112 = n1715 & n17111 ;
  assign n17113 = n17112 ^ n5469 ^ 1'b0 ;
  assign n17114 = n8203 & n8332 ;
  assign n17115 = n3359 & n7545 ;
  assign n17116 = n17115 ^ n7706 ^ 1'b0 ;
  assign n17117 = n14075 | n17116 ;
  assign n17118 = n17114 | n17117 ;
  assign n17119 = ( ~n2393 & n10949 ) | ( ~n2393 & n11796 ) | ( n10949 & n11796 ) ;
  assign n17120 = n17119 ^ n7872 ^ 1'b0 ;
  assign n17121 = n991 | n17120 ;
  assign n17123 = n3853 ^ n252 ^ 1'b0 ;
  assign n17122 = n1720 ^ n518 ^ 1'b0 ;
  assign n17124 = n17123 ^ n17122 ^ 1'b0 ;
  assign n17125 = n6167 & ~n17124 ;
  assign n17127 = n1990 & ~n6366 ;
  assign n17128 = n17127 ^ n8789 ^ 1'b0 ;
  assign n17126 = ~n895 & n8797 ;
  assign n17129 = n17128 ^ n17126 ^ 1'b0 ;
  assign n17130 = n5803 ^ n5545 ^ 1'b0 ;
  assign n17131 = ~n17129 & n17130 ;
  assign n17132 = ~n694 & n17131 ;
  assign n17133 = ~n9753 & n17132 ;
  assign n17134 = ~n4341 & n6413 ;
  assign n17135 = ( n8607 & n11213 ) | ( n8607 & ~n17134 ) | ( n11213 & ~n17134 ) ;
  assign n17136 = n885 & n12010 ;
  assign n17137 = n4327 | n17136 ;
  assign n17138 = n5946 & n6328 ;
  assign n17139 = n17138 ^ n14604 ^ n805 ;
  assign n17140 = n8071 & ~n11769 ;
  assign n17141 = n15454 ^ n3609 ^ n1281 ;
  assign n17142 = n14845 & ~n17141 ;
  assign n17143 = n3051 ^ n2145 ^ 1'b0 ;
  assign n17144 = n7949 & ~n12507 ;
  assign n17145 = n17144 ^ n3155 ^ 1'b0 ;
  assign n17146 = n13854 ^ n6277 ^ n1167 ;
  assign n17147 = ~n637 & n4249 ;
  assign n17148 = n10406 ^ n553 ^ 1'b0 ;
  assign n17149 = n17147 & n17148 ;
  assign n17150 = ~n17146 & n17149 ;
  assign n17151 = n401 & n16783 ;
  assign n17152 = n8889 ^ n361 ^ 1'b0 ;
  assign n17153 = ( n5114 & n7977 ) | ( n5114 & n17152 ) | ( n7977 & n17152 ) ;
  assign n17154 = n7746 & n8086 ;
  assign n17155 = n17153 & n17154 ;
  assign n17156 = n16641 & n17155 ;
  assign n17157 = n17156 ^ n12727 ^ 1'b0 ;
  assign n17158 = ~n4544 & n17157 ;
  assign n17159 = ~n3259 & n7164 ;
  assign n17160 = n17159 ^ n11029 ^ 1'b0 ;
  assign n17161 = n1287 | n3790 ;
  assign n17162 = n882 & ~n17161 ;
  assign n17163 = n8158 | n17162 ;
  assign n17164 = n10820 & ~n17163 ;
  assign n17165 = ~n6071 & n17164 ;
  assign n17166 = ~n211 & n2561 ;
  assign n17167 = ~n8025 & n17166 ;
  assign n17168 = n10956 & n17167 ;
  assign n17169 = n1260 ^ n886 ^ 1'b0 ;
  assign n17170 = n17169 ^ n8938 ^ 1'b0 ;
  assign n17171 = n17170 ^ n13980 ^ 1'b0 ;
  assign n17173 = n16064 ^ n2340 ^ 1'b0 ;
  assign n17172 = n3056 | n3823 ;
  assign n17174 = n17173 ^ n17172 ^ 1'b0 ;
  assign n17175 = n14776 ^ n7696 ^ 1'b0 ;
  assign n17176 = n15112 ^ n12541 ^ 1'b0 ;
  assign n17177 = ~n13243 & n17176 ;
  assign n17178 = n7807 & ~n9075 ;
  assign n17179 = n17178 ^ n6743 ^ 1'b0 ;
  assign n17180 = n10824 ^ n57 ^ 1'b0 ;
  assign n17181 = ~n2486 & n13097 ;
  assign n17182 = n5691 ^ n4359 ^ n1300 ;
  assign n17185 = n1220 ^ n342 ^ 1'b0 ;
  assign n17183 = ~n6819 & n12049 ;
  assign n17184 = n14177 | n17183 ;
  assign n17186 = n17185 ^ n17184 ^ 1'b0 ;
  assign n17187 = n17186 ^ n8380 ^ 1'b0 ;
  assign n17188 = n16822 ^ n9775 ^ 1'b0 ;
  assign n17189 = n2679 & n17188 ;
  assign n17190 = n17189 ^ n2081 ^ n306 ;
  assign n17191 = n4315 | n12885 ;
  assign n17192 = n17190 & ~n17191 ;
  assign n17193 = n7449 & ~n10167 ;
  assign n17194 = n17193 ^ n4838 ^ 1'b0 ;
  assign n17195 = n17194 ^ n8709 ^ 1'b0 ;
  assign n17196 = n13890 & n17195 ;
  assign n17197 = ( n1694 & n6166 ) | ( n1694 & ~n10427 ) | ( n6166 & ~n10427 ) ;
  assign n17198 = ~n9713 & n17197 ;
  assign n17199 = n3245 & n17198 ;
  assign n17200 = ( n3975 & n14937 ) | ( n3975 & n17199 ) | ( n14937 & n17199 ) ;
  assign n17201 = n3184 | n17200 ;
  assign n17202 = ~n2885 & n8660 ;
  assign n17203 = n16738 ^ n957 ^ n260 ;
  assign n17204 = n17203 ^ n15824 ^ 1'b0 ;
  assign n17205 = n10185 | n17204 ;
  assign n17206 = n7049 | n17205 ;
  assign n17208 = n13315 ^ n6166 ^ n51 ;
  assign n17207 = n8098 ^ n5590 ^ 1'b0 ;
  assign n17209 = n17208 ^ n17207 ^ 1'b0 ;
  assign n17210 = n17206 & ~n17209 ;
  assign n17211 = ~n6482 & n17210 ;
  assign n17212 = n17211 ^ n12634 ^ 1'b0 ;
  assign n17213 = n6903 ^ n150 ^ 1'b0 ;
  assign n17214 = n2584 & n17213 ;
  assign n17215 = ~n65 & n17214 ;
  assign n17216 = n9752 & n17215 ;
  assign n17217 = n10088 ^ n4445 ^ 1'b0 ;
  assign n17218 = n15046 ^ n15031 ^ n13088 ;
  assign n17219 = n4435 | n11915 ;
  assign n17220 = n17219 ^ n1990 ^ 1'b0 ;
  assign n17221 = ~n4560 & n17220 ;
  assign n17222 = n16652 & n17221 ;
  assign n17223 = n9951 | n15238 ;
  assign n17225 = n2089 & ~n8014 ;
  assign n17226 = ~n7542 & n17225 ;
  assign n17227 = n411 & ~n17226 ;
  assign n17224 = n2130 & n5864 ;
  assign n17228 = n17227 ^ n17224 ^ n1656 ;
  assign n17229 = n8493 ^ n5016 ^ 1'b0 ;
  assign n17230 = n176 & ~n5667 ;
  assign n17231 = n17230 ^ n15593 ^ 1'b0 ;
  assign n17232 = n242 | n17231 ;
  assign n17233 = n17232 ^ n16628 ^ 1'b0 ;
  assign n17234 = n7749 ^ n809 ^ 1'b0 ;
  assign n17235 = n471 | n17234 ;
  assign n17236 = ~n4750 & n5231 ;
  assign n17237 = n17235 | n17236 ;
  assign n17238 = n9144 & n13208 ;
  assign n17239 = n17238 ^ n9748 ^ 1'b0 ;
  assign n17240 = n5321 & n6030 ;
  assign n17241 = n16294 ^ n9246 ^ n3134 ;
  assign n17242 = n17241 ^ n14506 ^ 1'b0 ;
  assign n17243 = n5495 ^ n336 ^ 1'b0 ;
  assign n17244 = n17243 ^ n122 ^ 1'b0 ;
  assign n17245 = ~n6430 & n13568 ;
  assign n17248 = n1083 & n7761 ;
  assign n17249 = n6275 & n17248 ;
  assign n17246 = n3858 & ~n3912 ;
  assign n17247 = n17246 ^ n3370 ^ 1'b0 ;
  assign n17250 = n17249 ^ n17247 ^ n6089 ;
  assign n17251 = n3387 ^ n2382 ^ n1745 ;
  assign n17252 = n4485 | n17251 ;
  assign n17253 = n3925 | n9656 ;
  assign n17254 = n2391 | n17253 ;
  assign n17255 = n17254 ^ n4359 ^ 1'b0 ;
  assign n17256 = n11626 & ~n17255 ;
  assign n17257 = n1263 ^ n609 ^ 1'b0 ;
  assign n17258 = n17257 ^ n918 ^ 1'b0 ;
  assign n17259 = n6420 | n11288 ;
  assign n17260 = n8857 | n11773 ;
  assign n17261 = n15928 | n17260 ;
  assign n17262 = n17261 ^ n7237 ^ 1'b0 ;
  assign n17263 = n3299 ^ n134 ^ 1'b0 ;
  assign n17264 = n10747 & n17263 ;
  assign n17265 = n11749 & ~n12372 ;
  assign n17266 = ~n3912 & n17265 ;
  assign n17267 = n680 & n2206 ;
  assign n17268 = n17267 ^ n4150 ^ 1'b0 ;
  assign n17269 = ~n25 & n17268 ;
  assign n17270 = ~n3977 & n17269 ;
  assign n17271 = n6890 & n11824 ;
  assign n17272 = n7242 | n17271 ;
  assign n17273 = n13396 ^ n1880 ^ 1'b0 ;
  assign n17274 = n17273 ^ n6924 ^ 1'b0 ;
  assign n17275 = n8590 & n9550 ;
  assign n17276 = ( n118 & ~n7523 ) | ( n118 & n9787 ) | ( ~n7523 & n9787 ) ;
  assign n17277 = ( n2320 & n14985 ) | ( n2320 & n17276 ) | ( n14985 & n17276 ) ;
  assign n17278 = n2397 & ~n3759 ;
  assign n17279 = n1694 & n17278 ;
  assign n17280 = n17279 ^ n2190 ^ 1'b0 ;
  assign n17281 = n1279 | n5764 ;
  assign n17282 = n17281 ^ n7363 ^ 1'b0 ;
  assign n17283 = ~n1097 & n4394 ;
  assign n17284 = n15597 | n17283 ;
  assign n17285 = n17284 ^ n195 ^ 1'b0 ;
  assign n17286 = n17285 ^ n6214 ^ 1'b0 ;
  assign n17287 = ~n17282 & n17286 ;
  assign n17288 = n17287 ^ n15800 ^ 1'b0 ;
  assign n17289 = n1606 & n17288 ;
  assign n17291 = n3081 ^ n2864 ^ 1'b0 ;
  assign n17290 = n2391 & ~n4668 ;
  assign n17292 = n17291 ^ n17290 ^ 1'b0 ;
  assign n17293 = n8780 & ~n17292 ;
  assign n17294 = ~n4990 & n10943 ;
  assign n17295 = ~n3084 & n17294 ;
  assign n17296 = ( n8615 & n17293 ) | ( n8615 & n17295 ) | ( n17293 & n17295 ) ;
  assign n17297 = n5529 ^ n4011 ^ 1'b0 ;
  assign n17298 = ~n6309 & n8020 ;
  assign n17299 = n548 & n17298 ;
  assign n17300 = n5301 | n8006 ;
  assign n17301 = n7740 | n17300 ;
  assign n17302 = n15674 ^ n1877 ^ 1'b0 ;
  assign n17303 = n8854 ^ n7631 ^ 1'b0 ;
  assign n17304 = n76 | n4719 ;
  assign n17305 = ~n13453 & n17304 ;
  assign n17306 = n11601 & n17305 ;
  assign n17307 = n17303 & n17306 ;
  assign n17308 = n7956 ^ n3030 ^ n601 ;
  assign n17309 = n3832 | n6896 ;
  assign n17310 = n1666 ^ n761 ^ 1'b0 ;
  assign n17311 = n17310 ^ n16461 ^ n14696 ;
  assign n17314 = x10 & ~n9667 ;
  assign n17315 = n4189 & n17314 ;
  assign n17312 = n7839 ^ n4512 ^ 1'b0 ;
  assign n17313 = ~n10695 & n17312 ;
  assign n17316 = n17315 ^ n17313 ^ 1'b0 ;
  assign n17317 = n10793 ^ n6659 ^ 1'b0 ;
  assign n17318 = ~n5740 & n15999 ;
  assign n17319 = ~n16034 & n17318 ;
  assign n17320 = n17319 ^ n1485 ^ 1'b0 ;
  assign n17321 = ( n7017 & n17317 ) | ( n7017 & ~n17320 ) | ( n17317 & ~n17320 ) ;
  assign n17322 = n17321 ^ n1278 ^ 1'b0 ;
  assign n17323 = ~n2101 & n17322 ;
  assign n17324 = n2012 & ~n13965 ;
  assign n17326 = ( n5391 & n12286 ) | ( n5391 & ~n13157 ) | ( n12286 & ~n13157 ) ;
  assign n17325 = n3381 | n8592 ;
  assign n17327 = n17326 ^ n17325 ^ 1'b0 ;
  assign n17328 = ~n10472 & n10795 ;
  assign n17329 = n17328 ^ n3354 ^ 1'b0 ;
  assign n17332 = n5352 ^ n3463 ^ n1699 ;
  assign n17330 = n4520 & n8199 ;
  assign n17331 = n17330 ^ n4053 ^ 1'b0 ;
  assign n17333 = n17332 ^ n17331 ^ n13467 ;
  assign n17334 = ~n9791 & n17333 ;
  assign n17335 = n17189 ^ n11766 ^ n7535 ;
  assign n17336 = n5973 | n13909 ;
  assign n17337 = n8195 & ~n17336 ;
  assign n17338 = n17337 ^ n3888 ^ 1'b0 ;
  assign n17340 = n4269 & n6743 ;
  assign n17341 = ~n853 & n17340 ;
  assign n17339 = n3199 ^ n1465 ^ 1'b0 ;
  assign n17342 = n17341 ^ n17339 ^ 1'b0 ;
  assign n17343 = n2154 | n12209 ;
  assign n17352 = n445 & n4595 ;
  assign n17344 = n440 | n13531 ;
  assign n17345 = n17344 ^ n3035 ^ 1'b0 ;
  assign n17346 = n1715 | n3706 ;
  assign n17347 = ~n1348 & n17346 ;
  assign n17348 = ~n6468 & n17347 ;
  assign n17349 = n17348 ^ n3640 ^ 1'b0 ;
  assign n17350 = n17349 ^ n688 ^ 1'b0 ;
  assign n17351 = n17345 & n17350 ;
  assign n17353 = n17352 ^ n17351 ^ 1'b0 ;
  assign n17354 = ~n7460 & n17353 ;
  assign n17355 = n3309 & ~n17354 ;
  assign n17356 = n8897 ^ n7672 ^ n3464 ;
  assign n17357 = ( n11083 & n11340 ) | ( n11083 & ~n15712 ) | ( n11340 & ~n15712 ) ;
  assign n17359 = n11815 ^ n5224 ^ 1'b0 ;
  assign n17358 = n1108 & n4460 ;
  assign n17360 = n17359 ^ n17358 ^ 1'b0 ;
  assign n17361 = ~n10337 & n14710 ;
  assign n17362 = n3997 & n17361 ;
  assign n17363 = n6076 | n16785 ;
  assign n17364 = n17362 & ~n17363 ;
  assign n17365 = n860 | n17364 ;
  assign n17366 = ~n3761 & n5227 ;
  assign n17367 = ~n7055 & n17366 ;
  assign n17368 = ~n2858 & n3432 ;
  assign n17369 = n17368 ^ n4993 ^ 1'b0 ;
  assign n17370 = n17369 ^ n11999 ^ 1'b0 ;
  assign n17371 = n2716 & n17370 ;
  assign n17372 = n17371 ^ n15909 ^ 1'b0 ;
  assign n17373 = n5353 & n17372 ;
  assign n17374 = n12618 & n13854 ;
  assign n17375 = n3295 ^ n786 ^ 1'b0 ;
  assign n17376 = ~n12852 & n17375 ;
  assign n17377 = n8832 ^ n7017 ^ n1294 ;
  assign n17378 = ( n6587 & n8918 ) | ( n6587 & n17377 ) | ( n8918 & n17377 ) ;
  assign n17379 = n4402 & ~n15568 ;
  assign n17380 = n320 & n17379 ;
  assign n17381 = n11241 | n17380 ;
  assign n17382 = n1189 & ~n17381 ;
  assign n17383 = n17382 ^ n8406 ^ 1'b0 ;
  assign n17384 = ( ~n6413 & n6852 ) | ( ~n6413 & n10094 ) | ( n6852 & n10094 ) ;
  assign n17385 = n17384 ^ n4888 ^ 1'b0 ;
  assign n17386 = n12658 | n17385 ;
  assign n17387 = ( ~n8807 & n15026 ) | ( ~n8807 & n17386 ) | ( n15026 & n17386 ) ;
  assign n17388 = ~n2926 & n3551 ;
  assign n17389 = n4627 & n17388 ;
  assign n17390 = ( ~n1748 & n8380 ) | ( ~n1748 & n17389 ) | ( n8380 & n17389 ) ;
  assign n17391 = n17390 ^ n6689 ^ 1'b0 ;
  assign n17392 = n4500 | n17391 ;
  assign n17394 = n12782 ^ n10692 ^ n5924 ;
  assign n17395 = n3997 & n17394 ;
  assign n17393 = n7864 & ~n12206 ;
  assign n17396 = n17395 ^ n17393 ^ 1'b0 ;
  assign n17397 = n7090 | n13165 ;
  assign n17398 = n2979 | n17397 ;
  assign n17399 = ~n3489 & n9330 ;
  assign n17400 = n17398 & n17399 ;
  assign n17401 = n15987 & n17400 ;
  assign n17402 = n3531 | n6569 ;
  assign n17403 = n1558 & ~n12658 ;
  assign n17404 = n5704 ^ n5363 ^ 1'b0 ;
  assign n17405 = n11345 ^ n5533 ^ n1859 ;
  assign n17406 = ( n10210 & n10297 ) | ( n10210 & ~n17405 ) | ( n10297 & ~n17405 ) ;
  assign n17407 = n9433 ^ n7234 ^ n572 ;
  assign n17408 = ~n12830 & n17407 ;
  assign n17409 = n11711 ^ n9975 ^ 1'b0 ;
  assign n17410 = n17408 | n17409 ;
  assign n17411 = n17406 | n17410 ;
  assign n17412 = n9524 | n9713 ;
  assign n17413 = n12443 & ~n17412 ;
  assign n17414 = n12856 & n17413 ;
  assign n17415 = n14565 & ~n17414 ;
  assign n17416 = n7776 ^ n7387 ^ 1'b0 ;
  assign n17417 = n4234 & n7711 ;
  assign n17418 = n9606 & n17417 ;
  assign n17419 = n8845 ^ n4002 ^ 1'b0 ;
  assign n17420 = ~n1712 & n17419 ;
  assign n17421 = n6564 ^ n4281 ^ 1'b0 ;
  assign n17422 = n3332 & n17421 ;
  assign n17423 = n2140 ^ n261 ^ 1'b0 ;
  assign n17424 = ~n401 & n17423 ;
  assign n17425 = n13086 & n17424 ;
  assign n17426 = n17425 ^ n945 ^ 1'b0 ;
  assign n17427 = n16922 | n17426 ;
  assign n17428 = n17422 | n17427 ;
  assign n17429 = n5809 & n11272 ;
  assign n17430 = n17429 ^ n14616 ^ 1'b0 ;
  assign n17431 = n1241 & n17430 ;
  assign n17432 = n7188 & n17431 ;
  assign n17433 = ~n9183 & n11220 ;
  assign n17434 = ~n3739 & n17433 ;
  assign n17438 = n2385 | n3573 ;
  assign n17439 = n3483 & ~n17438 ;
  assign n17435 = n51 | n8557 ;
  assign n17436 = n17435 ^ n1507 ^ 1'b0 ;
  assign n17437 = ~n5146 & n17436 ;
  assign n17440 = n17439 ^ n17437 ^ 1'b0 ;
  assign n17441 = n436 & ~n10825 ;
  assign n17442 = n15791 ^ n13151 ^ 1'b0 ;
  assign n17443 = ~n17441 & n17442 ;
  assign n17444 = n14690 ^ n14032 ^ 1'b0 ;
  assign n17445 = n17443 & ~n17444 ;
  assign n17446 = n10208 ^ n2441 ^ 1'b0 ;
  assign n17447 = n10333 & ~n17446 ;
  assign n17448 = ~n3409 & n17447 ;
  assign n17449 = ~n17445 & n17448 ;
  assign n17450 = ~n2493 & n6417 ;
  assign n17451 = n6229 & ~n17450 ;
  assign n17454 = n455 | n3475 ;
  assign n17455 = n17454 ^ n7254 ^ 1'b0 ;
  assign n17456 = n3647 ^ n3626 ^ 1'b0 ;
  assign n17457 = n17455 & n17456 ;
  assign n17458 = ~n4656 & n17457 ;
  assign n17459 = n1787 & n17458 ;
  assign n17460 = n12290 | n17459 ;
  assign n17452 = n6646 ^ n481 ^ 1'b0 ;
  assign n17453 = n8647 & n17452 ;
  assign n17461 = n17460 ^ n17453 ^ 1'b0 ;
  assign n17462 = ( n8840 & n12582 ) | ( n8840 & ~n17461 ) | ( n12582 & ~n17461 ) ;
  assign n17463 = n3173 | n5225 ;
  assign n17464 = n93 | n978 ;
  assign n17465 = n498 & ~n17464 ;
  assign n17466 = n17465 ^ n11014 ^ x3 ;
  assign n17467 = n3269 | n4951 ;
  assign n17468 = n2062 & n10594 ;
  assign n17469 = n3079 & ~n15949 ;
  assign n17470 = n10560 ^ n8936 ^ 1'b0 ;
  assign n17471 = n1522 | n17470 ;
  assign n17472 = ( n3803 & n13376 ) | ( n3803 & n17471 ) | ( n13376 & n17471 ) ;
  assign n17477 = n10402 & n14484 ;
  assign n17473 = n4315 | n6205 ;
  assign n17474 = ~n6495 & n9760 ;
  assign n17475 = n17473 & n17474 ;
  assign n17476 = n6817 | n17475 ;
  assign n17478 = n17477 ^ n17476 ^ 1'b0 ;
  assign n17481 = n4454 | n6819 ;
  assign n17482 = n17481 ^ n3406 ^ 1'b0 ;
  assign n17479 = n3201 | n15675 ;
  assign n17480 = n2440 & ~n17479 ;
  assign n17483 = n17482 ^ n17480 ^ 1'b0 ;
  assign n17484 = n17478 | n17483 ;
  assign n17485 = n10572 | n12168 ;
  assign n17486 = n6473 & ~n17485 ;
  assign n17487 = n17486 ^ n9308 ^ n4120 ;
  assign n17488 = ( ~n1214 & n7490 ) | ( ~n1214 & n9929 ) | ( n7490 & n9929 ) ;
  assign n17489 = n1247 & n8608 ;
  assign n17490 = n17489 ^ n1666 ^ 1'b0 ;
  assign n17491 = n12348 & n17490 ;
  assign n17492 = n854 & ~n8960 ;
  assign n17493 = n17492 ^ n9621 ^ 1'b0 ;
  assign n17494 = n4809 ^ n1617 ^ n152 ;
  assign n17495 = n7358 ^ n4570 ^ 1'b0 ;
  assign n17496 = ~n12259 & n17495 ;
  assign n17497 = n3890 & n17496 ;
  assign n17498 = n17497 ^ n10462 ^ 1'b0 ;
  assign n17499 = ~n12728 & n17498 ;
  assign n17500 = ( n4880 & n17494 ) | ( n4880 & n17499 ) | ( n17494 & n17499 ) ;
  assign n17501 = ( n364 & ~n556 ) | ( n364 & n884 ) | ( ~n556 & n884 ) ;
  assign n17502 = n12402 & ~n17501 ;
  assign n17503 = n9987 ^ n4675 ^ 1'b0 ;
  assign n17504 = n1181 & ~n17282 ;
  assign n17505 = n17504 ^ n15375 ^ n5678 ;
  assign n17507 = ( n1386 & ~n7989 ) | ( n1386 & n9460 ) | ( ~n7989 & n9460 ) ;
  assign n17506 = n3201 | n15739 ;
  assign n17508 = n17507 ^ n17506 ^ 1'b0 ;
  assign n17509 = n13078 ^ n2789 ^ 1'b0 ;
  assign n17510 = n13202 & ~n17509 ;
  assign n17511 = n17510 ^ n13279 ^ 1'b0 ;
  assign n17512 = n1189 & ~n12168 ;
  assign n17513 = n255 & n17512 ;
  assign n17514 = n9962 ^ n3647 ^ 1'b0 ;
  assign n17515 = n727 & n2266 ;
  assign n17516 = n4688 & n17515 ;
  assign n17517 = n14016 ^ n1192 ^ 1'b0 ;
  assign n17518 = n7237 | n17517 ;
  assign n17520 = n4461 ^ n1982 ^ 1'b0 ;
  assign n17519 = ~n744 & n14892 ;
  assign n17521 = n17520 ^ n17519 ^ 1'b0 ;
  assign n17522 = n17521 ^ n9981 ^ 1'b0 ;
  assign n17523 = ~n17518 & n17522 ;
  assign n17524 = n5683 & ~n17180 ;
  assign n17525 = ~n1182 & n7443 ;
  assign n17526 = n7489 & n17525 ;
  assign n17534 = n1848 ^ n332 ^ 1'b0 ;
  assign n17535 = n17534 ^ n15213 ^ n8113 ;
  assign n17527 = n8537 ^ n6275 ^ 1'b0 ;
  assign n17528 = ~n1135 & n17527 ;
  assign n17529 = n3593 | n3793 ;
  assign n17530 = n17528 | n17529 ;
  assign n17531 = ( n2879 & n13505 ) | ( n2879 & n17530 ) | ( n13505 & n17530 ) ;
  assign n17532 = n16017 ^ n10465 ^ n4287 ;
  assign n17533 = n17531 & n17532 ;
  assign n17536 = n17535 ^ n17533 ^ 1'b0 ;
  assign n17537 = n6049 ^ n4657 ^ 1'b0 ;
  assign n17538 = n4897 & ~n17537 ;
  assign n17539 = n7020 & n17538 ;
  assign n17540 = n1569 | n16753 ;
  assign n17541 = n17540 ^ n9138 ^ 1'b0 ;
  assign n17542 = n57 & n1933 ;
  assign n17543 = n12799 & ~n17542 ;
  assign n17544 = ( n1946 & n10176 ) | ( n1946 & n17543 ) | ( n10176 & n17543 ) ;
  assign n17545 = n16220 ^ n2836 ^ 1'b0 ;
  assign n17546 = n5131 | n17545 ;
  assign n17547 = ~n320 & n9105 ;
  assign n17548 = n17547 ^ n16457 ^ 1'b0 ;
  assign n17549 = n10091 | n14956 ;
  assign n17550 = n17549 ^ n2706 ^ 1'b0 ;
  assign n17551 = n14409 ^ n7545 ^ 1'b0 ;
  assign n17552 = n4260 & n4785 ;
  assign n17555 = n8712 ^ n8485 ^ 1'b0 ;
  assign n17556 = n8215 & ~n17555 ;
  assign n17557 = ~n369 & n17556 ;
  assign n17558 = n17557 ^ n4657 ^ 1'b0 ;
  assign n17553 = n471 | n2735 ;
  assign n17554 = n180 | n17553 ;
  assign n17559 = n17558 ^ n17554 ^ 1'b0 ;
  assign n17560 = n11320 & ~n17559 ;
  assign n17561 = n5987 & n17514 ;
  assign n17562 = n1305 & ~n5860 ;
  assign n17563 = n9866 & n17562 ;
  assign n17564 = n17563 ^ n14238 ^ n11560 ;
  assign n17565 = n448 & n14158 ;
  assign n17566 = n1443 & n3916 ;
  assign n17567 = n17566 ^ n8878 ^ 1'b0 ;
  assign n17568 = n7113 & n17567 ;
  assign n17569 = ~n14145 & n17568 ;
  assign n17570 = n12010 ^ n5800 ^ 1'b0 ;
  assign n17571 = ~n12283 & n17570 ;
  assign n17572 = n17571 ^ n11366 ^ 1'b0 ;
  assign n17573 = n13524 ^ n5380 ^ 1'b0 ;
  assign n17574 = n4903 & n17573 ;
  assign n17575 = n3115 & ~n3751 ;
  assign n17576 = n1410 & n17575 ;
  assign n17577 = n7401 & ~n17576 ;
  assign n17578 = n17577 ^ n1793 ^ 1'b0 ;
  assign n17579 = n4427 | n11510 ;
  assign n17580 = n17579 ^ n15672 ^ n10523 ;
  assign n17581 = n4180 ^ n876 ^ 1'b0 ;
  assign n17582 = ~n11249 & n17581 ;
  assign n17583 = ~n12684 & n17582 ;
  assign n17584 = n6067 ^ n3805 ^ 1'b0 ;
  assign n17585 = n14628 | n17584 ;
  assign n17586 = n15192 & n16738 ;
  assign n17587 = ( n369 & n1105 ) | ( n369 & n17586 ) | ( n1105 & n17586 ) ;
  assign n17588 = n3329 & n11901 ;
  assign n17589 = n15555 & n17588 ;
  assign n17591 = n2126 & ~n3238 ;
  assign n17592 = n7643 & n17591 ;
  assign n17590 = n5858 | n13143 ;
  assign n17593 = n17592 ^ n17590 ^ 1'b0 ;
  assign n17594 = ~n17589 & n17593 ;
  assign n17595 = n42 & n11898 ;
  assign n17605 = ~n1450 & n2441 ;
  assign n17596 = n4629 & ~n5855 ;
  assign n17597 = n17596 ^ n8854 ^ 1'b0 ;
  assign n17602 = n12290 ^ n5658 ^ 1'b0 ;
  assign n17598 = n16155 ^ n3953 ^ 1'b0 ;
  assign n17599 = n3991 & n17598 ;
  assign n17600 = ~n1243 & n17599 ;
  assign n17601 = n17600 ^ n6481 ^ 1'b0 ;
  assign n17603 = n17602 ^ n17601 ^ 1'b0 ;
  assign n17604 = ~n17597 & n17603 ;
  assign n17606 = n17605 ^ n17604 ^ 1'b0 ;
  assign n17607 = n17595 | n17606 ;
  assign n17608 = n11536 ^ n11185 ^ n157 ;
  assign n17609 = n11593 & n12857 ;
  assign n17610 = n17608 & n17609 ;
  assign n17611 = n131 | n7421 ;
  assign n17612 = n17611 ^ n9860 ^ 1'b0 ;
  assign n17613 = n17612 ^ n10245 ^ n8775 ;
  assign n17614 = n16738 ^ n3109 ^ n1105 ;
  assign n17615 = n2859 & ~n17614 ;
  assign n17616 = n17615 ^ n431 ^ 1'b0 ;
  assign n17617 = n17616 ^ n803 ^ 1'b0 ;
  assign n17620 = ~n852 & n2217 ;
  assign n17621 = n17620 ^ n4653 ^ 1'b0 ;
  assign n17618 = n8941 & n10887 ;
  assign n17619 = n17618 ^ n9404 ^ 1'b0 ;
  assign n17622 = n17621 ^ n17619 ^ 1'b0 ;
  assign n17623 = n5382 | n15624 ;
  assign n17624 = n8321 | n8678 ;
  assign n17625 = n14075 | n17624 ;
  assign n17626 = n17293 | n17625 ;
  assign n17627 = n17626 ^ n17110 ^ n10835 ;
  assign n17628 = n185 & n2481 ;
  assign n17629 = ( n4704 & ~n5535 ) | ( n4704 & n13576 ) | ( ~n5535 & n13576 ) ;
  assign n17630 = n5630 | n17629 ;
  assign n17631 = ~n2526 & n17630 ;
  assign n17632 = n17631 ^ n9126 ^ 1'b0 ;
  assign n17633 = n2056 & n7395 ;
  assign n17634 = n1463 | n15718 ;
  assign n17635 = n14286 & n15122 ;
  assign n17639 = n2951 ^ n259 ^ 1'b0 ;
  assign n17640 = n43 | n17639 ;
  assign n17636 = ~n4222 & n6785 ;
  assign n17637 = n1982 & n17636 ;
  assign n17638 = n17637 ^ n13539 ^ n12704 ;
  assign n17641 = n17640 ^ n17638 ^ n9315 ;
  assign n17642 = ~n1660 & n3064 ;
  assign n17643 = n17642 ^ n2242 ^ 1'b0 ;
  assign n17644 = ( n17238 & n17641 ) | ( n17238 & ~n17643 ) | ( n17641 & ~n17643 ) ;
  assign n17645 = n17034 ^ n12411 ^ 1'b0 ;
  assign n17646 = n17222 ^ n10323 ^ 1'b0 ;
  assign n17647 = n2531 & n4695 ;
  assign n17648 = n15495 & n17647 ;
  assign n17649 = ~n13684 & n15830 ;
  assign n17650 = ~n1655 & n2763 ;
  assign n17651 = n17650 ^ n10690 ^ 1'b0 ;
  assign n17652 = n108 & ~n17651 ;
  assign n17653 = n17418 | n17652 ;
  assign n17654 = n119 & n9493 ;
  assign n17655 = ~n351 & n17654 ;
  assign n17656 = ~n3290 & n11632 ;
  assign n17657 = ~n5329 & n6640 ;
  assign n17658 = n17657 ^ n7873 ^ 1'b0 ;
  assign n17659 = n7598 & ~n17658 ;
  assign n17660 = ~n1952 & n4620 ;
  assign n17661 = n17660 ^ n6593 ^ 1'b0 ;
  assign n17662 = ~n72 & n8549 ;
  assign n17663 = n1324 & n17662 ;
  assign n17664 = ( n17659 & ~n17661 ) | ( n17659 & n17663 ) | ( ~n17661 & n17663 ) ;
  assign n17665 = n4799 | n13291 ;
  assign n17666 = n4653 & n4671 ;
  assign n17667 = n17666 ^ n11283 ^ 1'b0 ;
  assign n17668 = n15690 ^ n9625 ^ 1'b0 ;
  assign n17669 = n14102 & ~n17668 ;
  assign n17670 = n2044 | n10436 ;
  assign n17671 = n17669 | n17670 ;
  assign n17672 = n17671 ^ n7541 ^ 1'b0 ;
  assign n17673 = n17667 | n17672 ;
  assign n17674 = n962 | n6088 ;
  assign n17675 = ~n1589 & n15282 ;
  assign n17676 = n17675 ^ n15266 ^ n14476 ;
  assign n17677 = n8443 & ~n9917 ;
  assign n17678 = n2485 & n17677 ;
  assign n17679 = n17678 ^ n5286 ^ 1'b0 ;
  assign n17681 = n3753 ^ n953 ^ 1'b0 ;
  assign n17680 = n17325 ^ n15191 ^ 1'b0 ;
  assign n17682 = n17681 ^ n17680 ^ 1'b0 ;
  assign n17683 = n1521 & n17313 ;
  assign n17684 = n5350 & n12742 ;
  assign n17685 = ~n17683 & n17684 ;
  assign n17686 = n14606 ^ n7186 ^ 1'b0 ;
  assign n17687 = ~n10436 & n17686 ;
  assign n17688 = n13157 & ~n15267 ;
  assign n17689 = ~n8152 & n17688 ;
  assign n17690 = ( n711 & ~n17687 ) | ( n711 & n17689 ) | ( ~n17687 & n17689 ) ;
  assign n17691 = n3214 | n16705 ;
  assign n17692 = n17691 ^ n12973 ^ 1'b0 ;
  assign n17693 = ( ~n887 & n1357 ) | ( ~n887 & n3407 ) | ( n1357 & n3407 ) ;
  assign n17694 = n7678 | n17693 ;
  assign n17695 = ~n16804 & n17694 ;
  assign n17696 = n17692 & n17695 ;
  assign n17697 = n17386 | n17696 ;
  assign n17698 = n17697 ^ n15661 ^ 1'b0 ;
  assign n17699 = n2984 | n4376 ;
  assign n17700 = n17699 ^ n3844 ^ 1'b0 ;
  assign n17701 = n10260 ^ n9904 ^ 1'b0 ;
  assign n17702 = n14580 & n17701 ;
  assign n17703 = n17012 ^ n12096 ^ 1'b0 ;
  assign n17704 = n17702 & ~n17703 ;
  assign n17705 = n17603 ^ n2734 ^ 1'b0 ;
  assign n17706 = n14360 & ~n17705 ;
  assign n17707 = n7278 | n16901 ;
  assign n17708 = n17707 ^ n14030 ^ 1'b0 ;
  assign n17709 = n12131 ^ n3435 ^ 1'b0 ;
  assign n17710 = n17709 ^ n5102 ^ 1'b0 ;
  assign n17711 = ~n4834 & n11516 ;
  assign n17712 = n17711 ^ n3773 ^ 1'b0 ;
  assign n17713 = n17712 ^ n8079 ^ 1'b0 ;
  assign n17714 = n17710 & ~n17713 ;
  assign n17715 = n8938 ^ n7141 ^ 1'b0 ;
  assign n17716 = n1122 & n17715 ;
  assign n17717 = n17716 ^ n7284 ^ 1'b0 ;
  assign n17718 = ( n7173 & ~n10098 ) | ( n7173 & n15191 ) | ( ~n10098 & n15191 ) ;
  assign n17719 = n12803 ^ n8115 ^ 1'b0 ;
  assign n17720 = n17718 & n17719 ;
  assign n17721 = ( ~n384 & n5892 ) | ( ~n384 & n6924 ) | ( n5892 & n6924 ) ;
  assign n17722 = ( n2381 & n8683 ) | ( n2381 & ~n17721 ) | ( n8683 & ~n17721 ) ;
  assign n17723 = n1573 | n3581 ;
  assign n17724 = n12490 | n17723 ;
  assign n17725 = n5253 ^ n3842 ^ 1'b0 ;
  assign n17726 = n2471 | n2645 ;
  assign n17727 = n17726 ^ n648 ^ 1'b0 ;
  assign n17728 = n17725 & n17727 ;
  assign n17729 = ~n1672 & n17728 ;
  assign n17730 = n14903 ^ n9147 ^ 1'b0 ;
  assign n17731 = n9011 | n17730 ;
  assign n17732 = n17731 ^ n4278 ^ 1'b0 ;
  assign n17733 = n5845 ^ n648 ^ 1'b0 ;
  assign n17734 = n2098 & n17733 ;
  assign n17735 = n17424 ^ n5817 ^ 1'b0 ;
  assign n17736 = n17734 & n17735 ;
  assign n17737 = n17736 ^ n4156 ^ 1'b0 ;
  assign n17738 = ~n17732 & n17737 ;
  assign n17739 = n15643 ^ n5961 ^ 1'b0 ;
  assign n17740 = n169 & ~n16197 ;
  assign n17741 = n17740 ^ n1740 ^ 1'b0 ;
  assign n17743 = n10256 ^ n2760 ^ 1'b0 ;
  assign n17742 = n6229 ^ n865 ^ 1'b0 ;
  assign n17744 = n17743 ^ n17742 ^ n4071 ;
  assign n17751 = n10511 ^ n8249 ^ 1'b0 ;
  assign n17745 = n12445 ^ n6774 ^ 1'b0 ;
  assign n17746 = n2705 & ~n17745 ;
  assign n17747 = n962 & ~n17746 ;
  assign n17748 = n14213 ^ n10849 ^ 1'b0 ;
  assign n17749 = n17748 ^ n4118 ^ n2625 ;
  assign n17750 = n17747 | n17749 ;
  assign n17752 = n17751 ^ n17750 ^ 1'b0 ;
  assign n17754 = n139 & n6437 ;
  assign n17753 = n41 & ~n12091 ;
  assign n17755 = n17754 ^ n17753 ^ n33 ;
  assign n17756 = n17755 ^ n15383 ^ n32 ;
  assign n17757 = ~n6188 & n6743 ;
  assign n17758 = n191 & n17757 ;
  assign n17759 = n17758 ^ n11253 ^ 1'b0 ;
  assign n17760 = n12642 & n17759 ;
  assign n17761 = n6197 & ~n10380 ;
  assign n17762 = ~n8681 & n17761 ;
  assign n17763 = ( n8198 & ~n17760 ) | ( n8198 & n17762 ) | ( ~n17760 & n17762 ) ;
  assign n17764 = n1767 & ~n3647 ;
  assign n17765 = n17764 ^ n2144 ^ 1'b0 ;
  assign n17766 = ( n1612 & n4340 ) | ( n1612 & ~n5042 ) | ( n4340 & ~n5042 ) ;
  assign n17767 = n17766 ^ n14413 ^ 1'b0 ;
  assign n17768 = n150 & ~n2695 ;
  assign n17769 = ( n795 & ~n6274 ) | ( n795 & n12799 ) | ( ~n6274 & n12799 ) ;
  assign n17770 = n691 | n16709 ;
  assign n17771 = ~n41 & n3412 ;
  assign n17772 = n17771 ^ n4987 ^ n3740 ;
  assign n17773 = n2670 & n17772 ;
  assign n17774 = n1783 & n17773 ;
  assign n17775 = n17774 ^ n11730 ^ 1'b0 ;
  assign n17776 = n15111 & ~n17775 ;
  assign n17777 = n530 & ~n10153 ;
  assign n17778 = n17777 ^ n15708 ^ 1'b0 ;
  assign n17779 = n601 | n11271 ;
  assign n17780 = n2745 & ~n17779 ;
  assign n17781 = n17780 ^ n13903 ^ 1'b0 ;
  assign n17782 = n17781 ^ n11907 ^ n4562 ;
  assign n17783 = n5979 ^ n5264 ^ 1'b0 ;
  assign n17789 = n2551 & n4356 ;
  assign n17787 = n3663 & n5587 ;
  assign n17784 = ~n2160 & n4765 ;
  assign n17785 = n3581 & ~n11222 ;
  assign n17786 = ~n17784 & n17785 ;
  assign n17788 = n17787 ^ n17786 ^ 1'b0 ;
  assign n17790 = n17789 ^ n17788 ^ 1'b0 ;
  assign n17791 = n1746 & ~n17790 ;
  assign n17792 = n2261 & ~n15702 ;
  assign n17793 = n1751 | n4544 ;
  assign n17794 = n1502 | n17793 ;
  assign n17795 = n17792 | n17794 ;
  assign n17796 = n17795 ^ n12965 ^ 1'b0 ;
  assign n17797 = ~n4773 & n17796 ;
  assign n17798 = ~n567 & n4543 ;
  assign n17800 = n2078 | n2259 ;
  assign n17801 = ( n4941 & n7927 ) | ( n4941 & ~n17800 ) | ( n7927 & ~n17800 ) ;
  assign n17799 = n13939 ^ n838 ^ 1'b0 ;
  assign n17802 = n17801 ^ n17799 ^ 1'b0 ;
  assign n17803 = n10333 ^ n2302 ^ 1'b0 ;
  assign n17804 = n12184 ^ n3257 ^ n1932 ;
  assign n17805 = n17804 ^ n601 ^ 1'b0 ;
  assign n17806 = n17805 ^ n7069 ^ 1'b0 ;
  assign n17807 = ~n17803 & n17806 ;
  assign n17808 = n5535 ^ n5011 ^ 1'b0 ;
  assign n17809 = n14041 & ~n17808 ;
  assign n17810 = n7957 | n9435 ;
  assign n17811 = n17809 | n17810 ;
  assign n17812 = n11387 ^ n6614 ^ 1'b0 ;
  assign n17813 = n7481 ^ n1934 ^ n57 ;
  assign n17814 = ( n7574 & n16709 ) | ( n7574 & n17813 ) | ( n16709 & n17813 ) ;
  assign n17815 = n4197 & ~n13725 ;
  assign n17816 = n1029 & n5006 ;
  assign n17817 = n10812 & n17816 ;
  assign n17822 = n17164 ^ n2177 ^ 1'b0 ;
  assign n17818 = n2044 & n13676 ;
  assign n17819 = ~n1412 & n17818 ;
  assign n17820 = n6711 & n17819 ;
  assign n17821 = ( n216 & ~n11507 ) | ( n216 & n17820 ) | ( ~n11507 & n17820 ) ;
  assign n17823 = n17822 ^ n17821 ^ 1'b0 ;
  assign n17824 = n17817 | n17823 ;
  assign n17825 = n17815 & n17824 ;
  assign n17826 = n9345 & n17825 ;
  assign n17827 = x10 & n17826 ;
  assign n17828 = n2399 & n6579 ;
  assign n17829 = n10145 ^ n6230 ^ 1'b0 ;
  assign n17830 = ~n17828 & n17829 ;
  assign n17831 = n2960 ^ n1348 ^ 1'b0 ;
  assign n17832 = n17831 ^ n2622 ^ 1'b0 ;
  assign n17833 = ( n889 & n5392 ) | ( n889 & ~n11585 ) | ( n5392 & ~n11585 ) ;
  assign n17834 = ~n10939 & n14703 ;
  assign n17835 = n5285 & ~n9240 ;
  assign n17836 = n17249 ^ n12842 ^ n10868 ;
  assign n17837 = n6829 | n17836 ;
  assign n17838 = ~n5843 & n6477 ;
  assign n17839 = ~n355 & n17838 ;
  assign n17842 = n15254 ^ n14781 ^ n72 ;
  assign n17840 = n8964 ^ n7650 ^ n36 ;
  assign n17841 = n17840 ^ n14366 ^ n3953 ;
  assign n17843 = n17842 ^ n17841 ^ 1'b0 ;
  assign n17844 = n12221 ^ n9769 ^ n5604 ;
  assign n17845 = n9848 ^ n4012 ^ 1'b0 ;
  assign n17846 = n322 & ~n2322 ;
  assign n17847 = n10543 ^ n9210 ^ 1'b0 ;
  assign n17848 = n11103 & ~n17847 ;
  assign n17854 = n15824 ^ n2213 ^ 1'b0 ;
  assign n17853 = ~n6394 & n7374 ;
  assign n17855 = n17854 ^ n17853 ^ 1'b0 ;
  assign n17849 = n850 & n8625 ;
  assign n17850 = n259 & n17849 ;
  assign n17851 = n17850 ^ n8624 ^ n276 ;
  assign n17852 = n6698 & n17851 ;
  assign n17856 = n17855 ^ n17852 ^ n8371 ;
  assign n17857 = ~n6670 & n17856 ;
  assign n17858 = n7540 & n12517 ;
  assign n17859 = n8054 & n17858 ;
  assign n17860 = n1400 & n6623 ;
  assign n17861 = n8453 | n17860 ;
  assign n17862 = n17861 ^ n1894 ^ 1'b0 ;
  assign n17863 = ~n7081 & n11004 ;
  assign n17864 = n6766 & n17863 ;
  assign n17865 = n9032 ^ n5878 ^ 1'b0 ;
  assign n17866 = n7844 ^ n7279 ^ 1'b0 ;
  assign n17867 = n1078 | n2107 ;
  assign n17868 = n17866 & ~n17867 ;
  assign n17869 = n13221 ^ n6978 ^ n2635 ;
  assign n17870 = ~n448 & n2144 ;
  assign n17871 = n17869 & ~n17870 ;
  assign n17872 = n11119 & n17871 ;
  assign n17873 = ( n3473 & n4045 ) | ( n3473 & n17872 ) | ( n4045 & n17872 ) ;
  assign n17874 = ~n10255 & n10279 ;
  assign n17875 = n17874 ^ n12185 ^ 1'b0 ;
  assign n17876 = ~n6738 & n14004 ;
  assign n17877 = n11204 ^ n421 ^ 1'b0 ;
  assign n17878 = n3203 & n17877 ;
  assign n17879 = n6599 & ~n6787 ;
  assign n17880 = n7230 & n17879 ;
  assign n17881 = n17878 | n17880 ;
  assign n17882 = n13583 & n17881 ;
  assign n17883 = ~n17876 & n17882 ;
  assign n17884 = n7788 ^ n4977 ^ n784 ;
  assign n17885 = n16489 & n17884 ;
  assign n17886 = n17885 ^ n5363 ^ 1'b0 ;
  assign n17887 = n249 & ~n1039 ;
  assign n17888 = n17887 ^ n2667 ^ 1'b0 ;
  assign n17889 = n17888 ^ n4787 ^ n183 ;
  assign n17890 = n2130 & n17889 ;
  assign n17891 = n17890 ^ n8337 ^ n63 ;
  assign n17892 = n315 | n3812 ;
  assign n17893 = n7977 & ~n17892 ;
  assign n17894 = n17893 ^ n839 ^ n423 ;
  assign n17895 = n3019 ^ n2864 ^ 1'b0 ;
  assign n17896 = ~n10311 & n17895 ;
  assign n17897 = ~n17894 & n17896 ;
  assign n17898 = n619 & n13585 ;
  assign n17899 = n16158 ^ n10093 ^ 1'b0 ;
  assign n17900 = n2895 & ~n8269 ;
  assign n17901 = ( n3962 & n5396 ) | ( n3962 & n17900 ) | ( n5396 & n17900 ) ;
  assign n17902 = n202 & ~n9522 ;
  assign n17903 = n17902 ^ n8745 ^ 1'b0 ;
  assign n17904 = n5280 & ~n14292 ;
  assign n17905 = n1554 ^ n582 ^ 1'b0 ;
  assign n17906 = n1249 & n17905 ;
  assign n17907 = n16611 ^ n9462 ^ 1'b0 ;
  assign n17908 = n8420 ^ n5507 ^ 1'b0 ;
  assign n17909 = n10520 | n17908 ;
  assign n17910 = n17909 ^ n11064 ^ 1'b0 ;
  assign n17911 = n16153 ^ n3673 ^ 1'b0 ;
  assign n17912 = n1131 & ~n17911 ;
  assign n17913 = n1927 & n6546 ;
  assign n17914 = n1898 | n9411 ;
  assign n17915 = n17913 & ~n17914 ;
  assign n17916 = n17915 ^ n15043 ^ n14555 ;
  assign n17917 = n6076 | n17128 ;
  assign n17919 = n5930 ^ n4769 ^ n3177 ;
  assign n17920 = ~n2190 & n12519 ;
  assign n17921 = n17920 ^ n6813 ^ 1'b0 ;
  assign n17922 = n17919 | n17921 ;
  assign n17918 = ~n1851 & n7205 ;
  assign n17923 = n17922 ^ n17918 ^ 1'b0 ;
  assign n17924 = n5484 ^ n3644 ^ 1'b0 ;
  assign n17925 = ~n2177 & n17924 ;
  assign n17926 = n1364 & ~n6351 ;
  assign n17927 = ~n17925 & n17926 ;
  assign n17928 = n15197 ^ n11593 ^ 1'b0 ;
  assign n17929 = ( n4974 & n17402 ) | ( n4974 & ~n17405 ) | ( n17402 & ~n17405 ) ;
  assign n17930 = n3898 ^ n3461 ^ 1'b0 ;
  assign n17931 = n7398 ^ n326 ^ 1'b0 ;
  assign n17932 = n7542 & n17931 ;
  assign n17933 = n4115 | n17932 ;
  assign n17934 = ( n162 & n3062 ) | ( n162 & ~n4574 ) | ( n3062 & ~n4574 ) ;
  assign n17935 = n17934 ^ n16940 ^ n1600 ;
  assign n17936 = n17935 ^ n17388 ^ n3370 ;
  assign n17937 = n17936 ^ n12503 ^ 1'b0 ;
  assign n17938 = n17933 & n17937 ;
  assign n17939 = n6477 ^ n825 ^ 1'b0 ;
  assign n17941 = n4019 & n5679 ;
  assign n17942 = n17941 ^ n5227 ^ 1'b0 ;
  assign n17940 = ( ~n2733 & n3546 ) | ( ~n2733 & n6793 ) | ( n3546 & n6793 ) ;
  assign n17943 = n17942 ^ n17940 ^ 1'b0 ;
  assign n17944 = n3019 & n17943 ;
  assign n17945 = n17939 & n17944 ;
  assign n17946 = n7378 ^ n6217 ^ 1'b0 ;
  assign n17947 = n7076 | n17592 ;
  assign n17948 = n2316 & n5131 ;
  assign n17949 = n4486 ^ n1868 ^ 1'b0 ;
  assign n17950 = n3064 ^ n211 ^ 1'b0 ;
  assign n17951 = n1709 ^ n1110 ^ 1'b0 ;
  assign n17952 = n2246 & n17951 ;
  assign n17953 = n15114 ^ n11218 ^ 1'b0 ;
  assign n17954 = n13975 & n17953 ;
  assign n17955 = n17954 ^ n4383 ^ 1'b0 ;
  assign n17956 = n17952 | n17955 ;
  assign n17957 = ( n1578 & n3755 ) | ( n1578 & n12260 ) | ( n3755 & n12260 ) ;
  assign n17958 = ~n17956 & n17957 ;
  assign n17959 = n17958 ^ n7147 ^ 1'b0 ;
  assign n17960 = n109 & ~n6789 ;
  assign n17961 = n17960 ^ n6293 ^ 1'b0 ;
  assign n17962 = ~n3788 & n17961 ;
  assign n17963 = ~n3414 & n17962 ;
  assign n17964 = n5630 ^ n108 ^ 1'b0 ;
  assign n17965 = ( n9085 & n16412 ) | ( n9085 & n17964 ) | ( n16412 & n17964 ) ;
  assign n17975 = n201 & n6717 ;
  assign n17976 = ~n3888 & n17975 ;
  assign n17972 = n3043 | n5895 ;
  assign n17973 = n17972 ^ n4153 ^ 1'b0 ;
  assign n17974 = n17973 ^ n1131 ^ 1'b0 ;
  assign n17969 = n4914 ^ n4671 ^ 1'b0 ;
  assign n17966 = n5912 ^ n1107 ^ 1'b0 ;
  assign n17967 = ~n7034 & n17966 ;
  assign n17968 = ~n2732 & n17967 ;
  assign n17970 = n17969 ^ n17968 ^ 1'b0 ;
  assign n17971 = n4419 | n17970 ;
  assign n17977 = n17976 ^ n17974 ^ n17971 ;
  assign n17978 = ~n2986 & n4112 ;
  assign n17979 = n17978 ^ n16804 ^ 1'b0 ;
  assign n17980 = ~n2824 & n5507 ;
  assign n17981 = n6983 & n10277 ;
  assign n17982 = n9702 ^ n853 ^ 1'b0 ;
  assign n17983 = n17982 ^ n5895 ^ n1363 ;
  assign n17984 = n8279 & ~n12638 ;
  assign n17985 = ~n11935 & n17984 ;
  assign n17986 = ~n9500 & n10786 ;
  assign n17987 = ~n7661 & n17986 ;
  assign n17988 = n7363 & n17987 ;
  assign n17989 = n17988 ^ n11437 ^ 1'b0 ;
  assign n17990 = ~n8467 & n11120 ;
  assign n17991 = n7767 ^ n4317 ^ 1'b0 ;
  assign n17992 = n12247 & n17991 ;
  assign n17993 = n9939 & n17992 ;
  assign n17994 = n15402 & ~n17993 ;
  assign n17995 = ~n11175 & n17994 ;
  assign n17996 = ( n7231 & n16605 ) | ( n7231 & n17939 ) | ( n16605 & n17939 ) ;
  assign n17997 = n6116 & n16973 ;
  assign n17998 = ~n10795 & n16876 ;
  assign n17999 = n5958 & n10120 ;
  assign n18000 = n17999 ^ n5090 ^ n4863 ;
  assign n18001 = n8820 | n15627 ;
  assign n18002 = ~n6122 & n13023 ;
  assign n18003 = n4862 & ~n18002 ;
  assign n18004 = n6304 ^ n293 ^ 1'b0 ;
  assign n18005 = n18003 & ~n18004 ;
  assign n18006 = ~n5111 & n9493 ;
  assign n18007 = n1033 | n1681 ;
  assign n18008 = n18007 ^ n5495 ^ 1'b0 ;
  assign n18009 = n1596 & ~n18008 ;
  assign n18010 = n18009 ^ n15827 ^ 1'b0 ;
  assign n18011 = n10899 | n18010 ;
  assign n18012 = n18011 ^ n12421 ^ 1'b0 ;
  assign n18013 = n15714 ^ n7620 ^ n1346 ;
  assign n18014 = n480 | n18013 ;
  assign n18015 = n7128 & n17842 ;
  assign n18016 = n4622 & n15248 ;
  assign n18017 = n18016 ^ n241 ^ 1'b0 ;
  assign n18019 = ( n6304 & ~n11791 ) | ( n6304 & n14354 ) | ( ~n11791 & n14354 ) ;
  assign n18020 = n1822 & n18019 ;
  assign n18021 = ~n9009 & n18020 ;
  assign n18018 = ( n601 & ~n8174 ) | ( n601 & n10066 ) | ( ~n8174 & n10066 ) ;
  assign n18022 = n18021 ^ n18018 ^ 1'b0 ;
  assign n18023 = n18022 ^ n9147 ^ 1'b0 ;
  assign n18024 = n11154 ^ n8585 ^ n3590 ;
  assign n18025 = n5803 & n18024 ;
  assign n18026 = n12510 & n15976 ;
  assign n18027 = n937 & n18026 ;
  assign n18028 = n12787 ^ n11041 ^ 1'b0 ;
  assign n18029 = ~n10917 & n18028 ;
  assign n18030 = n744 & n15317 ;
  assign n18031 = n2118 ^ n2072 ^ 1'b0 ;
  assign n18032 = n8874 & n14375 ;
  assign n18033 = n18031 & n18032 ;
  assign n18034 = n874 & n6554 ;
  assign n18043 = n4373 | n5193 ;
  assign n18044 = n18043 ^ n12771 ^ 1'b0 ;
  assign n18045 = n6924 & n18044 ;
  assign n18046 = n5100 & n18045 ;
  assign n18035 = n12003 ^ n2179 ^ 1'b0 ;
  assign n18036 = n14706 & ~n18035 ;
  assign n18037 = n536 & n863 ;
  assign n18038 = n315 & n18037 ;
  assign n18039 = ~n619 & n7680 ;
  assign n18040 = n18038 | n18039 ;
  assign n18041 = n12020 | n18040 ;
  assign n18042 = n18036 & n18041 ;
  assign n18047 = n18046 ^ n18042 ^ 1'b0 ;
  assign n18048 = n4911 & ~n9276 ;
  assign n18049 = n10210 ^ n991 ^ 1'b0 ;
  assign n18050 = n18048 | n18049 ;
  assign n18051 = n13228 | n18050 ;
  assign n18052 = n6036 & n9393 ;
  assign n18053 = n13387 | n18052 ;
  assign n18054 = n8109 ^ n4508 ^ 1'b0 ;
  assign n18055 = n10277 & ~n17039 ;
  assign n18056 = n18055 ^ n13873 ^ 1'b0 ;
  assign n18057 = ~n18054 & n18056 ;
  assign n18058 = n15058 ^ n8301 ^ 1'b0 ;
  assign n18059 = n2313 & n18058 ;
  assign n18060 = n11708 ^ n10841 ^ 1'b0 ;
  assign n18061 = n5675 ^ n222 ^ 1'b0 ;
  assign n18062 = n9729 ^ n9420 ^ 1'b0 ;
  assign n18063 = n13979 ^ n11829 ^ 1'b0 ;
  assign n18064 = ~n4097 & n15140 ;
  assign n18065 = ~n811 & n18064 ;
  assign n18066 = n8141 ^ n5628 ^ n5329 ;
  assign n18067 = n718 ^ n649 ^ 1'b0 ;
  assign n18068 = n18067 ^ n6885 ^ 1'b0 ;
  assign n18069 = n8337 & ~n18068 ;
  assign n18070 = n14816 ^ n4645 ^ 1'b0 ;
  assign n18071 = n9286 & n18070 ;
  assign n18072 = n18071 ^ n11519 ^ 1'b0 ;
  assign n18073 = n1001 & n13433 ;
  assign n18075 = n2334 ^ n696 ^ 1'b0 ;
  assign n18074 = n4367 ^ n2642 ^ n1295 ;
  assign n18076 = n18075 ^ n18074 ^ 1'b0 ;
  assign n18077 = ( ~n614 & n9792 ) | ( ~n614 & n18076 ) | ( n9792 & n18076 ) ;
  assign n18078 = ~n3057 & n8199 ;
  assign n18079 = ~n18077 & n18078 ;
  assign n18080 = n3732 & ~n16691 ;
  assign n18081 = n18080 ^ n15114 ^ 1'b0 ;
  assign n18082 = ~n10057 & n18081 ;
  assign n18083 = n9644 | n18082 ;
  assign n18084 = n3819 | n18083 ;
  assign n18085 = n10767 & n11258 ;
  assign n18086 = n10714 ^ n5713 ^ 1'b0 ;
  assign n18087 = n18085 | n18086 ;
  assign n18088 = n13112 ^ n11976 ^ 1'b0 ;
  assign n18089 = ~n18087 & n18088 ;
  assign n18090 = n8067 & ~n18089 ;
  assign n18091 = n14815 ^ n9210 ^ 1'b0 ;
  assign n18092 = n14352 & n18091 ;
  assign n18093 = n711 | n6739 ;
  assign n18094 = n6924 & n17530 ;
  assign n18095 = n18094 ^ n7406 ^ 1'b0 ;
  assign n18096 = n7006 ^ n3225 ^ 1'b0 ;
  assign n18097 = n17449 ^ n13478 ^ n3184 ;
  assign n18098 = n3641 & ~n12707 ;
  assign n18101 = ( n7123 & n8327 ) | ( n7123 & ~n9686 ) | ( n8327 & ~n9686 ) ;
  assign n18099 = ~n409 & n12720 ;
  assign n18100 = n3686 | n18099 ;
  assign n18102 = n18101 ^ n18100 ^ 1'b0 ;
  assign n18103 = n641 | n15412 ;
  assign n18104 = n17945 | n18103 ;
  assign n18108 = n1841 | n14796 ;
  assign n18109 = n18108 ^ n16284 ^ 1'b0 ;
  assign n18106 = ( ~n426 & n1073 ) | ( ~n426 & n2696 ) | ( n1073 & n2696 ) ;
  assign n18105 = n6183 ^ n5486 ^ n5404 ;
  assign n18107 = n18106 ^ n18105 ^ 1'b0 ;
  assign n18110 = n18109 ^ n18107 ^ 1'b0 ;
  assign n18117 = n1081 & n4179 ;
  assign n18111 = ( ~n2402 & n6695 ) | ( ~n2402 & n12247 ) | ( n6695 & n12247 ) ;
  assign n18112 = n2825 ^ n1274 ^ 1'b0 ;
  assign n18113 = n2982 | n18112 ;
  assign n18114 = n18113 ^ n102 ^ 1'b0 ;
  assign n18115 = n8909 & n18114 ;
  assign n18116 = n18111 & n18115 ;
  assign n18118 = n18117 ^ n18116 ^ 1'b0 ;
  assign n18119 = n2086 & n6593 ;
  assign n18126 = n3931 & n6387 ;
  assign n18120 = n14778 ^ n4077 ^ 1'b0 ;
  assign n18121 = n7527 & ~n18120 ;
  assign n18122 = n7952 ^ n6105 ^ 1'b0 ;
  assign n18123 = ~n4964 & n18122 ;
  assign n18124 = ~x10 & n18123 ;
  assign n18125 = n18121 & ~n18124 ;
  assign n18127 = n18126 ^ n18125 ^ 1'b0 ;
  assign n18128 = n6962 & ~n13658 ;
  assign n18129 = n14802 & n18128 ;
  assign n18130 = n965 | n4823 ;
  assign n18131 = n18130 ^ n10034 ^ 1'b0 ;
  assign n18132 = ~n2447 & n18131 ;
  assign n18133 = n59 & n2745 ;
  assign n18134 = n15702 & n18133 ;
  assign n18135 = n14049 ^ n5117 ^ 1'b0 ;
  assign n18136 = n1909 & ~n18135 ;
  assign n18137 = ~n849 & n18136 ;
  assign n18138 = ~n8414 & n18137 ;
  assign n18139 = n7938 | n18138 ;
  assign n18140 = n4217 ^ n1400 ^ 1'b0 ;
  assign n18141 = n9683 | n18140 ;
  assign n18142 = n18139 & ~n18141 ;
  assign n18143 = n3245 & n17175 ;
  assign n18144 = n17859 ^ n5270 ^ 1'b0 ;
  assign n18145 = n18143 | n18144 ;
  assign n18146 = n15395 ^ n5406 ^ 1'b0 ;
  assign n18147 = ( n2885 & ~n2898 ) | ( n2885 & n18146 ) | ( ~n2898 & n18146 ) ;
  assign n18148 = n2519 & ~n2722 ;
  assign n18150 = n2022 & n9999 ;
  assign n18149 = ~n156 & n2566 ;
  assign n18151 = n18150 ^ n18149 ^ 1'b0 ;
  assign n18152 = n3551 & ~n14897 ;
  assign n18153 = n13541 ^ n3393 ^ 1'b0 ;
  assign n18154 = n12400 ^ n8211 ^ 1'b0 ;
  assign n18155 = n8738 & ~n14983 ;
  assign n18156 = n563 & n18155 ;
  assign n18157 = n18156 ^ n12327 ^ 1'b0 ;
  assign n18159 = n8995 ^ n7011 ^ n4219 ;
  assign n18158 = n6067 | n15169 ;
  assign n18160 = n18159 ^ n18158 ^ 1'b0 ;
  assign n18163 = n813 | n3307 ;
  assign n18164 = n18163 ^ n8790 ^ 1'b0 ;
  assign n18161 = ( n2280 & ~n2621 ) | ( n2280 & n5897 ) | ( ~n2621 & n5897 ) ;
  assign n18162 = n18161 ^ n8371 ^ 1'b0 ;
  assign n18165 = n18164 ^ n18162 ^ 1'b0 ;
  assign n18166 = n534 & ~n18165 ;
  assign n18167 = n8338 ^ n2294 ^ 1'b0 ;
  assign n18168 = ~n5008 & n18167 ;
  assign n18169 = n18168 ^ n6877 ^ n47 ;
  assign n18170 = n6019 | n7106 ;
  assign n18171 = n18170 ^ n11154 ^ 1'b0 ;
  assign n18172 = n2566 & ~n18171 ;
  assign n18173 = n13116 ^ n2606 ^ 1'b0 ;
  assign n18174 = n8536 & n18173 ;
  assign n18175 = n18174 ^ n9307 ^ 1'b0 ;
  assign n18178 = n8359 ^ n622 ^ 1'b0 ;
  assign n18179 = ~n4862 & n18178 ;
  assign n18176 = n6590 | n8365 ;
  assign n18177 = n3013 & n18176 ;
  assign n18180 = n18179 ^ n18177 ^ 1'b0 ;
  assign n18183 = n2316 & ~n3928 ;
  assign n18184 = ~n436 & n18183 ;
  assign n18185 = n4068 | n18048 ;
  assign n18186 = n18184 & ~n18185 ;
  assign n18181 = ~n2987 & n6392 ;
  assign n18182 = n18181 ^ n5802 ^ 1'b0 ;
  assign n18187 = n18186 ^ n18182 ^ 1'b0 ;
  assign n18188 = n1104 | n18187 ;
  assign n18189 = n3540 ^ n1803 ^ 1'b0 ;
  assign n18190 = n12834 | n18189 ;
  assign n18191 = n2551 & ~n9468 ;
  assign n18192 = n18190 & n18191 ;
  assign n18193 = n18192 ^ n11490 ^ n5482 ;
  assign n18194 = n4779 & ~n11124 ;
  assign n18195 = n18194 ^ n9011 ^ 1'b0 ;
  assign n18196 = n6008 | n7150 ;
  assign n18197 = n4489 | n18196 ;
  assign n18198 = n18197 ^ n6603 ^ 1'b0 ;
  assign n18199 = n3384 | n17887 ;
  assign n18200 = n18199 ^ n3566 ^ 1'b0 ;
  assign n18201 = n15999 & n18200 ;
  assign n18202 = ~n874 & n18201 ;
  assign n18203 = n4869 ^ n1836 ^ 1'b0 ;
  assign n18204 = n14586 | n18203 ;
  assign n18205 = n10296 & n18204 ;
  assign n18206 = n17089 ^ n6000 ^ 1'b0 ;
  assign n18207 = n7276 | n18206 ;
  assign n18208 = n13493 ^ n12945 ^ n3926 ;
  assign n18209 = ~n799 & n17349 ;
  assign n18210 = n18209 ^ n13627 ^ 1'b0 ;
  assign n18211 = ( ~n4118 & n7108 ) | ( ~n4118 & n18210 ) | ( n7108 & n18210 ) ;
  assign n18212 = ( ~n6227 & n9522 ) | ( ~n6227 & n13445 ) | ( n9522 & n13445 ) ;
  assign n18213 = n18212 ^ n8921 ^ 1'b0 ;
  assign n18214 = n15708 ^ n10125 ^ 1'b0 ;
  assign n18215 = n3803 & n18214 ;
  assign n18216 = ~n1525 & n6562 ;
  assign n18217 = ~n18215 & n18216 ;
  assign n18218 = n9939 | n18217 ;
  assign n18219 = n2958 & ~n5329 ;
  assign n18220 = n7707 & ~n18219 ;
  assign n18221 = n3244 | n5146 ;
  assign n18222 = ~n2321 & n4463 ;
  assign n18223 = n18221 & n18222 ;
  assign n18224 = n15448 ^ n686 ^ 1'b0 ;
  assign n18225 = n6537 ^ n5675 ^ n2126 ;
  assign n18226 = n18225 ^ n4294 ^ n4058 ;
  assign n18227 = n7792 & ~n9618 ;
  assign n18228 = n5408 & ~n11555 ;
  assign n18230 = n91 | n3170 ;
  assign n18229 = n1235 | n10741 ;
  assign n18231 = n18230 ^ n18229 ^ 1'b0 ;
  assign n18233 = ~n2418 & n3422 ;
  assign n18234 = ~n1698 & n18233 ;
  assign n18235 = n2859 ^ n2060 ^ 1'b0 ;
  assign n18236 = n18234 | n18235 ;
  assign n18232 = n6222 & n17138 ;
  assign n18237 = n18236 ^ n18232 ^ 1'b0 ;
  assign n18238 = n8780 ^ n1527 ^ n1234 ;
  assign n18239 = n3973 ^ n2071 ^ 1'b0 ;
  assign n18240 = n18239 ^ n9571 ^ n771 ;
  assign n18241 = ~n18238 & n18240 ;
  assign n18242 = ~n1503 & n2859 ;
  assign n18243 = ( ~n16153 & n16915 ) | ( ~n16153 & n18242 ) | ( n16915 & n18242 ) ;
  assign n18245 = n6511 & ~n6736 ;
  assign n18246 = ( n3517 & n4679 ) | ( n3517 & n18245 ) | ( n4679 & n18245 ) ;
  assign n18247 = ( ~n10408 & n11573 ) | ( ~n10408 & n18246 ) | ( n11573 & n18246 ) ;
  assign n18244 = n569 & n6340 ;
  assign n18248 = n18247 ^ n18244 ^ 1'b0 ;
  assign n18249 = n6269 ^ n2787 ^ 1'b0 ;
  assign n18250 = n18074 ^ n13963 ^ n12589 ;
  assign n18251 = n6639 ^ x3 ^ 1'b0 ;
  assign n18252 = ~n3833 & n18251 ;
  assign n18253 = n9605 ^ n6167 ^ 1'b0 ;
  assign n18254 = n18252 & ~n18253 ;
  assign n18255 = n4369 & ~n18254 ;
  assign n18256 = n2725 | n14119 ;
  assign n18257 = n5968 & ~n16556 ;
  assign n18258 = n5301 ^ n3567 ^ n1996 ;
  assign n18259 = ~n5318 & n18258 ;
  assign n18260 = ~n18257 & n18259 ;
  assign n18262 = ( ~n5440 & n7358 ) | ( ~n5440 & n9564 ) | ( n7358 & n9564 ) ;
  assign n18261 = n9173 & n9419 ;
  assign n18263 = n18262 ^ n18261 ^ 1'b0 ;
  assign n18264 = n7978 & ~n18263 ;
  assign n18265 = n6098 & ~n11594 ;
  assign n18266 = n10593 ^ n3792 ^ 1'b0 ;
  assign n18267 = n1009 | n4226 ;
  assign n18268 = n2248 & ~n18267 ;
  assign n18269 = n2801 & ~n18268 ;
  assign n18270 = n18269 ^ n8947 ^ 1'b0 ;
  assign n18271 = n2496 ^ n654 ^ 1'b0 ;
  assign n18272 = n18270 | n18271 ;
  assign n18273 = n2772 & n14593 ;
  assign n18274 = ~n5554 & n18273 ;
  assign n18276 = n8146 & n9658 ;
  assign n18277 = ~n8500 & n18276 ;
  assign n18275 = x7 & ~n830 ;
  assign n18278 = n18277 ^ n18275 ^ 1'b0 ;
  assign n18279 = n230 & ~n1666 ;
  assign n18280 = n18279 ^ n865 ^ 1'b0 ;
  assign n18281 = n13078 & n18280 ;
  assign n18282 = ~n18278 & n18281 ;
  assign n18283 = n3394 | n17809 ;
  assign n18284 = n18283 ^ n1848 ^ 1'b0 ;
  assign n18289 = n6482 ^ n4799 ^ 1'b0 ;
  assign n18288 = n13107 ^ n10484 ^ n5702 ;
  assign n18290 = n18289 ^ n18288 ^ n6625 ;
  assign n18285 = n12547 ^ n5167 ^ n3687 ;
  assign n18286 = ( n11073 & n11867 ) | ( n11073 & n18285 ) | ( n11867 & n18285 ) ;
  assign n18287 = n15692 & n18286 ;
  assign n18291 = n18290 ^ n18287 ^ 1'b0 ;
  assign n18292 = ( n1054 & ~n6833 ) | ( n1054 & n6887 ) | ( ~n6833 & n6887 ) ;
  assign n18294 = n9926 ^ n8281 ^ n416 ;
  assign n18293 = n2573 & ~n9724 ;
  assign n18295 = n18294 ^ n18293 ^ 1'b0 ;
  assign n18296 = ~n5512 & n15235 ;
  assign n18297 = n18296 ^ n957 ^ 1'b0 ;
  assign n18298 = n18297 ^ n10459 ^ 1'b0 ;
  assign n18299 = n18295 & ~n18298 ;
  assign n18300 = n1367 | n7062 ;
  assign n18301 = n18300 ^ n9541 ^ 1'b0 ;
  assign n18302 = n7433 & ~n12079 ;
  assign n18303 = n18302 ^ n11138 ^ 1'b0 ;
  assign n18304 = n18303 ^ n4231 ^ 1'b0 ;
  assign n18305 = n15233 ^ n12620 ^ n7866 ;
  assign n18306 = n17694 ^ n9700 ^ n9029 ;
  assign n18307 = ( ~n3894 & n5635 ) | ( ~n3894 & n18306 ) | ( n5635 & n18306 ) ;
  assign n18308 = n1779 ^ n1415 ^ 1'b0 ;
  assign n18309 = n3532 | n18308 ;
  assign n18310 = n949 | n18309 ;
  assign n18311 = n8275 & ~n18310 ;
  assign n18312 = n6000 | n18311 ;
  assign n18313 = ~n263 & n18312 ;
  assign n18314 = ~n18307 & n18313 ;
  assign n18315 = n2055 | n3563 ;
  assign n18316 = ( n1234 & n13862 ) | ( n1234 & ~n18315 ) | ( n13862 & ~n18315 ) ;
  assign n18317 = n2152 & ~n16777 ;
  assign n18318 = ~n11119 & n12750 ;
  assign n18319 = n18317 & n18318 ;
  assign n18320 = n18319 ^ n11724 ^ 1'b0 ;
  assign n18321 = n1069 | n4346 ;
  assign n18322 = ~n16499 & n18321 ;
  assign n18323 = n364 | n18322 ;
  assign n18324 = n8404 & ~n18323 ;
  assign n18325 = n7045 & n7935 ;
  assign n18326 = ~n2524 & n6745 ;
  assign n18327 = n15437 & ~n17038 ;
  assign n18330 = n5952 ^ n3824 ^ n2027 ;
  assign n18328 = n3029 ^ n2784 ^ 1'b0 ;
  assign n18329 = n12255 & ~n18328 ;
  assign n18331 = n18330 ^ n18329 ^ 1'b0 ;
  assign n18332 = n2999 | n9620 ;
  assign n18333 = n18332 ^ n13069 ^ n9052 ;
  assign n18337 = n2352 & ~n15651 ;
  assign n18336 = ( n3696 & n10356 ) | ( n3696 & n13099 ) | ( n10356 & n13099 ) ;
  assign n18334 = n1000 & ~n17116 ;
  assign n18335 = n1822 | n18334 ;
  assign n18338 = n18337 ^ n18336 ^ n18335 ;
  assign n18339 = n3610 ^ n1818 ^ 1'b0 ;
  assign n18340 = n3416 & ~n18339 ;
  assign n18341 = n18340 ^ n55 ^ 1'b0 ;
  assign n18342 = n6908 ^ n1754 ^ 1'b0 ;
  assign n18343 = n18342 ^ n9452 ^ 1'b0 ;
  assign n18344 = n6115 & n18343 ;
  assign n18345 = n7775 & n7870 ;
  assign n18346 = ~n18344 & n18345 ;
  assign n18347 = n570 | n7271 ;
  assign n18348 = n1709 | n11605 ;
  assign n18349 = n4769 ^ n1527 ^ 1'b0 ;
  assign n18350 = n11267 & n15003 ;
  assign n18351 = n9623 ^ n6139 ^ 1'b0 ;
  assign n18352 = n18351 ^ n23 ^ 1'b0 ;
  assign n18353 = n2886 & n18352 ;
  assign n18354 = n6609 ^ n5457 ^ 1'b0 ;
  assign n18355 = n18353 & ~n18354 ;
  assign n18356 = n15267 & n18355 ;
  assign n18357 = ( ~n10206 & n10380 ) | ( ~n10206 & n13002 ) | ( n10380 & n13002 ) ;
  assign n18358 = n11145 & n18357 ;
  assign n18359 = n15145 & n18358 ;
  assign n18360 = ( n5397 & n8385 ) | ( n5397 & ~n10090 ) | ( n8385 & ~n10090 ) ;
  assign n18361 = n6565 & ~n13627 ;
  assign n18362 = ~n11674 & n17989 ;
  assign n18363 = n18362 ^ n13230 ^ 1'b0 ;
  assign n18364 = n16467 ^ n15803 ^ 1'b0 ;
  assign n18365 = n2179 & ~n18364 ;
  assign n18366 = n6490 & ~n15801 ;
  assign n18367 = n18366 ^ n117 ^ 1'b0 ;
  assign n18368 = n4624 | n18367 ;
  assign n18369 = n18368 ^ n8994 ^ 1'b0 ;
  assign n18370 = n3584 & ~n13755 ;
  assign n18371 = n2807 & n18370 ;
  assign n18372 = n18371 ^ n1490 ^ 1'b0 ;
  assign n18373 = n16228 | n18372 ;
  assign n18374 = ~n9513 & n10404 ;
  assign n18375 = n13514 ^ n6564 ^ 1'b0 ;
  assign n18377 = ~n5195 & n7542 ;
  assign n18376 = n4976 & n5997 ;
  assign n18378 = n18377 ^ n18376 ^ 1'b0 ;
  assign n18382 = n7518 & n9753 ;
  assign n18381 = n4179 & n6431 ;
  assign n18379 = n4626 & n15715 ;
  assign n18380 = n18379 ^ n6277 ^ 1'b0 ;
  assign n18383 = n18382 ^ n18381 ^ n18380 ;
  assign n18384 = n17106 ^ n617 ^ 1'b0 ;
  assign n18385 = n17438 ^ n5969 ^ 1'b0 ;
  assign n18386 = n12084 & n18385 ;
  assign n18387 = n7021 & n11424 ;
  assign n18388 = n18387 ^ n6322 ^ 1'b0 ;
  assign n18389 = n521 & ~n13686 ;
  assign n18390 = n18389 ^ n11853 ^ 1'b0 ;
  assign n18391 = ( n3397 & ~n8891 ) | ( n3397 & n14170 ) | ( ~n8891 & n14170 ) ;
  assign n18392 = n11406 | n12214 ;
  assign n18393 = ( ~n249 & n9471 ) | ( ~n249 & n18392 ) | ( n9471 & n18392 ) ;
  assign n18394 = n18393 ^ n14632 ^ n2784 ;
  assign n18395 = n4884 | n15807 ;
  assign n18396 = n15631 ^ n3306 ^ n1561 ;
  assign n18397 = ~n2225 & n6527 ;
  assign n18398 = ~n15389 & n18397 ;
  assign n18399 = n5814 | n18398 ;
  assign n18400 = ~n1164 & n2825 ;
  assign n18401 = n14136 & n18400 ;
  assign n18402 = n18399 & ~n18401 ;
  assign n18403 = ( n2734 & n3128 ) | ( n2734 & ~n4300 ) | ( n3128 & ~n4300 ) ;
  assign n18404 = n11318 ^ n8654 ^ 1'b0 ;
  assign n18405 = n18404 ^ n17702 ^ 1'b0 ;
  assign n18406 = n6087 & ~n18405 ;
  assign n18407 = n18406 ^ n7785 ^ 1'b0 ;
  assign n18408 = n18403 & ~n18407 ;
  assign n18409 = n6186 & ~n9227 ;
  assign n18410 = n17449 & n18409 ;
  assign n18411 = n8026 ^ n6628 ^ 1'b0 ;
  assign n18412 = n788 & ~n18411 ;
  assign n18413 = ~n6457 & n18412 ;
  assign n18414 = ~n3473 & n18413 ;
  assign n18415 = ~n11119 & n14682 ;
  assign n18416 = n18415 ^ n16352 ^ n1825 ;
  assign n18417 = ~n10001 & n15009 ;
  assign n18418 = n2592 & n4002 ;
  assign n18419 = n18418 ^ n18272 ^ 1'b0 ;
  assign n18420 = n11053 & ~n13417 ;
  assign n18421 = n4458 & ~n7406 ;
  assign n18422 = n5280 & ~n6363 ;
  assign n18423 = n670 & n18422 ;
  assign n18424 = n3473 & ~n18423 ;
  assign n18425 = ~n566 & n18424 ;
  assign n18426 = n18421 & n18425 ;
  assign n18427 = n8074 & n17457 ;
  assign n18428 = ~n16231 & n18427 ;
  assign n18429 = n3871 ^ n2569 ^ 1'b0 ;
  assign n18430 = n18428 | n18429 ;
  assign n18431 = ~n2747 & n17995 ;
  assign n18432 = n1861 & ~n5601 ;
  assign n18433 = n612 | n7101 ;
  assign n18434 = n18432 & ~n18433 ;
  assign n18435 = ~n3271 & n18434 ;
  assign n18436 = n8191 & n15769 ;
  assign n18446 = n983 | n2587 ;
  assign n18437 = ~n7285 & n13844 ;
  assign n18438 = n12213 & n18437 ;
  assign n18442 = n3973 ^ n3483 ^ 1'b0 ;
  assign n18443 = n3084 & n18442 ;
  assign n18439 = n17035 ^ n5715 ^ 1'b0 ;
  assign n18440 = n17268 & ~n18439 ;
  assign n18441 = n2484 & n18440 ;
  assign n18444 = n18443 ^ n18441 ^ 1'b0 ;
  assign n18445 = n18438 | n18444 ;
  assign n18447 = n18446 ^ n18445 ^ 1'b0 ;
  assign n18448 = n8004 ^ n3299 ^ n1317 ;
  assign n18449 = ( ~n108 & n1645 ) | ( ~n108 & n18448 ) | ( n1645 & n18448 ) ;
  assign n18450 = n4480 & n18449 ;
  assign n18451 = ~n9919 & n18450 ;
  assign n18452 = n11632 | n18451 ;
  assign n18453 = n18452 ^ n10488 ^ 1'b0 ;
  assign n18454 = n7316 & n18453 ;
  assign n18455 = ( n664 & n8755 ) | ( n664 & ~n12918 ) | ( n8755 & ~n12918 ) ;
  assign n18456 = n18454 | n18455 ;
  assign n18457 = n14258 & ~n18456 ;
  assign n18458 = n18136 ^ n3238 ^ n107 ;
  assign n18459 = n18457 | n18458 ;
  assign n18460 = n13795 & ~n15819 ;
  assign n18461 = n3127 & n18460 ;
  assign n18462 = n601 | n2926 ;
  assign n18463 = ~n4014 & n18462 ;
  assign n18464 = n18463 ^ n10563 ^ 1'b0 ;
  assign n18465 = ~n18461 & n18464 ;
  assign n18466 = n7332 ^ n4138 ^ n1193 ;
  assign n18467 = n12708 & ~n18466 ;
  assign n18468 = n4086 | n17260 ;
  assign n18469 = n18468 ^ n3812 ^ 1'b0 ;
  assign n18470 = n7140 | n14604 ;
  assign n18471 = n5166 & n18470 ;
  assign n18472 = ~n6948 & n18471 ;
  assign n18473 = n18472 ^ n3223 ^ 1'b0 ;
  assign n18474 = n11041 ^ n965 ^ 1'b0 ;
  assign n18475 = n18474 ^ n7510 ^ 1'b0 ;
  assign n18476 = ~n13658 & n14555 ;
  assign n18477 = n1361 & n2662 ;
  assign n18478 = n18477 ^ n772 ^ 1'b0 ;
  assign n18479 = ( n6743 & n10884 ) | ( n6743 & n18478 ) | ( n10884 & n18478 ) ;
  assign n18480 = n11349 ^ n3393 ^ n1312 ;
  assign n18484 = n14126 ^ n9463 ^ n7060 ;
  assign n18481 = ~n557 & n680 ;
  assign n18482 = n18481 ^ n8994 ^ 1'b0 ;
  assign n18483 = n10059 & ~n18482 ;
  assign n18485 = n18484 ^ n18483 ^ 1'b0 ;
  assign n18486 = n7850 & ~n15163 ;
  assign n18487 = n18486 ^ n694 ^ 1'b0 ;
  assign n18488 = n3984 ^ n3688 ^ n517 ;
  assign n18489 = ~n9215 & n9388 ;
  assign n18490 = n18489 ^ n7228 ^ 1'b0 ;
  assign n18491 = n18490 ^ n3229 ^ 1'b0 ;
  assign n18492 = ~n18488 & n18491 ;
  assign n18493 = n12936 ^ n1374 ^ 1'b0 ;
  assign n18494 = n1448 & n3740 ;
  assign n18495 = n18494 ^ n8333 ^ 1'b0 ;
  assign n18496 = ~n15267 & n16671 ;
  assign n18497 = n12076 | n15138 ;
  assign n18498 = n17934 ^ n8206 ^ 1'b0 ;
  assign n18499 = n18498 ^ n4574 ^ n2148 ;
  assign n18500 = n18499 ^ n9005 ^ 1'b0 ;
  assign n18501 = n18500 ^ n15597 ^ n3227 ;
  assign n18502 = n2294 | n6743 ;
  assign n18503 = n18502 ^ n7103 ^ 1'b0 ;
  assign n18504 = n6050 & ~n15872 ;
  assign n18505 = n8182 | n18504 ;
  assign n18506 = n6161 & ~n18505 ;
  assign n18507 = ~n18503 & n18506 ;
  assign n18508 = ~n9222 & n18507 ;
  assign n18509 = ( n2218 & n4160 ) | ( n2218 & n8830 ) | ( n4160 & n8830 ) ;
  assign n18510 = ~n2303 & n2841 ;
  assign n18511 = n18510 ^ n7058 ^ n5006 ;
  assign n18512 = n18509 | n18511 ;
  assign n18513 = n18508 & ~n18512 ;
  assign n18514 = n811 & ~n15404 ;
  assign n18515 = ( ~n4270 & n13638 ) | ( ~n4270 & n17719 ) | ( n13638 & n17719 ) ;
  assign n18516 = ( ~n204 & n8356 ) | ( ~n204 & n15485 ) | ( n8356 & n15485 ) ;
  assign n18517 = n3867 | n18516 ;
  assign n18518 = n18515 | n18517 ;
  assign n18519 = n1950 | n5151 ;
  assign n18520 = n5793 & n18519 ;
  assign n18521 = n811 & n916 ;
  assign n18522 = n4889 ^ n2617 ^ 1'b0 ;
  assign n18523 = ~n15114 & n18522 ;
  assign n18524 = ~n18521 & n18523 ;
  assign n18525 = n18524 ^ n15238 ^ 1'b0 ;
  assign n18530 = n6899 & ~n8576 ;
  assign n18526 = n4144 | n7440 ;
  assign n18527 = n11535 | n18526 ;
  assign n18528 = n18527 ^ n3201 ^ 1'b0 ;
  assign n18529 = n5740 | n18528 ;
  assign n18531 = n18530 ^ n18529 ^ 1'b0 ;
  assign n18532 = n2199 | n6022 ;
  assign n18533 = n5534 & ~n18532 ;
  assign n18534 = n18533 ^ n2339 ^ 1'b0 ;
  assign n18535 = n18534 ^ n3660 ^ 1'b0 ;
  assign n18536 = n12133 | n18535 ;
  assign n18537 = n9746 | n16301 ;
  assign n18538 = n18537 ^ n3214 ^ 1'b0 ;
  assign n18539 = ( n6927 & n15330 ) | ( n6927 & n15874 ) | ( n15330 & n15874 ) ;
  assign n18540 = n17430 ^ n3163 ^ 1'b0 ;
  assign n18541 = n12375 & n18540 ;
  assign n18542 = n10674 | n18541 ;
  assign n18543 = n5856 | n8813 ;
  assign n18544 = n14354 | n18543 ;
  assign n18545 = n18544 ^ n6187 ^ 1'b0 ;
  assign n18546 = ~n8429 & n18545 ;
  assign n18547 = n11196 | n18546 ;
  assign n18548 = n2810 | n8633 ;
  assign n18549 = n2328 | n18548 ;
  assign n18550 = n18549 ^ n398 ^ 1'b0 ;
  assign n18551 = n1809 & n11999 ;
  assign n18552 = n18551 ^ n14534 ^ 1'b0 ;
  assign n18553 = n5715 ^ n3586 ^ 1'b0 ;
  assign n18554 = n18553 ^ n8533 ^ n2049 ;
  assign n18555 = ( ~n10052 & n18148 ) | ( ~n10052 & n18554 ) | ( n18148 & n18554 ) ;
  assign n18558 = n10576 ^ n7678 ^ 1'b0 ;
  assign n18559 = n14145 & n18558 ;
  assign n18556 = n7360 ^ n6585 ^ 1'b0 ;
  assign n18557 = n11316 & ~n18556 ;
  assign n18560 = n18559 ^ n18557 ^ 1'b0 ;
  assign n18561 = n12184 ^ n12180 ^ 1'b0 ;
  assign n18562 = n15712 & n18561 ;
  assign n18563 = n18562 ^ n11993 ^ n9616 ;
  assign n18564 = n961 | n4817 ;
  assign n18565 = n18564 ^ n5361 ^ 1'b0 ;
  assign n18566 = n18565 ^ n14125 ^ 1'b0 ;
  assign n18567 = n8895 ^ n6346 ^ 1'b0 ;
  assign n18568 = n1995 & n18567 ;
  assign n18569 = ~n760 & n3710 ;
  assign n18570 = ( ~n10106 & n18568 ) | ( ~n10106 & n18569 ) | ( n18568 & n18569 ) ;
  assign n18571 = n17251 ^ n1433 ^ 1'b0 ;
  assign n18572 = n5970 | n18571 ;
  assign n18573 = n18024 ^ n16883 ^ n12785 ;
  assign n18574 = n7071 | n18573 ;
  assign n18575 = n18572 | n18574 ;
  assign n18576 = ~n18570 & n18575 ;
  assign n18577 = ~n2190 & n18576 ;
  assign n18578 = ( n3847 & ~n6935 ) | ( n3847 & n18577 ) | ( ~n6935 & n18577 ) ;
  assign n18579 = n12167 ^ n3866 ^ 1'b0 ;
  assign n18580 = n1037 & ~n18579 ;
  assign n18581 = n1105 & n18580 ;
  assign n18582 = n5704 | n6743 ;
  assign n18583 = n18582 ^ n3737 ^ 1'b0 ;
  assign n18584 = n8472 | n18583 ;
  assign n18585 = n12751 | n18584 ;
  assign n18586 = ( n14084 & n18581 ) | ( n14084 & n18585 ) | ( n18581 & n18585 ) ;
  assign n18587 = n3214 ^ n2765 ^ 1'b0 ;
  assign n18588 = n8846 & n10628 ;
  assign n18589 = n18587 & n18588 ;
  assign n18590 = n8852 & n18589 ;
  assign n18591 = ~n17204 & n18590 ;
  assign n18592 = n706 & ~n11111 ;
  assign n18593 = n18592 ^ n11040 ^ n3687 ;
  assign n18594 = n15774 | n16409 ;
  assign n18595 = n8068 ^ n7634 ^ n7194 ;
  assign n18596 = n5292 & n18595 ;
  assign n18597 = ~n7500 & n13997 ;
  assign n18599 = n1862 & ~n5869 ;
  assign n18600 = n2984 & n18599 ;
  assign n18601 = n2170 | n18600 ;
  assign n18598 = n10131 ^ n5376 ^ n2571 ;
  assign n18602 = n18601 ^ n18598 ^ n2591 ;
  assign n18603 = n767 & ~n13056 ;
  assign n18604 = n18603 ^ n3703 ^ 1'b0 ;
  assign n18605 = n18604 ^ n4972 ^ 1'b0 ;
  assign n18606 = ~n12269 & n18605 ;
  assign n18607 = ~n9353 & n18606 ;
  assign n18608 = n18607 ^ n7657 ^ 1'b0 ;
  assign n18609 = n8882 ^ n7898 ^ 1'b0 ;
  assign n18611 = ~n1571 & n13899 ;
  assign n18612 = n18611 ^ n5625 ^ 1'b0 ;
  assign n18610 = n8389 | n8960 ;
  assign n18613 = n18612 ^ n18610 ^ 1'b0 ;
  assign n18614 = n6262 & ~n7167 ;
  assign n18615 = ~n2268 & n7587 ;
  assign n18616 = n18615 ^ n2980 ^ 1'b0 ;
  assign n18617 = n18616 ^ n8061 ^ n5043 ;
  assign n18618 = ~n4034 & n4156 ;
  assign n18619 = n18618 ^ n2870 ^ 1'b0 ;
  assign n18620 = n18619 ^ n3222 ^ 1'b0 ;
  assign n18621 = n18620 ^ n2768 ^ 1'b0 ;
  assign n18622 = n9824 ^ n6042 ^ n3930 ;
  assign n18623 = n1112 | n18622 ;
  assign n18624 = n18621 & n18623 ;
  assign n18625 = ~n18617 & n18624 ;
  assign n18626 = n13270 & n18625 ;
  assign n18627 = n13410 & ~n17827 ;
  assign n18628 = n18626 & n18627 ;
  assign n18629 = n4154 ^ n985 ^ 1'b0 ;
  assign n18630 = n17062 & ~n18629 ;
  assign n18631 = n3477 ^ n2344 ^ 1'b0 ;
  assign n18632 = n14299 ^ n12175 ^ 1'b0 ;
  assign n18633 = n18631 | n18632 ;
  assign n18634 = n13307 | n18633 ;
  assign n18635 = ~n15238 & n18634 ;
  assign n18636 = n18635 ^ n5028 ^ 1'b0 ;
  assign n18637 = n18630 & ~n18636 ;
  assign n18638 = ~n6282 & n13854 ;
  assign n18639 = n5325 ^ n556 ^ 1'b0 ;
  assign n18640 = n18639 ^ n4057 ^ 1'b0 ;
  assign n18641 = ~n592 & n11542 ;
  assign n18642 = n3158 & n18641 ;
  assign n18643 = n13890 ^ n5036 ^ n313 ;
  assign n18644 = n10500 & n18643 ;
  assign n18645 = ~n6705 & n18644 ;
  assign n18646 = n18255 ^ n6437 ^ 1'b0 ;
  assign n18647 = n10072 & ~n10224 ;
  assign n18648 = n18647 ^ n1439 ^ 1'b0 ;
  assign n18649 = ~n2080 & n9805 ;
  assign n18650 = n18648 & n18649 ;
  assign n18651 = n18650 ^ n3054 ^ 1'b0 ;
  assign n18652 = n9244 & ~n13109 ;
  assign n18653 = n16853 ^ n8772 ^ 1'b0 ;
  assign n18654 = n18652 & ~n18653 ;
  assign n18655 = ( n8567 & ~n12457 ) | ( n8567 & n12817 ) | ( ~n12457 & n12817 ) ;
  assign n18656 = ( n3853 & ~n7185 ) | ( n3853 & n15444 ) | ( ~n7185 & n15444 ) ;
  assign n18657 = n11243 ^ n8259 ^ 1'b0 ;
  assign n18658 = n18656 | n18657 ;
  assign n18659 = ~n6082 & n13520 ;
  assign n18660 = n10361 & n18659 ;
  assign n18661 = ~n9866 & n15184 ;
  assign n18662 = n6009 & n18661 ;
  assign n18663 = n13270 ^ n10129 ^ 1'b0 ;
  assign n18664 = ~n18662 & n18663 ;
  assign n18665 = ~n1311 & n6245 ;
  assign n18666 = ~n8824 & n18665 ;
  assign n18667 = n18666 ^ n7841 ^ 1'b0 ;
  assign n18668 = n527 & ~n17203 ;
  assign n18669 = n3193 & ~n12373 ;
  assign n18670 = ~n5022 & n18669 ;
  assign n18671 = n18670 ^ n1940 ^ 1'b0 ;
  assign n18672 = n1854 | n15870 ;
  assign n18673 = n16064 ^ n1000 ^ 1'b0 ;
  assign n18674 = ~n5175 & n18673 ;
  assign n18675 = n12296 ^ n9788 ^ n9245 ;
  assign n18676 = n16260 & ~n18675 ;
  assign n18677 = ~n9783 & n18676 ;
  assign n18678 = n368 & n5095 ;
  assign n18679 = n933 & n18678 ;
  assign n18680 = n18679 ^ n15075 ^ n8980 ;
  assign n18681 = n8889 & ~n14148 ;
  assign n18682 = n18680 & ~n18681 ;
  assign n18683 = n18682 ^ n18485 ^ 1'b0 ;
  assign n18684 = n14893 ^ n2090 ^ n1656 ;
  assign n18685 = n4009 | n18684 ;
  assign n18686 = n7763 | n18685 ;
  assign n18687 = n8490 | n18686 ;
  assign n18688 = n4116 ^ n2289 ^ n1108 ;
  assign n18689 = ( n6750 & n8644 ) | ( n6750 & ~n11311 ) | ( n8644 & ~n11311 ) ;
  assign n18698 = ~n890 & n2324 ;
  assign n18699 = ~n8185 & n18698 ;
  assign n18690 = ~n132 & n4745 ;
  assign n18691 = n8054 ^ n7790 ^ 1'b0 ;
  assign n18692 = n12252 & n18691 ;
  assign n18693 = ~n1752 & n7680 ;
  assign n18694 = n18693 ^ n7449 ^ 1'b0 ;
  assign n18695 = n18694 ^ n16534 ^ n2844 ;
  assign n18696 = n18692 & ~n18695 ;
  assign n18697 = ~n18690 & n18696 ;
  assign n18700 = n18699 ^ n18697 ^ 1'b0 ;
  assign n18701 = n12441 & n18700 ;
  assign n18705 = ~n498 & n7659 ;
  assign n18702 = ( n695 & n4228 ) | ( n695 & n15112 ) | ( n4228 & n15112 ) ;
  assign n18703 = n6638 & n18702 ;
  assign n18704 = n18703 ^ n15697 ^ 1'b0 ;
  assign n18706 = n18705 ^ n18704 ^ 1'b0 ;
  assign n18707 = n12249 & n15405 ;
  assign n18708 = ~n5233 & n9041 ;
  assign n18709 = n18708 ^ n711 ^ 1'b0 ;
  assign n18710 = ~n716 & n18709 ;
  assign n18711 = n15610 ^ n1748 ^ 1'b0 ;
  assign n18712 = ( n6889 & n11511 ) | ( n6889 & n18711 ) | ( n11511 & n18711 ) ;
  assign n18714 = n4058 | n6018 ;
  assign n18715 = n7373 | n18714 ;
  assign n18716 = n18715 ^ n4426 ^ n3307 ;
  assign n18713 = n1201 & ~n4900 ;
  assign n18717 = n18716 ^ n18713 ^ 1'b0 ;
  assign n18718 = n945 & ~n11986 ;
  assign n18719 = n3581 & n18718 ;
  assign n18720 = ( n2673 & ~n16648 ) | ( n2673 & n18719 ) | ( ~n16648 & n18719 ) ;
  assign n18721 = n15638 | n18720 ;
  assign n18722 = n9441 & ~n17836 ;
  assign n18723 = ( ~n358 & n2607 ) | ( ~n358 & n6692 ) | ( n2607 & n6692 ) ;
  assign n18724 = n18722 & ~n18723 ;
  assign n18725 = ~n1969 & n18724 ;
  assign n18726 = ( n4941 & n4959 ) | ( n4941 & n16758 ) | ( n4959 & n16758 ) ;
  assign n18727 = n3137 | n10265 ;
  assign n18728 = n7707 & n17638 ;
  assign n18729 = ~n3069 & n11117 ;
  assign n18730 = ( n11902 & ~n18728 ) | ( n11902 & n18729 ) | ( ~n18728 & n18729 ) ;
  assign n18731 = n18727 | n18730 ;
  assign n18732 = n12060 | n12573 ;
  assign n18733 = n14603 ^ n9091 ^ 1'b0 ;
  assign n18734 = n12379 ^ n2760 ^ 1'b0 ;
  assign n18735 = n18733 | n18734 ;
  assign n18736 = n18735 ^ n14587 ^ n784 ;
  assign n18748 = n6557 | n12033 ;
  assign n18749 = ~n3780 & n4147 ;
  assign n18750 = n18749 ^ n4114 ^ 1'b0 ;
  assign n18751 = ~n18748 & n18750 ;
  assign n18752 = n741 & n18751 ;
  assign n18753 = n18752 ^ n13733 ^ 1'b0 ;
  assign n18754 = n9902 ^ n1789 ^ 1'b0 ;
  assign n18755 = ~n818 & n18754 ;
  assign n18756 = n18753 & n18755 ;
  assign n18742 = ( n462 & n1033 ) | ( n462 & n5153 ) | ( n1033 & n5153 ) ;
  assign n18738 = ~n2485 & n9716 ;
  assign n18739 = n6104 & n18738 ;
  assign n18740 = n2382 | n18739 ;
  assign n18741 = n7307 | n18740 ;
  assign n18743 = n18742 ^ n18741 ^ 1'b0 ;
  assign n18737 = n13172 & ~n18733 ;
  assign n18744 = n18743 ^ n18737 ^ 1'b0 ;
  assign n18745 = n12632 | n18744 ;
  assign n18746 = n18745 ^ n3392 ^ 1'b0 ;
  assign n18747 = n14228 & n18746 ;
  assign n18757 = n18756 ^ n18747 ^ 1'b0 ;
  assign n18758 = n3694 ^ n2492 ^ 1'b0 ;
  assign n18759 = n741 & ~n895 ;
  assign n18760 = n11084 ^ n2256 ^ 1'b0 ;
  assign n18761 = n5366 | n18760 ;
  assign n18762 = n18761 ^ n4429 ^ 1'b0 ;
  assign n18763 = n17855 | n18762 ;
  assign n18764 = n1817 & ~n14706 ;
  assign n18765 = ( n145 & n10775 ) | ( n145 & ~n13216 ) | ( n10775 & ~n13216 ) ;
  assign n18766 = n14049 ^ n1568 ^ 1'b0 ;
  assign n18767 = n6301 ^ n5259 ^ 1'b0 ;
  assign n18768 = n3329 & ~n18767 ;
  assign n18769 = ~n299 & n2723 ;
  assign n18770 = ~n3040 & n18769 ;
  assign n18771 = ~n30 & n18770 ;
  assign n18772 = ~n2845 & n7925 ;
  assign n18773 = n18772 ^ n5799 ^ 1'b0 ;
  assign n18774 = n256 & n1281 ;
  assign n18775 = ~n4497 & n18774 ;
  assign n18776 = n18181 & ~n18775 ;
  assign n18777 = n18773 & n18776 ;
  assign n18784 = n1771 & ~n1896 ;
  assign n18785 = n680 | n18784 ;
  assign n18786 = n6110 | n18785 ;
  assign n18780 = n8349 & ~n11184 ;
  assign n18781 = ~n14677 & n16816 ;
  assign n18782 = n18781 ^ n13463 ^ 1'b0 ;
  assign n18783 = n18780 & n18782 ;
  assign n18778 = n18008 ^ n6345 ^ 1'b0 ;
  assign n18779 = n1245 | n18778 ;
  assign n18787 = n18786 ^ n18783 ^ n18779 ;
  assign n18788 = n14409 ^ n6475 ^ 1'b0 ;
  assign n18789 = n7264 ^ n5628 ^ 1'b0 ;
  assign n18790 = n3314 | n16836 ;
  assign n18791 = n13232 & ~n18790 ;
  assign n18792 = n9401 ^ n5587 ^ 1'b0 ;
  assign n18793 = n8733 & n13660 ;
  assign n18794 = n15857 ^ n12432 ^ 1'b0 ;
  assign n18795 = ~n5601 & n11254 ;
  assign n18796 = n18794 & n18795 ;
  assign n18797 = n10852 ^ n7121 ^ 1'b0 ;
  assign n18798 = n7994 & ~n16588 ;
  assign n18799 = n18798 ^ n1962 ^ 1'b0 ;
  assign n18800 = n18799 ^ n13008 ^ 1'b0 ;
  assign n18801 = n6842 ^ n6245 ^ 1'b0 ;
  assign n18802 = n16510 | n18801 ;
  assign n18803 = n3964 & n11642 ;
  assign n18804 = n4053 & n12017 ;
  assign n18805 = n15334 ^ n11219 ^ 1'b0 ;
  assign n18806 = n17748 | n18805 ;
  assign n18807 = n18804 | n18806 ;
  assign n18808 = n2209 & ~n18807 ;
  assign n18810 = n1529 & ~n1630 ;
  assign n18811 = ~n6175 & n18810 ;
  assign n18809 = n8362 & ~n9462 ;
  assign n18812 = n18811 ^ n18809 ^ 1'b0 ;
  assign n18813 = n3236 & ~n5458 ;
  assign n18814 = n18692 ^ n9371 ^ 1'b0 ;
  assign n18815 = n5189 & ~n18814 ;
  assign n18816 = n18813 | n18815 ;
  assign n18817 = ~n6607 & n18816 ;
  assign n18818 = ~n18812 & n18817 ;
  assign n18819 = n237 & ~n2858 ;
  assign n18820 = n15056 & ~n18819 ;
  assign n18821 = n8304 ^ n7134 ^ 1'b0 ;
  assign n18822 = n18820 & n18821 ;
  assign n18823 = n8239 & n17264 ;
  assign n18824 = n12463 ^ n5692 ^ 1'b0 ;
  assign n18827 = n7956 ^ n3872 ^ 1'b0 ;
  assign n18828 = n8106 & ~n18827 ;
  assign n18825 = n13546 ^ n975 ^ 1'b0 ;
  assign n18826 = ( ~n324 & n11372 ) | ( ~n324 & n18825 ) | ( n11372 & n18825 ) ;
  assign n18829 = n18828 ^ n18826 ^ 1'b0 ;
  assign n18834 = n8684 ^ n8023 ^ n6520 ;
  assign n18831 = n1796 ^ x7 ^ 1'b0 ;
  assign n18830 = n5766 | n8441 ;
  assign n18832 = n18831 ^ n18830 ^ 1'b0 ;
  assign n18833 = n6383 & n18832 ;
  assign n18835 = n18834 ^ n18833 ^ 1'b0 ;
  assign n18836 = n18289 ^ n859 ^ 1'b0 ;
  assign n18837 = ( n3309 & n12433 ) | ( n3309 & n18836 ) | ( n12433 & n18836 ) ;
  assign n18838 = n10428 & n18837 ;
  assign n18839 = n18838 ^ n4381 ^ 1'b0 ;
  assign n18840 = n18835 & n18839 ;
  assign n18844 = n12017 ^ n8852 ^ 1'b0 ;
  assign n18845 = n5080 & n18844 ;
  assign n18841 = n6917 & n9966 ;
  assign n18842 = ~n13990 & n18841 ;
  assign n18843 = n18842 ^ n7613 ^ 1'b0 ;
  assign n18846 = n18845 ^ n18843 ^ n12191 ;
  assign n18847 = n394 & n5432 ;
  assign n18848 = n18847 ^ n12129 ^ 1'b0 ;
  assign n18849 = n888 & ~n14202 ;
  assign n18854 = n8608 & ~n8972 ;
  assign n18855 = n969 & n18854 ;
  assign n18856 = n2854 | n18855 ;
  assign n18857 = n10475 | n18856 ;
  assign n18852 = n3002 ^ n1197 ^ 1'b0 ;
  assign n18853 = n9605 & ~n18852 ;
  assign n18850 = n12553 ^ n9012 ^ 1'b0 ;
  assign n18851 = n7414 & n18850 ;
  assign n18858 = n18857 ^ n18853 ^ n18851 ;
  assign n18859 = n10500 ^ n191 ^ 1'b0 ;
  assign n18860 = n18859 ^ n11184 ^ n6210 ;
  assign n18861 = n18860 ^ n3350 ^ 1'b0 ;
  assign n18862 = n10451 & n18861 ;
  assign n18863 = n4313 ^ n1462 ^ 1'b0 ;
  assign n18864 = ~n6193 & n11155 ;
  assign n18865 = n11258 ^ n6758 ^ 1'b0 ;
  assign n18866 = n18864 | n18865 ;
  assign n18867 = n7607 ^ n4322 ^ 1'b0 ;
  assign n18868 = n18866 | n18867 ;
  assign n18869 = n18868 ^ n10527 ^ 1'b0 ;
  assign n18870 = ( n16260 & ~n18863 ) | ( n16260 & n18869 ) | ( ~n18863 & n18869 ) ;
  assign n18872 = ( ~n415 & n6221 ) | ( ~n415 & n9085 ) | ( n6221 & n9085 ) ;
  assign n18871 = n10790 & n13522 ;
  assign n18873 = n18872 ^ n18871 ^ 1'b0 ;
  assign n18874 = n4212 & n9845 ;
  assign n18875 = n8697 ^ n1010 ^ 1'b0 ;
  assign n18876 = n18875 ^ n3833 ^ 1'b0 ;
  assign n18877 = n18876 ^ n12275 ^ 1'b0 ;
  assign n18878 = n18877 ^ n14999 ^ 1'b0 ;
  assign n18879 = n1931 & ~n18878 ;
  assign n18880 = ~n665 & n5806 ;
  assign n18881 = ~n271 & n4269 ;
  assign n18882 = n18881 ^ n4385 ^ 1'b0 ;
  assign n18883 = n13252 & n18882 ;
  assign n18884 = ~n12080 & n15868 ;
  assign n18885 = n18883 | n18884 ;
  assign n18888 = ( n590 & n11128 ) | ( n590 & ~n17257 ) | ( n11128 & ~n17257 ) ;
  assign n18886 = n6234 & n18620 ;
  assign n18887 = ~n7387 & n18886 ;
  assign n18889 = n18888 ^ n18887 ^ 1'b0 ;
  assign n18890 = n18889 ^ n3843 ^ n82 ;
  assign n18891 = n1319 | n5258 ;
  assign n18892 = n17951 & ~n18891 ;
  assign n18893 = n18892 ^ n6186 ^ 1'b0 ;
  assign n18894 = n5014 ^ n2041 ^ 1'b0 ;
  assign n18895 = n13748 ^ n548 ^ 1'b0 ;
  assign n18896 = ~n10118 & n17860 ;
  assign n18897 = n15410 ^ n6919 ^ 1'b0 ;
  assign n18898 = n5001 & n18897 ;
  assign n18899 = n1766 & n18898 ;
  assign n18901 = n12680 ^ n5958 ^ 1'b0 ;
  assign n18902 = n9903 & ~n18901 ;
  assign n18903 = n13427 & n18902 ;
  assign n18904 = n18903 ^ n5626 ^ 1'b0 ;
  assign n18900 = n4972 & ~n11275 ;
  assign n18905 = n18904 ^ n18900 ^ 1'b0 ;
  assign n18906 = ~n2230 & n4712 ;
  assign n18907 = n18906 ^ n2695 ^ 1'b0 ;
  assign n18908 = n688 & n18907 ;
  assign n18909 = ~n913 & n18908 ;
  assign n18910 = n8008 & n18909 ;
  assign n18911 = ~n5298 & n8635 ;
  assign n18912 = n2541 & ~n18911 ;
  assign n18913 = n18912 ^ n11865 ^ 1'b0 ;
  assign n18914 = n17100 ^ n3519 ^ 1'b0 ;
  assign n18915 = n10854 ^ n5098 ^ 1'b0 ;
  assign n18916 = n5534 & ~n18915 ;
  assign n18917 = n12002 | n18916 ;
  assign n18919 = n1979 & n9519 ;
  assign n18918 = n11213 & n13812 ;
  assign n18920 = n18919 ^ n18918 ^ 1'b0 ;
  assign n18921 = n18920 ^ n14202 ^ 1'b0 ;
  assign n18923 = n17800 ^ n5281 ^ n1525 ;
  assign n18922 = n3867 & n4485 ;
  assign n18924 = n18923 ^ n18922 ^ 1'b0 ;
  assign n18925 = n2955 | n18924 ;
  assign n18926 = n4701 | n18925 ;
  assign n18927 = n401 & ~n10319 ;
  assign n18928 = n18926 | n18927 ;
  assign n18929 = n18928 ^ n10815 ^ 1'b0 ;
  assign n18930 = n6115 ^ n1861 ^ 1'b0 ;
  assign n18931 = n5149 | n11871 ;
  assign n18932 = n14437 ^ n9947 ^ 1'b0 ;
  assign n18933 = ( n6811 & n7344 ) | ( n6811 & ~n13676 ) | ( n7344 & ~n13676 ) ;
  assign n18934 = n1150 & ~n1186 ;
  assign n18935 = ~n2841 & n8766 ;
  assign n18936 = ~n18745 & n18935 ;
  assign n18937 = n18934 & n18936 ;
  assign n18938 = ( n7680 & ~n12608 ) | ( n7680 & n18937 ) | ( ~n12608 & n18937 ) ;
  assign n18939 = n18192 | n18938 ;
  assign n18940 = n18470 | n18939 ;
  assign n18941 = ( n2493 & n11044 ) | ( n2493 & n18940 ) | ( n11044 & n18940 ) ;
  assign n18942 = n13782 | n18899 ;
  assign n18943 = n18942 ^ n14580 ^ 1'b0 ;
  assign n18944 = n10428 & ~n15517 ;
  assign n18945 = n16282 ^ n14699 ^ 1'b0 ;
  assign n18946 = n18945 ^ n2138 ^ 1'b0 ;
  assign n18947 = n12874 & n18946 ;
  assign n18948 = n12439 & ~n13202 ;
  assign n18949 = n14547 ^ n5123 ^ 1'b0 ;
  assign n18950 = n11977 | n18949 ;
  assign n18951 = n18950 ^ n5324 ^ 1'b0 ;
  assign n18952 = ( n11769 & ~n18948 ) | ( n11769 & n18951 ) | ( ~n18948 & n18951 ) ;
  assign n18953 = ~n500 & n7705 ;
  assign n18954 = n18953 ^ n10025 ^ 1'b0 ;
  assign n18955 = n18954 ^ n8549 ^ n897 ;
  assign n18956 = ~n12233 & n18955 ;
  assign n18957 = n14694 & n18956 ;
  assign n18958 = n4627 & ~n15636 ;
  assign n18959 = ( ~n4986 & n12525 ) | ( ~n4986 & n18958 ) | ( n12525 & n18958 ) ;
  assign n18960 = n11529 ^ n6047 ^ 1'b0 ;
  assign n18961 = ~n5156 & n18960 ;
  assign n18962 = n2452 ^ n2044 ^ 1'b0 ;
  assign n18963 = ~n2044 & n18962 ;
  assign n18964 = n98 & ~n1052 ;
  assign n18965 = n18963 & ~n18964 ;
  assign n18966 = ~n18961 & n18965 ;
  assign n18967 = n153 | n8061 ;
  assign n18968 = n18716 ^ n4685 ^ 1'b0 ;
  assign n18969 = ~n18967 & n18968 ;
  assign n18971 = n2479 | n13123 ;
  assign n18972 = ( ~n8441 & n9868 ) | ( ~n8441 & n18971 ) | ( n9868 & n18971 ) ;
  assign n18970 = n41 | n11276 ;
  assign n18973 = n18972 ^ n18970 ^ 1'b0 ;
  assign n18974 = n18973 ^ n8135 ^ 1'b0 ;
  assign n18975 = n8735 ^ n6829 ^ 1'b0 ;
  assign n18976 = n15214 ^ n3581 ^ 1'b0 ;
  assign n18977 = n13546 ^ n3585 ^ 1'b0 ;
  assign n18978 = n8857 ^ n3027 ^ 1'b0 ;
  assign n18979 = n18977 & n18978 ;
  assign n18980 = n18979 ^ n530 ^ 1'b0 ;
  assign n18981 = n7978 & n18980 ;
  assign n18982 = ~n5289 & n5339 ;
  assign n18983 = n18982 ^ n14057 ^ 1'b0 ;
  assign n18984 = n7694 & n18983 ;
  assign n18985 = ( n3309 & n4275 ) | ( n3309 & ~n5218 ) | ( n4275 & ~n5218 ) ;
  assign n18986 = ( n8014 & n18984 ) | ( n8014 & ~n18985 ) | ( n18984 & ~n18985 ) ;
  assign n18987 = ( n5517 & n18981 ) | ( n5517 & ~n18986 ) | ( n18981 & ~n18986 ) ;
  assign n18988 = n829 & n5175 ;
  assign n18989 = ~n18987 & n18988 ;
  assign n18990 = n1545 & ~n7943 ;
  assign n18991 = n18059 ^ n16158 ^ n3633 ;
  assign n18992 = n9032 ^ n1370 ^ 1'b0 ;
  assign n18995 = n13902 ^ n8201 ^ 1'b0 ;
  assign n18996 = n8014 | n18995 ;
  assign n18993 = n8226 & n17272 ;
  assign n18994 = n18993 ^ n7543 ^ 1'b0 ;
  assign n18997 = n18996 ^ n18994 ^ n1893 ;
  assign n18998 = n7218 ^ n3897 ^ 1'b0 ;
  assign n18999 = n18998 ^ n18904 ^ 1'b0 ;
  assign n19000 = n533 & ~n11283 ;
  assign n19001 = n5794 | n19000 ;
  assign n19002 = n19001 ^ n4684 ^ 1'b0 ;
  assign n19003 = n2542 | n19002 ;
  assign n19004 = n19003 ^ n8885 ^ 1'b0 ;
  assign n19007 = n7307 | n11446 ;
  assign n19005 = n7178 ^ n6639 ^ n2644 ;
  assign n19006 = n19005 ^ n17789 ^ n14188 ;
  assign n19008 = n19007 ^ n19006 ^ 1'b0 ;
  assign n19009 = n19004 | n19008 ;
  assign n19010 = ~n99 & n8480 ;
  assign n19011 = ~n139 & n2751 ;
  assign n19012 = n19011 ^ n10098 ^ 1'b0 ;
  assign n19013 = n19012 ^ n14885 ^ 1'b0 ;
  assign n19014 = n19013 ^ n2984 ^ 1'b0 ;
  assign n19015 = n7182 ^ n2251 ^ 1'b0 ;
  assign n19016 = ~n19014 & n19015 ;
  assign n19017 = ~n9158 & n16593 ;
  assign n19018 = n7741 ^ n1642 ^ 1'b0 ;
  assign n19019 = n2662 | n6985 ;
  assign n19020 = n11372 & n19019 ;
  assign n19021 = ~n5253 & n19020 ;
  assign n19022 = n5845 ^ n2176 ^ 1'b0 ;
  assign n19023 = n12140 ^ n8907 ^ n7210 ;
  assign n19024 = n5095 | n8813 ;
  assign n19025 = ( n158 & n2456 ) | ( n158 & ~n5832 ) | ( n2456 & ~n5832 ) ;
  assign n19026 = n3717 | n19025 ;
  assign n19027 = n2416 & n9755 ;
  assign n19028 = ~n15336 & n19027 ;
  assign n19029 = n18899 ^ n12405 ^ 1'b0 ;
  assign n19030 = n17128 ^ n13708 ^ 1'b0 ;
  assign n19031 = ~n1276 & n14170 ;
  assign n19032 = n19031 ^ n7069 ^ 1'b0 ;
  assign n19033 = n19030 | n19032 ;
  assign n19034 = n19033 ^ n16500 ^ 1'b0 ;
  assign n19037 = ~n1414 & n2867 ;
  assign n19038 = n19037 ^ n2280 ^ 1'b0 ;
  assign n19035 = ~n2216 & n10734 ;
  assign n19036 = n7575 & ~n19035 ;
  assign n19039 = n19038 ^ n19036 ^ 1'b0 ;
  assign n19041 = x10 & ~n5640 ;
  assign n19040 = n5122 | n6306 ;
  assign n19042 = n19041 ^ n19040 ^ 1'b0 ;
  assign n19044 = ( ~n3867 & n4304 ) | ( ~n3867 & n6638 ) | ( n4304 & n6638 ) ;
  assign n19043 = ~n3971 & n9887 ;
  assign n19045 = n19044 ^ n19043 ^ 1'b0 ;
  assign n19046 = n13393 & ~n13764 ;
  assign n19047 = n19046 ^ n5665 ^ 1'b0 ;
  assign n19049 = ~n7361 & n16212 ;
  assign n19050 = ~n388 & n19049 ;
  assign n19048 = ~n4543 & n5666 ;
  assign n19051 = n19050 ^ n19048 ^ 1'b0 ;
  assign n19052 = n6762 ^ n3658 ^ n3127 ;
  assign n19053 = n16402 | n19052 ;
  assign n19054 = n11712 ^ n10078 ^ 1'b0 ;
  assign n19055 = ~n11064 & n19054 ;
  assign n19056 = ~n478 & n6374 ;
  assign n19057 = ~n9432 & n19056 ;
  assign n19058 = n16551 ^ n181 ^ 1'b0 ;
  assign n19059 = n1988 | n5086 ;
  assign n19060 = n19059 ^ n10416 ^ 1'b0 ;
  assign n19061 = n19060 ^ n13157 ^ 1'b0 ;
  assign n19062 = n19058 & ~n19061 ;
  assign n19063 = ~n126 & n14042 ;
  assign n19064 = n19063 ^ n14692 ^ 1'b0 ;
  assign n19065 = n2432 | n6813 ;
  assign n19066 = n3607 ^ n2942 ^ 1'b0 ;
  assign n19067 = ~n2588 & n4127 ;
  assign n19068 = ~n4455 & n19067 ;
  assign n19069 = n15739 ^ n1656 ^ 1'b0 ;
  assign n19070 = n3357 & n19069 ;
  assign n19071 = ( n5716 & n12368 ) | ( n5716 & n19070 ) | ( n12368 & n19070 ) ;
  assign n19072 = n5003 & n12725 ;
  assign n19073 = n5333 & n7092 ;
  assign n19074 = n9905 & n19073 ;
  assign n19076 = n299 & ~n7265 ;
  assign n19075 = n7449 & n9592 ;
  assign n19077 = n19076 ^ n19075 ^ 1'b0 ;
  assign n19078 = ~n2693 & n16628 ;
  assign n19079 = n19078 ^ n10311 ^ n9855 ;
  assign n19080 = n19079 ^ n7886 ^ 1'b0 ;
  assign n19081 = n6305 & n8460 ;
  assign n19082 = n6561 & n19081 ;
  assign n19083 = ~n8625 & n19082 ;
  assign n19084 = n16850 ^ n11420 ^ 1'b0 ;
  assign n19085 = n3241 ^ n3158 ^ 1'b0 ;
  assign n19086 = n11741 | n19085 ;
  assign n19087 = n698 & ~n5909 ;
  assign n19088 = n19087 ^ n3250 ^ 1'b0 ;
  assign n19089 = n16648 & n19088 ;
  assign n19090 = ~n12697 & n19089 ;
  assign n19091 = n13345 | n18688 ;
  assign n19092 = n6287 & n19091 ;
  assign n19093 = n9741 | n19092 ;
  assign n19094 = n19093 ^ n9423 ^ 1'b0 ;
  assign n19095 = n12183 | n13558 ;
  assign n19096 = n11182 | n16739 ;
  assign n19097 = n942 & ~n2583 ;
  assign n19098 = n15224 | n19097 ;
  assign n19099 = n6387 & n7150 ;
  assign n19100 = n14220 ^ n8027 ^ 1'b0 ;
  assign n19101 = n11439 ^ n5520 ^ 1'b0 ;
  assign n19102 = n7802 & ~n7996 ;
  assign n19103 = n13683 ^ n7477 ^ 1'b0 ;
  assign n19104 = n19102 | n19103 ;
  assign n19105 = ( n10955 & ~n11254 ) | ( n10955 & n18200 ) | ( ~n11254 & n18200 ) ;
  assign n19106 = n10280 ^ n8114 ^ 1'b0 ;
  assign n19107 = n1600 & ~n10222 ;
  assign n19108 = n19107 ^ n14887 ^ 1'b0 ;
  assign n19109 = ( n12071 & n19106 ) | ( n12071 & ~n19108 ) | ( n19106 & ~n19108 ) ;
  assign n19110 = ~n926 & n2785 ;
  assign n19111 = ~n2785 & n19110 ;
  assign n19112 = x4 & ~n453 ;
  assign n19113 = ~x4 & n19112 ;
  assign n19114 = n472 | n19113 ;
  assign n19115 = n472 & ~n19114 ;
  assign n19116 = n453 | n19115 ;
  assign n19117 = n453 & ~n19116 ;
  assign n19118 = n19111 | n19117 ;
  assign n19119 = n19111 & ~n19118 ;
  assign n19120 = n913 & n19119 ;
  assign n19121 = ~n1437 & n19120 ;
  assign n19122 = n1437 & n19121 ;
  assign n19134 = n940 & n5106 ;
  assign n19135 = ~n9457 & n19134 ;
  assign n19123 = n887 & ~n1502 ;
  assign n19124 = ~n887 & n19123 ;
  assign n19125 = n3120 & n14097 ;
  assign n19126 = ~n3120 & n19125 ;
  assign n19127 = n13366 | n19126 ;
  assign n19128 = n13366 & ~n19127 ;
  assign n19129 = n19128 ^ n8443 ^ 1'b0 ;
  assign n19130 = n2055 & n5010 ;
  assign n19131 = ~n2055 & n19130 ;
  assign n19132 = n19129 & ~n19131 ;
  assign n19133 = n19124 & n19132 ;
  assign n19136 = n19135 ^ n19133 ^ 1'b0 ;
  assign n19137 = ~n19122 & n19136 ;
  assign n19138 = n17964 & n19137 ;
  assign n19139 = ~n19137 & n19138 ;
  assign n19140 = n569 | n14386 ;
  assign n19141 = n10724 ^ n7646 ^ 1'b0 ;
  assign n19142 = n5924 & ~n16909 ;
  assign n19143 = ~n5596 & n19142 ;
  assign n19144 = n5098 ^ n1526 ^ 1'b0 ;
  assign n19146 = ~n4648 & n9999 ;
  assign n19145 = n9805 ^ n2144 ^ 1'b0 ;
  assign n19147 = n19146 ^ n19145 ^ 1'b0 ;
  assign n19148 = n7064 ^ n6860 ^ 1'b0 ;
  assign n19149 = n19148 ^ n8820 ^ n772 ;
  assign n19150 = n13103 ^ n8408 ^ 1'b0 ;
  assign n19151 = n19150 ^ n6539 ^ 1'b0 ;
  assign n19152 = n19149 & n19151 ;
  assign n19153 = n1572 & ~n11660 ;
  assign n19154 = n4588 | n5554 ;
  assign n19155 = n19153 & ~n19154 ;
  assign n19156 = n11487 ^ n1737 ^ 1'b0 ;
  assign n19157 = ~n156 & n17390 ;
  assign n19158 = ~n19156 & n19157 ;
  assign n19159 = n12463 ^ n9801 ^ n44 ;
  assign n19160 = n19159 ^ n13266 ^ 1'b0 ;
  assign n19161 = n16035 & ~n19160 ;
  assign n19162 = n16443 ^ n11708 ^ 1'b0 ;
  assign n19163 = n11964 & ~n19162 ;
  assign n19164 = n1684 & n5303 ;
  assign n19165 = n18679 ^ n4153 ^ 1'b0 ;
  assign n19166 = n19164 | n19165 ;
  assign n19167 = n19166 ^ n16155 ^ 1'b0 ;
  assign n19168 = ~n5786 & n15172 ;
  assign n19169 = n11833 & n19168 ;
  assign n19170 = n953 & ~n1248 ;
  assign n19171 = n19170 ^ n2068 ^ 1'b0 ;
  assign n19172 = ~n3737 & n19171 ;
  assign n19173 = ~n9455 & n19172 ;
  assign n19174 = n19173 ^ n2813 ^ 1'b0 ;
  assign n19175 = ~n19169 & n19174 ;
  assign n19176 = n1185 & n2635 ;
  assign n19177 = n16411 ^ n13423 ^ 1'b0 ;
  assign n19178 = n5106 & n19177 ;
  assign n19179 = ~n3066 & n19178 ;
  assign n19180 = n19176 & n19179 ;
  assign n19181 = n11720 | n19180 ;
  assign n19182 = n18516 ^ n7559 ^ n4930 ;
  assign n19183 = n11958 ^ n8953 ^ x2 ;
  assign n19184 = n2089 ^ n957 ^ 1'b0 ;
  assign n19185 = x3 & ~n19184 ;
  assign n19188 = n14680 ^ n14206 ^ n9832 ;
  assign n19186 = n19035 ^ n7129 ^ 1'b0 ;
  assign n19187 = n887 & n19186 ;
  assign n19189 = n19188 ^ n19187 ^ 1'b0 ;
  assign n19190 = n7643 & ~n19189 ;
  assign n19191 = n6800 & n12562 ;
  assign n19192 = n10380 ^ n5966 ^ 1'b0 ;
  assign n19193 = ( n1314 & n19191 ) | ( n1314 & n19192 ) | ( n19191 & n19192 ) ;
  assign n19194 = n11157 ^ n10035 ^ 1'b0 ;
  assign n19195 = n9137 & ~n18438 ;
  assign n19196 = ( n1880 & ~n3313 ) | ( n1880 & n17817 ) | ( ~n3313 & n17817 ) ;
  assign n19197 = n1055 & n15592 ;
  assign n19198 = n19196 & n19197 ;
  assign n19199 = n3524 ^ n1540 ^ 1'b0 ;
  assign n19200 = n8615 & ~n11605 ;
  assign n19201 = ( n844 & n3299 ) | ( n844 & ~n8291 ) | ( n3299 & ~n8291 ) ;
  assign n19202 = n838 | n19201 ;
  assign n19203 = n20 & ~n19202 ;
  assign n19204 = n10924 ^ n9217 ^ n5716 ;
  assign n19205 = ~n19203 & n19204 ;
  assign n19206 = n6205 ^ n2911 ^ 1'b0 ;
  assign n19207 = n7471 & ~n19206 ;
  assign n19208 = ~n12696 & n19207 ;
  assign n19209 = n11095 & n19208 ;
  assign n19210 = n1175 ^ n1082 ^ 1'b0 ;
  assign n19211 = n19210 ^ n5392 ^ 1'b0 ;
  assign n19212 = n8211 | n19211 ;
  assign n19213 = ( n982 & n19209 ) | ( n982 & ~n19212 ) | ( n19209 & ~n19212 ) ;
  assign n19214 = n16295 & n19213 ;
  assign n19215 = n3102 | n11204 ;
  assign n19216 = n19215 ^ n2778 ^ 1'b0 ;
  assign n19217 = n11282 & ~n19216 ;
  assign n19218 = ~n8936 & n19217 ;
  assign n19219 = n5273 ^ n316 ^ 1'b0 ;
  assign n19220 = n7245 & ~n19219 ;
  assign n19221 = n19220 ^ n2885 ^ 1'b0 ;
  assign n19222 = n12500 & ~n19221 ;
  assign n19223 = n19222 ^ n3090 ^ 1'b0 ;
  assign n19224 = n4243 | n8841 ;
  assign n19225 = ~n12036 & n19224 ;
  assign n19226 = ~n7713 & n19225 ;
  assign n19227 = n13509 ^ n8474 ^ 1'b0 ;
  assign n19228 = n5122 & n19227 ;
  assign n19229 = n19228 ^ n18150 ^ 1'b0 ;
  assign n19231 = n6695 ^ n4536 ^ 1'b0 ;
  assign n19230 = ( ~n1509 & n1956 ) | ( ~n1509 & n7523 ) | ( n1956 & n7523 ) ;
  assign n19232 = n19231 ^ n19230 ^ n4560 ;
  assign n19233 = n434 & n2845 ;
  assign n19234 = n19233 ^ n906 ^ 1'b0 ;
  assign n19235 = n5490 & ~n19234 ;
  assign n19236 = n317 | n2476 ;
  assign n19237 = n19236 ^ n5442 ^ 1'b0 ;
  assign n19239 = n1156 & ~n1688 ;
  assign n19240 = n5303 | n19239 ;
  assign n19238 = n2391 ^ n1894 ^ n235 ;
  assign n19241 = n19240 ^ n19238 ^ n12426 ;
  assign n19242 = ( n3929 & ~n19237 ) | ( n3929 & n19241 ) | ( ~n19237 & n19241 ) ;
  assign n19243 = n11617 & ~n12366 ;
  assign n19244 = ~n12175 & n19243 ;
  assign n19245 = n3398 & n4795 ;
  assign n19247 = n1988 | n14964 ;
  assign n19248 = n19247 ^ n10594 ^ 1'b0 ;
  assign n19246 = n11794 ^ n3514 ^ n845 ;
  assign n19249 = n19248 ^ n19246 ^ 1'b0 ;
  assign n19250 = n15092 & ~n19249 ;
  assign n19251 = n16000 ^ n1554 ^ 1'b0 ;
  assign n19252 = n10190 & n19251 ;
  assign n19256 = ( n6607 & n7912 ) | ( n6607 & n15037 ) | ( n7912 & n15037 ) ;
  assign n19253 = n4949 ^ n935 ^ 1'b0 ;
  assign n19254 = n14222 | n19253 ;
  assign n19255 = n9716 & ~n19254 ;
  assign n19257 = n19256 ^ n19255 ^ 1'b0 ;
  assign n19258 = n7738 & ~n19257 ;
  assign n19259 = n19258 ^ n312 ^ 1'b0 ;
  assign n19260 = n19252 & n19259 ;
  assign n19261 = n17977 ^ n7896 ^ 1'b0 ;
  assign n19262 = ~n5684 & n11570 ;
  assign n19263 = ~n2281 & n19262 ;
  assign n19264 = ( n7315 & ~n11053 ) | ( n7315 & n19263 ) | ( ~n11053 & n19263 ) ;
  assign n19265 = ~n10178 & n19264 ;
  assign n19266 = n1554 ^ n652 ^ 1'b0 ;
  assign n19267 = ~n10007 & n19266 ;
  assign n19268 = n19267 ^ n12752 ^ 1'b0 ;
  assign n19269 = n4999 ^ n3737 ^ 1'b0 ;
  assign n19270 = n2833 & n13143 ;
  assign n19271 = ( n5627 & n8018 ) | ( n5627 & ~n19270 ) | ( n8018 & ~n19270 ) ;
  assign n19272 = n1023 & ~n19271 ;
  assign n19273 = n2918 & ~n14711 ;
  assign n19279 = n7427 & n15024 ;
  assign n19280 = n19279 ^ n8228 ^ 1'b0 ;
  assign n19274 = n2930 & n9889 ;
  assign n19275 = ~n3125 & n19274 ;
  assign n19276 = n1154 | n19275 ;
  assign n19277 = n19276 ^ n4163 ^ 1'b0 ;
  assign n19278 = ~n587 & n19277 ;
  assign n19281 = n19280 ^ n19278 ^ 1'b0 ;
  assign n19282 = ~n1406 & n1848 ;
  assign n19283 = ( n3749 & n13559 ) | ( n3749 & n14623 ) | ( n13559 & n14623 ) ;
  assign n19284 = ~n9921 & n19283 ;
  assign n19285 = n19282 & n19284 ;
  assign n19286 = n1231 ^ n1007 ^ 1'b0 ;
  assign n19287 = n1124 & ~n19286 ;
  assign n19288 = n19287 ^ n15555 ^ 1'b0 ;
  assign n19289 = n6446 ^ n5578 ^ 1'b0 ;
  assign n19290 = n8055 & n9068 ;
  assign n19291 = n3324 & n19290 ;
  assign n19292 = n19289 & ~n19291 ;
  assign n19293 = n4909 & ~n16932 ;
  assign n19294 = ~n19292 & n19293 ;
  assign n19295 = n1858 & ~n19294 ;
  assign n19296 = n19295 ^ n7646 ^ 1'b0 ;
  assign n19297 = n10319 ^ n8941 ^ 1'b0 ;
  assign n19298 = n14204 ^ n6334 ^ n3414 ;
  assign n19299 = x0 & n2186 ;
  assign n19300 = n19299 ^ n6361 ^ n667 ;
  assign n19301 = n19300 ^ n15809 ^ 1'b0 ;
  assign n19302 = n16880 & n19301 ;
  assign n19303 = n405 & n5066 ;
  assign n19304 = n428 & ~n2514 ;
  assign n19305 = n10850 ^ n10221 ^ 1'b0 ;
  assign n19306 = ( n9409 & n19304 ) | ( n9409 & ~n19305 ) | ( n19304 & ~n19305 ) ;
  assign n19307 = n19303 & ~n19306 ;
  assign n19308 = ~n3505 & n19307 ;
  assign n19309 = n11827 ^ n10195 ^ 1'b0 ;
  assign n19313 = n5963 ^ n2173 ^ 1'b0 ;
  assign n19314 = n11227 | n19313 ;
  assign n19310 = n3256 & ~n7581 ;
  assign n19311 = n19310 ^ n11904 ^ 1'b0 ;
  assign n19312 = n17693 & n19311 ;
  assign n19315 = n19314 ^ n19312 ^ 1'b0 ;
  assign n19316 = n17511 ^ n16373 ^ 1'b0 ;
  assign n19317 = n6835 ^ n6339 ^ 1'b0 ;
  assign n19318 = n19317 ^ n13025 ^ 1'b0 ;
  assign n19319 = n12360 | n19318 ;
  assign n19320 = ( n4817 & n5301 ) | ( n4817 & n8474 ) | ( n5301 & n8474 ) ;
  assign n19321 = n10035 ^ n4241 ^ 1'b0 ;
  assign n19322 = n4505 ^ n2932 ^ 1'b0 ;
  assign n19323 = n6616 | n6813 ;
  assign n19324 = n10008 | n19323 ;
  assign n19325 = n19324 ^ n11038 ^ 1'b0 ;
  assign n19326 = ~n19322 & n19325 ;
  assign n19327 = n19326 ^ n4915 ^ 1'b0 ;
  assign n19328 = ~n12107 & n14195 ;
  assign n19329 = ~n13457 & n19328 ;
  assign n19330 = n19329 ^ n4889 ^ 1'b0 ;
  assign n19331 = n6443 | n9490 ;
  assign n19332 = n8994 | n19331 ;
  assign n19333 = ~n6045 & n8558 ;
  assign n19334 = n19333 ^ n3592 ^ 1'b0 ;
  assign n19335 = n19334 ^ n10850 ^ 1'b0 ;
  assign n19336 = n9363 & n17656 ;
  assign n19337 = n19335 & n19336 ;
  assign n19339 = ( n3647 & n12089 ) | ( n3647 & ~n14409 ) | ( n12089 & ~n14409 ) ;
  assign n19338 = n8333 & ~n9723 ;
  assign n19340 = n19339 ^ n19338 ^ 1'b0 ;
  assign n19341 = n7968 ^ n2595 ^ 1'b0 ;
  assign n19342 = n17487 ^ n8673 ^ 1'b0 ;
  assign n19343 = n3763 | n8961 ;
  assign n19344 = n19343 ^ n12896 ^ n11262 ;
  assign n19345 = ( ~n6368 & n15020 ) | ( ~n6368 & n19344 ) | ( n15020 & n19344 ) ;
  assign n19346 = n3985 & n4627 ;
  assign n19347 = n5113 & ~n19346 ;
  assign n19348 = n16049 | n19347 ;
  assign n19349 = n19348 ^ n5478 ^ 1'b0 ;
  assign n19350 = n8037 & n19349 ;
  assign n19351 = ( ~n3252 & n19345 ) | ( ~n3252 & n19350 ) | ( n19345 & n19350 ) ;
  assign n19352 = n10920 ^ n8577 ^ 1'b0 ;
  assign n19353 = n8143 & ~n14707 ;
  assign n19354 = ( n5944 & n7401 ) | ( n5944 & n16160 ) | ( n7401 & n16160 ) ;
  assign n19355 = ~n17240 & n19354 ;
  assign n19356 = n6973 ^ n5587 ^ 1'b0 ;
  assign n19357 = n2674 & n19356 ;
  assign n19358 = n19357 ^ n18420 ^ n8154 ;
  assign n19359 = n8441 ^ n949 ^ 1'b0 ;
  assign n19360 = n6076 ^ n4367 ^ n2321 ;
  assign n19361 = n420 | n4620 ;
  assign n19362 = n2977 & n19361 ;
  assign n19363 = ~n19360 & n19362 ;
  assign n19364 = n19363 ^ n15890 ^ 1'b0 ;
  assign n19365 = n19364 ^ n134 ^ 1'b0 ;
  assign n19366 = n10868 ^ n135 ^ 1'b0 ;
  assign n19367 = ~n8375 & n19366 ;
  assign n19368 = n9730 & ~n19367 ;
  assign n19369 = n597 ^ n247 ^ 1'b0 ;
  assign n19370 = ~n19368 & n19369 ;
  assign n19371 = n2154 | n5377 ;
  assign n19372 = n8700 ^ n7291 ^ 1'b0 ;
  assign n19373 = ( n959 & n5891 ) | ( n959 & ~n11378 ) | ( n5891 & ~n11378 ) ;
  assign n19374 = n1727 & ~n19373 ;
  assign n19375 = ~n19372 & n19374 ;
  assign n19376 = n411 | n5327 ;
  assign n19377 = n19376 ^ n3501 ^ 1'b0 ;
  assign n19378 = n18984 & ~n19377 ;
  assign n19379 = n19375 & n19378 ;
  assign n19380 = ~n500 & n7228 ;
  assign n19381 = n19380 ^ n8448 ^ 1'b0 ;
  assign n19382 = n624 & n19381 ;
  assign n19383 = n19382 ^ n1022 ^ 1'b0 ;
  assign n19384 = n12420 ^ n8359 ^ n6625 ;
  assign n19386 = n533 & ~n11080 ;
  assign n19387 = ~n5197 & n19386 ;
  assign n19388 = n2466 | n3993 ;
  assign n19389 = n19387 & ~n19388 ;
  assign n19385 = n13088 ^ n11615 ^ 1'b0 ;
  assign n19390 = n19389 ^ n19385 ^ n4275 ;
  assign n19391 = n13638 ^ n1932 ^ 1'b0 ;
  assign n19392 = n3384 | n19391 ;
  assign n19393 = n9861 | n19392 ;
  assign n19394 = n9560 ^ n6689 ^ 1'b0 ;
  assign n19395 = n2538 | n19394 ;
  assign n19396 = n12740 | n19395 ;
  assign n19397 = n4882 ^ n2770 ^ 1'b0 ;
  assign n19398 = ~n5048 & n19397 ;
  assign n19399 = n19398 ^ n716 ^ 1'b0 ;
  assign n19400 = n8648 | n19399 ;
  assign n19401 = n7544 | n11052 ;
  assign n19402 = n19400 | n19401 ;
  assign n19403 = n6272 | n15700 ;
  assign n19404 = n19403 ^ n6384 ^ 1'b0 ;
  assign n19405 = n14083 & ~n19404 ;
  assign n19406 = n13725 & ~n17024 ;
  assign n19407 = n3855 & ~n6571 ;
  assign n19408 = n13350 & n19407 ;
  assign n19409 = ~n19406 & n19408 ;
  assign n19410 = ( n2217 & ~n6625 ) | ( n2217 & n14381 ) | ( ~n6625 & n14381 ) ;
  assign n19411 = n63 & n19410 ;
  assign n19412 = n1400 | n8478 ;
  assign n19413 = n349 | n352 ;
  assign n19414 = n849 & ~n5175 ;
  assign n19415 = n14614 ^ n2758 ^ 1'b0 ;
  assign n19416 = n15065 | n19415 ;
  assign n19417 = n19108 & ~n19416 ;
  assign n19418 = ( ~n8987 & n10467 ) | ( ~n8987 & n12404 ) | ( n10467 & n12404 ) ;
  assign n19419 = n15317 & n19418 ;
  assign n19420 = ~n1913 & n19419 ;
  assign n19421 = n17954 | n19420 ;
  assign n19422 = n14239 & n17656 ;
  assign n19424 = n13338 ^ n6245 ^ 1'b0 ;
  assign n19423 = n842 & ~n5554 ;
  assign n19425 = n19424 ^ n19423 ^ 1'b0 ;
  assign n19426 = n2909 & n3625 ;
  assign n19427 = n19426 ^ n7395 ^ 1'b0 ;
  assign n19428 = n4806 ^ n2429 ^ 1'b0 ;
  assign n19429 = n2920 & ~n19428 ;
  assign n19430 = n15192 ^ n14962 ^ 1'b0 ;
  assign n19431 = n19429 & ~n19430 ;
  assign n19432 = n2828 & ~n6058 ;
  assign n19433 = n82 & n19432 ;
  assign n19434 = n19433 ^ n14784 ^ 1'b0 ;
  assign n19435 = n19434 ^ n1380 ^ 1'b0 ;
  assign n19436 = n17530 ^ n8975 ^ n6262 ;
  assign n19437 = n873 | n18389 ;
  assign n19438 = n1009 & ~n19437 ;
  assign n19439 = ( n13486 & n16527 ) | ( n13486 & ~n19438 ) | ( n16527 & ~n19438 ) ;
  assign n19440 = ~n19436 & n19439 ;
  assign n19441 = n19440 ^ n15949 ^ 1'b0 ;
  assign n19442 = n11781 ^ n8508 ^ 1'b0 ;
  assign n19443 = n17346 | n19442 ;
  assign n19444 = x3 & n19443 ;
  assign n19445 = n5880 & n11045 ;
  assign n19446 = n19445 ^ n13325 ^ 1'b0 ;
  assign n19447 = n44 & n5692 ;
  assign n19448 = ~n17378 & n19447 ;
  assign n19449 = n230 | n4058 ;
  assign n19450 = n9799 | n19449 ;
  assign n19451 = n19450 ^ n10063 ^ 1'b0 ;
  assign n19452 = n13909 ^ n2047 ^ 1'b0 ;
  assign n19453 = n2523 & n19452 ;
  assign n19454 = n19453 ^ n6302 ^ 1'b0 ;
  assign n19455 = ~n4615 & n19454 ;
  assign n19458 = n8070 ^ n3199 ^ 1'b0 ;
  assign n19456 = n13854 ^ n4217 ^ 1'b0 ;
  assign n19457 = n6255 | n19456 ;
  assign n19459 = n19458 ^ n19457 ^ 1'b0 ;
  assign n19460 = n19455 & ~n19459 ;
  assign n19461 = ~n12765 & n19460 ;
  assign n19462 = n890 | n7659 ;
  assign n19463 = n12991 | n19462 ;
  assign n19464 = n2589 & n19463 ;
  assign n19465 = n19464 ^ n4574 ^ 1'b0 ;
  assign n19466 = n101 | n19465 ;
  assign n19467 = n19466 ^ n15376 ^ 1'b0 ;
  assign n19468 = n12248 ^ n2436 ^ 1'b0 ;
  assign n19469 = n13707 ^ n12204 ^ 1'b0 ;
  assign n19470 = n2612 & n19469 ;
  assign n19471 = n6402 | n6883 ;
  assign n19472 = n19471 ^ n15103 ^ 1'b0 ;
  assign n19475 = n11498 ^ n44 ^ 1'b0 ;
  assign n19476 = n16865 | n19475 ;
  assign n19473 = n117 | n6010 ;
  assign n19474 = n8625 & n19473 ;
  assign n19477 = n19476 ^ n19474 ^ 1'b0 ;
  assign n19478 = n5090 ^ n222 ^ 1'b0 ;
  assign n19479 = ( ~n1965 & n5110 ) | ( ~n1965 & n6753 ) | ( n5110 & n6753 ) ;
  assign n19480 = n19479 ^ n16663 ^ 1'b0 ;
  assign n19481 = n3833 ^ n2156 ^ 1'b0 ;
  assign n19482 = n1630 | n19481 ;
  assign n19483 = n19482 ^ n2556 ^ 1'b0 ;
  assign n19484 = n7287 & ~n18602 ;
  assign n19485 = n19484 ^ n12041 ^ 1'b0 ;
  assign n19486 = n12931 ^ n5782 ^ 1'b0 ;
  assign n19487 = n19485 & n19486 ;
  assign n19488 = n2004 & ~n5883 ;
  assign n19489 = ~n9345 & n19488 ;
  assign n19490 = n6440 ^ n2246 ^ 1'b0 ;
  assign n19491 = n3294 & n19490 ;
  assign n19492 = n10568 & ~n19491 ;
  assign n19493 = n19492 ^ n14738 ^ 1'b0 ;
  assign n19494 = n9566 ^ n5348 ^ n4463 ;
  assign n19495 = n8532 | n9796 ;
  assign n19496 = n19495 ^ n3578 ^ 1'b0 ;
  assign n19497 = ~n12271 & n15600 ;
  assign n19498 = n11152 & ~n19497 ;
  assign n19499 = n19498 ^ n8457 ^ 1'b0 ;
  assign n19504 = n590 & ~n5048 ;
  assign n19505 = ~n18136 & n19504 ;
  assign n19500 = ~n411 & n5919 ;
  assign n19501 = ~n7147 & n19500 ;
  assign n19502 = n15677 ^ n8509 ^ 1'b0 ;
  assign n19503 = n19501 | n19502 ;
  assign n19506 = n19505 ^ n19503 ^ n10527 ;
  assign n19507 = x0 & n7190 ;
  assign n19508 = n459 & n1231 ;
  assign n19509 = n12599 & n19508 ;
  assign n19510 = n19509 ^ n263 ^ 1'b0 ;
  assign n19511 = n9680 | n12436 ;
  assign n19512 = n19511 ^ n16650 ^ 1'b0 ;
  assign n19513 = n18929 | n19512 ;
  assign n19514 = n3818 & ~n17564 ;
  assign n19515 = n19514 ^ n10874 ^ 1'b0 ;
  assign n19517 = n6334 | n7081 ;
  assign n19518 = n19517 ^ n1448 ^ 1'b0 ;
  assign n19519 = n19518 ^ n11019 ^ 1'b0 ;
  assign n19520 = n965 & ~n19519 ;
  assign n19516 = ~n5986 & n13522 ;
  assign n19521 = n19520 ^ n19516 ^ 1'b0 ;
  assign n19522 = n15208 ^ n11111 ^ 1'b0 ;
  assign n19523 = ~n3134 & n19522 ;
  assign n19524 = x0 & n1500 ;
  assign n19525 = n2048 & ~n7128 ;
  assign n19526 = ( n8998 & n11051 ) | ( n8998 & ~n15690 ) | ( n11051 & ~n15690 ) ;
  assign n19527 = n19526 ^ n18494 ^ 1'b0 ;
  assign n19528 = ( ~n15208 & n19525 ) | ( ~n15208 & n19527 ) | ( n19525 & n19527 ) ;
  assign n19529 = n11915 ^ n7608 ^ 1'b0 ;
  assign n19530 = n1677 ^ n1001 ^ 1'b0 ;
  assign n19531 = n19530 ^ n8692 ^ 1'b0 ;
  assign n19532 = n19529 | n19531 ;
  assign n19536 = n3007 ^ n2443 ^ 1'b0 ;
  assign n19533 = n9224 ^ n5973 ^ n3753 ;
  assign n19534 = n8500 & ~n19533 ;
  assign n19535 = n19534 ^ n3983 ^ 1'b0 ;
  assign n19537 = n19536 ^ n19535 ^ 1'b0 ;
  assign n19538 = n16594 & ~n19537 ;
  assign n19539 = ( n4378 & ~n5077 ) | ( n4378 & n17994 ) | ( ~n5077 & n17994 ) ;
  assign n19540 = n19539 ^ n11428 ^ 1'b0 ;
  assign n19541 = n19538 & n19540 ;
  assign n19542 = n7738 ^ n491 ^ 1'b0 ;
  assign n19543 = n19541 & n19542 ;
  assign n19544 = n2209 ^ n806 ^ 1'b0 ;
  assign n19545 = n19544 ^ n14345 ^ n879 ;
  assign n19546 = n19545 ^ n11867 ^ 1'b0 ;
  assign n19547 = n67 & n19546 ;
  assign n19548 = n2958 & ~n4240 ;
  assign n19549 = ~n3119 & n5159 ;
  assign n19550 = n8016 ^ n6609 ^ n5791 ;
  assign n19551 = n19549 | n19550 ;
  assign n19552 = n9312 ^ n4660 ^ 1'b0 ;
  assign n19553 = n5531 & n19552 ;
  assign n19554 = n19553 ^ n10999 ^ 1'b0 ;
  assign n19555 = ~n10597 & n19554 ;
  assign n19557 = n360 | n797 ;
  assign n19558 = n5268 & ~n19557 ;
  assign n19556 = n5169 | n5732 ;
  assign n19559 = n19558 ^ n19556 ^ 1'b0 ;
  assign n19562 = n54 & ~n1064 ;
  assign n19563 = n11967 | n19562 ;
  assign n19564 = n19563 ^ n11424 ^ 1'b0 ;
  assign n19560 = n4704 ^ n2686 ^ 1'b0 ;
  assign n19561 = n19560 ^ n17131 ^ 1'b0 ;
  assign n19565 = n19564 ^ n19561 ^ n16730 ;
  assign n19566 = n11003 ^ n411 ^ 1'b0 ;
  assign n19567 = n7357 & n19566 ;
  assign n19568 = ( n5969 & ~n6623 ) | ( n5969 & n12821 ) | ( ~n6623 & n12821 ) ;
  assign n19569 = n1160 & ~n8907 ;
  assign n19570 = n19569 ^ n9532 ^ n5694 ;
  assign n19571 = n1861 & n9332 ;
  assign n19572 = n19571 ^ n5567 ^ 1'b0 ;
  assign n19573 = n19570 & n19572 ;
  assign n19574 = ~n3508 & n19573 ;
  assign n19575 = ( ~n2558 & n5290 ) | ( ~n2558 & n9683 ) | ( n5290 & n9683 ) ;
  assign n19576 = n3256 & ~n19575 ;
  assign n19577 = n19574 & n19576 ;
  assign n19578 = ( n10444 & n19568 ) | ( n10444 & n19577 ) | ( n19568 & n19577 ) ;
  assign n19579 = ~n17897 & n19315 ;
  assign n19581 = n67 | n4411 ;
  assign n19582 = n67 & ~n19581 ;
  assign n19583 = n13621 | n19582 ;
  assign n19584 = n19582 & ~n19583 ;
  assign n19585 = n13237 & ~n19584 ;
  assign n19586 = ~n13237 & n19585 ;
  assign n19580 = ( n1329 & n9141 ) | ( n1329 & n13107 ) | ( n9141 & n13107 ) ;
  assign n19587 = n19586 ^ n19580 ^ n11618 ;
  assign n19588 = n99 & n3825 ;
  assign n19589 = n18631 ^ n7357 ^ 1'b0 ;
  assign n19590 = n764 & ~n19589 ;
  assign n19591 = n2797 & ~n19590 ;
  assign n19592 = n5006 & n9341 ;
  assign n19593 = n4713 ^ n1247 ^ 1'b0 ;
  assign n19594 = n14338 ^ n6278 ^ 1'b0 ;
  assign n19595 = n10477 ^ n6611 ^ 1'b0 ;
  assign n19596 = n242 | n19595 ;
  assign n19597 = n19596 ^ n14338 ^ 1'b0 ;
  assign n19602 = ~n1945 & n4503 ;
  assign n19603 = n9208 | n19602 ;
  assign n19604 = n19603 ^ n11658 ^ 1'b0 ;
  assign n19598 = n5486 & ~n8938 ;
  assign n19599 = ( n3361 & n6168 ) | ( n3361 & n7507 ) | ( n6168 & n7507 ) ;
  assign n19600 = ~n5279 & n19599 ;
  assign n19601 = ~n19598 & n19600 ;
  assign n19605 = n19604 ^ n19601 ^ 1'b0 ;
  assign n19606 = n4703 & n8995 ;
  assign n19607 = ( n3308 & ~n12081 ) | ( n3308 & n19606 ) | ( ~n12081 & n19606 ) ;
  assign n19608 = n9172 ^ n5169 ^ 1'b0 ;
  assign n19609 = n17957 & n19608 ;
  assign n19610 = n18612 & n19609 ;
  assign n19611 = n17761 ^ n13580 ^ 1'b0 ;
  assign n19612 = n1137 | n8569 ;
  assign n19613 = n6596 | n19612 ;
  assign n19614 = n3883 & n19613 ;
  assign n19615 = ( n14571 & n19372 ) | ( n14571 & n19614 ) | ( n19372 & n19614 ) ;
  assign n19616 = n6648 ^ n5310 ^ 1'b0 ;
  assign n19617 = n19616 ^ n8597 ^ 1'b0 ;
  assign n19618 = ~n13188 & n19617 ;
  assign n19619 = n9721 | n19618 ;
  assign n19620 = n15007 ^ n7136 ^ 1'b0 ;
  assign n19621 = n19620 ^ n7402 ^ 1'b0 ;
  assign n19622 = n19621 ^ n13567 ^ 1'b0 ;
  assign n19623 = n12687 | n19622 ;
  assign n19624 = n13258 ^ n2810 ^ 1'b0 ;
  assign n19625 = n3195 & n19624 ;
  assign n19626 = n7554 | n9984 ;
  assign n19627 = n9984 & ~n19626 ;
  assign n19628 = n6643 | n19627 ;
  assign n19629 = n6643 & ~n19628 ;
  assign n19630 = ~n269 & n3713 ;
  assign n19631 = n3122 | n19630 ;
  assign n19632 = n19631 ^ n16079 ^ 1'b0 ;
  assign n19633 = n6551 & ~n6630 ;
  assign n19634 = ~n813 & n7730 ;
  assign n19635 = n13546 ^ n5281 ^ 1'b0 ;
  assign n19636 = ~n4544 & n19635 ;
  assign n19637 = n9148 & n19636 ;
  assign n19638 = n19637 ^ n14766 ^ 1'b0 ;
  assign n19639 = n3312 ^ n2196 ^ 1'b0 ;
  assign n19640 = n19639 ^ n14197 ^ 1'b0 ;
  assign n19641 = n1382 & n19640 ;
  assign n19642 = n9098 & n19641 ;
  assign n19643 = n13972 ^ n2725 ^ 1'b0 ;
  assign n19644 = n3789 & ~n19643 ;
  assign n19645 = ( ~n7350 & n12404 ) | ( ~n7350 & n19644 ) | ( n12404 & n19644 ) ;
  assign n19646 = n16954 ^ n14201 ^ n5852 ;
  assign n19647 = n6958 & n19646 ;
  assign n19648 = ~n19645 & n19647 ;
  assign n19649 = ~n734 & n3370 ;
  assign n19650 = ~n10569 & n19649 ;
  assign n19651 = n4673 | n19650 ;
  assign n19652 = n19651 ^ n2234 ^ 1'b0 ;
  assign n19653 = n15014 ^ n3079 ^ n2297 ;
  assign n19654 = ( ~n5466 & n6821 ) | ( ~n5466 & n19653 ) | ( n6821 & n19653 ) ;
  assign n19655 = n19654 ^ n8625 ^ n1139 ;
  assign n19656 = n1787 | n5564 ;
  assign n19664 = n10183 & ~n10559 ;
  assign n19657 = ~n5949 & n6816 ;
  assign n19658 = n397 ^ n63 ^ 1'b0 ;
  assign n19659 = n4044 | n13500 ;
  assign n19660 = n19658 & ~n19659 ;
  assign n19661 = n8390 | n19660 ;
  assign n19662 = n19657 | n19661 ;
  assign n19663 = ~n1213 & n19662 ;
  assign n19665 = n19664 ^ n19663 ^ 1'b0 ;
  assign n19666 = n12952 & n19665 ;
  assign n19667 = ~n3308 & n18381 ;
  assign n19668 = n2879 & n15100 ;
  assign n19669 = n5715 & n9833 ;
  assign n19670 = ~n3180 & n19669 ;
  assign n19671 = n1151 & ~n4987 ;
  assign n19672 = n19671 ^ n2736 ^ 1'b0 ;
  assign n19673 = n9776 | n19672 ;
  assign n19674 = n5176 | n18039 ;
  assign n19675 = n220 & ~n19674 ;
  assign n19676 = n1666 ^ n517 ^ 1'b0 ;
  assign n19677 = ( n1946 & n10488 ) | ( n1946 & n19676 ) | ( n10488 & n19676 ) ;
  assign n19678 = ~n8597 & n19677 ;
  assign n19679 = n18077 & n19678 ;
  assign n19680 = n2523 ^ n974 ^ 1'b0 ;
  assign n19681 = ~n5449 & n19680 ;
  assign n19682 = n19681 ^ n18971 ^ 1'b0 ;
  assign n19683 = n7462 | n19682 ;
  assign n19684 = n9039 & n19683 ;
  assign n19694 = n1502 ^ n1457 ^ 1'b0 ;
  assign n19695 = n2832 | n19694 ;
  assign n19696 = n19695 ^ n11302 ^ 1'b0 ;
  assign n19685 = ( n2729 & n4591 ) | ( n2729 & n7728 ) | ( n4591 & n7728 ) ;
  assign n19686 = ~n3304 & n15308 ;
  assign n19687 = n19686 ^ n5254 ^ 1'b0 ;
  assign n19688 = n3540 | n6116 ;
  assign n19689 = n19688 ^ n2869 ^ 1'b0 ;
  assign n19690 = n19689 ^ n6435 ^ 1'b0 ;
  assign n19691 = n13221 & n19690 ;
  assign n19692 = n19687 & n19691 ;
  assign n19693 = ~n19685 & n19692 ;
  assign n19697 = n19696 ^ n19693 ^ 1'b0 ;
  assign n19698 = n5686 ^ n3430 ^ 1'b0 ;
  assign n19699 = n780 & ~n19698 ;
  assign n19700 = n19699 ^ n14285 ^ 1'b0 ;
  assign n19702 = n14850 ^ n4147 ^ 1'b0 ;
  assign n19703 = n1489 & n19702 ;
  assign n19701 = n7312 & ~n14124 ;
  assign n19704 = n19703 ^ n19701 ^ 1'b0 ;
  assign n19705 = ~n656 & n19704 ;
  assign n19706 = n12293 & n13442 ;
  assign n19707 = n1348 & n1623 ;
  assign n19708 = n5936 & n19707 ;
  assign n19709 = n4271 | n19708 ;
  assign n19710 = n9857 ^ n9507 ^ 1'b0 ;
  assign n19711 = ~n8215 & n19710 ;
  assign n19712 = n19711 ^ n4287 ^ 1'b0 ;
  assign n19713 = n8508 & ~n18032 ;
  assign n19714 = n6142 ^ n3038 ^ n2408 ;
  assign n19715 = n15821 & ~n19714 ;
  assign n19716 = n4404 ^ n2170 ^ n1461 ;
  assign n19717 = ~n5627 & n19716 ;
  assign n19718 = n8713 & n19717 ;
  assign n19719 = n19718 ^ n4485 ^ 1'b0 ;
  assign n19720 = n3108 & n19277 ;
  assign n19721 = ~n10393 & n19720 ;
  assign n19722 = n9110 ^ n1280 ^ 1'b0 ;
  assign n19723 = ~n2655 & n19722 ;
  assign n19724 = n118 & n12782 ;
  assign n19725 = ~n19723 & n19724 ;
  assign n19726 = n19721 | n19725 ;
  assign n19727 = n9004 ^ n6647 ^ 1'b0 ;
  assign n19728 = n3202 & n15364 ;
  assign n19729 = n15189 & n19728 ;
  assign n19730 = n19729 ^ n11247 ^ 1'b0 ;
  assign n19731 = ~n5048 & n19730 ;
  assign n19732 = ~n19727 & n19731 ;
  assign n19733 = n18237 ^ n12827 ^ n2037 ;
  assign n19734 = ~n4252 & n13046 ;
  assign n19735 = n19347 ^ n14211 ^ 1'b0 ;
  assign n19736 = n14766 & ~n19735 ;
  assign n19737 = n19736 ^ n2556 ^ 1'b0 ;
  assign n19738 = n2083 & n8654 ;
  assign n19739 = n19738 ^ n5691 ^ 1'b0 ;
  assign n19745 = ( n4931 & ~n12498 ) | ( n4931 & n17326 ) | ( ~n12498 & n17326 ) ;
  assign n19740 = n14978 ^ n1878 ^ 1'b0 ;
  assign n19741 = n4195 & n19740 ;
  assign n19742 = ~n2237 & n12042 ;
  assign n19743 = ( n19092 & n19741 ) | ( n19092 & ~n19742 ) | ( n19741 & ~n19742 ) ;
  assign n19744 = n19743 ^ n8020 ^ 1'b0 ;
  assign n19746 = n19745 ^ n19744 ^ 1'b0 ;
  assign n19747 = ~n7395 & n19746 ;
  assign n19748 = n19747 ^ n10958 ^ 1'b0 ;
  assign n19749 = n15607 ^ n11901 ^ 1'b0 ;
  assign n19750 = n9311 ^ n1642 ^ n1082 ;
  assign n19751 = n15614 ^ n9115 ^ 1'b0 ;
  assign n19752 = ~n210 & n19751 ;
  assign n19753 = ~n1932 & n19752 ;
  assign n19754 = n19753 ^ n10258 ^ 1'b0 ;
  assign n19755 = ~n4684 & n19754 ;
  assign n19756 = n19755 ^ n18067 ^ 1'b0 ;
  assign n19757 = n3317 & n6595 ;
  assign n19758 = n19757 ^ n5302 ^ 1'b0 ;
  assign n19759 = n3482 & ~n5131 ;
  assign n19760 = n19759 ^ n12549 ^ 1'b0 ;
  assign n19761 = n16899 & ~n19760 ;
  assign n19762 = n13179 & n19761 ;
  assign n19763 = n19758 & n19762 ;
  assign n19764 = n5128 & ~n6495 ;
  assign n19765 = n19764 ^ n2274 ^ 1'b0 ;
  assign n19766 = n19765 ^ n9681 ^ 1'b0 ;
  assign n19767 = ~n7182 & n19766 ;
  assign n19768 = n2652 & ~n4313 ;
  assign n19769 = n19768 ^ n5354 ^ 1'b0 ;
  assign n19770 = n19769 ^ n7248 ^ 1'b0 ;
  assign n19771 = n19770 ^ n17133 ^ 1'b0 ;
  assign n19772 = n3061 & n10301 ;
  assign n19775 = n3892 ^ n1031 ^ 1'b0 ;
  assign n19773 = ~n3737 & n19625 ;
  assign n19774 = n19773 ^ n16573 ^ 1'b0 ;
  assign n19776 = n19775 ^ n19774 ^ 1'b0 ;
  assign n19777 = n19220 ^ n3521 ^ x3 ;
  assign n19778 = n10124 ^ n6890 ^ 1'b0 ;
  assign n19779 = n19778 ^ n3945 ^ 1'b0 ;
  assign n19780 = ~n19777 & n19779 ;
  assign n19781 = n19780 ^ n6922 ^ 1'b0 ;
  assign n19782 = ( ~n5651 & n8701 ) | ( ~n5651 & n10541 ) | ( n8701 & n10541 ) ;
  assign n19783 = n7836 & n9929 ;
  assign n19784 = n18637 ^ n9402 ^ 1'b0 ;
  assign n19785 = n149 & ~n19784 ;
  assign n19787 = ( n982 & n7927 ) | ( n982 & ~n12005 ) | ( n7927 & ~n12005 ) ;
  assign n19786 = n18283 & ~n19529 ;
  assign n19788 = n19787 ^ n19786 ^ 1'b0 ;
  assign n19789 = n6273 ^ n5237 ^ 1'b0 ;
  assign n19790 = ~n40 & n19789 ;
  assign n19791 = ~n3855 & n5175 ;
  assign n19792 = ~n3870 & n19791 ;
  assign n19793 = n3158 & ~n5864 ;
  assign n19794 = ~n7089 & n19793 ;
  assign n19795 = n19794 ^ n12418 ^ 1'b0 ;
  assign n19796 = n2080 | n3953 ;
  assign n19797 = ( ~n2960 & n6135 ) | ( ~n2960 & n17534 ) | ( n6135 & n17534 ) ;
  assign n19798 = ( n2733 & n19796 ) | ( n2733 & ~n19797 ) | ( n19796 & ~n19797 ) ;
  assign n19799 = n8483 & ~n19798 ;
  assign n19800 = ( n5415 & n7498 ) | ( n5415 & n19799 ) | ( n7498 & n19799 ) ;
  assign n19801 = ~n989 & n11231 ;
  assign n19802 = n19801 ^ n3131 ^ 1'b0 ;
  assign n19803 = n15194 & n19802 ;
  assign n19804 = n7590 & ~n11132 ;
  assign n19805 = n19804 ^ n4455 ^ 1'b0 ;
  assign n19806 = n6612 & ~n13943 ;
  assign n19807 = n19806 ^ n3824 ^ 1'b0 ;
  assign n19808 = n19807 ^ n12439 ^ 1'b0 ;
  assign n19809 = n11809 & ~n19808 ;
  assign n19810 = n19809 ^ n3620 ^ 1'b0 ;
  assign n19811 = ~n12575 & n19810 ;
  assign n19812 = n15076 ^ n7077 ^ n4262 ;
  assign n19813 = n91 & ~n2588 ;
  assign n19814 = n8438 ^ n4298 ^ 1'b0 ;
  assign n19815 = n9821 | n19814 ;
  assign n19816 = n9363 & n19815 ;
  assign n19817 = n1630 & n19816 ;
  assign n19818 = n2129 & ~n3722 ;
  assign n19819 = n10441 & n19818 ;
  assign n19823 = ~n15382 & n18262 ;
  assign n19820 = n8821 ^ n2492 ^ 1'b0 ;
  assign n19821 = n12101 & n19820 ;
  assign n19822 = n12145 & n19821 ;
  assign n19824 = n19823 ^ n19822 ^ 1'b0 ;
  assign n19825 = n11664 ^ n1684 ^ n1305 ;
  assign n19826 = n19825 ^ n8542 ^ 1'b0 ;
  assign n19827 = n3039 ^ n923 ^ 1'b0 ;
  assign n19828 = n19826 & n19827 ;
  assign n19829 = ~n8727 & n16762 ;
  assign n19832 = n1240 | n10504 ;
  assign n19833 = n19832 ^ n7802 ^ 1'b0 ;
  assign n19830 = n10345 & n18486 ;
  assign n19831 = n6941 & n19830 ;
  assign n19834 = n19833 ^ n19831 ^ 1'b0 ;
  assign n19835 = n12478 | n19834 ;
  assign n19836 = n11325 ^ n8801 ^ 1'b0 ;
  assign n19837 = n6792 & n19836 ;
  assign n19838 = n3655 & n19837 ;
  assign n19839 = ~n178 & n19838 ;
  assign n19840 = ( n3106 & n4982 ) | ( n3106 & n14716 ) | ( n4982 & n14716 ) ;
  assign n19841 = n14813 & ~n15588 ;
  assign n19842 = n19841 ^ n1888 ^ 1'b0 ;
  assign n19843 = n4126 ^ n45 ^ 1'b0 ;
  assign n19844 = n13680 ^ n5496 ^ 1'b0 ;
  assign n19845 = n19844 ^ n3260 ^ 1'b0 ;
  assign n19846 = ~n7071 & n12753 ;
  assign n19847 = n19845 | n19846 ;
  assign n19848 = n19335 ^ n6004 ^ n839 ;
  assign n19849 = ~n383 & n18641 ;
  assign n19850 = n19849 ^ n7327 ^ 1'b0 ;
  assign n19851 = n2102 | n3184 ;
  assign n19852 = n575 | n19851 ;
  assign n19853 = ~n1290 & n19852 ;
  assign n19854 = n11690 & n19853 ;
  assign n19855 = n10452 ^ n6564 ^ 1'b0 ;
  assign n19856 = ( n9792 & ~n19854 ) | ( n9792 & n19855 ) | ( ~n19854 & n19855 ) ;
  assign n19857 = n3040 & n19856 ;
  assign n19858 = n191 & n8950 ;
  assign n19859 = n19858 ^ n7363 ^ 1'b0 ;
  assign n19860 = n10291 & n19859 ;
  assign n19861 = n1076 | n5466 ;
  assign n19862 = n3313 | n6161 ;
  assign n19863 = n19745 ^ n15823 ^ 1'b0 ;
  assign n19864 = ~n1638 & n19863 ;
  assign n19865 = ~n17078 & n19864 ;
  assign n19867 = n3787 & n4495 ;
  assign n19868 = n10270 & n19867 ;
  assign n19866 = n543 & n11708 ;
  assign n19869 = n19868 ^ n19866 ^ 1'b0 ;
  assign n19870 = n8348 | n8644 ;
  assign n19871 = n7386 & n19870 ;
  assign n19872 = n16790 ^ n3156 ^ n1320 ;
  assign n19873 = ~n1367 & n19872 ;
  assign n19874 = ( n14475 & n19871 ) | ( n14475 & n19873 ) | ( n19871 & n19873 ) ;
  assign n19875 = n5774 | n7017 ;
  assign n19876 = n19875 ^ n18539 ^ 1'b0 ;
  assign n19877 = ( ~n5037 & n10059 ) | ( ~n5037 & n10777 ) | ( n10059 & n10777 ) ;
  assign n19878 = n7832 & ~n10665 ;
  assign n19879 = ( ~n16798 & n19877 ) | ( ~n16798 & n19878 ) | ( n19877 & n19878 ) ;
  assign n19880 = n6904 | n10073 ;
  assign n19881 = n19880 ^ n5020 ^ 1'b0 ;
  assign n19882 = n16935 ^ n14273 ^ 1'b0 ;
  assign n19883 = ~n7190 & n19882 ;
  assign n19884 = n9986 ^ n1412 ^ 1'b0 ;
  assign n19885 = n1563 & ~n2408 ;
  assign n19886 = n19885 ^ n16557 ^ 1'b0 ;
  assign n19887 = n19886 ^ n1770 ^ 1'b0 ;
  assign n19888 = n10941 | n19887 ;
  assign n19889 = n19884 | n19888 ;
  assign n19890 = n2898 ^ n1472 ^ 1'b0 ;
  assign n19891 = ~n126 & n2650 ;
  assign n19892 = n19891 ^ n3581 ^ 1'b0 ;
  assign n19894 = n11592 ^ n3246 ^ 1'b0 ;
  assign n19895 = ~n2665 & n19894 ;
  assign n19893 = n5458 ^ n5149 ^ 1'b0 ;
  assign n19896 = n19895 ^ n19893 ^ 1'b0 ;
  assign n19897 = n14816 | n19896 ;
  assign n19898 = n17873 ^ n3410 ^ 1'b0 ;
  assign n19899 = n9036 ^ n4543 ^ 1'b0 ;
  assign n19900 = n4735 & n4884 ;
  assign n19901 = n11766 ^ n1623 ^ 1'b0 ;
  assign n19902 = n19900 & n19901 ;
  assign n19903 = n15373 ^ n12281 ^ n1315 ;
  assign n19904 = n249 & ~n19903 ;
  assign n19905 = n19902 | n19904 ;
  assign n19906 = ( n6152 & n13167 ) | ( n6152 & ~n17718 ) | ( n13167 & ~n17718 ) ;
  assign n19907 = n2483 & n9757 ;
  assign n19908 = ~n14048 & n19907 ;
  assign n19909 = ~n19906 & n19908 ;
  assign n19910 = n6848 & ~n19909 ;
  assign n19911 = n19910 ^ n15226 ^ 1'b0 ;
  assign n19912 = ~n3988 & n5415 ;
  assign n19913 = n19912 ^ n7976 ^ 1'b0 ;
  assign n19914 = ~n11301 & n16331 ;
  assign n19915 = n19914 ^ n6199 ^ 1'b0 ;
  assign n19916 = ~n734 & n4983 ;
  assign n19917 = ~n1647 & n19916 ;
  assign n19920 = ~n3313 & n4134 ;
  assign n19918 = n8426 | n16234 ;
  assign n19919 = n7130 | n19918 ;
  assign n19921 = n19920 ^ n19919 ^ 1'b0 ;
  assign n19922 = ~n19917 & n19921 ;
  assign n19923 = n445 & n2677 ;
  assign n19924 = ( ~n7147 & n7468 ) | ( ~n7147 & n19923 ) | ( n7468 & n19923 ) ;
  assign n19925 = ~n2658 & n10826 ;
  assign n19926 = n16890 | n19925 ;
  assign n19927 = n17903 | n19926 ;
  assign n19930 = n5725 & n14475 ;
  assign n19928 = n10488 & ~n17455 ;
  assign n19929 = ( n57 & ~n13876 ) | ( n57 & n19928 ) | ( ~n13876 & n19928 ) ;
  assign n19931 = n19930 ^ n19929 ^ n1026 ;
  assign n19934 = n2370 & ~n13391 ;
  assign n19935 = ~n5921 & n19934 ;
  assign n19932 = n10393 ^ n432 ^ 1'b0 ;
  assign n19933 = n784 & ~n19932 ;
  assign n19936 = n19935 ^ n19933 ^ n14175 ;
  assign n19937 = n15574 & n19936 ;
  assign n19938 = n19931 & n19937 ;
  assign n19939 = n9208 ^ n2581 ^ 1'b0 ;
  assign n19940 = n19312 & ~n19939 ;
  assign n19941 = ( ~n8962 & n11910 ) | ( ~n8962 & n19940 ) | ( n11910 & n19940 ) ;
  assign n19942 = n4258 | n19941 ;
  assign n19943 = n1945 & ~n19942 ;
  assign n19945 = n9506 ^ n51 ^ 1'b0 ;
  assign n19946 = n3477 & n19945 ;
  assign n19947 = ~n5837 & n19946 ;
  assign n19944 = n19858 ^ n3189 ^ 1'b0 ;
  assign n19948 = n19947 ^ n19944 ^ n17116 ;
  assign n19949 = n6546 & n9228 ;
  assign n19950 = n19949 ^ n3870 ^ 1'b0 ;
  assign n19951 = n12220 ^ n6568 ^ 1'b0 ;
  assign n19952 = ~n12482 & n19951 ;
  assign n19953 = n19952 ^ n9962 ^ 1'b0 ;
  assign n19954 = n18921 | n19953 ;
  assign n19955 = n5891 ^ n3784 ^ 1'b0 ;
  assign n19956 = n4305 | n13766 ;
  assign n19957 = n19956 ^ n1824 ^ 1'b0 ;
  assign n19958 = ~n4602 & n9267 ;
  assign n19966 = ~n6766 & n15832 ;
  assign n19967 = n6890 & n19966 ;
  assign n19968 = n15401 & n19967 ;
  assign n19959 = n2552 ^ n496 ^ n490 ;
  assign n19960 = n19959 ^ n7342 ^ 1'b0 ;
  assign n19961 = n1013 | n19960 ;
  assign n19962 = n19961 ^ n13500 ^ 1'b0 ;
  assign n19963 = n1108 & ~n19962 ;
  assign n19964 = ~n8958 & n19963 ;
  assign n19965 = n13642 & n19964 ;
  assign n19969 = n19968 ^ n19965 ^ 1'b0 ;
  assign n19971 = n4408 & n17106 ;
  assign n19970 = n4247 | n15729 ;
  assign n19972 = n19971 ^ n19970 ^ 1'b0 ;
  assign n19973 = n11975 & n19972 ;
  assign n19974 = ( n218 & n2677 ) | ( n218 & n6128 ) | ( n2677 & n6128 ) ;
  assign n19975 = n19974 ^ n5898 ^ 1'b0 ;
  assign n19976 = n19973 & ~n19975 ;
  assign n19977 = n13972 & ~n17034 ;
  assign n19978 = n19977 ^ n9369 ^ 1'b0 ;
  assign n19979 = ( n2561 & ~n8978 ) | ( n2561 & n19978 ) | ( ~n8978 & n19978 ) ;
  assign n19980 = n16505 & n19979 ;
  assign n19981 = n10007 & n19980 ;
  assign n19982 = n2878 & ~n7322 ;
  assign n19983 = n15978 ^ n469 ^ 1'b0 ;
  assign n19984 = n19983 ^ n12008 ^ n779 ;
  assign n19985 = n9580 ^ n9322 ^ 1'b0 ;
  assign n19986 = n12403 & ~n19985 ;
  assign n19987 = n19354 ^ n10946 ^ 1'b0 ;
  assign n19988 = n19987 ^ n1804 ^ 1'b0 ;
  assign n19989 = ( ~n4637 & n19986 ) | ( ~n4637 & n19988 ) | ( n19986 & n19988 ) ;
  assign n19990 = ~n1201 & n2289 ;
  assign n19991 = n19990 ^ n10943 ^ 1'b0 ;
  assign n19992 = n7979 | n10850 ;
  assign n19993 = n2704 & ~n19992 ;
  assign n19994 = n5273 & ~n19993 ;
  assign n19995 = n2623 | n16228 ;
  assign n19996 = n510 & n14833 ;
  assign n19997 = ~n473 & n19996 ;
  assign n19998 = n4394 & n12591 ;
  assign n19999 = n18711 & n19998 ;
  assign n20000 = n19999 ^ n17653 ^ n426 ;
  assign n20001 = n524 | n6462 ;
  assign n20002 = n5012 | n10963 ;
  assign n20003 = ( ~n9813 & n13113 ) | ( ~n9813 & n17351 ) | ( n13113 & n17351 ) ;
  assign n20004 = n10836 | n20003 ;
  assign n20005 = n20002 & ~n20004 ;
  assign n20006 = n16781 | n17770 ;
  assign n20007 = n20006 ^ n6638 ^ 1'b0 ;
  assign n20008 = n7904 & ~n9998 ;
  assign n20012 = n4368 ^ n401 ^ 1'b0 ;
  assign n20013 = n2539 & n20012 ;
  assign n20009 = n3192 ^ n1612 ^ n168 ;
  assign n20010 = n20009 ^ n9909 ^ 1'b0 ;
  assign n20011 = ~n9029 & n20010 ;
  assign n20014 = n20013 ^ n20011 ^ n5400 ;
  assign n20015 = n20014 ^ n12484 ^ 1'b0 ;
  assign n20016 = n11123 | n20015 ;
  assign n20017 = n20008 & ~n20016 ;
  assign n20018 = n5437 ^ n1581 ^ 1'b0 ;
  assign n20021 = n7742 & ~n16876 ;
  assign n20019 = n1346 & n2346 ;
  assign n20020 = n2723 & n20019 ;
  assign n20022 = n20021 ^ n20020 ^ 1'b0 ;
  assign n20023 = ~n15753 & n20022 ;
  assign n20024 = n14930 & n20023 ;
  assign n20025 = n20024 ^ n16136 ^ 1'b0 ;
  assign n20026 = n4679 & ~n20025 ;
  assign n20027 = n5888 | n18109 ;
  assign n20028 = n20027 ^ n12601 ^ 1'b0 ;
  assign n20029 = n7332 ^ n6249 ^ 1'b0 ;
  assign n20030 = n20028 & ~n20029 ;
  assign n20031 = n9984 ^ n2766 ^ 1'b0 ;
  assign n20032 = n20031 ^ n15470 ^ 1'b0 ;
  assign n20033 = n1677 | n20032 ;
  assign n20034 = ~n20002 & n20033 ;
  assign n20035 = ( ~n5706 & n6126 ) | ( ~n5706 & n20034 ) | ( n6126 & n20034 ) ;
  assign n20036 = ( n4260 & n13467 ) | ( n4260 & ~n15246 ) | ( n13467 & ~n15246 ) ;
  assign n20037 = n17748 ^ n15996 ^ n9727 ;
  assign n20038 = n20036 & ~n20037 ;
  assign n20039 = n20038 ^ n18236 ^ 1'b0 ;
  assign n20040 = ~n374 & n3119 ;
  assign n20041 = n20040 ^ n378 ^ 1'b0 ;
  assign n20043 = n5212 & ~n11724 ;
  assign n20044 = n20043 ^ n11090 ^ 1'b0 ;
  assign n20042 = ~n3923 & n7366 ;
  assign n20045 = n20044 ^ n20042 ^ n11438 ;
  assign n20046 = n12355 ^ n8052 ^ 1'b0 ;
  assign n20047 = n187 & ~n15804 ;
  assign n20048 = n19698 ^ n191 ^ 1'b0 ;
  assign n20049 = n2692 | n6217 ;
  assign n20050 = ~n3751 & n4948 ;
  assign n20051 = ( n82 & ~n5408 ) | ( n82 & n20050 ) | ( ~n5408 & n20050 ) ;
  assign n20052 = n20049 & ~n20051 ;
  assign n20053 = n16047 ^ n9013 ^ 1'b0 ;
  assign n20054 = n20053 ^ n2691 ^ 1'b0 ;
  assign n20055 = n14296 | n20054 ;
  assign n20056 = n5504 | n8446 ;
  assign n20057 = n20056 ^ n3782 ^ 1'b0 ;
  assign n20058 = n2504 ^ n2325 ^ 1'b0 ;
  assign n20059 = ~n8179 & n20058 ;
  assign n20060 = n5866 & n20059 ;
  assign n20061 = n2441 & ~n4067 ;
  assign n20062 = n20061 ^ n12396 ^ 1'b0 ;
  assign n20063 = n20062 ^ n15267 ^ 1'b0 ;
  assign n20064 = n18681 | n20063 ;
  assign n20065 = n10657 & ~n15785 ;
  assign n20066 = n20065 ^ n8400 ^ 1'b0 ;
  assign n20067 = n20066 ^ n19084 ^ 1'b0 ;
  assign n20068 = n17511 ^ n13795 ^ 1'b0 ;
  assign n20069 = n20068 ^ n9524 ^ 1'b0 ;
  assign n20070 = ~n3916 & n15359 ;
  assign n20071 = n4475 & n7089 ;
  assign n20072 = n16372 & n20071 ;
  assign n20073 = n20072 ^ n12472 ^ 1'b0 ;
  assign n20074 = n20070 | n20073 ;
  assign n20075 = ~n5397 & n8976 ;
  assign n20076 = ~n714 & n3098 ;
  assign n20077 = ~n3359 & n20076 ;
  assign n20078 = n20077 ^ n14947 ^ n14110 ;
  assign n20079 = n650 | n4285 ;
  assign n20080 = n2684 & ~n3667 ;
  assign n20081 = n20079 & n20080 ;
  assign n20082 = n604 ^ n322 ^ 1'b0 ;
  assign n20083 = n15513 ^ n10800 ^ 1'b0 ;
  assign n20084 = n20083 ^ n1550 ^ 1'b0 ;
  assign n20085 = n20082 & ~n20084 ;
  assign n20086 = ~n5864 & n16833 ;
  assign n20087 = n14428 | n17019 ;
  assign n20088 = n2350 | n15801 ;
  assign n20089 = n341 | n20088 ;
  assign n20090 = n6533 & n20089 ;
  assign n20091 = n3048 & n20090 ;
  assign n20092 = n20091 ^ n1542 ^ 1'b0 ;
  assign n20093 = n20092 ^ n13707 ^ 1'b0 ;
  assign n20094 = n10968 & n20093 ;
  assign n20095 = ~n4563 & n15535 ;
  assign n20096 = n13923 ^ n9824 ^ 1'b0 ;
  assign n20097 = n20096 ^ n18739 ^ 1'b0 ;
  assign n20098 = n20097 ^ n13594 ^ 1'b0 ;
  assign n20099 = n9799 & n20098 ;
  assign n20100 = ~n12460 & n14169 ;
  assign n20101 = n20100 ^ n15720 ^ n13684 ;
  assign n20102 = n16011 & ~n18346 ;
  assign n20103 = n20102 ^ n8777 ^ 1'b0 ;
  assign n20104 = n4699 ^ n53 ^ 1'b0 ;
  assign n20105 = n5363 & n20104 ;
  assign n20106 = n20105 ^ n5004 ^ 1'b0 ;
  assign n20107 = n18950 ^ n6074 ^ 1'b0 ;
  assign n20108 = n9448 ^ n3285 ^ 1'b0 ;
  assign n20109 = ~n4887 & n20108 ;
  assign n20110 = n16126 ^ n6743 ^ 1'b0 ;
  assign n20111 = ~n6326 & n6612 ;
  assign n20112 = n854 & n17736 ;
  assign n20113 = n20112 ^ n3277 ^ 1'b0 ;
  assign n20114 = n12066 | n20113 ;
  assign n20115 = n20114 ^ n645 ^ 1'b0 ;
  assign n20116 = n19830 & n20115 ;
  assign n20117 = ~n8807 & n20116 ;
  assign n20118 = n20111 & n20117 ;
  assign n20119 = n14848 ^ n8674 ^ 1'b0 ;
  assign n20120 = ~n3345 & n20119 ;
  assign n20121 = n20120 ^ n12036 ^ 1'b0 ;
  assign n20122 = ~n517 & n10718 ;
  assign n20123 = n1693 | n5156 ;
  assign n20124 = n20123 ^ n6380 ^ 1'b0 ;
  assign n20125 = ( n2391 & n17380 ) | ( n2391 & ~n20124 ) | ( n17380 & ~n20124 ) ;
  assign n20126 = n13037 ^ n11385 ^ 1'b0 ;
  assign n20127 = ~n8441 & n20126 ;
  assign n20128 = n2825 | n11704 ;
  assign n20129 = n3824 & ~n9373 ;
  assign n20130 = n557 & ~n3192 ;
  assign n20131 = n20129 & ~n20130 ;
  assign n20132 = n12460 & n20131 ;
  assign n20133 = n9439 ^ n3085 ^ 1'b0 ;
  assign n20134 = n19483 | n20133 ;
  assign n20135 = n20134 ^ n12520 ^ n7581 ;
  assign n20136 = n17057 ^ n7580 ^ 1'b0 ;
  assign n20137 = n16318 | n20136 ;
  assign n20138 = n319 | n8726 ;
  assign n20139 = n20138 ^ n13488 ^ 1'b0 ;
  assign n20140 = n1616 & n14479 ;
  assign n20141 = n20140 ^ n3833 ^ 1'b0 ;
  assign n20142 = n15395 & n20141 ;
  assign n20143 = n20142 ^ n4411 ^ 1'b0 ;
  assign n20144 = n4743 & n20143 ;
  assign n20145 = n10890 ^ n1099 ^ 1'b0 ;
  assign n20146 = n10088 & n20145 ;
  assign n20147 = n5785 ^ n2674 ^ 1'b0 ;
  assign n20148 = n8497 & n9727 ;
  assign n20149 = n194 | n20148 ;
  assign n20150 = n7428 ^ n7020 ^ 1'b0 ;
  assign n20151 = n7500 | n20150 ;
  assign n20152 = n11341 & n15969 ;
  assign n20153 = ~n19877 & n20152 ;
  assign n20154 = n1129 ^ n760 ^ 1'b0 ;
  assign n20155 = n4330 & ~n20154 ;
  assign n20156 = n20155 ^ n6976 ^ 1'b0 ;
  assign n20157 = ~n3273 & n20156 ;
  assign n20158 = ~n5690 & n20157 ;
  assign n20159 = n11033 & n16923 ;
  assign n20160 = n20159 ^ n8414 ^ 1'b0 ;
  assign n20161 = n15200 | n20160 ;
  assign n20162 = n8304 & ~n11465 ;
  assign n20163 = n20162 ^ n17710 ^ 1'b0 ;
  assign n20164 = ~n1800 & n4163 ;
  assign n20165 = n12986 ^ n8047 ^ 1'b0 ;
  assign n20166 = n20164 & n20165 ;
  assign n20167 = n9984 ^ n4565 ^ 1'b0 ;
  assign n20171 = ~n5749 & n10163 ;
  assign n20172 = n20171 ^ n7289 ^ 1'b0 ;
  assign n20168 = n4689 ^ n1182 ^ 1'b0 ;
  assign n20169 = n2757 & n20168 ;
  assign n20170 = ~n5800 & n20169 ;
  assign n20173 = n20172 ^ n20170 ^ 1'b0 ;
  assign n20174 = n7506 | n13461 ;
  assign n20175 = n20173 & ~n20174 ;
  assign n20176 = n3858 & ~n7915 ;
  assign n20177 = n788 | n3500 ;
  assign n20178 = n20177 ^ n1270 ^ 1'b0 ;
  assign n20179 = n20176 | n20178 ;
  assign n20180 = n20179 ^ n16703 ^ 1'b0 ;
  assign n20181 = n4577 | n20180 ;
  assign n20182 = n3575 | n20181 ;
  assign n20183 = n15423 | n20182 ;
  assign n20184 = n11577 ^ n1823 ^ 1'b0 ;
  assign n20185 = n20184 ^ n434 ^ 1'b0 ;
  assign n20186 = n1959 & ~n2054 ;
  assign n20187 = ( n3313 & ~n15464 ) | ( n3313 & n20186 ) | ( ~n15464 & n20186 ) ;
  assign n20188 = n20187 ^ n4715 ^ 1'b0 ;
  assign n20189 = n20188 ^ n13513 ^ n4310 ;
  assign n20190 = n10076 ^ n7665 ^ 1'b0 ;
  assign n20191 = n6366 | n20190 ;
  assign n20192 = n4156 & ~n20191 ;
  assign n20193 = n20192 ^ n4936 ^ 1'b0 ;
  assign n20194 = ~n3891 & n4376 ;
  assign n20195 = ~n10532 & n20194 ;
  assign n20196 = n15208 & ~n20195 ;
  assign n20197 = n13391 | n20196 ;
  assign n20198 = n14697 ^ n11480 ^ n2752 ;
  assign n20199 = n1402 | n1961 ;
  assign n20200 = n10856 | n20199 ;
  assign n20201 = n17520 ^ n1154 ^ 1'b0 ;
  assign n20202 = ~n20200 & n20201 ;
  assign n20203 = n20202 ^ n6740 ^ 1'b0 ;
  assign n20204 = n4397 ^ n1629 ^ 1'b0 ;
  assign n20205 = n12248 & ~n15161 ;
  assign n20206 = n20205 ^ n14047 ^ n2670 ;
  assign n20208 = n7598 ^ n5047 ^ 1'b0 ;
  assign n20209 = n8362 & n20208 ;
  assign n20207 = n5022 | n7988 ;
  assign n20210 = n20209 ^ n20207 ^ 1'b0 ;
  assign n20211 = n10087 ^ n8115 ^ 1'b0 ;
  assign n20212 = n11356 & n20211 ;
  assign n20213 = ( n5355 & ~n7694 ) | ( n5355 & n20212 ) | ( ~n7694 & n20212 ) ;
  assign n20214 = n15335 ^ n4681 ^ n4465 ;
  assign n20215 = ( ~n11697 & n13496 ) | ( ~n11697 & n20214 ) | ( n13496 & n20214 ) ;
  assign n20216 = ~n3313 & n5151 ;
  assign n20217 = n8029 ^ n3329 ^ 1'b0 ;
  assign n20218 = ~n499 & n20217 ;
  assign n20219 = ~n13552 & n20218 ;
  assign n20220 = n11406 & n20219 ;
  assign n20221 = n5444 ^ n3491 ^ 1'b0 ;
  assign n20222 = n20221 ^ n17336 ^ n8968 ;
  assign n20223 = n3158 & ~n16461 ;
  assign n20224 = ~n11063 & n20223 ;
  assign n20225 = n9003 | n11874 ;
  assign n20226 = ~n78 & n17619 ;
  assign n20227 = ~n7817 & n10163 ;
  assign n20228 = n20227 ^ n16056 ^ 1'b0 ;
  assign n20229 = n3159 ^ n3142 ^ 1'b0 ;
  assign n20230 = n4640 & n20229 ;
  assign n20231 = ~n8783 & n20230 ;
  assign n20232 = n7686 & n20231 ;
  assign n20233 = ~n2919 & n9981 ;
  assign n20234 = n41 & n2684 ;
  assign n20235 = ~n6762 & n20234 ;
  assign n20236 = n649 & n2405 ;
  assign n20237 = n20236 ^ n1531 ^ 1'b0 ;
  assign n20238 = ( n5806 & ~n16914 ) | ( n5806 & n20237 ) | ( ~n16914 & n20237 ) ;
  assign n20239 = n16060 & n20238 ;
  assign n20240 = n20235 & n20239 ;
  assign n20244 = n2723 & ~n8801 ;
  assign n20245 = n20244 ^ n3486 ^ 1'b0 ;
  assign n20243 = n7060 & n10675 ;
  assign n20246 = n20245 ^ n20243 ^ 1'b0 ;
  assign n20241 = n7122 & ~n12168 ;
  assign n20242 = n20241 ^ n1861 ^ 1'b0 ;
  assign n20247 = n20246 ^ n20242 ^ 1'b0 ;
  assign n20248 = n9687 ^ n9400 ^ 1'b0 ;
  assign n20249 = n205 | n6902 ;
  assign n20250 = n10215 & ~n20249 ;
  assign n20251 = n20248 | n20250 ;
  assign n20252 = ~n5618 & n7974 ;
  assign n20253 = n13275 ^ n2176 ^ 1'b0 ;
  assign n20254 = n2797 & n20253 ;
  assign n20255 = n12452 ^ n7527 ^ 1'b0 ;
  assign n20256 = n20255 ^ n18126 ^ n7357 ;
  assign n20257 = n5059 & n9109 ;
  assign n20258 = ~n4966 & n20257 ;
  assign n20259 = n8993 & ~n9884 ;
  assign n20260 = ~n16806 & n20259 ;
  assign n20261 = n17736 ^ n11542 ^ 1'b0 ;
  assign n20262 = n5231 & ~n20261 ;
  assign n20263 = n7624 & n20262 ;
  assign n20264 = n14745 ^ n1353 ^ 1'b0 ;
  assign n20265 = ~n177 & n5968 ;
  assign n20266 = n20265 ^ n19639 ^ 1'b0 ;
  assign n20267 = n15807 ^ n8812 ^ 1'b0 ;
  assign n20268 = n20266 & ~n20267 ;
  assign n20269 = ( n134 & ~n20264 ) | ( n134 & n20268 ) | ( ~n20264 & n20268 ) ;
  assign n20270 = n18377 ^ n4135 ^ 1'b0 ;
  assign n20271 = ~n9140 & n20270 ;
  assign n20272 = ( ~n2497 & n6021 ) | ( ~n2497 & n6247 ) | ( n6021 & n6247 ) ;
  assign n20273 = n3769 & n8621 ;
  assign n20274 = n19839 ^ n6922 ^ n1957 ;
  assign n20275 = ~n2292 & n3876 ;
  assign n20276 = n20275 ^ n17321 ^ 1'b0 ;
  assign n20277 = n4135 & n8856 ;
  assign n20278 = n7867 & ~n20277 ;
  assign n20279 = n20278 ^ n6411 ^ 1'b0 ;
  assign n20280 = n5585 | n8753 ;
  assign n20281 = n20280 ^ n1023 ^ n188 ;
  assign n20282 = n1794 & ~n20281 ;
  assign n20283 = n9666 & n15586 ;
  assign n20284 = n17586 ^ n2835 ^ 1'b0 ;
  assign n20285 = n5509 | n20284 ;
  assign n20286 = ( n6022 & n7016 ) | ( n6022 & n20285 ) | ( n7016 & n20285 ) ;
  assign n20287 = ~n1168 & n2667 ;
  assign n20288 = ~n11361 & n20287 ;
  assign n20289 = ( n6970 & ~n18454 ) | ( n6970 & n20288 ) | ( ~n18454 & n20288 ) ;
  assign n20290 = ( ~n18516 & n20286 ) | ( ~n18516 & n20289 ) | ( n20286 & n20289 ) ;
  assign n20291 = ( n7751 & ~n11606 ) | ( n7751 & n20290 ) | ( ~n11606 & n20290 ) ;
  assign n20294 = n12413 ^ n4512 ^ 1'b0 ;
  assign n20292 = n139 & ~n11460 ;
  assign n20293 = n19150 | n20292 ;
  assign n20295 = n20294 ^ n20293 ^ 1'b0 ;
  assign n20296 = n20295 ^ n10744 ^ 1'b0 ;
  assign n20297 = n4195 & ~n20296 ;
  assign n20298 = n2482 | n18062 ;
  assign n20299 = n9506 & n11339 ;
  assign n20300 = n1280 ^ n51 ^ 1'b0 ;
  assign n20301 = n20299 & ~n20300 ;
  assign n20302 = n20301 ^ n10559 ^ 1'b0 ;
  assign n20303 = ( ~n6911 & n12576 ) | ( ~n6911 & n18719 ) | ( n12576 & n18719 ) ;
  assign n20304 = n18006 & ~n20303 ;
  assign n20305 = n20304 ^ n8610 ^ 1'b0 ;
  assign n20316 = ~n678 & n11609 ;
  assign n20306 = n7751 ^ n5874 ^ 1'b0 ;
  assign n20307 = ( n10206 & n11374 ) | ( n10206 & n20306 ) | ( n11374 & n20306 ) ;
  assign n20308 = n20307 ^ n7404 ^ 1'b0 ;
  assign n20309 = ~n14644 & n20308 ;
  assign n20310 = n3636 ^ n2949 ^ 1'b0 ;
  assign n20311 = n10079 ^ n8025 ^ n434 ;
  assign n20312 = n20310 | n20311 ;
  assign n20313 = n8547 | n20312 ;
  assign n20314 = n20309 | n20313 ;
  assign n20315 = n14612 & n20314 ;
  assign n20317 = n20316 ^ n20315 ^ 1'b0 ;
  assign n20318 = n1681 | n8033 ;
  assign n20319 = n20318 ^ n2488 ^ 1'b0 ;
  assign n20320 = ( n2510 & n7323 ) | ( n2510 & n20319 ) | ( n7323 & n20319 ) ;
  assign n20321 = ~n12457 & n15159 ;
  assign n20322 = n17913 ^ n5265 ^ 1'b0 ;
  assign n20323 = n6221 & ~n20322 ;
  assign n20324 = n19505 & n20323 ;
  assign n20325 = ~n5864 & n8986 ;
  assign n20326 = n369 & n20325 ;
  assign n20327 = n4959 & ~n18849 ;
  assign n20328 = n20327 ^ n12431 ^ 1'b0 ;
  assign n20329 = ( n3517 & ~n13221 ) | ( n3517 & n13943 ) | ( ~n13221 & n13943 ) ;
  assign n20333 = n132 | n11266 ;
  assign n20334 = n20333 ^ n2857 ^ 1'b0 ;
  assign n20331 = n9996 ^ n3581 ^ 1'b0 ;
  assign n20332 = n14715 & ~n20331 ;
  assign n20330 = n8268 & n9335 ;
  assign n20335 = n20334 ^ n20332 ^ n20330 ;
  assign n20336 = n4327 | n9746 ;
  assign n20337 = n20336 ^ n16799 ^ n12457 ;
  assign n20338 = n17605 ^ n13366 ^ 1'b0 ;
  assign n20339 = n1168 | n20338 ;
  assign n20340 = ( n3709 & n15195 ) | ( n3709 & n20339 ) | ( n15195 & n20339 ) ;
  assign n20341 = n17107 ^ n6013 ^ 1'b0 ;
  assign n20342 = n2324 & ~n19695 ;
  assign n20343 = n20342 ^ n4140 ^ 1'b0 ;
  assign n20344 = ~n67 & n20343 ;
  assign n20345 = n1081 | n20344 ;
  assign n20346 = ~n1142 & n14885 ;
  assign n20347 = n20346 ^ n15746 ^ 1'b0 ;
  assign n20348 = n17900 & ~n20347 ;
  assign n20349 = n11829 & n20348 ;
  assign n20350 = n14057 | n20349 ;
  assign n20351 = ( n1596 & ~n10862 ) | ( n1596 & n12071 ) | ( ~n10862 & n12071 ) ;
  assign n20352 = n20351 ^ n14409 ^ n4114 ;
  assign n20353 = ~n9942 & n20352 ;
  assign n20356 = n6478 ^ n3790 ^ 1'b0 ;
  assign n20354 = ~n2261 & n4322 ;
  assign n20355 = ( x3 & ~n44 ) | ( x3 & n20354 ) | ( ~n44 & n20354 ) ;
  assign n20357 = n20356 ^ n20355 ^ 1'b0 ;
  assign n20358 = n20357 ^ n11766 ^ n7567 ;
  assign n20359 = n2942 & n17267 ;
  assign n20360 = n20359 ^ n11188 ^ 1'b0 ;
  assign n20361 = n523 & ~n16346 ;
  assign n20362 = n3908 & n20361 ;
  assign n20363 = ( n1218 & n8472 ) | ( n1218 & ~n8527 ) | ( n8472 & ~n8527 ) ;
  assign n20364 = ( ~n5441 & n13178 ) | ( ~n5441 & n14824 ) | ( n13178 & n14824 ) ;
  assign n20365 = n20364 ^ n2335 ^ 1'b0 ;
  assign n20366 = n20363 | n20365 ;
  assign n20367 = n7864 & n13975 ;
  assign n20368 = n20367 ^ n1897 ^ 1'b0 ;
  assign n20369 = n13684 ^ n11378 ^ n8569 ;
  assign n20370 = n20368 | n20369 ;
  assign n20371 = n3563 ^ n3207 ^ n221 ;
  assign n20372 = ~n3662 & n20371 ;
  assign n20373 = n7799 | n10319 ;
  assign n20374 = n20373 ^ n1000 ^ 1'b0 ;
  assign n20375 = n20374 ^ n7704 ^ 1'b0 ;
  assign n20376 = n1552 & ~n9535 ;
  assign n20377 = ~n1552 & n20376 ;
  assign n20378 = n16942 ^ n15031 ^ 1'b0 ;
  assign n20379 = n20377 | n20378 ;
  assign n20380 = n10870 & ~n20379 ;
  assign n20381 = ~n5473 & n20380 ;
  assign n20382 = n5355 ^ n2515 ^ 1'b0 ;
  assign n20383 = ~n3302 & n4434 ;
  assign n20384 = n20383 ^ n3962 ^ 1'b0 ;
  assign n20385 = ~n20382 & n20384 ;
  assign n20386 = n19931 ^ n278 ^ 1'b0 ;
  assign n20387 = ~n4520 & n15800 ;
  assign n20388 = n4330 ^ n2330 ^ 1'b0 ;
  assign n20389 = ~n20387 & n20388 ;
  assign n20391 = ~n139 & n4283 ;
  assign n20392 = n20391 ^ n3932 ^ 1'b0 ;
  assign n20393 = n8567 & n13881 ;
  assign n20394 = n20392 & n20393 ;
  assign n20390 = n4383 | n9519 ;
  assign n20395 = n20394 ^ n20390 ^ 1'b0 ;
  assign n20396 = n332 & ~n20395 ;
  assign n20397 = ~n1001 & n9596 ;
  assign n20398 = ~n14868 & n20397 ;
  assign n20399 = n20396 & n20398 ;
  assign n20400 = n14255 ^ n1702 ^ 1'b0 ;
  assign n20401 = ~n20399 & n20400 ;
  assign n20402 = ~n20389 & n20401 ;
  assign n20403 = n20402 ^ n44 ^ 1'b0 ;
  assign n20404 = n10456 ^ n9457 ^ n8656 ;
  assign n20405 = n10727 & ~n15779 ;
  assign n20406 = n15194 | n15863 ;
  assign n20407 = n9242 ^ n8269 ^ 1'b0 ;
  assign n20408 = n20407 ^ n17718 ^ 1'b0 ;
  assign n20409 = ~n4549 & n20408 ;
  assign n20410 = ~n3773 & n9557 ;
  assign n20411 = n20410 ^ n11920 ^ 1'b0 ;
  assign n20412 = n20411 ^ n157 ^ 1'b0 ;
  assign n20413 = n11768 ^ n2745 ^ 1'b0 ;
  assign n20414 = n12963 & n15330 ;
  assign n20415 = ~n20413 & n20414 ;
  assign n20416 = n11053 & ~n20415 ;
  assign n20417 = ( n36 & ~n6363 ) | ( n36 & n8750 ) | ( ~n6363 & n8750 ) ;
  assign n20418 = n6806 & ~n20417 ;
  assign n20419 = n20418 ^ n4633 ^ 1'b0 ;
  assign n20420 = n3408 & ~n20419 ;
  assign n20421 = n20420 ^ n645 ^ 1'b0 ;
  assign n20422 = n1125 & ~n10254 ;
  assign n20426 = n6093 ^ n5086 ^ 1'b0 ;
  assign n20423 = n5361 ^ n3508 ^ 1'b0 ;
  assign n20424 = ~n9936 & n20423 ;
  assign n20425 = n20424 ^ n1684 ^ 1'b0 ;
  assign n20427 = n20426 ^ n20425 ^ 1'b0 ;
  assign n20428 = ~n1180 & n20427 ;
  assign n20429 = n15070 ^ n1084 ^ 1'b0 ;
  assign n20430 = n20428 & ~n20429 ;
  assign n20431 = n2250 & n5866 ;
  assign n20432 = n20431 ^ n12276 ^ 1'b0 ;
  assign n20433 = ~n12211 & n20432 ;
  assign n20434 = n278 & n8435 ;
  assign n20435 = n20434 ^ n10197 ^ 1'b0 ;
  assign n20436 = n10385 & ~n20435 ;
  assign n20437 = n7692 & n20436 ;
  assign n20438 = n6852 ^ n2369 ^ 1'b0 ;
  assign n20439 = ( ~n14697 & n20086 ) | ( ~n14697 & n20438 ) | ( n20086 & n20438 ) ;
  assign n20440 = n6510 & n10125 ;
  assign n20441 = n20440 ^ n7329 ^ 1'b0 ;
  assign n20442 = ~n1412 & n4717 ;
  assign n20443 = ~n5352 & n20442 ;
  assign n20444 = n20443 ^ n10031 ^ 1'b0 ;
  assign n20445 = n947 & n15946 ;
  assign n20446 = n20444 & n20445 ;
  assign n20447 = n10838 | n20446 ;
  assign n20448 = n20447 ^ n4916 ^ 1'b0 ;
  assign n20449 = n12520 ^ n525 ^ 1'b0 ;
  assign n20450 = n8733 & n10350 ;
  assign n20451 = n16625 ^ n14033 ^ 1'b0 ;
  assign n20452 = n1768 | n20451 ;
  assign n20453 = n20452 ^ n19068 ^ n16200 ;
  assign n20454 = ~n249 & n18174 ;
  assign n20455 = ~n6696 & n20454 ;
  assign n20456 = ( ~n1918 & n10404 ) | ( ~n1918 & n19005 ) | ( n10404 & n19005 ) ;
  assign n20457 = n8896 ^ n4544 ^ n544 ;
  assign n20458 = ( n1156 & ~n1865 ) | ( n1156 & n20457 ) | ( ~n1865 & n20457 ) ;
  assign n20459 = n3192 & ~n12003 ;
  assign n20460 = n20459 ^ n15347 ^ 1'b0 ;
  assign n20461 = n20460 ^ n15980 ^ 1'b0 ;
  assign n20462 = n1071 & n20461 ;
  assign n20463 = n835 & ~n18711 ;
  assign n20464 = n20463 ^ n8896 ^ 1'b0 ;
  assign n20465 = n9699 ^ n2541 ^ 1'b0 ;
  assign n20466 = n3628 & n20465 ;
  assign n20467 = ~n3552 & n20062 ;
  assign n20468 = ~n6743 & n20467 ;
  assign n20469 = ~n7231 & n20468 ;
  assign n20470 = n20469 ^ n9344 ^ 1'b0 ;
  assign n20471 = n6292 ^ n3590 ^ 1'b0 ;
  assign n20472 = ~n3104 & n15677 ;
  assign n20473 = n20471 & n20472 ;
  assign n20474 = n4235 & n6005 ;
  assign n20475 = n14622 & n20474 ;
  assign n20476 = n20475 ^ n9879 ^ n8678 ;
  assign n20477 = n2419 ^ n1822 ^ 1'b0 ;
  assign n20485 = n3489 ^ n1023 ^ 1'b0 ;
  assign n20486 = n649 | n20485 ;
  assign n20483 = ~n1905 & n11794 ;
  assign n20484 = n18662 & n20483 ;
  assign n20487 = n20486 ^ n20484 ^ n17173 ;
  assign n20488 = ~n790 & n20487 ;
  assign n20489 = n6306 & n20488 ;
  assign n20478 = n2445 | n2873 ;
  assign n20479 = n2873 & ~n20478 ;
  assign n20480 = n1638 | n20479 ;
  assign n20481 = n20479 & ~n20480 ;
  assign n20482 = n11120 & ~n20481 ;
  assign n20490 = n20489 ^ n20482 ^ 1'b0 ;
  assign n20491 = n5704 ^ n13 ^ 1'b0 ;
  assign n20493 = n2999 & ~n6866 ;
  assign n20494 = n20493 ^ n923 ^ 1'b0 ;
  assign n20495 = n2684 & n12292 ;
  assign n20496 = n20494 & n20495 ;
  assign n20497 = ~n8682 & n20496 ;
  assign n20492 = n3637 & n6249 ;
  assign n20498 = n20497 ^ n20492 ^ 1'b0 ;
  assign n20499 = n20498 ^ n2132 ^ 1'b0 ;
  assign n20500 = ~n16038 & n20499 ;
  assign n20501 = n20491 & n20500 ;
  assign n20502 = ( n6491 & n12558 ) | ( n6491 & ~n17077 ) | ( n12558 & ~n17077 ) ;
  assign n20503 = ( n1455 & n12271 ) | ( n1455 & n13338 ) | ( n12271 & n13338 ) ;
  assign n20504 = ~n15310 & n20503 ;
  assign n20505 = ~n20502 & n20504 ;
  assign n20506 = ~n8937 & n20272 ;
  assign n20507 = n20506 ^ n8493 ^ 1'b0 ;
  assign n20508 = n10793 ^ n890 ^ 1'b0 ;
  assign n20509 = ~n3936 & n20508 ;
  assign n20510 = n20509 ^ n10379 ^ 1'b0 ;
  assign n20511 = n13032 ^ n7737 ^ 1'b0 ;
  assign n20512 = ~n4222 & n14141 ;
  assign n20513 = n8045 & ~n20512 ;
  assign n20514 = ~n1370 & n9208 ;
  assign n20515 = n14443 ^ n7505 ^ n4066 ;
  assign n20516 = n126 | n13789 ;
  assign n20517 = n20516 ^ n18103 ^ 1'b0 ;
  assign n20518 = n1312 | n7789 ;
  assign n20520 = ~n6284 & n19372 ;
  assign n20521 = n20520 ^ n17147 ^ 1'b0 ;
  assign n20519 = n9942 | n15114 ;
  assign n20522 = n20521 ^ n20519 ^ 1'b0 ;
  assign n20525 = n437 & ~n5502 ;
  assign n20526 = n1253 & n20525 ;
  assign n20523 = ~n6582 & n7868 ;
  assign n20524 = n20523 ^ n10992 ^ 1'b0 ;
  assign n20527 = n20526 ^ n20524 ^ 1'b0 ;
  assign n20528 = ~n5533 & n20527 ;
  assign n20529 = n12438 ^ n5484 ^ 1'b0 ;
  assign n20530 = n11059 ^ n4237 ^ n2073 ;
  assign n20531 = n20529 & n20530 ;
  assign n20532 = n4195 & ~n14373 ;
  assign n20533 = n10867 & ~n20532 ;
  assign n20534 = n9755 ^ n4109 ^ n241 ;
  assign n20535 = ~n7226 & n20534 ;
  assign n20536 = ( n2976 & ~n6683 ) | ( n2976 & n20535 ) | ( ~n6683 & n20535 ) ;
  assign n20537 = n10379 ^ n2176 ^ 1'b0 ;
  assign n20538 = n16561 ^ n2804 ^ 1'b0 ;
  assign n20542 = n8333 ^ n8172 ^ 1'b0 ;
  assign n20543 = n7701 ^ n2229 ^ 1'b0 ;
  assign n20544 = n2904 & n20543 ;
  assign n20545 = n20542 & n20544 ;
  assign n20539 = n17194 ^ n11433 ^ 1'b0 ;
  assign n20540 = n3376 & n20539 ;
  assign n20541 = n20540 ^ n10210 ^ 1'b0 ;
  assign n20546 = n20545 ^ n20541 ^ 1'b0 ;
  assign n20547 = n70 & n2242 ;
  assign n20548 = n20547 ^ n19213 ^ 1'b0 ;
  assign n20549 = n11676 & n18458 ;
  assign n20550 = n12879 | n20549 ;
  assign n20551 = n13114 ^ n8476 ^ n900 ;
  assign n20552 = n15774 ^ n7022 ^ 1'b0 ;
  assign n20553 = n20552 ^ n6421 ^ 1'b0 ;
  assign n20554 = n10405 & n20553 ;
  assign n20555 = n20105 ^ n79 ^ 1'b0 ;
  assign n20556 = ~n601 & n20555 ;
  assign n20557 = ~n10748 & n20556 ;
  assign n20558 = n1731 & ~n3807 ;
  assign n20559 = n20558 ^ n816 ^ 1'b0 ;
  assign n20560 = n11135 & ~n20559 ;
  assign n20561 = ( n523 & n8874 ) | ( n523 & n20560 ) | ( n8874 & n20560 ) ;
  assign n20562 = n14557 & ~n20042 ;
  assign n20563 = n20562 ^ n10812 ^ 1'b0 ;
  assign n20564 = n12423 ^ n11480 ^ n8987 ;
  assign n20565 = n10241 ^ n1784 ^ 1'b0 ;
  assign n20566 = ( n20563 & n20564 ) | ( n20563 & n20565 ) | ( n20564 & n20565 ) ;
  assign n20570 = n7881 ^ n5556 ^ 1'b0 ;
  assign n20567 = n4021 | n16293 ;
  assign n20568 = ~n3229 & n20567 ;
  assign n20569 = n10632 & ~n20568 ;
  assign n20571 = n20570 ^ n20569 ^ 1'b0 ;
  assign n20572 = n379 | n3564 ;
  assign n20573 = n1056 | n20572 ;
  assign n20574 = n20248 ^ n5594 ^ n4854 ;
  assign n20575 = n4840 & ~n20574 ;
  assign n20576 = ~n20573 & n20575 ;
  assign n20577 = ~n4058 & n18133 ;
  assign n20578 = ~n19640 & n20577 ;
  assign n20582 = n20446 ^ n3654 ^ n2942 ;
  assign n20579 = n11772 & ~n20009 ;
  assign n20580 = n20579 ^ n5083 ^ 1'b0 ;
  assign n20581 = n4582 & ~n20580 ;
  assign n20583 = n20582 ^ n20581 ^ 1'b0 ;
  assign n20584 = n20112 ^ n6670 ^ 1'b0 ;
  assign n20585 = n12262 | n20584 ;
  assign n20586 = n7698 ^ n3776 ^ n3008 ;
  assign n20587 = n508 | n2569 ;
  assign n20588 = n20587 ^ n3008 ^ 1'b0 ;
  assign n20589 = n9295 | n16939 ;
  assign n20590 = ( n2786 & ~n20588 ) | ( n2786 & n20589 ) | ( ~n20588 & n20589 ) ;
  assign n20591 = n15341 ^ n12495 ^ 1'b0 ;
  assign n20592 = n694 | n20591 ;
  assign n20593 = n12059 ^ n5876 ^ n5389 ;
  assign n20594 = n1109 | n20593 ;
  assign n20595 = n1022 & n2867 ;
  assign n20596 = n20595 ^ n5428 ^ 1'b0 ;
  assign n20597 = n20596 ^ n6864 ^ 1'b0 ;
  assign n20598 = n4427 & n20597 ;
  assign n20599 = ~n6016 & n20598 ;
  assign n20600 = ( n99 & n7796 ) | ( n99 & n20599 ) | ( n7796 & n20599 ) ;
  assign n20602 = ~n285 & n1841 ;
  assign n20601 = ~n2004 & n19191 ;
  assign n20603 = n20602 ^ n20601 ^ n7699 ;
  assign n20604 = n3087 | n20603 ;
  assign n20605 = n20600 | n20604 ;
  assign n20606 = ~n15005 & n16118 ;
  assign n20607 = n18516 & n20606 ;
  assign n20608 = ~n360 & n20607 ;
  assign n20609 = ~n17700 & n20608 ;
  assign n20610 = n10583 ^ n6890 ^ 1'b0 ;
  assign n20611 = n20610 ^ n13057 ^ 1'b0 ;
  assign n20612 = n10708 ^ n10677 ^ 1'b0 ;
  assign n20613 = n3372 ^ n2580 ^ 1'b0 ;
  assign n20614 = n20612 & ~n20613 ;
  assign n20615 = n20614 ^ n8888 ^ 1'b0 ;
  assign n20616 = n19637 | n20615 ;
  assign n20617 = n17860 ^ n9615 ^ n441 ;
  assign n20618 = n10989 & n20617 ;
  assign n20619 = n4482 & n20618 ;
  assign n20620 = n17659 ^ n9984 ^ 1'b0 ;
  assign n20621 = n20619 | n20620 ;
  assign n20622 = n8142 ^ n2695 ^ 1'b0 ;
  assign n20623 = n20621 & n20622 ;
  assign n20624 = n1071 & ~n3463 ;
  assign n20625 = n20624 ^ n1979 ^ 1'b0 ;
  assign n20626 = ( ~n1568 & n9486 ) | ( ~n1568 & n20625 ) | ( n9486 & n20625 ) ;
  assign n20627 = n2867 & ~n20626 ;
  assign n20628 = n14298 ^ n9901 ^ 1'b0 ;
  assign n20629 = n20627 | n20628 ;
  assign n20630 = n20629 ^ n11403 ^ 1'b0 ;
  assign n20631 = ( n8915 & n14405 ) | ( n8915 & n15006 ) | ( n14405 & n15006 ) ;
  assign n20632 = n15265 ^ n10594 ^ n9690 ;
  assign n20633 = n2230 ^ n527 ^ 1'b0 ;
  assign n20634 = ~n1533 & n20633 ;
  assign n20635 = n20634 ^ n3179 ^ 1'b0 ;
  assign n20636 = ( n5830 & ~n14603 ) | ( n5830 & n14857 ) | ( ~n14603 & n14857 ) ;
  assign n20637 = n3040 & n5818 ;
  assign n20638 = n408 & n20637 ;
  assign n20639 = n12083 & ~n20638 ;
  assign n20640 = n20639 ^ n7151 ^ 1'b0 ;
  assign n20641 = n20640 ^ n19983 ^ 1'b0 ;
  assign n20642 = n18778 ^ n937 ^ 1'b0 ;
  assign n20643 = n20641 | n20642 ;
  assign n20644 = n20636 & ~n20643 ;
  assign n20646 = n472 | n885 ;
  assign n20645 = n3157 ^ n388 ^ 1'b0 ;
  assign n20647 = n20646 ^ n20645 ^ 1'b0 ;
  assign n20648 = n20647 ^ n16919 ^ 1'b0 ;
  assign n20649 = ~n12681 & n17450 ;
  assign n20650 = n13296 ^ n5188 ^ 1'b0 ;
  assign n20651 = n3449 | n6987 ;
  assign n20652 = n14101 & ~n20651 ;
  assign n20653 = n20650 & ~n20652 ;
  assign n20654 = ~n2670 & n4677 ;
  assign n20655 = n11983 | n20252 ;
  assign n20656 = n12682 ^ n9496 ^ 1'b0 ;
  assign n20657 = n16647 ^ n236 ^ 1'b0 ;
  assign n20658 = n5173 & ~n20657 ;
  assign n20659 = ( ~n1295 & n10527 ) | ( ~n1295 & n20658 ) | ( n10527 & n20658 ) ;
  assign n20660 = ( n6320 & n19610 ) | ( n6320 & ~n20659 ) | ( n19610 & ~n20659 ) ;
  assign n20661 = n13326 ^ n592 ^ 1'b0 ;
  assign n20664 = n5957 ^ n2184 ^ n164 ;
  assign n20663 = n15729 | n16597 ;
  assign n20665 = n20664 ^ n20663 ^ 1'b0 ;
  assign n20662 = n1606 & ~n4126 ;
  assign n20666 = n20665 ^ n20662 ^ n16189 ;
  assign n20667 = n13558 & ~n20666 ;
  assign n20668 = n11961 ^ n6129 ^ 1'b0 ;
  assign n20669 = ( n465 & n7708 ) | ( n465 & ~n20668 ) | ( n7708 & ~n20668 ) ;
  assign n20670 = n2858 | n19399 ;
  assign n20671 = n18123 | n20670 ;
  assign n20672 = n10481 ^ n3025 ^ 1'b0 ;
  assign n20673 = n188 & n20672 ;
  assign n20674 = ~n20671 & n20673 ;
  assign n20675 = n2008 ^ n873 ^ 1'b0 ;
  assign n20676 = n5370 & n17693 ;
  assign n20677 = n20675 & n20676 ;
  assign n20678 = n8894 ^ n3998 ^ 1'b0 ;
  assign n20680 = n15260 ^ n6356 ^ n471 ;
  assign n20679 = ~n9649 & n17099 ;
  assign n20681 = n20680 ^ n20679 ^ 1'b0 ;
  assign n20682 = n18522 ^ n9395 ^ 1'b0 ;
  assign n20683 = ~n8597 & n9702 ;
  assign n20684 = n3603 & n20683 ;
  assign n20685 = ~n10638 & n15382 ;
  assign n20686 = n570 | n20685 ;
  assign n20687 = ~n6754 & n7545 ;
  assign n20688 = n20687 ^ n12519 ^ 1'b0 ;
  assign n20689 = ~n1362 & n17628 ;
  assign n20690 = ~n961 & n8206 ;
  assign n20691 = n20690 ^ n811 ^ 1'b0 ;
  assign n20692 = n7195 ^ n5321 ^ 1'b0 ;
  assign n20693 = n11648 | n20692 ;
  assign n20694 = n57 & n784 ;
  assign n20695 = n20694 ^ n15787 ^ 1'b0 ;
  assign n20696 = ( n12576 & n13346 ) | ( n12576 & n13986 ) | ( n13346 & n13986 ) ;
  assign n20697 = n13133 ^ n8684 ^ 1'b0 ;
  assign n20698 = ~n20696 & n20697 ;
  assign n20699 = n2677 ^ n1798 ^ 1'b0 ;
  assign n20700 = ( n20695 & n20698 ) | ( n20695 & n20699 ) | ( n20698 & n20699 ) ;
  assign n20701 = n19875 ^ n2408 ^ 1'b0 ;
  assign n20702 = ~n16370 & n20701 ;
  assign n20703 = n1809 & ~n4889 ;
  assign n20704 = n20703 ^ n16345 ^ 1'b0 ;
  assign n20705 = n20704 ^ n401 ^ 1'b0 ;
  assign n20706 = n16923 ^ n6470 ^ n3546 ;
  assign n20707 = n6658 ^ n1419 ^ 1'b0 ;
  assign n20708 = n6736 | n20707 ;
  assign n20709 = n20708 ^ n4540 ^ 1'b0 ;
  assign n20710 = ~n10406 & n20709 ;
  assign n20711 = ( ~n14353 & n20706 ) | ( ~n14353 & n20710 ) | ( n20706 & n20710 ) ;
  assign n20712 = n10004 ^ n6522 ^ 1'b0 ;
  assign n20713 = ~n7825 & n17098 ;
  assign n20714 = n20452 ^ n4412 ^ 1'b0 ;
  assign n20715 = ( n361 & n20096 ) | ( n361 & ~n20714 ) | ( n20096 & ~n20714 ) ;
  assign n20716 = n7880 ^ n2149 ^ n990 ;
  assign n20717 = n16150 & n20716 ;
  assign n20718 = ~n2358 & n7315 ;
  assign n20719 = n19038 & ~n20718 ;
  assign n20720 = ~n2217 & n9905 ;
  assign n20721 = n3919 ^ n3115 ^ 1'b0 ;
  assign n20722 = ( n5415 & n14724 ) | ( n5415 & ~n20721 ) | ( n14724 & ~n20721 ) ;
  assign n20724 = ~n539 & n16021 ;
  assign n20725 = n20724 ^ n18819 ^ n2984 ;
  assign n20723 = ~n11750 & n19058 ;
  assign n20726 = n20725 ^ n20723 ^ 1'b0 ;
  assign n20727 = ( ~n973 & n1857 ) | ( ~n973 & n8543 ) | ( n1857 & n8543 ) ;
  assign n20728 = n20727 ^ n9721 ^ 1'b0 ;
  assign n20729 = ~n10594 & n20728 ;
  assign n20730 = n20729 ^ n6159 ^ 1'b0 ;
  assign n20731 = n20726 | n20730 ;
  assign n20732 = n15554 ^ n7690 ^ 1'b0 ;
  assign n20733 = n3789 & n20732 ;
  assign n20734 = n4271 ^ n1311 ^ 1'b0 ;
  assign n20735 = n20734 ^ n523 ^ 1'b0 ;
  assign n20736 = n18032 & n20735 ;
  assign n20737 = ( ~n1800 & n13737 ) | ( ~n1800 & n16492 ) | ( n13737 & n16492 ) ;
  assign n20738 = n20737 ^ n7864 ^ 1'b0 ;
  assign n20739 = ~n551 & n12480 ;
  assign n20740 = ( n1877 & ~n7813 ) | ( n1877 & n17576 ) | ( ~n7813 & n17576 ) ;
  assign n20741 = n20740 ^ n15467 ^ 1'b0 ;
  assign n20742 = ~n20739 & n20741 ;
  assign n20743 = n15348 ^ n811 ^ 1'b0 ;
  assign n20744 = n10523 & n20743 ;
  assign n20745 = ~n7545 & n20744 ;
  assign n20746 = n5492 & n7778 ;
  assign n20747 = n20746 ^ n3832 ^ 1'b0 ;
  assign n20748 = n11574 & n17381 ;
  assign n20749 = n17763 ^ n6211 ^ 1'b0 ;
  assign n20750 = ~n20748 & n20749 ;
  assign n20751 = ~n1787 & n20196 ;
  assign n20752 = n892 & n923 ;
  assign n20753 = ~n15674 & n20752 ;
  assign n20754 = n1766 & n2521 ;
  assign n20755 = n8549 & n19988 ;
  assign n20756 = ( n5534 & ~n7077 ) | ( n5534 & n8622 ) | ( ~n7077 & n8622 ) ;
  assign n20758 = n2314 | n3787 ;
  assign n20759 = n7736 & ~n20758 ;
  assign n20757 = ~n2393 & n16356 ;
  assign n20760 = n20759 ^ n20757 ^ 1'b0 ;
  assign n20761 = ~n10862 & n14628 ;
  assign n20762 = n18602 | n20761 ;
  assign n20763 = n10773 & n15189 ;
  assign n20764 = ( ~n9999 & n16917 ) | ( ~n9999 & n19283 ) | ( n16917 & n19283 ) ;
  assign n20765 = n676 & ~n5289 ;
  assign n20766 = ~n2114 & n12569 ;
  assign n20767 = ( n7421 & n9685 ) | ( n7421 & n11805 ) | ( n9685 & n11805 ) ;
  assign n20768 = n7404 ^ n1031 ^ 1'b0 ;
  assign n20769 = n20768 ^ n12852 ^ n9397 ;
  assign n20772 = ( n1365 & ~n5156 ) | ( n1365 & n6537 ) | ( ~n5156 & n6537 ) ;
  assign n20773 = ~n5022 & n20772 ;
  assign n20770 = n7954 & ~n10130 ;
  assign n20771 = ~n13457 & n20770 ;
  assign n20774 = n20773 ^ n20771 ^ 1'b0 ;
  assign n20775 = n20774 ^ n16547 ^ 1'b0 ;
  assign n20781 = n3622 & n9944 ;
  assign n20782 = n20781 ^ n13654 ^ 1'b0 ;
  assign n20776 = n2857 ^ n2056 ^ 1'b0 ;
  assign n20777 = n14500 ^ n8176 ^ 1'b0 ;
  assign n20778 = n20776 & ~n20777 ;
  assign n20779 = n20778 ^ n6632 ^ 1'b0 ;
  assign n20780 = n19292 & ~n20779 ;
  assign n20783 = n20782 ^ n20780 ^ 1'b0 ;
  assign n20784 = n15729 ^ n3113 ^ 1'b0 ;
  assign n20785 = n953 & n4144 ;
  assign n20786 = n3892 & n20785 ;
  assign n20787 = n20786 ^ n14664 ^ 1'b0 ;
  assign n20788 = ~n20784 & n20787 ;
  assign n20789 = n8780 ^ n929 ^ 1'b0 ;
  assign n20790 = n5144 & n20789 ;
  assign n20791 = ~n14426 & n20790 ;
  assign n20792 = ( ~n5195 & n9481 ) | ( ~n5195 & n20791 ) | ( n9481 & n20791 ) ;
  assign n20793 = n1367 & ~n2160 ;
  assign n20794 = n5237 & n12793 ;
  assign n20795 = ~n20793 & n20794 ;
  assign n20796 = n10967 ^ n4830 ^ 1'b0 ;
  assign n20797 = n17285 ^ n15700 ^ 1'b0 ;
  assign n20798 = n20796 | n20797 ;
  assign n20799 = n12903 & ~n20798 ;
  assign n20800 = ~n2566 & n14967 ;
  assign n20801 = n20800 ^ n8165 ^ 1'b0 ;
  assign n20802 = n1523 & ~n9713 ;
  assign n20803 = ~n20801 & n20802 ;
  assign n20804 = ~n78 & n3371 ;
  assign n20805 = n20804 ^ n2064 ^ 1'b0 ;
  assign n20806 = n19607 ^ n17480 ^ 1'b0 ;
  assign n20807 = n20805 & ~n20806 ;
  assign n20808 = n20227 ^ n6455 ^ 1'b0 ;
  assign n20809 = n7900 & ~n20808 ;
  assign n20810 = n11002 ^ n1397 ^ 1'b0 ;
  assign n20811 = n13584 ^ n2050 ^ 1'b0 ;
  assign n20812 = n20811 ^ n14226 ^ n10318 ;
  assign n20813 = n20812 ^ n7694 ^ 1'b0 ;
  assign n20814 = n5377 ^ n1332 ^ 1'b0 ;
  assign n20815 = n10412 | n20814 ;
  assign n20816 = n20815 ^ n20027 ^ n3995 ;
  assign n20817 = n4662 ^ n541 ^ 1'b0 ;
  assign n20818 = n9392 ^ n4467 ^ 1'b0 ;
  assign n20819 = n11258 | n20818 ;
  assign n20820 = n20817 & ~n20819 ;
  assign n20821 = ~n20816 & n20820 ;
  assign n20822 = n7468 & ~n8441 ;
  assign n20823 = ~n13297 & n15130 ;
  assign n20824 = ~n15552 & n20823 ;
  assign n20825 = n12677 & n14848 ;
  assign n20826 = ~n11654 & n20825 ;
  assign n20827 = ( n8712 & n13514 ) | ( n8712 & ~n20826 ) | ( n13514 & ~n20826 ) ;
  assign n20828 = n5285 ^ n5047 ^ 1'b0 ;
  assign n20829 = n115 | n20828 ;
  assign n20830 = ( ~n13690 & n18252 ) | ( ~n13690 & n20829 ) | ( n18252 & n20829 ) ;
  assign n20831 = n11804 & n20830 ;
  assign n20832 = n6118 & ~n20831 ;
  assign n20833 = n1201 | n18590 ;
  assign n20834 = n1102 | n20833 ;
  assign n20835 = ~n6305 & n7540 ;
  assign n20836 = n3515 & ~n20835 ;
  assign n20837 = n165 & ~n1328 ;
  assign n20838 = n4978 & n20837 ;
  assign n20839 = n9895 & n20838 ;
  assign n20840 = n13825 ^ n8009 ^ 1'b0 ;
  assign n20846 = n12879 | n13703 ;
  assign n20847 = n7387 & ~n20846 ;
  assign n20848 = n2216 | n20847 ;
  assign n20841 = n18770 ^ n1816 ^ 1'b0 ;
  assign n20842 = n1078 | n20841 ;
  assign n20843 = n20842 ^ n11479 ^ n5781 ;
  assign n20844 = n12937 & n20843 ;
  assign n20845 = ( n10459 & n10934 ) | ( n10459 & ~n20844 ) | ( n10934 & ~n20844 ) ;
  assign n20849 = n20848 ^ n20845 ^ n15683 ;
  assign n20850 = n9493 ^ n1179 ^ 1'b0 ;
  assign n20851 = n2524 & n18813 ;
  assign n20852 = n11573 & n20851 ;
  assign n20853 = ~n1104 & n9799 ;
  assign n20854 = n20853 ^ n4768 ^ 1'b0 ;
  assign n20855 = n20854 ^ n441 ^ 1'b0 ;
  assign n20856 = ~n237 & n5631 ;
  assign n20857 = n11422 & ~n20856 ;
  assign n20858 = n10303 & n20857 ;
  assign n20859 = n4271 ^ n1276 ^ 1'b0 ;
  assign n20860 = n16666 & n20859 ;
  assign n20861 = n8764 & n20860 ;
  assign n20862 = n12243 & ~n20861 ;
  assign n20863 = n20858 & n20862 ;
  assign n20865 = n6415 ^ n2172 ^ 1'b0 ;
  assign n20866 = ~n17315 & n20865 ;
  assign n20864 = n682 & n11157 ;
  assign n20867 = n20866 ^ n20864 ^ 1'b0 ;
  assign n20876 = n142 & n5662 ;
  assign n20868 = n499 | n10091 ;
  assign n20869 = n20868 ^ n20497 ^ 1'b0 ;
  assign n20870 = n984 | n6654 ;
  assign n20871 = n10239 & ~n16896 ;
  assign n20872 = n20870 | n20871 ;
  assign n20873 = ( ~n3071 & n19426 ) | ( ~n3071 & n20872 ) | ( n19426 & n20872 ) ;
  assign n20874 = ~n989 & n20873 ;
  assign n20875 = n20869 | n20874 ;
  assign n20877 = n20876 ^ n20875 ^ 1'b0 ;
  assign n20878 = ~n475 & n17766 ;
  assign n20879 = n8170 & n9288 ;
  assign n20880 = n10846 ^ n2152 ^ 1'b0 ;
  assign n20881 = n20880 ^ n19693 ^ 1'b0 ;
  assign n20882 = n17548 & ~n20881 ;
  assign n20883 = n670 | n14973 ;
  assign n20884 = n285 & ~n20883 ;
  assign n20885 = n11565 ^ n8761 ^ 1'b0 ;
  assign n20886 = ~n17627 & n20885 ;
  assign n20887 = n35 | n19341 ;
  assign n20888 = ~n2346 & n8241 ;
  assign n20889 = ~n2712 & n17658 ;
  assign n20890 = ~n9109 & n20889 ;
  assign n20891 = n20890 ^ n7981 ^ 1'b0 ;
  assign n20892 = n20891 ^ n20827 ^ 1'b0 ;
  assign n20893 = n2926 ^ n732 ^ 1'b0 ;
  assign n20894 = n12089 ^ n1597 ^ 1'b0 ;
  assign n20895 = n14462 & n20894 ;
  assign n20896 = ( n5589 & n7684 ) | ( n5589 & ~n9597 ) | ( n7684 & ~n9597 ) ;
  assign n20897 = n7008 ^ n5997 ^ 1'b0 ;
  assign n20898 = ~n11902 & n19058 ;
  assign n20899 = n3650 ^ n2341 ^ 1'b0 ;
  assign n20901 = n966 | n8360 ;
  assign n20902 = n3725 | n20901 ;
  assign n20900 = n6727 | n14953 ;
  assign n20903 = n20902 ^ n20900 ^ 1'b0 ;
  assign n20904 = n20903 ^ n13455 ^ 1'b0 ;
  assign n20905 = n11846 ^ n5638 ^ 1'b0 ;
  assign n20906 = ~n9532 & n18595 ;
  assign n20907 = ( n885 & n7040 ) | ( n885 & ~n12987 ) | ( n7040 & ~n12987 ) ;
  assign n20908 = n16846 | n20907 ;
  assign n20909 = n20908 ^ n11472 ^ n2471 ;
  assign n20910 = n11195 & n15396 ;
  assign n20911 = n8664 | n19210 ;
  assign n20912 = n20911 ^ n20885 ^ 1'b0 ;
  assign n20913 = ~n20910 & n20912 ;
  assign n20914 = n14371 ^ n1704 ^ 1'b0 ;
  assign n20915 = n6864 | n20914 ;
  assign n20916 = n1311 | n3447 ;
  assign n20917 = n2070 | n20916 ;
  assign n20918 = n20917 ^ n7648 ^ 1'b0 ;
  assign n20919 = n2377 & n20918 ;
  assign n20924 = ~n4021 & n5427 ;
  assign n20920 = n4497 & ~n9274 ;
  assign n20921 = n14674 & n20920 ;
  assign n20922 = n13041 ^ n4258 ^ 1'b0 ;
  assign n20923 = ~n20921 & n20922 ;
  assign n20925 = n20924 ^ n20923 ^ 1'b0 ;
  assign n20926 = n8033 ^ n2995 ^ 1'b0 ;
  assign n20927 = ( n4092 & ~n4769 ) | ( n4092 & n12147 ) | ( ~n4769 & n12147 ) ;
  assign n20928 = n20927 ^ n4390 ^ 1'b0 ;
  assign n20929 = n20926 & ~n20928 ;
  assign n20930 = n7428 ^ n2158 ^ 1'b0 ;
  assign n20931 = n10534 & n20930 ;
  assign n20932 = ~n20537 & n20931 ;
  assign n20933 = n20932 ^ n12440 ^ 1'b0 ;
  assign n20936 = n6503 ^ n874 ^ 1'b0 ;
  assign n20937 = n10254 & ~n20936 ;
  assign n20934 = n1024 & ~n3426 ;
  assign n20935 = n5272 & ~n20934 ;
  assign n20938 = n20937 ^ n20935 ^ 1'b0 ;
  assign n20939 = ~n1105 & n1744 ;
  assign n20940 = n20939 ^ n9471 ^ 1'b0 ;
  assign n20941 = n20940 ^ n2758 ^ 1'b0 ;
  assign n20942 = n10879 & ~n20941 ;
  assign n20948 = n12812 ^ n3109 ^ 1'b0 ;
  assign n20946 = n5610 & ~n13356 ;
  assign n20947 = n5913 & ~n20946 ;
  assign n20949 = n20948 ^ n20947 ^ 1'b0 ;
  assign n20945 = n545 & ~n11549 ;
  assign n20950 = n20949 ^ n20945 ^ 1'b0 ;
  assign n20943 = ( n2170 & n6298 ) | ( n2170 & ~n8674 ) | ( n6298 & ~n8674 ) ;
  assign n20944 = n7009 | n20943 ;
  assign n20951 = n20950 ^ n20944 ^ 1'b0 ;
  assign n20952 = n18330 | n20564 ;
  assign n20953 = n20952 ^ n6991 ^ 1'b0 ;
  assign n20954 = n8736 ^ n4754 ^ 1'b0 ;
  assign n20955 = ( ~n453 & n5054 ) | ( ~n453 & n6983 ) | ( n5054 & n6983 ) ;
  assign n20956 = n8447 ^ n1658 ^ 1'b0 ;
  assign n20957 = ~n10781 & n13139 ;
  assign n20959 = n2161 & n8271 ;
  assign n20958 = n213 | n17774 ;
  assign n20960 = n20959 ^ n20958 ^ 1'b0 ;
  assign n20961 = n15210 | n20960 ;
  assign n20962 = n8960 ^ n4161 ^ n1380 ;
  assign n20963 = n20962 ^ n141 ^ 1'b0 ;
  assign n20964 = ~n8903 & n20963 ;
  assign n20965 = n18387 & n20964 ;
  assign n20966 = n14403 ^ n7449 ^ 1'b0 ;
  assign n20967 = n1046 & ~n20966 ;
  assign n20968 = n6500 & ~n14211 ;
  assign n20969 = n12954 ^ n5551 ^ 1'b0 ;
  assign n20970 = n6635 | n12690 ;
  assign n20971 = n10491 & ~n20970 ;
  assign n20976 = n2367 ^ n2216 ^ 1'b0 ;
  assign n20977 = n9813 | n20976 ;
  assign n20972 = n5122 ^ n1035 ^ 1'b0 ;
  assign n20973 = ~n17380 & n20972 ;
  assign n20974 = n13124 & n20973 ;
  assign n20975 = n19656 | n20974 ;
  assign n20978 = n20977 ^ n20975 ^ 1'b0 ;
  assign n20979 = n7275 ^ n3112 ^ n1346 ;
  assign n20980 = n20979 ^ n2640 ^ 1'b0 ;
  assign n20981 = n15591 | n20980 ;
  assign n20982 = n20981 ^ n14906 ^ 1'b0 ;
  assign n20983 = n12028 & ~n20982 ;
  assign n20984 = n10851 ^ n10835 ^ 1'b0 ;
  assign n20985 = n10131 & n16738 ;
  assign n20986 = ~n2987 & n9178 ;
  assign n20987 = n20986 ^ n15079 ^ 1'b0 ;
  assign n20988 = n5876 & n17906 ;
  assign n20989 = n14688 ^ n3558 ^ n710 ;
  assign n20990 = n3894 ^ n1320 ^ n450 ;
  assign n20991 = n7636 ^ n7165 ^ 1'b0 ;
  assign n20992 = n7087 | n20121 ;
  assign n20993 = n20991 | n20992 ;
  assign n20994 = n8055 & n16641 ;
  assign n20995 = n670 & n20994 ;
  assign n20996 = n20995 ^ n2638 ^ 1'b0 ;
  assign n20997 = n8945 | n20996 ;
  assign n20998 = n10568 & ~n19828 ;
  assign n21010 = n15 | n6008 ;
  assign n21011 = n9453 ^ n9264 ^ 1'b0 ;
  assign n21012 = n21010 | n21011 ;
  assign n21000 = n2967 | n5284 ;
  assign n20999 = n514 & ~n3093 ;
  assign n21001 = n21000 ^ n20999 ^ 1'b0 ;
  assign n21002 = ~n5475 & n21001 ;
  assign n21003 = n14305 & n21002 ;
  assign n21004 = n18605 & ~n21003 ;
  assign n21005 = n21004 ^ n16132 ^ 1'b0 ;
  assign n21006 = n7795 ^ n5227 ^ 1'b0 ;
  assign n21007 = n12481 & ~n21006 ;
  assign n21008 = ~n9713 & n21007 ;
  assign n21009 = n21005 & n21008 ;
  assign n21013 = n21012 ^ n21009 ^ 1'b0 ;
  assign n21014 = n2048 & n4377 ;
  assign n21015 = n21014 ^ n15127 ^ 1'b0 ;
  assign n21016 = n13740 ^ n10939 ^ 1'b0 ;
  assign n21019 = n10731 ^ n4339 ^ n3734 ;
  assign n21020 = n16169 ^ n15736 ^ 1'b0 ;
  assign n21021 = n21019 & n21020 ;
  assign n21017 = n3837 | n10576 ;
  assign n21018 = n19621 & n21017 ;
  assign n21022 = n21021 ^ n21018 ^ 1'b0 ;
  assign n21023 = n14312 ^ n1932 ^ 1'b0 ;
  assign n21024 = ~n8821 & n21023 ;
  assign n21025 = n21024 ^ n3803 ^ 1'b0 ;
  assign n21028 = n4869 & ~n9055 ;
  assign n21029 = ~n909 & n21028 ;
  assign n21026 = ~x10 & n3644 ;
  assign n21027 = ~n6801 & n21026 ;
  assign n21030 = n21029 ^ n21027 ^ 1'b0 ;
  assign n21031 = ( n10008 & n10900 ) | ( n10008 & ~n13574 ) | ( n10900 & ~n13574 ) ;
  assign n21032 = n4394 & ~n14373 ;
  assign n21033 = n21032 ^ n11142 ^ 1'b0 ;
  assign n21035 = ( n4911 & ~n14912 ) | ( n4911 & n15736 ) | ( ~n14912 & n15736 ) ;
  assign n21036 = n570 | n21035 ;
  assign n21037 = n21036 ^ n6602 ^ 1'b0 ;
  assign n21034 = n10170 & ~n15320 ;
  assign n21038 = n21037 ^ n21034 ^ 1'b0 ;
  assign n21039 = n617 | n19503 ;
  assign n21040 = n21038 | n21039 ;
  assign n21041 = n11756 ^ n2510 ^ 1'b0 ;
  assign n21046 = n769 | n4701 ;
  assign n21042 = n4354 ^ n437 ^ 1'b0 ;
  assign n21043 = n18404 | n21042 ;
  assign n21044 = n3386 | n21043 ;
  assign n21045 = n7680 | n21044 ;
  assign n21047 = n21046 ^ n21045 ^ 1'b0 ;
  assign n21048 = ~n15173 & n21047 ;
  assign n21049 = n11347 ^ n6196 ^ 1'b0 ;
  assign n21050 = ~n15323 & n21049 ;
  assign n21051 = n21048 & n21050 ;
  assign n21052 = n21041 & n21051 ;
  assign n21053 = n1339 & n9373 ;
  assign n21054 = n21053 ^ n336 ^ 1'b0 ;
  assign n21055 = n21054 ^ n14865 ^ 1'b0 ;
  assign n21056 = n2257 & ~n21055 ;
  assign n21057 = n304 & n452 ;
  assign n21058 = ~n153 & n21057 ;
  assign n21059 = n1786 | n6681 ;
  assign n21060 = n21059 ^ n12815 ^ 1'b0 ;
  assign n21061 = n21060 ^ n20971 ^ n10325 ;
  assign n21062 = n2768 & n8215 ;
  assign n21063 = n668 | n14239 ;
  assign n21064 = n21062 | n21063 ;
  assign n21065 = n5279 & n21064 ;
  assign n21066 = ( n224 & n551 ) | ( n224 & ~n1414 ) | ( n551 & ~n1414 ) ;
  assign n21068 = n4818 & ~n16940 ;
  assign n21069 = ~n9285 & n21068 ;
  assign n21067 = ( ~n11205 & n11731 ) | ( ~n11205 & n14714 ) | ( n11731 & n14714 ) ;
  assign n21070 = n21069 ^ n21067 ^ 1'b0 ;
  assign n21071 = n12934 ^ n1817 ^ 1'b0 ;
  assign n21072 = n14848 & ~n21071 ;
  assign n21073 = n10794 ^ n1348 ^ n1121 ;
  assign n21074 = n100 & ~n7765 ;
  assign n21075 = n6447 ^ n5066 ^ n3398 ;
  assign n21076 = n9964 & ~n21075 ;
  assign n21077 = n3295 & n10870 ;
  assign n21078 = n15317 ^ n7710 ^ n782 ;
  assign n21079 = ~n12712 & n21078 ;
  assign n21080 = n11088 ^ n9520 ^ 1'b0 ;
  assign n21081 = n4144 & ~n21080 ;
  assign n21082 = n2895 & ~n16642 ;
  assign n21083 = n21082 ^ n13362 ^ 1'b0 ;
  assign n21084 = n21081 & n21083 ;
  assign n21085 = n14170 & n17496 ;
  assign n21086 = n13327 ^ n9104 ^ 1'b0 ;
  assign n21087 = n21085 & ~n21086 ;
  assign n21088 = n3881 | n18410 ;
  assign n21089 = n12355 | n21088 ;
  assign n21090 = ~n706 & n21089 ;
  assign n21091 = n17792 & n18146 ;
  assign n21092 = n6306 & n21091 ;
  assign n21096 = n132 | n772 ;
  assign n21097 = n132 & ~n21096 ;
  assign n21098 = n557 | n21097 ;
  assign n21099 = n557 & ~n21098 ;
  assign n21100 = n1859 | n21099 ;
  assign n21101 = n1859 & ~n21100 ;
  assign n21102 = n1724 & ~n21101 ;
  assign n21103 = ~n1724 & n21102 ;
  assign n21104 = n446 | n21103 ;
  assign n21105 = n446 & ~n21104 ;
  assign n21106 = n1032 | n6867 ;
  assign n21107 = n1032 & ~n21106 ;
  assign n21108 = n21105 | n21107 ;
  assign n21109 = n21105 & ~n21108 ;
  assign n21110 = n3327 | n5006 ;
  assign n21111 = ~n21109 & n21110 ;
  assign n21112 = n21109 & n21111 ;
  assign n21093 = n4317 & ~n6322 ;
  assign n21094 = n6322 & n21093 ;
  assign n21095 = n2357 & ~n21094 ;
  assign n21113 = n21112 ^ n21095 ^ 1'b0 ;
  assign n21114 = n4710 ^ n4272 ^ n4072 ;
  assign n21115 = n2805 | n21114 ;
  assign n21116 = n491 | n21115 ;
  assign n21117 = n5324 & n21116 ;
  assign n21118 = n1633 & ~n4140 ;
  assign n21119 = n15730 & n21118 ;
  assign n21120 = n7138 & n21119 ;
  assign n21122 = n59 | n19928 ;
  assign n21123 = n63 & ~n21122 ;
  assign n21121 = n5182 & ~n9274 ;
  assign n21124 = n21123 ^ n21121 ^ 1'b0 ;
  assign n21127 = n7914 ^ n5815 ^ 1'b0 ;
  assign n21125 = n7867 & n9332 ;
  assign n21126 = ~n17872 & n21125 ;
  assign n21128 = n21127 ^ n21126 ^ 1'b0 ;
  assign n21129 = ~n135 & n940 ;
  assign n21130 = ~n2999 & n21129 ;
  assign n21131 = n21130 ^ n13258 ^ 1'b0 ;
  assign n21132 = ~n4251 & n10965 ;
  assign n21133 = n2432 | n2720 ;
  assign n21134 = n21132 & ~n21133 ;
  assign n21135 = n1596 | n21134 ;
  assign n21136 = n10478 ^ n8826 ^ n7836 ;
  assign n21137 = n3537 ^ n776 ^ 1'b0 ;
  assign n21138 = n435 & n21137 ;
  assign n21139 = n13752 & n21138 ;
  assign n21140 = n7529 & ~n21139 ;
  assign n21141 = n3432 & ~n6073 ;
  assign n21142 = n21140 & n21141 ;
  assign n21143 = n14852 & ~n16313 ;
  assign n21144 = n21143 ^ n6526 ^ 1'b0 ;
  assign n21145 = n355 | n21144 ;
  assign n21146 = n8418 ^ n7128 ^ n1084 ;
  assign n21147 = n139 | n11829 ;
  assign n21148 = ~n7039 & n17952 ;
  assign n21149 = n21148 ^ n4767 ^ 1'b0 ;
  assign n21150 = n12828 ^ n78 ^ 1'b0 ;
  assign n21151 = ~n5773 & n21150 ;
  assign n21152 = ~n11196 & n21151 ;
  assign n21153 = n10436 & n21152 ;
  assign n21154 = n10186 & n13945 ;
  assign n21155 = n21154 ^ n1805 ^ 1'b0 ;
  assign n21156 = n21155 ^ n11989 ^ 1'b0 ;
  assign n21157 = ~n2923 & n4196 ;
  assign n21158 = n21157 ^ n17013 ^ 1'b0 ;
  assign n21159 = n3341 | n5725 ;
  assign n21160 = n2667 & ~n21159 ;
  assign n21161 = n21160 ^ n12860 ^ 1'b0 ;
  assign n21162 = ~n4297 & n10213 ;
  assign n21165 = n2162 ^ n1047 ^ 1'b0 ;
  assign n21163 = n10720 ^ n4596 ^ 1'b0 ;
  assign n21164 = n5124 | n21163 ;
  assign n21166 = n21165 ^ n21164 ^ 1'b0 ;
  assign n21167 = n8395 ^ n2836 ^ 1'b0 ;
  assign n21168 = n11544 ^ n2449 ^ n225 ;
  assign n21169 = n1310 | n2332 ;
  assign n21170 = n21169 ^ n12882 ^ 1'b0 ;
  assign n21171 = n21168 | n21170 ;
  assign n21172 = n21171 ^ n17974 ^ n12925 ;
  assign n21173 = n9134 & ~n21172 ;
  assign n21174 = n13406 & n21173 ;
  assign n21175 = n13560 | n19660 ;
  assign n21176 = n2216 & ~n3912 ;
  assign n21177 = n10883 ^ n3517 ^ 1'b0 ;
  assign n21178 = n21176 | n21177 ;
  assign n21179 = n10183 | n15145 ;
  assign n21180 = n21179 ^ n18285 ^ 1'b0 ;
  assign n21181 = ~n5244 & n5841 ;
  assign n21182 = n691 | n5589 ;
  assign n21187 = n12562 ^ n2144 ^ 1'b0 ;
  assign n21188 = n5088 & ~n21187 ;
  assign n21189 = n5042 | n7011 ;
  assign n21190 = n21188 | n21189 ;
  assign n21183 = ~n1461 & n3890 ;
  assign n21184 = n13243 ^ n6027 ^ n853 ;
  assign n21185 = n21184 ^ n9722 ^ n37 ;
  assign n21186 = n21183 & ~n21185 ;
  assign n21191 = n21190 ^ n21186 ^ 1'b0 ;
  assign n21192 = n14049 ^ n10192 ^ 1'b0 ;
  assign n21193 = n1092 & n21192 ;
  assign n21194 = ~n1921 & n11446 ;
  assign n21195 = ~n21193 & n21194 ;
  assign n21196 = n12079 ^ n7599 ^ n710 ;
  assign n21200 = n1456 & n10647 ;
  assign n21201 = n21200 ^ n6241 ^ 1'b0 ;
  assign n21197 = n5660 & n12951 ;
  assign n21198 = n21197 ^ n8872 ^ 1'b0 ;
  assign n21199 = n9063 & ~n21198 ;
  assign n21202 = n21201 ^ n21199 ^ 1'b0 ;
  assign n21203 = n2028 | n5337 ;
  assign n21204 = n15781 | n21203 ;
  assign n21205 = n670 & ~n5037 ;
  assign n21206 = n13673 ^ n8122 ^ 1'b0 ;
  assign n21207 = n21206 ^ n20189 ^ 1'b0 ;
  assign n21208 = n2531 & n21207 ;
  assign n21209 = n1231 ^ n676 ^ 1'b0 ;
  assign n21210 = n20471 | n21209 ;
  assign n21211 = ~n157 & n1909 ;
  assign n21212 = n21211 ^ n3676 ^ 1'b0 ;
  assign n21213 = ( n1550 & n10624 ) | ( n1550 & n21212 ) | ( n10624 & n21212 ) ;
  assign n21214 = n21210 & n21213 ;
  assign n21215 = n2452 | n5630 ;
  assign n21216 = n1746 | n21215 ;
  assign n21217 = ~n786 & n21216 ;
  assign n21218 = n20638 ^ n1267 ^ 1'b0 ;
  assign n21219 = n5912 | n21218 ;
  assign n21220 = n20339 & ~n21219 ;
  assign n21221 = n2027 & ~n21220 ;
  assign n21222 = ~n17776 & n20299 ;
  assign n21223 = ( n2365 & n13946 ) | ( n2365 & ~n19660 ) | ( n13946 & ~n19660 ) ;
  assign n21224 = n11201 & n20736 ;
  assign n21230 = n448 & n17278 ;
  assign n21228 = ( ~n5173 & n8919 ) | ( ~n5173 & n14347 ) | ( n8919 & n14347 ) ;
  assign n21229 = n2621 | n21228 ;
  assign n21231 = n21230 ^ n21229 ^ 1'b0 ;
  assign n21225 = n3079 & n8082 ;
  assign n21226 = n17993 ^ n15794 ^ n10425 ;
  assign n21227 = n21225 | n21226 ;
  assign n21232 = n21231 ^ n21227 ^ 1'b0 ;
  assign n21233 = n13990 ^ n9369 ^ 1'b0 ;
  assign n21234 = n7634 ^ n7614 ^ 1'b0 ;
  assign n21235 = n12536 ^ n9286 ^ 1'b0 ;
  assign n21236 = n9096 & n21235 ;
  assign n21237 = ~n991 & n8323 ;
  assign n21238 = n21237 ^ n13136 ^ 1'b0 ;
  assign n21239 = n21238 ^ n7477 ^ 1'b0 ;
  assign n21240 = ~n7137 & n21239 ;
  assign n21241 = n1723 | n2569 ;
  assign n21242 = n7261 ^ n1632 ^ 1'b0 ;
  assign n21243 = n8085 | n18482 ;
  assign n21244 = n21242 | n21243 ;
  assign n21245 = ( ~n16998 & n21241 ) | ( ~n16998 & n21244 ) | ( n21241 & n21244 ) ;
  assign n21246 = ~n2217 & n10667 ;
  assign n21247 = n11000 ^ x3 ^ 1'b0 ;
  assign n21248 = n12519 & n21247 ;
  assign n21249 = ~n15046 & n21248 ;
  assign n21250 = n21249 ^ n6497 ^ 1'b0 ;
  assign n21260 = n7488 ^ n5076 ^ n3089 ;
  assign n21251 = n8954 & n10790 ;
  assign n21252 = n7943 ^ n6508 ^ 1'b0 ;
  assign n21253 = ~n2469 & n21252 ;
  assign n21254 = n9130 | n21253 ;
  assign n21255 = n7587 & n7701 ;
  assign n21256 = n21255 ^ n1856 ^ 1'b0 ;
  assign n21257 = ( ~n5595 & n7255 ) | ( ~n5595 & n21256 ) | ( n7255 & n21256 ) ;
  assign n21258 = n21257 ^ n6990 ^ 1'b0 ;
  assign n21259 = ( n21251 & n21254 ) | ( n21251 & n21258 ) | ( n21254 & n21258 ) ;
  assign n21261 = n21260 ^ n21259 ^ n868 ;
  assign n21262 = n14484 ^ n1035 ^ 1'b0 ;
  assign n21263 = ~n14889 & n14980 ;
  assign n21264 = n9431 & n21263 ;
  assign n21265 = n2510 & ~n21264 ;
  assign n21266 = n21262 & n21265 ;
  assign n21267 = n21266 ^ n9416 ^ 1'b0 ;
  assign n21268 = n12288 ^ n6479 ^ 1'b0 ;
  assign n21269 = ~n9947 & n21268 ;
  assign n21270 = ~n1362 & n2176 ;
  assign n21271 = n21270 ^ n1024 ^ 1'b0 ;
  assign n21272 = ~n6201 & n21271 ;
  assign n21273 = n6201 & n21272 ;
  assign n21274 = n484 | n1013 ;
  assign n21275 = n1013 & ~n21274 ;
  assign n21276 = n1787 | n21275 ;
  assign n21277 = n21275 & ~n21276 ;
  assign n21278 = n8114 | n21277 ;
  assign n21279 = n57 & n1210 ;
  assign n21280 = ~n1210 & n21279 ;
  assign n21281 = n21278 | n21280 ;
  assign n21282 = n21278 & ~n21281 ;
  assign n21283 = n2422 | n21282 ;
  assign n21284 = n21282 & ~n21283 ;
  assign n21285 = n5359 & ~n21284 ;
  assign n21286 = ~n5359 & n21285 ;
  assign n21287 = ( n19510 & n21273 ) | ( n19510 & n21286 ) | ( n21273 & n21286 ) ;
  assign n21288 = ~n5796 & n16483 ;
  assign n21289 = n364 & n21288 ;
  assign n21290 = n8485 & n9027 ;
  assign n21291 = n14825 | n21290 ;
  assign n21292 = n21291 ^ n10862 ^ 1'b0 ;
  assign n21293 = n5159 & n14067 ;
  assign n21294 = n21293 ^ n7558 ^ 1'b0 ;
  assign n21295 = n21294 ^ n5024 ^ 1'b0 ;
  assign n21296 = n14644 ^ n11330 ^ 1'b0 ;
  assign n21297 = ~n1676 & n14291 ;
  assign n21298 = n15 & n772 ;
  assign n21299 = n8355 & n21298 ;
  assign n21300 = n21299 ^ n8258 ^ 1'b0 ;
  assign n21301 = n10044 | n21300 ;
  assign n21302 = n571 & n21301 ;
  assign n21303 = n800 & ~n7234 ;
  assign n21304 = n21303 ^ x5 ^ 1'b0 ;
  assign n21305 = n21304 ^ n1332 ^ 1'b0 ;
  assign n21306 = n20430 ^ n2476 ^ 1'b0 ;
  assign n21307 = n5373 | n21306 ;
  assign n21311 = n6271 ^ n5864 ^ n586 ;
  assign n21312 = n7214 ^ n2513 ^ 1'b0 ;
  assign n21313 = n5227 & ~n21312 ;
  assign n21314 = n7043 & ~n21313 ;
  assign n21315 = n21311 & n21314 ;
  assign n21316 = ( ~n255 & n1641 ) | ( ~n255 & n8618 ) | ( n1641 & n8618 ) ;
  assign n21317 = ~n21315 & n21316 ;
  assign n21308 = n16223 ^ n848 ^ 1'b0 ;
  assign n21309 = ~n7448 & n21308 ;
  assign n21310 = n18839 & n21309 ;
  assign n21318 = n21317 ^ n21310 ^ 1'b0 ;
  assign n21319 = n976 & ~n13246 ;
  assign n21326 = n7705 ^ n5225 ^ 1'b0 ;
  assign n21327 = n21326 ^ n15439 ^ 1'b0 ;
  assign n21328 = x10 & n21327 ;
  assign n21323 = n7003 & ~n9078 ;
  assign n21324 = n12327 ^ n12322 ^ 1'b0 ;
  assign n21325 = n21323 & ~n21324 ;
  assign n21320 = n4658 ^ n2791 ^ 1'b0 ;
  assign n21321 = n6670 & n21320 ;
  assign n21322 = n21321 ^ n7158 ^ 1'b0 ;
  assign n21329 = n21328 ^ n21325 ^ n21322 ;
  assign n21334 = ~n790 & n5325 ;
  assign n21335 = n21334 ^ n16368 ^ 1'b0 ;
  assign n21336 = ( n3138 & n3885 ) | ( n3138 & ~n21335 ) | ( n3885 & ~n21335 ) ;
  assign n21337 = n10533 & n12906 ;
  assign n21338 = n17954 & n21337 ;
  assign n21339 = n21336 & n21338 ;
  assign n21330 = n11596 ^ n4773 ^ 1'b0 ;
  assign n21331 = n9199 | n21330 ;
  assign n21332 = n21331 ^ n6705 ^ n356 ;
  assign n21333 = ~n17685 & n21332 ;
  assign n21340 = n21339 ^ n21333 ^ 1'b0 ;
  assign n21341 = n3484 | n18099 ;
  assign n21342 = n5380 & ~n21341 ;
  assign n21343 = n6625 & ~n12022 ;
  assign n21344 = n7642 & ~n13643 ;
  assign n21347 = n5466 ^ n4204 ^ 1'b0 ;
  assign n21348 = n21347 ^ n7115 ^ 1'b0 ;
  assign n21349 = ( ~n3079 & n13175 ) | ( ~n3079 & n21348 ) | ( n13175 & n21348 ) ;
  assign n21345 = n5337 | n5693 ;
  assign n21346 = n362 | n21345 ;
  assign n21350 = n21349 ^ n21346 ^ 1'b0 ;
  assign n21351 = n6153 & n6935 ;
  assign n21352 = ~n4399 & n21351 ;
  assign n21353 = n21352 ^ n5339 ^ 1'b0 ;
  assign n21354 = n18258 ^ n6473 ^ 1'b0 ;
  assign n21355 = n3467 | n14898 ;
  assign n21356 = n4520 ^ n3742 ^ 1'b0 ;
  assign n21357 = n21355 & n21356 ;
  assign n21358 = n16917 & n18230 ;
  assign n21359 = n829 & ~n16215 ;
  assign n21360 = n21359 ^ n19455 ^ 1'b0 ;
  assign n21361 = ( ~n3082 & n4110 ) | ( ~n3082 & n16799 ) | ( n4110 & n16799 ) ;
  assign n21362 = n6277 ^ n3665 ^ 1'b0 ;
  assign n21363 = ~n8470 & n21362 ;
  assign n21364 = n21363 ^ n5576 ^ 1'b0 ;
  assign n21365 = n2859 | n21364 ;
  assign n21366 = ( n688 & n15926 ) | ( n688 & ~n21365 ) | ( n15926 & ~n21365 ) ;
  assign n21367 = n21361 & n21366 ;
  assign n21368 = n11360 & n15632 ;
  assign n21369 = n21368 ^ n4004 ^ 1'b0 ;
  assign n21370 = ~n21367 & n21369 ;
  assign n21371 = n5309 ^ n1666 ^ n1312 ;
  assign n21372 = n13737 & n21371 ;
  assign n21373 = n21372 ^ n1694 ^ 1'b0 ;
  assign n21374 = n21373 ^ n4659 ^ 1'b0 ;
  assign n21375 = ~n19526 & n21374 ;
  assign n21376 = n712 ^ x6 ^ 1'b0 ;
  assign n21377 = ( n1944 & ~n2819 ) | ( n1944 & n21376 ) | ( ~n2819 & n21376 ) ;
  assign n21378 = n829 ^ n543 ^ 1'b0 ;
  assign n21379 = n11321 & n21378 ;
  assign n21380 = n18867 & n21379 ;
  assign n21381 = n5741 & n12119 ;
  assign n21382 = n17222 ^ n15013 ^ 1'b0 ;
  assign n21383 = n20160 ^ n17916 ^ n6227 ;
  assign n21384 = n18085 ^ n6940 ^ 1'b0 ;
  assign n21385 = n3566 & n21384 ;
  assign n21386 = n5873 ^ n3295 ^ 1'b0 ;
  assign n21387 = ~n263 & n21386 ;
  assign n21388 = ( n1350 & ~n12219 ) | ( n1350 & n21387 ) | ( ~n12219 & n21387 ) ;
  assign n21389 = n18169 ^ n2335 ^ 1'b0 ;
  assign n21390 = n21388 | n21389 ;
  assign n21391 = ( n1063 & n8824 ) | ( n1063 & n13567 ) | ( n8824 & n13567 ) ;
  assign n21392 = n21391 ^ n3738 ^ 1'b0 ;
  assign n21393 = n4665 ^ n3071 ^ 1'b0 ;
  assign n21394 = n21393 ^ n14167 ^ n8688 ;
  assign n21395 = n4797 & n13312 ;
  assign n21396 = ( n8154 & n21394 ) | ( n8154 & ~n21395 ) | ( n21394 & ~n21395 ) ;
  assign n21397 = n18401 ^ n11102 ^ n7531 ;
  assign n21398 = n17407 ^ n4057 ^ 1'b0 ;
  assign n21399 = n21398 ^ n3870 ^ 1'b0 ;
  assign n21400 = n19698 | n21399 ;
  assign n21401 = n764 ^ n115 ^ 1'b0 ;
  assign n21402 = n14936 ^ n6696 ^ 1'b0 ;
  assign n21403 = n20352 | n21402 ;
  assign n21404 = n21403 ^ n5997 ^ 1'b0 ;
  assign n21405 = n21401 & ~n21404 ;
  assign n21406 = n11666 ^ n3010 ^ 1'b0 ;
  assign n21407 = ~n7280 & n21406 ;
  assign n21408 = n11331 | n12393 ;
  assign n21410 = n14700 ^ n1082 ^ 1'b0 ;
  assign n21409 = n17640 ^ n3785 ^ 1'b0 ;
  assign n21411 = n21410 ^ n21409 ^ 1'b0 ;
  assign n21412 = ( ~n2636 & n4789 ) | ( ~n2636 & n21411 ) | ( n4789 & n21411 ) ;
  assign n21413 = n18519 ^ n40 ^ 1'b0 ;
  assign n21414 = n12915 ^ n6937 ^ 1'b0 ;
  assign n21415 = n7253 ^ n4916 ^ 1'b0 ;
  assign n21416 = n21414 | n21415 ;
  assign n21417 = n9211 | n12153 ;
  assign n21418 = n2650 ^ n2100 ^ 1'b0 ;
  assign n21419 = ( n2190 & n9144 ) | ( n2190 & n21418 ) | ( n9144 & n21418 ) ;
  assign n21420 = n11809 & ~n21419 ;
  assign n21421 = n21420 ^ n16409 ^ 1'b0 ;
  assign n21422 = n10402 | n11844 ;
  assign n21423 = n21422 ^ n9902 ^ 1'b0 ;
  assign n21424 = ~n151 & n639 ;
  assign n21425 = n12197 & ~n17640 ;
  assign n21426 = n21424 | n21425 ;
  assign n21427 = n17424 | n21426 ;
  assign n21429 = n15367 & ~n19303 ;
  assign n21430 = n4259 ^ n3475 ^ 1'b0 ;
  assign n21431 = ~n21429 & n21430 ;
  assign n21428 = n8778 & n16965 ;
  assign n21432 = n21431 ^ n21428 ^ 1'b0 ;
  assign n21433 = n15982 ^ n5682 ^ 1'b0 ;
  assign n21434 = ( n2745 & n4025 ) | ( n2745 & n4745 ) | ( n4025 & n4745 ) ;
  assign n21435 = ( n3428 & n10949 ) | ( n3428 & ~n21434 ) | ( n10949 & ~n21434 ) ;
  assign n21436 = n16295 & n21435 ;
  assign n21437 = ~n21433 & n21436 ;
  assign n21438 = n21437 ^ n16811 ^ 1'b0 ;
  assign n21439 = ~n3582 & n21438 ;
  assign n21444 = n4376 & ~n7830 ;
  assign n21445 = ( n10093 & n12966 ) | ( n10093 & ~n21444 ) | ( n12966 & ~n21444 ) ;
  assign n21440 = n3181 ^ n1061 ^ 1'b0 ;
  assign n21441 = n1320 & n21440 ;
  assign n21442 = ~n16149 & n21441 ;
  assign n21443 = n21442 ^ n1267 ^ 1'b0 ;
  assign n21446 = n21445 ^ n21443 ^ 1'b0 ;
  assign n21447 = n12123 | n16115 ;
  assign n21448 = ~n1603 & n11314 ;
  assign n21449 = n5125 ^ n1633 ^ n654 ;
  assign n21454 = n734 & n1281 ;
  assign n21450 = n2186 ^ n498 ^ 1'b0 ;
  assign n21451 = n3687 & ~n21450 ;
  assign n21452 = n21451 ^ n483 ^ 1'b0 ;
  assign n21453 = n9589 & n21452 ;
  assign n21455 = n21454 ^ n21453 ^ n8485 ;
  assign n21456 = n21455 ^ n2670 ^ 1'b0 ;
  assign n21457 = n21449 & ~n21456 ;
  assign n21458 = n21457 ^ n14106 ^ 1'b0 ;
  assign n21459 = ~n5255 & n21458 ;
  assign n21460 = n15498 | n19296 ;
  assign n21461 = n21460 ^ n1064 ^ 1'b0 ;
  assign n21462 = ~n8159 & n21461 ;
  assign n21463 = n7976 ^ n5028 ^ n373 ;
  assign n21464 = n21463 ^ n6485 ^ 1'b0 ;
  assign n21465 = n15937 | n21464 ;
  assign n21466 = n11443 ^ n2666 ^ 1'b0 ;
  assign n21467 = ~n12683 & n21466 ;
  assign n21475 = n11511 ^ n11389 ^ 1'b0 ;
  assign n21472 = n1856 ^ n1605 ^ 1'b0 ;
  assign n21473 = n5069 | n21472 ;
  assign n21468 = n17855 ^ n7739 ^ 1'b0 ;
  assign n21469 = ~n5866 & n21468 ;
  assign n21470 = n5582 & n21469 ;
  assign n21471 = n5696 & n21470 ;
  assign n21474 = n21473 ^ n21471 ^ 1'b0 ;
  assign n21476 = n21475 ^ n21474 ^ 1'b0 ;
  assign n21477 = n21476 ^ n17275 ^ 1'b0 ;
  assign n21478 = n10939 | n21477 ;
  assign n21479 = n17643 | n21182 ;
  assign n21480 = n21479 ^ n8041 ^ 1'b0 ;
  assign n21481 = n14131 ^ n3016 ^ 1'b0 ;
  assign n21482 = n9487 & ~n21481 ;
  assign n21483 = n3053 & n21482 ;
  assign n21486 = ( ~n5576 & n9330 ) | ( ~n5576 & n18423 ) | ( n9330 & n18423 ) ;
  assign n21487 = n21486 ^ n7316 ^ 1'b0 ;
  assign n21488 = n11282 & n21487 ;
  assign n21484 = n4807 | n4957 ;
  assign n21485 = n21484 ^ n12124 ^ 1'b0 ;
  assign n21489 = n21488 ^ n21485 ^ n6426 ;
  assign n21490 = n8847 | n14041 ;
  assign n21491 = n1489 & n14524 ;
  assign n21492 = n21491 ^ x6 ^ 1'b0 ;
  assign n21493 = n6817 & ~n17601 ;
  assign n21494 = ~n2765 & n21493 ;
  assign n21495 = ~n21492 & n21494 ;
  assign n21496 = n18660 ^ n11827 ^ 1'b0 ;
  assign n21497 = n21495 & ~n21496 ;
  assign n21498 = n16597 ^ n10063 ^ n3495 ;
  assign n21499 = ~n16730 & n21498 ;
  assign n21500 = ~n15237 & n21499 ;
  assign n21501 = n289 & n21500 ;
  assign n21502 = n6956 ^ n5026 ^ 1'b0 ;
  assign n21503 = ~n3211 & n21502 ;
  assign n21504 = n145 & n882 ;
  assign n21505 = n1290 | n21504 ;
  assign n21506 = n21505 ^ n14163 ^ 1'b0 ;
  assign n21507 = n6045 & ~n7188 ;
  assign n21508 = n2960 & n21507 ;
  assign n21509 = n21506 & ~n21508 ;
  assign n21510 = n7337 & n21509 ;
  assign n21511 = n4835 ^ n36 ^ 1'b0 ;
  assign n21512 = ~n21510 & n21511 ;
  assign n21513 = ( n5095 & ~n14423 ) | ( n5095 & n21512 ) | ( ~n14423 & n21512 ) ;
  assign n21514 = n21513 ^ n14007 ^ 1'b0 ;
  assign n21515 = n5009 | n9555 ;
  assign n21516 = n1080 | n21515 ;
  assign n21517 = n21516 ^ n10233 ^ 1'b0 ;
  assign n21518 = ( n825 & n3435 ) | ( n825 & n3704 ) | ( n3435 & n3704 ) ;
  assign n21519 = n19677 & n21518 ;
  assign n21520 = n6039 ^ n2312 ^ 1'b0 ;
  assign n21521 = n21519 | n21520 ;
  assign n21522 = n15718 ^ n3334 ^ 1'b0 ;
  assign n21523 = n17650 ^ n16793 ^ 1'b0 ;
  assign n21524 = n11795 ^ n4772 ^ 1'b0 ;
  assign n21525 = n21523 & ~n21524 ;
  assign n21526 = n11323 ^ n10210 ^ 1'b0 ;
  assign n21527 = n14129 ^ n12166 ^ 1'b0 ;
  assign n21528 = n4796 | n21527 ;
  assign n21529 = n21528 ^ n10668 ^ 1'b0 ;
  assign n21530 = n16950 ^ n6878 ^ 1'b0 ;
  assign n21534 = n10295 ^ n9498 ^ n5975 ;
  assign n21531 = n3114 & ~n7251 ;
  assign n21532 = ~n6839 & n21531 ;
  assign n21533 = n10209 | n21532 ;
  assign n21535 = n21534 ^ n21533 ^ 1'b0 ;
  assign n21536 = n4894 & n9848 ;
  assign n21537 = ~n4894 & n21536 ;
  assign n21538 = n21537 ^ n11120 ^ 1'b0 ;
  assign n21539 = n21538 ^ n12418 ^ n10689 ;
  assign n21540 = n3154 & n3637 ;
  assign n21541 = n2784 | n2995 ;
  assign n21542 = n16145 ^ n14386 ^ 1'b0 ;
  assign n21543 = n609 & n21542 ;
  assign n21544 = n4339 & n9248 ;
  assign n21545 = n12371 ^ n8684 ^ 1'b0 ;
  assign n21546 = n9890 | n21545 ;
  assign n21551 = n2620 & n5219 ;
  assign n21552 = n21551 ^ n818 ^ 1'b0 ;
  assign n21549 = n3574 ^ n2330 ^ 1'b0 ;
  assign n21550 = n21549 ^ n1649 ^ 1'b0 ;
  assign n21553 = n21552 ^ n21550 ^ 1'b0 ;
  assign n21554 = n11014 | n21553 ;
  assign n21555 = n11117 | n21554 ;
  assign n21547 = n11904 ^ n788 ^ 1'b0 ;
  assign n21548 = ~n10311 & n21547 ;
  assign n21556 = n21555 ^ n21548 ^ n7221 ;
  assign n21557 = n7248 | n21556 ;
  assign n21559 = n5344 & ~n14024 ;
  assign n21558 = n4851 | n20181 ;
  assign n21560 = n21559 ^ n21558 ^ 1'b0 ;
  assign n21561 = ~n1509 & n21560 ;
  assign n21562 = n7128 ^ n1617 ^ 1'b0 ;
  assign n21563 = ~n11153 & n21562 ;
  assign n21564 = ~n3314 & n21563 ;
  assign n21565 = n1762 ^ n1749 ^ 1'b0 ;
  assign n21566 = n6302 ^ n181 ^ 1'b0 ;
  assign n21567 = ~n1350 & n21566 ;
  assign n21568 = n21567 ^ n1713 ^ 1'b0 ;
  assign n21570 = n929 & ~n7527 ;
  assign n21569 = n563 & n15490 ;
  assign n21571 = n21570 ^ n21569 ^ n13558 ;
  assign n21572 = n21568 & n21571 ;
  assign n21573 = n10187 & n21572 ;
  assign n21574 = n9921 ^ n4761 ^ 1'b0 ;
  assign n21575 = n19399 ^ n7112 ^ 1'b0 ;
  assign n21576 = n10940 & n12748 ;
  assign n21577 = n18656 | n21365 ;
  assign n21578 = n18897 ^ n1408 ^ 1'b0 ;
  assign n21579 = n830 | n5219 ;
  assign n21580 = n5645 & n14023 ;
  assign n21581 = n21580 ^ n8896 ^ 1'b0 ;
  assign n21582 = n6455 & n16058 ;
  assign n21583 = ~n21581 & n21582 ;
  assign n21584 = n3591 | n18169 ;
  assign n21585 = n6846 & n8043 ;
  assign n21586 = n10290 & n21585 ;
  assign n21587 = n19805 | n20164 ;
  assign n21588 = ~n10034 & n21587 ;
  assign n21589 = n21588 ^ n1694 ^ 1'b0 ;
  assign n21590 = n7756 | n16957 ;
  assign n21591 = n2211 | n21590 ;
  assign n21592 = n15493 ^ n13366 ^ 1'b0 ;
  assign n21593 = n13695 | n21592 ;
  assign n21594 = n14350 | n15972 ;
  assign n21595 = n7240 ^ n823 ^ 1'b0 ;
  assign n21599 = ~n864 & n4205 ;
  assign n21600 = n2418 & n21599 ;
  assign n21596 = n6093 & n8669 ;
  assign n21597 = n13046 & n21596 ;
  assign n21598 = ~n6020 & n21597 ;
  assign n21601 = n21600 ^ n21598 ^ 1'b0 ;
  assign n21602 = n965 & n15335 ;
  assign n21603 = n21602 ^ n8646 ^ 1'b0 ;
  assign n21604 = n1247 | n3782 ;
  assign n21605 = ~n21603 & n21604 ;
  assign n21606 = ~n615 & n7912 ;
  assign n21607 = n21606 ^ n1579 ^ 1'b0 ;
  assign n21608 = n21607 ^ n15433 ^ 1'b0 ;
  assign n21609 = n3506 | n21608 ;
  assign n21610 = n2391 | n21609 ;
  assign n21611 = ~n6787 & n21610 ;
  assign n21612 = ~n5896 & n17559 ;
  assign n21613 = n11396 ^ n332 ^ n245 ;
  assign n21614 = n21613 ^ n9230 ^ 1'b0 ;
  assign n21615 = n11347 & ~n21614 ;
  assign n21616 = ( n2174 & ~n9830 ) | ( n2174 & n21615 ) | ( ~n9830 & n21615 ) ;
  assign n21617 = ( n5352 & n12827 ) | ( n5352 & ~n14619 ) | ( n12827 & ~n14619 ) ;
  assign n21618 = ~n3041 & n10118 ;
  assign n21619 = ~n7280 & n21618 ;
  assign n21620 = ( n2137 & ~n14805 ) | ( n2137 & n21619 ) | ( ~n14805 & n21619 ) ;
  assign n21621 = n9150 ^ n3826 ^ 1'b0 ;
  assign n21622 = n3650 & ~n21621 ;
  assign n21623 = n7864 & n8576 ;
  assign n21624 = n2722 & n21623 ;
  assign n21625 = n21622 & n21624 ;
  assign n21626 = n6948 & ~n17608 ;
  assign n21627 = n3097 & n21626 ;
  assign n21628 = n8927 & ~n9134 ;
  assign n21629 = n6667 ^ n6406 ^ 1'b0 ;
  assign n21630 = n7256 | n21629 ;
  assign n21631 = n3544 & ~n6129 ;
  assign n21632 = n241 & n21631 ;
  assign n21633 = n21632 ^ n19971 ^ n1312 ;
  assign n21634 = n6628 & ~n14520 ;
  assign n21635 = ~n9253 & n21634 ;
  assign n21636 = n6988 & n21635 ;
  assign n21637 = n1542 & ~n7484 ;
  assign n21638 = n309 & n21637 ;
  assign n21639 = ~n16731 & n21638 ;
  assign n21640 = n16110 ^ n9437 ^ n8181 ;
  assign n21641 = n21640 ^ n14531 ^ n6249 ;
  assign n21642 = n771 & n21641 ;
  assign n21643 = n21639 & n21642 ;
  assign n21644 = n3372 & ~n12050 ;
  assign n21645 = n9950 & ~n21644 ;
  assign n21646 = n21645 ^ n5828 ^ 1'b0 ;
  assign n21647 = n11429 ^ n8406 ^ 1'b0 ;
  assign n21651 = n6386 ^ n4813 ^ n4712 ;
  assign n21650 = ~n73 & n5151 ;
  assign n21652 = n21651 ^ n21650 ^ 1'b0 ;
  assign n21648 = n6043 ^ n2882 ^ 1'b0 ;
  assign n21649 = n6887 & n21648 ;
  assign n21653 = n21652 ^ n21649 ^ 1'b0 ;
  assign n21654 = n13732 & n21653 ;
  assign n21655 = n21654 ^ n15285 ^ n3604 ;
  assign n21656 = n3514 & n12138 ;
  assign n21657 = n20540 ^ n10427 ^ 1'b0 ;
  assign n21658 = n21656 & n21657 ;
  assign n21659 = n9983 & ~n15732 ;
  assign n21660 = ~n8787 & n21659 ;
  assign n21661 = n926 | n2658 ;
  assign n21662 = n21661 ^ n10939 ^ 1'b0 ;
  assign n21663 = n1085 | n6804 ;
  assign n21664 = ( ~n7288 & n12449 ) | ( ~n7288 & n13754 ) | ( n12449 & n13754 ) ;
  assign n21665 = n21664 ^ n17283 ^ n9434 ;
  assign n21666 = n13261 & n18366 ;
  assign n21667 = n21666 ^ n4497 ^ 1'b0 ;
  assign n21668 = n7180 ^ n2901 ^ 1'b0 ;
  assign n21669 = ( ~n6947 & n21667 ) | ( ~n6947 & n21668 ) | ( n21667 & n21668 ) ;
  assign n21670 = n6648 ^ n2461 ^ 1'b0 ;
  assign n21671 = n4803 ^ n220 ^ 1'b0 ;
  assign n21672 = n21671 ^ n1545 ^ 1'b0 ;
  assign n21673 = n15640 & ~n19660 ;
  assign n21674 = n21673 ^ n20737 ^ 1'b0 ;
  assign n21675 = n13938 ^ n10192 ^ 1'b0 ;
  assign n21676 = n13378 | n21675 ;
  assign n21677 = ( ~n7087 & n12127 ) | ( ~n7087 & n21676 ) | ( n12127 & n21676 ) ;
  assign n21678 = n169 & n9919 ;
  assign n21679 = ~n15330 & n21678 ;
  assign n21680 = n21679 ^ n4944 ^ 1'b0 ;
  assign n21681 = n21680 ^ n8030 ^ n2677 ;
  assign n21682 = n5856 ^ n4388 ^ n2405 ;
  assign n21683 = n18393 ^ n4233 ^ 1'b0 ;
  assign n21684 = n7804 & ~n21683 ;
  assign n21685 = ~n21682 & n21684 ;
  assign n21686 = n76 | n3195 ;
  assign n21687 = n21686 ^ n1656 ^ 1'b0 ;
  assign n21688 = n4048 & n21687 ;
  assign n21689 = n8606 & ~n21688 ;
  assign n21690 = n21689 ^ n1538 ^ 1'b0 ;
  assign n21691 = n12923 ^ n10230 ^ n8485 ;
  assign n21693 = n10451 ^ n6060 ^ 1'b0 ;
  assign n21694 = n4038 & ~n21693 ;
  assign n21692 = n1962 & ~n19300 ;
  assign n21695 = n21694 ^ n21692 ^ 1'b0 ;
  assign n21696 = n9933 ^ n2664 ^ 1'b0 ;
  assign n21697 = n20526 ^ n15569 ^ 1'b0 ;
  assign n21698 = ~n2340 & n3329 ;
  assign n21699 = ~n7575 & n21698 ;
  assign n21700 = n10576 ^ n195 ^ 1'b0 ;
  assign n21701 = n850 & n11642 ;
  assign n21702 = n7670 | n11095 ;
  assign n21703 = n21701 | n21702 ;
  assign n21707 = n7828 ^ n2100 ^ 1'b0 ;
  assign n21704 = n7367 ^ n4890 ^ 1'b0 ;
  assign n21705 = n3762 | n21704 ;
  assign n21706 = n21705 ^ n4469 ^ 1'b0 ;
  assign n21708 = n21707 ^ n21706 ^ 1'b0 ;
  assign n21709 = n21703 & ~n21708 ;
  assign n21710 = ( n890 & n15912 ) | ( n890 & ~n21709 ) | ( n15912 & ~n21709 ) ;
  assign n21711 = n475 & ~n4544 ;
  assign n21712 = n21711 ^ n4804 ^ 1'b0 ;
  assign n21713 = n9444 ^ n9108 ^ 1'b0 ;
  assign n21714 = n21713 ^ n18940 ^ n6683 ;
  assign n21716 = n2001 & n6182 ;
  assign n21715 = n4706 | n17199 ;
  assign n21717 = n21716 ^ n21715 ^ 1'b0 ;
  assign n21718 = n4796 & n21717 ;
  assign n21719 = n8745 & n10270 ;
  assign n21720 = n21719 ^ n6278 ^ 1'b0 ;
  assign n21721 = ( n6406 & n13761 ) | ( n6406 & n21720 ) | ( n13761 & n21720 ) ;
  assign n21722 = n4873 ^ n4857 ^ 1'b0 ;
  assign n21723 = n10181 | n21722 ;
  assign n21724 = n21723 ^ n14972 ^ n2566 ;
  assign n21725 = n21724 ^ n20612 ^ 1'b0 ;
  assign n21726 = ~n3983 & n7976 ;
  assign n21727 = n9274 ^ n7219 ^ 1'b0 ;
  assign n21728 = n21726 & n21727 ;
  assign n21735 = n5968 & ~n8695 ;
  assign n21736 = n4436 & n21735 ;
  assign n21732 = ~n2853 & n9018 ;
  assign n21733 = ( n4812 & n9490 ) | ( n4812 & n21732 ) | ( n9490 & n21732 ) ;
  assign n21729 = n8015 ^ n6262 ^ 1'b0 ;
  assign n21730 = n2531 & ~n21729 ;
  assign n21731 = n4272 & n21730 ;
  assign n21734 = n21733 ^ n21731 ^ 1'b0 ;
  assign n21737 = n21736 ^ n21734 ^ 1'b0 ;
  assign n21738 = n7985 | n8089 ;
  assign n21739 = n11773 ^ n4096 ^ n2176 ;
  assign n21740 = ( n3638 & ~n10393 ) | ( n3638 & n11589 ) | ( ~n10393 & n11589 ) ;
  assign n21741 = n11942 & ~n16457 ;
  assign n21742 = n3951 & ~n21741 ;
  assign n21743 = n21608 & ~n21688 ;
  assign n21744 = ~n3225 & n15040 ;
  assign n21745 = n9452 & n20570 ;
  assign n21746 = ~n1693 & n21745 ;
  assign n21747 = ~n17741 & n21746 ;
  assign n21748 = n20371 ^ n8618 ^ 1'b0 ;
  assign n21749 = n8765 & ~n12918 ;
  assign n21750 = n21749 ^ n10353 ^ 1'b0 ;
  assign n21751 = ~n2089 & n21750 ;
  assign n21752 = ~n11128 & n21751 ;
  assign n21753 = n21752 ^ n14711 ^ 1'b0 ;
  assign n21754 = n16925 ^ n4032 ^ 1'b0 ;
  assign n21755 = n3439 & n5561 ;
  assign n21756 = n21755 ^ n6093 ^ 1'b0 ;
  assign n21757 = n21756 ^ n18069 ^ 1'b0 ;
  assign n21758 = n11378 & ~n16345 ;
  assign n21759 = n13932 & n21758 ;
  assign n21760 = ~n20628 & n21759 ;
  assign n21761 = n5057 ^ n3359 ^ n1543 ;
  assign n21762 = n6517 & n9072 ;
  assign n21763 = n21762 ^ n2667 ^ 1'b0 ;
  assign n21764 = ( n2597 & ~n16450 ) | ( n2597 & n17388 ) | ( ~n16450 & n17388 ) ;
  assign n21765 = n9372 ^ n2355 ^ 1'b0 ;
  assign n21766 = n8964 & ~n21765 ;
  assign n21767 = n4968 & n11806 ;
  assign n21768 = n21767 ^ n15714 ^ 1'b0 ;
  assign n21769 = ~n787 & n17332 ;
  assign n21770 = n21769 ^ n18704 ^ 1'b0 ;
  assign n21771 = n21770 ^ n20960 ^ 1'b0 ;
  assign n21772 = n11219 | n11811 ;
  assign n21773 = n21772 ^ n6815 ^ 1'b0 ;
  assign n21774 = n124 | n2958 ;
  assign n21775 = n8143 & ~n21774 ;
  assign n21776 = n5223 & ~n21775 ;
  assign n21777 = n19097 & n19439 ;
  assign n21778 = n21777 ^ n5940 ^ 1'b0 ;
  assign n21779 = n21778 ^ n8958 ^ 1'b0 ;
  assign n21780 = n21776 & ~n21779 ;
  assign n21781 = ~n1322 & n2836 ;
  assign n21782 = n21781 ^ n15306 ^ 1'b0 ;
  assign n21783 = n10802 | n12586 ;
  assign n21784 = n9057 | n21783 ;
  assign n21785 = ~n16950 & n21784 ;
  assign n21786 = n1495 & n19280 ;
  assign n21787 = n8597 & n21786 ;
  assign n21788 = n17990 | n21787 ;
  assign n21789 = n9151 ^ n3214 ^ 1'b0 ;
  assign n21790 = n21789 ^ n9487 ^ n4428 ;
  assign n21792 = n5228 & n7468 ;
  assign n21793 = ( n6888 & n11500 ) | ( n6888 & ~n21792 ) | ( n11500 & ~n21792 ) ;
  assign n21794 = ~n7276 & n21793 ;
  assign n21791 = n14131 ^ n7785 ^ 1'b0 ;
  assign n21795 = n21794 ^ n21791 ^ 1'b0 ;
  assign n21796 = n2797 & n13235 ;
  assign n21797 = n6034 & n21796 ;
  assign n21798 = n1784 ^ n201 ^ 1'b0 ;
  assign n21799 = n18078 ^ n9999 ^ 1'b0 ;
  assign n21800 = n21798 & ~n21799 ;
  assign n21801 = n19327 | n19928 ;
  assign n21802 = n17339 | n21801 ;
  assign n21803 = ~n14865 & n17118 ;
  assign n21804 = n4698 & ~n14721 ;
  assign n21807 = n13116 ^ n10143 ^ 1'b0 ;
  assign n21808 = n21807 ^ n15321 ^ n13491 ;
  assign n21809 = x10 & ~n10726 ;
  assign n21810 = n21808 & n21809 ;
  assign n21805 = ~n5396 & n11033 ;
  assign n21806 = ~n223 & n21805 ;
  assign n21811 = n21810 ^ n21806 ^ 1'b0 ;
  assign n21813 = n11389 ^ n5778 ^ 1'b0 ;
  assign n21812 = n2174 & ~n13714 ;
  assign n21814 = n21813 ^ n21812 ^ 1'b0 ;
  assign n21815 = n11846 ^ n7988 ^ n6675 ;
  assign n21816 = n14651 & n21815 ;
  assign n21824 = n15092 ^ n6601 ^ n5134 ;
  assign n21817 = n17906 ^ n5473 ^ n3973 ;
  assign n21818 = n21817 ^ n13775 ^ n9061 ;
  assign n21819 = n5054 | n15799 ;
  assign n21820 = n21819 ^ n181 ^ 1'b0 ;
  assign n21821 = n21818 & n21820 ;
  assign n21822 = n21821 ^ n4563 ^ 1'b0 ;
  assign n21823 = n21822 ^ n765 ^ 1'b0 ;
  assign n21825 = n21824 ^ n21823 ^ n11600 ;
  assign n21826 = n19727 ^ n14752 ^ n3049 ;
  assign n21827 = n9416 ^ n4143 ^ 1'b0 ;
  assign n21828 = ~n3571 & n21827 ;
  assign n21829 = ( ~n4538 & n12470 ) | ( ~n4538 & n21518 ) | ( n12470 & n21518 ) ;
  assign n21830 = n15338 ^ n5679 ^ 1'b0 ;
  assign n21831 = n19538 ^ n3906 ^ 1'b0 ;
  assign n21832 = n4221 & ~n21831 ;
  assign n21833 = ~n2148 & n21832 ;
  assign n21834 = ~n14777 & n21833 ;
  assign n21835 = ~n21830 & n21834 ;
  assign n21836 = n6466 | n18786 ;
  assign n21837 = ~n2589 & n13363 ;
  assign n21838 = n9986 & n21837 ;
  assign n21840 = ( n617 & n2214 ) | ( n617 & n4413 ) | ( n2214 & n4413 ) ;
  assign n21839 = n1786 | n6186 ;
  assign n21841 = n21840 ^ n21839 ^ 1'b0 ;
  assign n21842 = n21838 | n21841 ;
  assign n21843 = n15136 ^ n9485 ^ n6948 ;
  assign n21844 = n18824 ^ n10968 ^ n10070 ;
  assign n21845 = n3282 | n8638 ;
  assign n21846 = n6825 & ~n21845 ;
  assign n21847 = n21846 ^ n19483 ^ 1'b0 ;
  assign n21848 = n5864 ^ n1906 ^ n1320 ;
  assign n21849 = n21848 ^ n4588 ^ 1'b0 ;
  assign n21850 = n21849 ^ n945 ^ 1'b0 ;
  assign n21851 = ( n14422 & n18458 ) | ( n14422 & n18565 ) | ( n18458 & n18565 ) ;
  assign n21852 = n14600 & n19385 ;
  assign n21853 = n16632 & n21852 ;
  assign n21854 = n18089 & ~n21853 ;
  assign n21855 = n1543 & n6040 ;
  assign n21856 = ~n4882 & n21855 ;
  assign n21857 = n15733 ^ n5912 ^ n2436 ;
  assign n21858 = n21857 ^ n12457 ^ 1'b0 ;
  assign n21859 = n8201 ^ n4845 ^ 1'b0 ;
  assign n21860 = n21859 ^ n19443 ^ 1'b0 ;
  assign n21861 = ~n4210 & n21860 ;
  assign n21862 = n21861 ^ n14566 ^ n11566 ;
  assign n21863 = n10774 | n11967 ;
  assign n21864 = n21862 & n21863 ;
  assign n21865 = n9384 ^ n5583 ^ 1'b0 ;
  assign n21866 = n1134 ^ n593 ^ 1'b0 ;
  assign n21867 = n656 & n21866 ;
  assign n21868 = n10780 & ~n21867 ;
  assign n21869 = n21865 & ~n21868 ;
  assign n21870 = n16771 ^ n12963 ^ 1'b0 ;
  assign n21871 = n252 | n21870 ;
  assign n21872 = n5654 & ~n21871 ;
  assign n21873 = n7499 ^ n3154 ^ 1'b0 ;
  assign n21874 = n9563 ^ n8801 ^ 1'b0 ;
  assign n21875 = ( n8398 & ~n10527 ) | ( n8398 & n13412 ) | ( ~n10527 & n13412 ) ;
  assign n21876 = n21874 & ~n21875 ;
  assign n21877 = n4251 & n5795 ;
  assign n21878 = ( n3088 & n5562 ) | ( n3088 & ~n15999 ) | ( n5562 & ~n15999 ) ;
  assign n21880 = n707 | n10845 ;
  assign n21879 = ~n20716 & n21818 ;
  assign n21881 = n21880 ^ n21879 ^ 1'b0 ;
  assign n21882 = n17938 & n21323 ;
  assign n21883 = ~n3257 & n21882 ;
  assign n21884 = n21883 ^ n19292 ^ 1'b0 ;
  assign n21885 = ~n1360 & n4584 ;
  assign n21886 = n12421 & n21885 ;
  assign n21887 = ( n1189 & n6259 ) | ( n1189 & n21886 ) | ( n6259 & n21886 ) ;
  assign n21888 = n8941 & n15865 ;
  assign n21889 = n21888 ^ n15618 ^ n4724 ;
  assign n21890 = n21652 ^ n19941 ^ 1'b0 ;
  assign n21891 = ( n705 & n4354 ) | ( n705 & n20042 ) | ( n4354 & n20042 ) ;
  assign n21892 = n9244 & ~n21891 ;
  assign n21893 = n10863 ^ n4330 ^ 1'b0 ;
  assign n21894 = n3294 & ~n10240 ;
  assign n21895 = ~n2989 & n21894 ;
  assign n21896 = n2134 & ~n12347 ;
  assign n21897 = n19096 & ~n21896 ;
  assign n21898 = n21897 ^ n10339 ^ 1'b0 ;
  assign n21899 = ( n15468 & n21895 ) | ( n15468 & ~n21898 ) | ( n21895 & ~n21898 ) ;
  assign n21900 = n17447 ^ n16959 ^ 1'b0 ;
  assign n21901 = n8980 ^ n6345 ^ 1'b0 ;
  assign n21902 = n1591 | n21901 ;
  assign n21903 = n1251 & ~n21902 ;
  assign n21904 = n17576 ^ n6970 ^ 1'b0 ;
  assign n21905 = n3392 & n21904 ;
  assign n21906 = n5309 & n21905 ;
  assign n21907 = n21906 ^ n8443 ^ 1'b0 ;
  assign n21908 = ~n21903 & n21907 ;
  assign n21909 = ~n1367 & n3898 ;
  assign n21910 = n11844 & n21909 ;
  assign n21911 = n16716 & n21651 ;
  assign n21912 = n16328 ^ n15370 ^ 1'b0 ;
  assign n21913 = n12556 ^ n9425 ^ 1'b0 ;
  assign n21914 = n8770 & ~n21913 ;
  assign n21915 = n21914 ^ n8008 ^ n6587 ;
  assign n21916 = n14619 | n19536 ;
  assign n21917 = n19753 ^ n13134 ^ 1'b0 ;
  assign n21918 = ~n17283 & n21917 ;
  assign n21919 = n21918 ^ n18280 ^ n15907 ;
  assign n21920 = n12541 ^ n10134 ^ 1'b0 ;
  assign n21921 = n13942 & ~n21920 ;
  assign n21922 = n12147 & n21921 ;
  assign n21923 = n21922 ^ n7047 ^ 1'b0 ;
  assign n21924 = n305 & n366 ;
  assign n21925 = n21924 ^ n16835 ^ 1'b0 ;
  assign n21926 = n6059 & ~n20230 ;
  assign n21927 = n13461 ^ n6478 ^ n4706 ;
  assign n21928 = ~n2722 & n6229 ;
  assign n21929 = n21928 ^ n14915 ^ 1'b0 ;
  assign n21930 = n21927 & n21929 ;
  assign n21931 = n1930 & n21930 ;
  assign n21932 = n3914 ^ n1022 ^ 1'b0 ;
  assign n21933 = n21932 ^ n19544 ^ 1'b0 ;
  assign n21935 = ~n2028 & n3651 ;
  assign n21934 = n7854 & ~n12988 ;
  assign n21936 = n21935 ^ n21934 ^ 1'b0 ;
  assign n21937 = n15184 & n21936 ;
  assign n21938 = n21937 ^ n5492 ^ 1'b0 ;
  assign n21939 = n3457 & n13547 ;
  assign n21940 = n21939 ^ n396 ^ 1'b0 ;
  assign n21947 = ~n726 & n1904 ;
  assign n21948 = ~n4463 & n21947 ;
  assign n21949 = n21948 ^ n11272 ^ 1'b0 ;
  assign n21941 = n11609 ^ n2160 ^ 1'b0 ;
  assign n21943 = n7989 | n13052 ;
  assign n21944 = ~n21679 & n21943 ;
  assign n21942 = n5958 & n19192 ;
  assign n21945 = n21944 ^ n21942 ^ 1'b0 ;
  assign n21946 = ( ~n2221 & n21941 ) | ( ~n2221 & n21945 ) | ( n21941 & n21945 ) ;
  assign n21950 = n21949 ^ n21946 ^ 1'b0 ;
  assign n21951 = n21940 & n21950 ;
  assign n21952 = n9108 & ~n10017 ;
  assign n21953 = n7925 & n8119 ;
  assign n21954 = n21953 ^ n15797 ^ n8635 ;
  assign n21955 = ( n9707 & ~n19701 ) | ( n9707 & n21954 ) | ( ~n19701 & n21954 ) ;
  assign n21956 = ~n7902 & n8842 ;
  assign n21957 = n21956 ^ n1956 ^ 1'b0 ;
  assign n21958 = n7893 ^ n627 ^ 1'b0 ;
  assign n21959 = n2150 & n11393 ;
  assign n21960 = n1093 & n21959 ;
  assign n21961 = n994 & n4897 ;
  assign n21962 = n672 & n21961 ;
  assign n21963 = n7713 & ~n21962 ;
  assign n21966 = n4294 ^ n488 ^ 1'b0 ;
  assign n21967 = n6691 & n21966 ;
  assign n21968 = n16694 & n21967 ;
  assign n21964 = n1031 | n16984 ;
  assign n21965 = n21964 ^ n4387 ^ 1'b0 ;
  assign n21969 = n21968 ^ n21965 ^ n20805 ;
  assign n21971 = ~n10722 & n19564 ;
  assign n21972 = n21971 ^ n13486 ^ 1'b0 ;
  assign n21970 = n5572 & n6776 ;
  assign n21973 = n21972 ^ n21970 ^ 1'b0 ;
  assign n21974 = ( n6709 & n8206 ) | ( n6709 & n20031 ) | ( n8206 & n20031 ) ;
  assign n21975 = n21552 ^ n16382 ^ n10594 ;
  assign n21976 = n4867 | n21975 ;
  assign n21977 = n21976 ^ n14657 ^ 1'b0 ;
  assign n21978 = n6352 & n17578 ;
  assign n21979 = n2940 & n3899 ;
  assign n21980 = ~n772 & n21979 ;
  assign n21981 = n20206 ^ n1104 ^ 1'b0 ;
  assign n21982 = n13215 ^ n10449 ^ 1'b0 ;
  assign n21983 = ~n11097 & n21982 ;
  assign n21985 = ( ~n1929 & n5331 ) | ( ~n1929 & n19191 ) | ( n5331 & n19191 ) ;
  assign n21984 = n20281 & ~n20462 ;
  assign n21986 = n21985 ^ n21984 ^ n18927 ;
  assign n21987 = ( n2012 & n9983 ) | ( n2012 & n13107 ) | ( n9983 & n13107 ) ;
  assign n21988 = n16298 ^ n11569 ^ 1'b0 ;
  assign n21989 = n5786 ^ n5468 ^ 1'b0 ;
  assign n21991 = ~n1569 & n14964 ;
  assign n21990 = n2471 & ~n9997 ;
  assign n21992 = n21991 ^ n21990 ^ 1'b0 ;
  assign n21993 = n10177 ^ n6722 ^ 1'b0 ;
  assign n21994 = n21992 & ~n21993 ;
  assign n21997 = ~n11513 & n19606 ;
  assign n21995 = n12080 & n13211 ;
  assign n21996 = n8168 & n21995 ;
  assign n21998 = n21997 ^ n21996 ^ n9563 ;
  assign n21999 = n10741 ^ n8025 ^ 1'b0 ;
  assign n22000 = n3131 | n21999 ;
  assign n22001 = n22000 ^ n2385 ^ 1'b0 ;
  assign n22003 = n5139 | n7306 ;
  assign n22002 = ~n5749 & n9026 ;
  assign n22004 = n22003 ^ n22002 ^ 1'b0 ;
  assign n22005 = n12555 | n22004 ;
  assign n22006 = n22005 ^ n1085 ^ 1'b0 ;
  assign n22007 = ~n1003 & n22006 ;
  assign n22008 = n8731 ^ n914 ^ 1'b0 ;
  assign n22011 = n10669 ^ n919 ^ 1'b0 ;
  assign n22012 = ~n7772 & n22011 ;
  assign n22009 = n780 & n9402 ;
  assign n22010 = n22009 ^ n2044 ^ 1'b0 ;
  assign n22013 = n22012 ^ n22010 ^ 1'b0 ;
  assign n22014 = ~n15061 & n22013 ;
  assign n22016 = ( n3329 & n3941 ) | ( n3329 & ~n7357 ) | ( n3941 & ~n7357 ) ;
  assign n22015 = n12937 & n13972 ;
  assign n22017 = n22016 ^ n22015 ^ 1'b0 ;
  assign n22018 = n1322 | n3810 ;
  assign n22019 = n10556 & n22018 ;
  assign n22020 = ( n9314 & n9620 ) | ( n9314 & ~n17985 ) | ( n9620 & ~n17985 ) ;
  assign n22021 = n14361 & ~n22020 ;
  assign n22022 = ( n2482 & ~n6762 ) | ( n2482 & n7062 ) | ( ~n6762 & n7062 ) ;
  assign n22023 = n4854 & n19105 ;
  assign n22024 = n13133 ^ n9748 ^ n835 ;
  assign n22025 = n22024 ^ n5908 ^ 1'b0 ;
  assign n22026 = n9815 ^ n5924 ^ 1'b0 ;
  assign n22027 = n5838 | n8919 ;
  assign n22028 = n17183 ^ n13814 ^ 1'b0 ;
  assign n22029 = ( n8726 & n12088 ) | ( n8726 & n22028 ) | ( n12088 & n22028 ) ;
  assign n22030 = n3199 & ~n9411 ;
  assign n22031 = ~n16477 & n22030 ;
  assign n22032 = n22031 ^ n8816 ^ 1'b0 ;
  assign n22033 = ( n6136 & n21471 ) | ( n6136 & ~n22032 ) | ( n21471 & ~n22032 ) ;
  assign n22034 = n3760 & n12416 ;
  assign n22035 = ~n11365 & n13597 ;
  assign n22036 = ~n22034 & n22035 ;
  assign n22037 = n22036 ^ n1079 ^ 1'b0 ;
  assign n22038 = n20856 ^ n18728 ^ 1'b0 ;
  assign n22039 = n3807 & ~n22038 ;
  assign n22040 = n15 & n21492 ;
  assign n22041 = ( n8037 & ~n8610 ) | ( n8037 & n15987 ) | ( ~n8610 & n15987 ) ;
  assign n22042 = n270 | n22041 ;
  assign n22043 = ( n411 & n2943 ) | ( n411 & n11991 ) | ( n2943 & n11991 ) ;
  assign n22044 = n22043 ^ n2048 ^ 1'b0 ;
  assign n22045 = n21435 ^ n14809 ^ 1'b0 ;
  assign n22046 = n6875 | n22045 ;
  assign n22047 = n4275 & n22046 ;
  assign n22048 = ~n1084 & n18059 ;
  assign n22049 = n17886 ^ n6560 ^ 1'b0 ;
  assign n22050 = n8088 | n14497 ;
  assign n22051 = n22050 ^ n2048 ^ 1'b0 ;
  assign n22052 = n3508 ^ n1965 ^ 1'b0 ;
  assign n22053 = n22052 ^ n7005 ^ 1'b0 ;
  assign n22054 = n22051 & ~n22053 ;
  assign n22055 = n16006 ^ n5161 ^ 1'b0 ;
  assign n22056 = n22055 ^ n4602 ^ 1'b0 ;
  assign n22057 = n6383 & ~n22056 ;
  assign n22058 = n2588 ^ n2414 ^ 1'b0 ;
  assign n22059 = n19782 | n22058 ;
  assign n22060 = n3713 & n13947 ;
  assign n22061 = n22060 ^ n3234 ^ 1'b0 ;
  assign n22062 = ( ~n1827 & n6844 ) | ( ~n1827 & n22061 ) | ( n6844 & n22061 ) ;
  assign n22063 = ( n164 & ~n4777 ) | ( n164 & n10760 ) | ( ~n4777 & n10760 ) ;
  assign n22064 = ~n5533 & n22063 ;
  assign n22065 = n19237 ^ n17372 ^ 1'b0 ;
  assign n22066 = n12788 | n22065 ;
  assign n22067 = n774 ^ n529 ^ 1'b0 ;
  assign n22068 = n21269 & ~n22067 ;
  assign n22069 = n19719 ^ n2966 ^ 1'b0 ;
  assign n22070 = ~n12570 & n22069 ;
  assign n22071 = ( ~n6622 & n9264 ) | ( ~n6622 & n10917 ) | ( n9264 & n10917 ) ;
  assign n22072 = n19007 | n22071 ;
  assign n22073 = n11508 | n22072 ;
  assign n22074 = ( n8480 & n14665 ) | ( n8480 & n19002 ) | ( n14665 & n19002 ) ;
  assign n22075 = n1272 & ~n12586 ;
  assign n22076 = n2529 & n5033 ;
  assign n22077 = n22076 ^ n2074 ^ 1'b0 ;
  assign n22078 = n1577 & n3133 ;
  assign n22079 = n4981 & ~n22078 ;
  assign n22080 = n22077 | n22079 ;
  assign n22081 = n19770 ^ n14522 ^ n11264 ;
  assign n22082 = n8881 | n22081 ;
  assign n22083 = n22080 & ~n22082 ;
  assign n22084 = n530 & ~n1182 ;
  assign n22085 = n5490 & ~n22084 ;
  assign n22086 = ~n3550 & n22085 ;
  assign n22087 = ~n3128 & n22086 ;
  assign n22088 = n22087 ^ n17932 ^ n884 ;
  assign n22089 = n8268 & ~n22088 ;
  assign n22090 = n16212 & n22089 ;
  assign n22091 = n22090 ^ n9538 ^ 1'b0 ;
  assign n22092 = n7561 & n22091 ;
  assign n22093 = n11832 ^ n3123 ^ 1'b0 ;
  assign n22094 = n4048 & ~n22093 ;
  assign n22095 = ~n2896 & n22094 ;
  assign n22097 = n213 & ~n8397 ;
  assign n22098 = n12555 ^ n108 ^ 1'b0 ;
  assign n22099 = n22097 & n22098 ;
  assign n22096 = n13629 & n20646 ;
  assign n22100 = n22099 ^ n22096 ^ n10328 ;
  assign n22104 = n41 | n315 ;
  assign n22105 = n3469 & ~n22104 ;
  assign n22101 = n4569 & ~n12401 ;
  assign n22102 = n22101 ^ n5608 ^ 1'b0 ;
  assign n22103 = n5062 | n22102 ;
  assign n22106 = n22105 ^ n22103 ^ n12510 ;
  assign n22107 = n14778 ^ n411 ^ 1'b0 ;
  assign n22108 = n12259 ^ n4043 ^ n1427 ;
  assign n22109 = n19511 ^ n732 ^ 1'b0 ;
  assign n22110 = ~n22108 & n22109 ;
  assign n22111 = n22110 ^ n216 ^ 1'b0 ;
  assign n22112 = n22107 & ~n22111 ;
  assign n22113 = n3337 ^ n1367 ^ 1'b0 ;
  assign n22114 = n12482 | n21827 ;
  assign n22115 = n1131 ^ n719 ^ n483 ;
  assign n22116 = n22115 ^ n4851 ^ 1'b0 ;
  assign n22117 = n9201 | n22116 ;
  assign n22118 = n16302 | n22117 ;
  assign n22119 = n1021 | n1389 ;
  assign n22120 = ( n2428 & ~n19277 ) | ( n2428 & n22119 ) | ( ~n19277 & n22119 ) ;
  assign n22121 = n22120 ^ n20874 ^ 1'b0 ;
  assign n22122 = n412 & ~n21508 ;
  assign n22123 = n20471 & n22122 ;
  assign n22124 = n283 | n2722 ;
  assign n22125 = n10273 & n22124 ;
  assign n22126 = n2094 & ~n6646 ;
  assign n22127 = n22126 ^ n265 ^ 1'b0 ;
  assign n22128 = n15979 & ~n22127 ;
  assign n22129 = n5040 & n22128 ;
  assign n22130 = n3540 ^ n1403 ^ 1'b0 ;
  assign n22131 = n3217 | n7020 ;
  assign n22132 = ( n1443 & ~n22130 ) | ( n1443 & n22131 ) | ( ~n22130 & n22131 ) ;
  assign n22133 = n2190 & n3799 ;
  assign n22134 = ~n2618 & n22133 ;
  assign n22135 = n10095 & ~n22134 ;
  assign n22136 = ~n3902 & n22135 ;
  assign n22137 = n13151 & n22136 ;
  assign n22138 = n14285 ^ n1849 ^ 1'b0 ;
  assign n22139 = n19923 | n22138 ;
  assign n22140 = n17906 & n22139 ;
  assign n22141 = n11396 & n22140 ;
  assign n22142 = n4733 & ~n19192 ;
  assign n22143 = n22077 ^ n12853 ^ 1'b0 ;
  assign n22144 = n20112 ^ n105 ^ 1'b0 ;
  assign n22145 = n19642 ^ n3662 ^ 1'b0 ;
  assign n22146 = n9959 & ~n18728 ;
  assign n22147 = n20650 ^ n17107 ^ n4001 ;
  assign n22148 = n4925 ^ n351 ^ 1'b0 ;
  assign n22149 = n6091 & n22148 ;
  assign n22150 = n21010 | n22149 ;
  assign n22151 = n5262 & ~n13817 ;
  assign n22152 = n2281 & n7254 ;
  assign n22153 = ~n6382 & n22152 ;
  assign n22154 = n7268 ^ n639 ^ 1'b0 ;
  assign n22155 = ~n17801 & n22154 ;
  assign n22156 = ~n2095 & n12547 ;
  assign n22157 = ~n6352 & n22156 ;
  assign n22158 = n21498 | n22157 ;
  assign n22159 = n848 & ~n22158 ;
  assign n22160 = ~n22155 & n22159 ;
  assign n22161 = ~n1139 & n8891 ;
  assign n22162 = n13932 | n22161 ;
  assign n22163 = n15981 | n22162 ;
  assign n22164 = n1694 & ~n19846 ;
  assign n22165 = n21418 ^ n15228 ^ 1'b0 ;
  assign n22166 = n9208 & n21765 ;
  assign n22167 = n5109 & ~n22166 ;
  assign n22168 = n22167 ^ n12270 ^ 1'b0 ;
  assign n22173 = n8962 ^ n2721 ^ 1'b0 ;
  assign n22169 = n9232 ^ n1226 ^ 1'b0 ;
  assign n22170 = n13428 & ~n22169 ;
  assign n22171 = ( ~n11733 & n15944 ) | ( ~n11733 & n15977 ) | ( n15944 & n15977 ) ;
  assign n22172 = n22170 & n22171 ;
  assign n22174 = n22173 ^ n22172 ^ 1'b0 ;
  assign n22175 = n7713 & ~n16247 ;
  assign n22176 = n299 & ~n6451 ;
  assign n22177 = n4777 & ~n18592 ;
  assign n22178 = n22176 | n22177 ;
  assign n22180 = n7988 ^ n1437 ^ 1'b0 ;
  assign n22179 = n12090 | n12687 ;
  assign n22181 = n22180 ^ n22179 ^ 1'b0 ;
  assign n22182 = n13958 & ~n22181 ;
  assign n22184 = ~n17122 & n17574 ;
  assign n22185 = n22184 ^ n7218 ^ 1'b0 ;
  assign n22186 = n11626 & n22185 ;
  assign n22183 = ~n3696 & n20773 ;
  assign n22187 = n22186 ^ n22183 ^ 1'b0 ;
  assign n22188 = n5222 & ~n20574 ;
  assign n22189 = ~n6414 & n22188 ;
  assign n22190 = n306 & n4733 ;
  assign n22191 = ~n15167 & n22190 ;
  assign n22192 = n164 & n6551 ;
  assign n22193 = ~n1825 & n22192 ;
  assign n22194 = n22193 ^ n21069 ^ 1'b0 ;
  assign n22195 = n8008 & ~n22194 ;
  assign n22196 = n22195 ^ n21453 ^ 1'b0 ;
  assign n22197 = n22196 ^ n17174 ^ 1'b0 ;
  assign n22198 = ~n22191 & n22197 ;
  assign n22199 = n12619 & n18530 ;
  assign n22200 = n12491 & n22199 ;
  assign n22201 = n17986 & n18863 ;
  assign n22202 = ~n8192 & n22201 ;
  assign n22203 = ~n3365 & n4972 ;
  assign n22204 = n22203 ^ n7013 ^ 1'b0 ;
  assign n22205 = n405 | n22204 ;
  assign n22206 = ( n8827 & n11147 ) | ( n8827 & n22205 ) | ( n11147 & n22205 ) ;
  assign n22207 = n22206 ^ n13117 ^ 1'b0 ;
  assign n22208 = ~n22202 & n22207 ;
  assign n22209 = ~n22200 & n22208 ;
  assign n22210 = n14957 ^ n11154 ^ n7794 ;
  assign n22211 = n7073 & ~n12791 ;
  assign n22212 = n11104 & ~n22211 ;
  assign n22213 = n2566 & n22212 ;
  assign n22214 = n22213 ^ n13743 ^ 1'b0 ;
  assign n22215 = ~n22210 & n22214 ;
  assign n22216 = n813 & ~n20688 ;
  assign n22219 = n2497 ^ n645 ^ 1'b0 ;
  assign n22220 = n6288 & n22219 ;
  assign n22217 = n12611 & n14172 ;
  assign n22218 = n22217 ^ n10326 ^ 1'b0 ;
  assign n22221 = n22220 ^ n22218 ^ 1'b0 ;
  assign n22222 = n12060 & ~n22221 ;
  assign n22223 = n352 | n2561 ;
  assign n22224 = n8794 & n22223 ;
  assign n22225 = n3488 & ~n22224 ;
  assign n22226 = n6240 | n19974 ;
  assign n22227 = n22226 ^ n4077 ^ 1'b0 ;
  assign n22228 = n9732 & ~n22227 ;
  assign n22229 = n22228 ^ n11124 ^ 1'b0 ;
  assign n22230 = ~n1350 & n22229 ;
  assign n22231 = n9679 & ~n9683 ;
  assign n22232 = ~n22230 & n22231 ;
  assign n22233 = n6036 & ~n7326 ;
  assign n22234 = n18896 ^ n7571 ^ 1'b0 ;
  assign n22235 = ~n22233 & n22234 ;
  assign n22236 = n22235 ^ n12400 ^ 1'b0 ;
  assign n22237 = ~n2676 & n22236 ;
  assign n22238 = n13032 ^ n2729 ^ 1'b0 ;
  assign n22239 = n2306 | n22238 ;
  assign n22240 = n22239 ^ n12574 ^ 1'b0 ;
  assign n22241 = n21679 ^ n12044 ^ n9522 ;
  assign n22242 = n711 & n1698 ;
  assign n22243 = n22242 ^ n13680 ^ 1'b0 ;
  assign n22244 = n20970 ^ n7649 ^ 1'b0 ;
  assign n22250 = n19755 ^ n8337 ^ 1'b0 ;
  assign n22245 = n20444 ^ n19254 ^ 1'b0 ;
  assign n22246 = n10053 & n22245 ;
  assign n22247 = n16596 & n22246 ;
  assign n22248 = n16411 | n22247 ;
  assign n22249 = n22248 ^ n11777 ^ 1'b0 ;
  assign n22251 = n22250 ^ n22249 ^ 1'b0 ;
  assign n22252 = ~n22244 & n22251 ;
  assign n22253 = n4482 | n18715 ;
  assign n22254 = ~n13797 & n22253 ;
  assign n22255 = n5410 & n22254 ;
  assign n22256 = n7069 ^ n3615 ^ n3137 ;
  assign n22257 = ~n18008 & n22256 ;
  assign n22258 = n398 & n22257 ;
  assign n22259 = ~n13707 & n14502 ;
  assign n22260 = ( n3901 & n22258 ) | ( n3901 & n22259 ) | ( n22258 & n22259 ) ;
  assign n22261 = n13248 ^ n3580 ^ 1'b0 ;
  assign n22262 = n1668 | n12844 ;
  assign n22263 = n22261 & ~n22262 ;
  assign n22264 = n22263 ^ n20081 ^ 1'b0 ;
  assign n22265 = n55 & n22264 ;
  assign n22266 = n16129 & n17948 ;
  assign n22267 = n22266 ^ n2986 ^ 1'b0 ;
  assign n22268 = ~n6121 & n22267 ;
  assign n22269 = n22268 ^ n17151 ^ 1'b0 ;
  assign n22270 = n18601 ^ n3329 ^ 1'b0 ;
  assign n22271 = n17872 ^ n8470 ^ n1243 ;
  assign n22272 = n9701 | n18454 ;
  assign n22273 = ~n427 & n16282 ;
  assign n22274 = n22273 ^ n7312 ^ 1'b0 ;
  assign n22275 = ~n3469 & n19172 ;
  assign n22276 = n17308 ^ n4608 ^ 1'b0 ;
  assign n22277 = n6360 ^ n5848 ^ 1'b0 ;
  assign n22278 = n5856 | n22277 ;
  assign n22279 = ~n5146 & n9412 ;
  assign n22280 = n16771 & n22279 ;
  assign n22281 = n2266 & n22280 ;
  assign n22282 = n4737 & ~n22281 ;
  assign n22283 = n6242 & ~n21991 ;
  assign n22284 = n22283 ^ n19034 ^ n18621 ;
  assign n22285 = n22284 ^ n9362 ^ 1'b0 ;
  assign n22286 = n22282 | n22285 ;
  assign n22287 = ~n576 & n21385 ;
  assign n22288 = ~n1105 & n7495 ;
  assign n22289 = n22288 ^ n12311 ^ n9460 ;
  assign n22290 = n16169 | n22289 ;
  assign n22291 = n22290 ^ n10714 ^ n1193 ;
  assign n22292 = n1468 & ~n10591 ;
  assign n22293 = n22292 ^ n9743 ^ n3734 ;
  assign n22294 = n913 & ~n7106 ;
  assign n22295 = n6908 | n22294 ;
  assign n22296 = n22295 ^ n10511 ^ 1'b0 ;
  assign n22297 = ~n694 & n5284 ;
  assign n22298 = n22297 ^ n1263 ^ 1'b0 ;
  assign n22299 = n19518 & ~n22298 ;
  assign n22300 = ~n5057 & n22299 ;
  assign n22301 = n13766 & n22300 ;
  assign n22302 = n6356 & ~n22301 ;
  assign n22303 = n22302 ^ n5337 ^ 1'b0 ;
  assign n22304 = ~n4030 & n18143 ;
  assign n22306 = n7747 & ~n15744 ;
  assign n22307 = n5853 & n22306 ;
  assign n22308 = n14425 | n22307 ;
  assign n22309 = n22308 ^ n8262 ^ 1'b0 ;
  assign n22305 = n10411 | n14964 ;
  assign n22310 = n22309 ^ n22305 ^ 1'b0 ;
  assign n22311 = n328 & n764 ;
  assign n22312 = n22311 ^ n2327 ^ 1'b0 ;
  assign n22313 = n63 | n7199 ;
  assign n22314 = n22313 ^ n2176 ^ n68 ;
  assign n22315 = n1340 & n5891 ;
  assign n22316 = n22314 & n22315 ;
  assign n22317 = n22316 ^ n5864 ^ 1'b0 ;
  assign n22318 = n15830 & n22317 ;
  assign n22319 = n7763 ^ n5811 ^ n1650 ;
  assign n22320 = n21749 & n22319 ;
  assign n22321 = n7218 & n22320 ;
  assign n22322 = n22321 ^ n829 ^ 1'b0 ;
  assign n22323 = n6215 | n22322 ;
  assign n22324 = n221 | n14893 ;
  assign n22325 = n22324 ^ n11925 ^ 1'b0 ;
  assign n22326 = n18462 ^ n366 ^ 1'b0 ;
  assign n22327 = n11901 & n22326 ;
  assign n22328 = ~n2222 & n22327 ;
  assign n22329 = n22328 ^ n4394 ^ 1'b0 ;
  assign n22330 = n16263 & ~n22329 ;
  assign n22331 = n8058 & n13682 ;
  assign n22332 = n22331 ^ n811 ^ 1'b0 ;
  assign n22333 = n9830 & ~n22332 ;
  assign n22334 = n1625 | n8063 ;
  assign n22335 = ( n749 & ~n10804 ) | ( n749 & n22334 ) | ( ~n10804 & n22334 ) ;
  assign n22336 = n22335 ^ n5162 ^ n3824 ;
  assign n22337 = n1603 | n2832 ;
  assign n22338 = n1603 & ~n22337 ;
  assign n22339 = n1400 | n22338 ;
  assign n22340 = ~n953 & n9874 ;
  assign n22341 = n22339 & n22340 ;
  assign n22342 = n22336 & n22341 ;
  assign n22343 = n5078 | n5279 ;
  assign n22344 = n19180 ^ n6654 ^ 1'b0 ;
  assign n22345 = ~n1248 & n22344 ;
  assign n22346 = n13477 ^ n1058 ^ 1'b0 ;
  assign n22347 = ~n5876 & n6670 ;
  assign n22348 = n19297 & n22347 ;
  assign n22349 = x1 & n15944 ;
  assign n22350 = n4187 & n22349 ;
  assign n22351 = n10726 | n22350 ;
  assign n22352 = n411 & ~n22351 ;
  assign n22353 = n14258 ^ n5673 ^ 1'b0 ;
  assign n22354 = n11654 ^ n2804 ^ 1'b0 ;
  assign n22355 = n22353 & n22354 ;
  assign n22356 = ~n51 & n7532 ;
  assign n22357 = n22356 ^ n2958 ^ 1'b0 ;
  assign n22358 = ( ~n3776 & n4622 ) | ( ~n3776 & n22357 ) | ( n4622 & n22357 ) ;
  assign n22359 = n7010 & ~n22358 ;
  assign n22360 = n22359 ^ n19465 ^ 1'b0 ;
  assign n22362 = n4588 | n21506 ;
  assign n22361 = n12484 ^ n11292 ^ 1'b0 ;
  assign n22363 = n22362 ^ n22361 ^ n5572 ;
  assign n22364 = n17035 | n22363 ;
  assign n22365 = n22360 | n22364 ;
  assign n22366 = ~n7485 & n17046 ;
  assign n22367 = n22366 ^ n11356 ^ 1'b0 ;
  assign n22368 = n22367 ^ n498 ^ 1'b0 ;
  assign n22372 = n7876 ^ n6501 ^ n4186 ;
  assign n22369 = n4608 ^ n1043 ^ 1'b0 ;
  assign n22370 = ( n5132 & n19936 ) | ( n5132 & ~n22369 ) | ( n19936 & ~n22369 ) ;
  assign n22371 = n14817 & ~n22370 ;
  assign n22373 = n22372 ^ n22371 ^ 1'b0 ;
  assign n22374 = n22223 ^ n987 ^ 1'b0 ;
  assign n22375 = n17134 & ~n22374 ;
  assign n22376 = n22375 ^ n5537 ^ 1'b0 ;
  assign n22377 = n16378 ^ n9504 ^ 1'b0 ;
  assign n22378 = n13603 & n22377 ;
  assign n22379 = n15159 & n22378 ;
  assign n22380 = n1003 & n11345 ;
  assign n22381 = n22380 ^ n19558 ^ n16850 ;
  assign n22382 = n14204 | n22381 ;
  assign n22383 = n22382 ^ n12619 ^ 1'b0 ;
  assign n22384 = ( n2177 & n12260 ) | ( n2177 & n16132 ) | ( n12260 & n16132 ) ;
  assign n22385 = n22384 ^ n7150 ^ 1'b0 ;
  assign n22386 = n2129 & n22385 ;
  assign n22387 = n16278 ^ n5400 ^ 1'b0 ;
  assign n22388 = n6415 ^ n4177 ^ 1'b0 ;
  assign n22389 = ~n13895 & n19741 ;
  assign n22390 = n22389 ^ n1515 ^ 1'b0 ;
  assign n22391 = n10229 ^ n5150 ^ 1'b0 ;
  assign n22392 = n22391 ^ n6089 ^ 1'b0 ;
  assign n22393 = n68 | n10943 ;
  assign n22394 = n22393 ^ n2101 ^ 1'b0 ;
  assign n22395 = n3581 & ~n11144 ;
  assign n22396 = n18077 ^ n13426 ^ n4534 ;
  assign n22397 = n835 & ~n14737 ;
  assign n22398 = ~n14208 & n22397 ;
  assign n22399 = n22398 ^ n20426 ^ n7345 ;
  assign n22400 = n21815 ^ n20096 ^ 1'b0 ;
  assign n22401 = n14279 ^ n291 ^ 1'b0 ;
  assign n22402 = n1412 | n22401 ;
  assign n22403 = n22402 ^ n4970 ^ 1'b0 ;
  assign n22404 = n22403 ^ n13238 ^ n4819 ;
  assign n22405 = n22404 ^ n18055 ^ 1'b0 ;
  assign n22406 = ~n972 & n7120 ;
  assign n22407 = n22406 ^ n20737 ^ 1'b0 ;
  assign n22408 = ( n8709 & n15310 ) | ( n8709 & n19147 ) | ( n15310 & n19147 ) ;
  assign n22413 = n1330 | n5111 ;
  assign n22414 = n22413 ^ n1245 ^ 1'b0 ;
  assign n22415 = n8028 & n22414 ;
  assign n22416 = ~n13537 & n22415 ;
  assign n22409 = n11769 ^ n1400 ^ 1'b0 ;
  assign n22410 = n269 | n22409 ;
  assign n22411 = n22410 ^ n4128 ^ 1'b0 ;
  assign n22412 = n18816 & n22411 ;
  assign n22417 = n22416 ^ n22412 ^ 1'b0 ;
  assign n22418 = n8926 | n16998 ;
  assign n22419 = n22418 ^ n17380 ^ 1'b0 ;
  assign n22423 = n4093 & ~n11459 ;
  assign n22424 = n22423 ^ n717 ^ 1'b0 ;
  assign n22425 = n4014 & n16175 ;
  assign n22426 = n22424 & n22425 ;
  assign n22420 = n2355 & ~n2877 ;
  assign n22421 = ~n17801 & n22420 ;
  assign n22422 = n10083 & n22421 ;
  assign n22427 = n22426 ^ n22422 ^ 1'b0 ;
  assign n22428 = n22419 | n22427 ;
  assign n22429 = n22099 ^ n6292 ^ 1'b0 ;
  assign n22434 = n15009 ^ n2825 ^ 1'b0 ;
  assign n22435 = n3302 & n22434 ;
  assign n22432 = n2288 | n6973 ;
  assign n22433 = n7119 | n22432 ;
  assign n22430 = n19203 ^ n8696 ^ 1'b0 ;
  assign n22431 = n8882 | n22430 ;
  assign n22436 = n22435 ^ n22433 ^ n22431 ;
  assign n22437 = ( n1697 & ~n2126 ) | ( n1697 & n7791 ) | ( ~n2126 & n7791 ) ;
  assign n22438 = n22437 ^ n530 ^ 1'b0 ;
  assign n22439 = n10528 & n17012 ;
  assign n22440 = n22439 ^ n18410 ^ n15855 ;
  assign n22441 = n7649 ^ n3038 ^ 1'b0 ;
  assign n22442 = n22441 ^ n9514 ^ 1'b0 ;
  assign n22443 = n12979 & n22442 ;
  assign n22444 = n22443 ^ n3314 ^ 1'b0 ;
  assign n22445 = n892 & n15364 ;
  assign n22446 = n11626 | n12431 ;
  assign n22447 = ~n6569 & n16475 ;
  assign n22448 = n22447 ^ n16077 ^ n3774 ;
  assign n22450 = n14219 ^ n2413 ^ 1'b0 ;
  assign n22449 = n5036 & ~n12439 ;
  assign n22451 = n22450 ^ n22449 ^ 1'b0 ;
  assign n22452 = n1039 & ~n2356 ;
  assign n22453 = n7364 | n13356 ;
  assign n22454 = n22453 ^ n10883 ^ n7335 ;
  assign n22455 = n3702 | n8629 ;
  assign n22456 = n22455 ^ n8537 ^ 1'b0 ;
  assign n22457 = n22456 ^ n8172 ^ 1'b0 ;
  assign n22458 = n22457 ^ n11698 ^ 1'b0 ;
  assign n22459 = ( n3761 & n7739 ) | ( n3761 & ~n22458 ) | ( n7739 & ~n22458 ) ;
  assign n22460 = n22454 & ~n22459 ;
  assign n22461 = ~n13426 & n22460 ;
  assign n22462 = n18432 & n22461 ;
  assign n22463 = ~n5834 & n10452 ;
  assign n22464 = n18867 & n22463 ;
  assign n22465 = ( ~n6091 & n7895 ) | ( ~n6091 & n22464 ) | ( n7895 & n22464 ) ;
  assign n22466 = n22391 ^ n10739 ^ n2195 ;
  assign n22467 = n22466 ^ n4091 ^ 1'b0 ;
  assign n22468 = n9244 & n22467 ;
  assign n22469 = n17887 ^ n4693 ^ n1864 ;
  assign n22470 = ( n4447 & n12597 ) | ( n4447 & ~n22469 ) | ( n12597 & ~n22469 ) ;
  assign n22471 = n1600 & n22470 ;
  assign n22472 = ~n22468 & n22471 ;
  assign n22473 = n8498 & ~n12044 ;
  assign n22474 = n6490 ^ n102 ^ 1'b0 ;
  assign n22475 = n22473 & ~n22474 ;
  assign n22477 = n11318 ^ n9271 ^ 1'b0 ;
  assign n22476 = n6245 & ~n14987 ;
  assign n22478 = n22477 ^ n22476 ^ 1'b0 ;
  assign n22479 = n22478 ^ n13845 ^ 1'b0 ;
  assign n22480 = ~n6181 & n22479 ;
  assign n22481 = ~n8972 & n13198 ;
  assign n22482 = n19904 ^ n355 ^ 1'b0 ;
  assign n22483 = n704 & n3505 ;
  assign n22484 = n2004 & ~n5607 ;
  assign n22485 = n22483 & n22484 ;
  assign n22486 = n1838 | n9075 ;
  assign n22487 = n22486 ^ n15824 ^ 1'b0 ;
  assign n22488 = n15299 ^ n346 ^ 1'b0 ;
  assign n22489 = n7687 | n22488 ;
  assign n22490 = n3508 | n22489 ;
  assign n22491 = n7473 ^ n3330 ^ 1'b0 ;
  assign n22492 = ~n8712 & n22491 ;
  assign n22493 = n9213 ^ n3031 ^ x7 ;
  assign n22494 = ~n2365 & n22493 ;
  assign n22495 = n22494 ^ n1204 ^ 1'b0 ;
  assign n22496 = ( n2339 & ~n14499 ) | ( n2339 & n22495 ) | ( ~n14499 & n22495 ) ;
  assign n22497 = ~n9374 & n22496 ;
  assign n22498 = n22497 ^ n15744 ^ 1'b0 ;
  assign n22499 = n22492 & n22498 ;
  assign n22500 = n16913 ^ n3713 ^ 1'b0 ;
  assign n22501 = ~n2321 & n22500 ;
  assign n22502 = ( ~n3236 & n4993 ) | ( ~n3236 & n9145 ) | ( n4993 & n9145 ) ;
  assign n22508 = ( n3625 & ~n6844 ) | ( n3625 & n7358 ) | ( ~n6844 & n7358 ) ;
  assign n22507 = n10093 & n12328 ;
  assign n22503 = n968 | n1100 ;
  assign n22504 = ~n11938 & n22503 ;
  assign n22505 = n17834 ^ n4404 ^ 1'b0 ;
  assign n22506 = n22504 & ~n22505 ;
  assign n22509 = n22508 ^ n22507 ^ n22506 ;
  assign n22510 = n11006 & n22509 ;
  assign n22511 = ~n20761 & n22510 ;
  assign n22512 = n19959 ^ n3840 ^ 1'b0 ;
  assign n22513 = n6678 & ~n11288 ;
  assign n22514 = n22513 ^ n15690 ^ 1'b0 ;
  assign n22515 = n6360 ^ n6118 ^ n505 ;
  assign n22516 = ~n1040 & n22515 ;
  assign n22517 = n8076 & n22516 ;
  assign n22518 = n22517 ^ n18294 ^ 1'b0 ;
  assign n22519 = n13245 ^ n8353 ^ 1'b0 ;
  assign n22520 = n4622 & ~n22519 ;
  assign n22521 = ( n5188 & ~n13881 ) | ( n5188 & n22520 ) | ( ~n13881 & n22520 ) ;
  assign n22522 = n16381 | n22521 ;
  assign n22523 = n22518 | n22522 ;
  assign n22524 = n14949 ^ n10594 ^ 1'b0 ;
  assign n22525 = n4751 | n5696 ;
  assign n22526 = ( ~n17891 & n19098 ) | ( ~n17891 & n22525 ) | ( n19098 & n22525 ) ;
  assign n22527 = ~n4694 & n8665 ;
  assign n22528 = n3011 & ~n7219 ;
  assign n22529 = n14082 ^ n8544 ^ 1'b0 ;
  assign n22530 = n8684 | n8750 ;
  assign n22531 = n15411 ^ n6660 ^ 1'b0 ;
  assign n22532 = n134 & ~n22531 ;
  assign n22533 = n22532 ^ n10873 ^ 1'b0 ;
  assign n22534 = n22530 & n22533 ;
  assign n22535 = n22534 ^ n20405 ^ 1'b0 ;
  assign n22536 = ~n22529 & n22535 ;
  assign n22537 = ~n22528 & n22536 ;
  assign n22538 = n408 & n22537 ;
  assign n22539 = n2433 ^ n1726 ^ 1'b0 ;
  assign n22540 = n13969 | n22539 ;
  assign n22541 = ( ~n4054 & n8826 ) | ( ~n4054 & n10939 ) | ( n8826 & n10939 ) ;
  assign n22542 = n21376 ^ n8711 ^ 1'b0 ;
  assign n22543 = ~n18294 & n22542 ;
  assign n22544 = n22541 & n22543 ;
  assign n22545 = ( n1387 & ~n12491 ) | ( n1387 & n21499 ) | ( ~n12491 & n21499 ) ;
  assign n22546 = n22544 | n22545 ;
  assign n22548 = n2674 & n4485 ;
  assign n22549 = ~n543 & n22548 ;
  assign n22550 = n22549 ^ n7915 ^ n6951 ;
  assign n22547 = n10890 & ~n14294 ;
  assign n22551 = n22550 ^ n22547 ^ 1'b0 ;
  assign n22552 = n12711 ^ n8655 ^ n4180 ;
  assign n22553 = n22552 ^ n9937 ^ n2139 ;
  assign n22554 = ~n17589 & n17932 ;
  assign n22556 = ~n350 & n10357 ;
  assign n22555 = n6664 & ~n10344 ;
  assign n22557 = n22556 ^ n22555 ^ 1'b0 ;
  assign n22558 = n7080 ^ n3561 ^ 1'b0 ;
  assign n22559 = n9144 ^ n4943 ^ 1'b0 ;
  assign n22560 = ~n9969 & n22559 ;
  assign n22561 = n22558 & n22560 ;
  assign n22562 = ( ~n2294 & n8625 ) | ( ~n2294 & n9414 ) | ( n8625 & n9414 ) ;
  assign n22563 = n5085 | n9936 ;
  assign n22564 = n5047 | n22563 ;
  assign n22565 = ~n7979 & n22564 ;
  assign n22566 = n15785 & n22565 ;
  assign n22567 = n22566 ^ n12163 ^ 1'b0 ;
  assign n22568 = n22562 & ~n22567 ;
  assign n22569 = n1745 & ~n6958 ;
  assign n22570 = n11178 & ~n22569 ;
  assign n22571 = ~n15229 & n22570 ;
  assign n22572 = n14421 ^ n3483 ^ 1'b0 ;
  assign n22573 = ~n10448 & n22572 ;
  assign n22574 = n9119 & ~n20245 ;
  assign n22575 = n22574 ^ n6805 ^ 1'b0 ;
  assign n22576 = n6299 & n22575 ;
  assign n22577 = n22573 & n22576 ;
  assign n22578 = n20498 ^ n8838 ^ 1'b0 ;
  assign n22579 = n3357 & ~n4004 ;
  assign n22580 = n22579 ^ n12235 ^ 1'b0 ;
  assign n22581 = n13030 | n19483 ;
  assign n22582 = n1162 & ~n22581 ;
  assign n22583 = n22582 ^ n4487 ^ 1'b0 ;
  assign n22584 = n6650 & ~n14920 ;
  assign n22585 = n12396 & n22584 ;
  assign n22586 = n9188 & ~n20114 ;
  assign n22587 = n14489 ^ n4055 ^ 1'b0 ;
  assign n22588 = ~n8697 & n22587 ;
  assign n22589 = n17460 ^ n12840 ^ n11009 ;
  assign n22590 = n9428 & ~n11448 ;
  assign n22591 = ~n4338 & n6396 ;
  assign n22592 = n22591 ^ n20985 ^ 1'b0 ;
  assign n22593 = ~n12408 & n19305 ;
  assign n22594 = n621 | n22593 ;
  assign n22595 = n1223 | n3059 ;
  assign n22596 = n1314 & ~n22595 ;
  assign n22597 = n655 | n2601 ;
  assign n22598 = n22596 | n22597 ;
  assign n22599 = n1951 ^ n1198 ^ 1'b0 ;
  assign n22600 = n14873 | n22599 ;
  assign n22601 = n22600 ^ n6957 ^ 1'b0 ;
  assign n22602 = ~n7549 & n22601 ;
  assign n22603 = n13754 ^ n10289 ^ 1'b0 ;
  assign n22604 = n13013 ^ n6275 ^ 1'b0 ;
  assign n22605 = ~n2207 & n20556 ;
  assign n22606 = n22604 & ~n22605 ;
  assign n22607 = n22603 & n22606 ;
  assign n22608 = n1492 & n8408 ;
  assign n22609 = n22608 ^ n22577 ^ 1'b0 ;
  assign n22610 = n22607 & ~n22609 ;
  assign n22611 = ~n11967 & n21050 ;
  assign n22612 = n6430 ^ n3202 ^ 1'b0 ;
  assign n22613 = n14531 ^ n11740 ^ 1'b0 ;
  assign n22614 = n22613 ^ n17763 ^ 1'b0 ;
  assign n22615 = n1875 | n22614 ;
  assign n22616 = n4628 & n13334 ;
  assign n22617 = ~n3916 & n22616 ;
  assign n22619 = n11503 ^ n10263 ^ n809 ;
  assign n22618 = ~n839 & n11329 ;
  assign n22620 = n22619 ^ n22618 ^ 1'b0 ;
  assign n22622 = n10562 ^ n1668 ^ 1'b0 ;
  assign n22621 = n7240 | n19236 ;
  assign n22623 = n22622 ^ n22621 ^ 1'b0 ;
  assign n22624 = n22564 ^ n12430 ^ n4216 ;
  assign n22625 = n22624 ^ n3092 ^ 1'b0 ;
  assign n22626 = n14041 & n22625 ;
  assign n22627 = ( n4331 & n6754 ) | ( n4331 & n22626 ) | ( n6754 & n22626 ) ;
  assign n22628 = n8030 & ~n21494 ;
  assign n22632 = ( n803 & ~n8917 ) | ( n803 & n15061 ) | ( ~n8917 & n15061 ) ;
  assign n22629 = n356 & ~n5580 ;
  assign n22630 = ~n9989 & n22629 ;
  assign n22631 = n22630 ^ n10481 ^ 1'b0 ;
  assign n22633 = n22632 ^ n22631 ^ 1'b0 ;
  assign n22634 = n8661 ^ n6440 ^ 1'b0 ;
  assign n22635 = n17811 & ~n19518 ;
  assign n22636 = n22635 ^ n10827 ^ 1'b0 ;
  assign n22637 = n15355 ^ n8143 ^ 1'b0 ;
  assign n22638 = ~n22224 & n22637 ;
  assign n22639 = ~n1412 & n10650 ;
  assign n22640 = ( n10199 & n12180 ) | ( n10199 & n22639 ) | ( n12180 & n22639 ) ;
  assign n22641 = ~n14249 & n21116 ;
  assign n22642 = n962 | n12421 ;
  assign n22643 = n17766 ^ n2499 ^ 1'b0 ;
  assign n22644 = n17714 & n22643 ;
  assign n22646 = n8738 | n22058 ;
  assign n22647 = n22646 ^ n2932 ^ 1'b0 ;
  assign n22648 = n15046 & n22647 ;
  assign n22645 = n17247 ^ n2440 ^ 1'b0 ;
  assign n22649 = n22648 ^ n22645 ^ 1'b0 ;
  assign n22650 = n19687 ^ n14066 ^ 1'b0 ;
  assign n22651 = n21651 | n22650 ;
  assign n22652 = ( n12402 & ~n15643 ) | ( n12402 & n22651 ) | ( ~n15643 & n22651 ) ;
  assign n22653 = n7900 ^ n5924 ^ 1'b0 ;
  assign n22654 = ( ~n1906 & n11908 ) | ( ~n1906 & n22653 ) | ( n11908 & n22653 ) ;
  assign n22655 = n10900 & ~n16580 ;
  assign n22656 = n22655 ^ n9835 ^ 1'b0 ;
  assign n22658 = n22435 ^ n14409 ^ 1'b0 ;
  assign n22659 = ( n9828 & ~n17809 ) | ( n9828 & n22658 ) | ( ~n17809 & n22658 ) ;
  assign n22657 = n19596 ^ n1803 ^ 1'b0 ;
  assign n22660 = n22659 ^ n22657 ^ 1'b0 ;
  assign n22661 = n4301 & n8172 ;
  assign n22662 = n12880 ^ n1399 ^ 1'b0 ;
  assign n22663 = n2945 & ~n3039 ;
  assign n22664 = ~n7763 & n22663 ;
  assign n22665 = n22664 ^ n16513 ^ 1'b0 ;
  assign n22666 = ~n22662 & n22665 ;
  assign n22667 = ~n2621 & n7099 ;
  assign n22668 = ~n4665 & n22667 ;
  assign n22669 = ( n957 & n6007 ) | ( n957 & n10986 ) | ( n6007 & n10986 ) ;
  assign n22670 = n12335 ^ n2135 ^ 1'b0 ;
  assign n22671 = ~n4961 & n22670 ;
  assign n22672 = n22671 ^ n4750 ^ 1'b0 ;
  assign n22673 = ~n10897 & n22672 ;
  assign n22674 = n15684 & n22673 ;
  assign n22675 = n3546 | n22674 ;
  assign n22676 = n2288 & ~n22675 ;
  assign n22677 = n1596 & n13879 ;
  assign n22678 = n13686 ^ n10960 ^ 1'b0 ;
  assign n22679 = n16398 & n22678 ;
  assign n22680 = n22677 | n22679 ;
  assign n22681 = n20856 & ~n22680 ;
  assign n22682 = n5880 & n8601 ;
  assign n22683 = n22682 ^ n6804 ^ n3767 ;
  assign n22684 = n8471 ^ n451 ^ 1'b0 ;
  assign n22685 = n18600 | n22684 ;
  assign n22686 = ~n201 & n22685 ;
  assign n22687 = n22686 ^ n3187 ^ 1'b0 ;
  assign n22688 = ~n6972 & n7045 ;
  assign n22689 = n2839 & ~n9716 ;
  assign n22690 = ~n19186 & n22689 ;
  assign n22691 = n22690 ^ n5661 ^ 1'b0 ;
  assign n22692 = n5507 & ~n22691 ;
  assign n22693 = ~x3 & n12771 ;
  assign n22694 = ~n7957 & n22693 ;
  assign n22696 = n3579 | n8509 ;
  assign n22697 = n22696 ^ n368 ^ 1'b0 ;
  assign n22698 = n22697 ^ n9245 ^ 1'b0 ;
  assign n22695 = n7506 ^ n5352 ^ 1'b0 ;
  assign n22699 = n22698 ^ n22695 ^ 1'b0 ;
  assign n22700 = n5817 & ~n14083 ;
  assign n22701 = n6471 ^ n4866 ^ 1'b0 ;
  assign n22702 = n22700 & n22701 ;
  assign n22703 = n2597 & n17576 ;
  assign n22704 = n4818 | n17000 ;
  assign n22705 = n14674 ^ n4543 ^ 1'b0 ;
  assign n22706 = n2983 ^ n533 ^ 1'b0 ;
  assign n22707 = n6924 & ~n22706 ;
  assign n22708 = n22707 ^ n1023 ^ 1'b0 ;
  assign n22709 = n9179 & ~n22708 ;
  assign n22710 = n22705 & n22709 ;
  assign n22711 = n5195 & n22710 ;
  assign n22712 = n2304 ^ n1155 ^ 1'b0 ;
  assign n22713 = n2874 | n6814 ;
  assign n22714 = n22712 | n22713 ;
  assign n22715 = n1026 | n1516 ;
  assign n22716 = n5440 | n22715 ;
  assign n22717 = n7272 & n22716 ;
  assign n22719 = n21017 ^ n15426 ^ 1'b0 ;
  assign n22720 = ~n17843 & n22719 ;
  assign n22718 = n3120 & n22186 ;
  assign n22721 = n22720 ^ n22718 ^ 1'b0 ;
  assign n22722 = ( ~n102 & n3785 ) | ( ~n102 & n3884 ) | ( n3785 & n3884 ) ;
  assign n22723 = ( ~n8220 & n13927 ) | ( ~n8220 & n22722 ) | ( n13927 & n22722 ) ;
  assign n22724 = n22723 ^ n16027 ^ n5706 ;
  assign n22725 = n16605 ^ n3560 ^ 1'b0 ;
  assign n22726 = n9246 | n22725 ;
  assign n22727 = n9073 ^ n1142 ^ 1'b0 ;
  assign n22728 = ( ~n16406 & n22726 ) | ( ~n16406 & n22727 ) | ( n22726 & n22727 ) ;
  assign n22729 = n18784 ^ n8272 ^ 1'b0 ;
  assign n22730 = n6202 & n22728 ;
  assign n22731 = n22729 & n22730 ;
  assign n22735 = n122 & ~n7631 ;
  assign n22732 = n12030 ^ n2496 ^ 1'b0 ;
  assign n22733 = ~n2725 & n22732 ;
  assign n22734 = n22733 ^ n13146 ^ n6574 ;
  assign n22736 = n22735 ^ n22734 ^ 1'b0 ;
  assign n22737 = n22736 ^ n20426 ^ 1'b0 ;
  assign n22738 = n10353 & n22737 ;
  assign n22739 = ( n940 & n17319 ) | ( n940 & ~n22123 ) | ( n17319 & ~n22123 ) ;
  assign n22740 = ~n4249 & n9614 ;
  assign n22741 = n36 & ~n22740 ;
  assign n22742 = n7771 & n17280 ;
  assign n22743 = n6752 & n22742 ;
  assign n22744 = n1052 & ~n5938 ;
  assign n22745 = n213 & ~n22744 ;
  assign n22749 = n19807 ^ n686 ^ 1'b0 ;
  assign n22750 = n22749 ^ n491 ^ 1'b0 ;
  assign n22746 = n1387 & ~n12512 ;
  assign n22747 = n22746 ^ n1773 ^ 1'b0 ;
  assign n22748 = n11033 & n22747 ;
  assign n22751 = n22750 ^ n22748 ^ 1'b0 ;
  assign n22752 = n22745 | n22751 ;
  assign n22753 = n22752 ^ n7283 ^ 1'b0 ;
  assign n22758 = n16641 ^ n8061 ^ 1'b0 ;
  assign n22754 = n8957 & n13457 ;
  assign n22755 = ~n8957 & n22754 ;
  assign n22756 = n22755 ^ n15794 ^ 1'b0 ;
  assign n22757 = ( n2101 & n10865 ) | ( n2101 & n22756 ) | ( n10865 & n22756 ) ;
  assign n22759 = n22758 ^ n22757 ^ n1959 ;
  assign n22760 = ~n3832 & n7147 ;
  assign n22761 = n22760 ^ n8296 ^ 1'b0 ;
  assign n22762 = n17932 ^ n14701 ^ 1'b0 ;
  assign n22763 = n22761 | n22762 ;
  assign n22764 = n9326 | n20419 ;
  assign n22765 = n22764 ^ n17842 ^ 1'b0 ;
  assign n22766 = ~n3406 & n10267 ;
  assign n22767 = n5761 ^ n787 ^ 1'b0 ;
  assign n22768 = n4763 & n22767 ;
  assign n22769 = n22768 ^ n17809 ^ 1'b0 ;
  assign n22770 = n2004 & n22769 ;
  assign n22771 = ~n9633 & n21054 ;
  assign n22772 = n22771 ^ n6915 ^ n2323 ;
  assign n22773 = n5457 & ~n22628 ;
  assign n22774 = n19660 ^ n17661 ^ n15864 ;
  assign n22775 = n6537 & ~n7020 ;
  assign n22776 = n22775 ^ n2412 ^ 1'b0 ;
  assign n22777 = ( ~n1950 & n5455 ) | ( ~n1950 & n22776 ) | ( n5455 & n22776 ) ;
  assign n22778 = n8471 & ~n11575 ;
  assign n22779 = n22777 & ~n22778 ;
  assign n22780 = n22779 ^ n5729 ^ 1'b0 ;
  assign n22781 = n4273 ^ n3544 ^ 1'b0 ;
  assign n22782 = n16419 ^ n16098 ^ 1'b0 ;
  assign n22783 = ~n1010 & n22782 ;
  assign n22784 = n17916 ^ n2565 ^ 1'b0 ;
  assign n22785 = n22783 & n22784 ;
  assign n22786 = n3785 | n11218 ;
  assign n22787 = n22786 ^ n8919 ^ 1'b0 ;
  assign n22788 = n9583 & ~n22787 ;
  assign n22789 = n16576 ^ n5963 ^ 1'b0 ;
  assign n22790 = n22788 & n22789 ;
  assign n22791 = n4559 ^ n122 ^ 1'b0 ;
  assign n22792 = n21183 ^ n7970 ^ 1'b0 ;
  assign n22793 = ~n804 & n18950 ;
  assign n22794 = n22793 ^ n4543 ^ 1'b0 ;
  assign n22795 = n7974 ^ n2008 ^ 1'b0 ;
  assign n22796 = n1387 & ~n22795 ;
  assign n22797 = ~n10304 & n22796 ;
  assign n22798 = n22797 ^ n7834 ^ 1'b0 ;
  assign n22799 = n982 & n12986 ;
  assign n22800 = ~n6609 & n22799 ;
  assign n22801 = n22800 ^ n7128 ^ n3020 ;
  assign n22802 = n19244 ^ n76 ^ 1'b0 ;
  assign n22807 = n8446 | n20419 ;
  assign n22808 = n1142 & ~n22807 ;
  assign n22803 = n7650 & ~n22695 ;
  assign n22804 = n13716 & n22803 ;
  assign n22805 = n22804 ^ n20186 ^ 1'b0 ;
  assign n22806 = ( n12006 & ~n16786 ) | ( n12006 & n22805 ) | ( ~n16786 & n22805 ) ;
  assign n22809 = n22808 ^ n22806 ^ 1'b0 ;
  assign n22810 = ( n3971 & ~n12855 ) | ( n3971 & n19677 ) | ( ~n12855 & n19677 ) ;
  assign n22817 = n4334 | n13388 ;
  assign n22811 = n12382 ^ n3508 ^ 1'b0 ;
  assign n22812 = n11041 & ~n22811 ;
  assign n22813 = n5099 ^ n4150 ^ 1'b0 ;
  assign n22814 = ~n22812 & n22813 ;
  assign n22815 = n14503 ^ n7028 ^ 1'b0 ;
  assign n22816 = ~n22814 & n22815 ;
  assign n22818 = n22817 ^ n22816 ^ 1'b0 ;
  assign n22819 = n14452 | n22818 ;
  assign n22820 = n22142 ^ n19169 ^ 1'b0 ;
  assign n22821 = ~n7102 & n22820 ;
  assign n22822 = n4160 | n16443 ;
  assign n22823 = n22196 & ~n22822 ;
  assign n22824 = n21001 ^ n11975 ^ 1'b0 ;
  assign n22825 = ~n22823 & n22824 ;
  assign n22826 = n17291 ^ n153 ^ 1'b0 ;
  assign n22827 = n9034 | n18825 ;
  assign n22828 = n22827 ^ n14997 ^ 1'b0 ;
  assign n22839 = n2421 & ~n17398 ;
  assign n22835 = n11790 ^ n10929 ^ 1'b0 ;
  assign n22836 = n488 ^ n412 ^ 1'b0 ;
  assign n22837 = n22836 ^ n17851 ^ 1'b0 ;
  assign n22838 = n22835 | n22837 ;
  assign n22840 = n22839 ^ n22838 ^ 1'b0 ;
  assign n22830 = n13983 ^ n4436 ^ 1'b0 ;
  assign n22831 = ~n4240 & n22830 ;
  assign n22832 = n8051 | n8177 ;
  assign n22833 = n22831 | n22832 ;
  assign n22829 = n11440 ^ n3620 ^ 1'b0 ;
  assign n22834 = n22833 ^ n22829 ^ n3241 ;
  assign n22841 = n22840 ^ n22834 ^ n3234 ;
  assign n22842 = n22135 ^ n19109 ^ 1'b0 ;
  assign n22843 = n15915 | n22842 ;
  assign n22844 = n1296 & n7275 ;
  assign n22845 = n16728 ^ n1811 ^ 1'b0 ;
  assign n22846 = ~n4030 & n22845 ;
  assign n22847 = ( ~n2631 & n2885 ) | ( ~n2631 & n22846 ) | ( n2885 & n22846 ) ;
  assign n22848 = n22847 ^ n19181 ^ n6098 ;
  assign n22849 = n6741 ^ n2078 ^ 1'b0 ;
  assign n22850 = n9296 & n22849 ;
  assign n22851 = n1198 & n22850 ;
  assign n22852 = n3946 & ~n11227 ;
  assign n22853 = n3518 & ~n22852 ;
  assign n22854 = n6549 & n22853 ;
  assign n22855 = n22851 & ~n22854 ;
  assign n22856 = n14210 ^ n2592 ^ 1'b0 ;
  assign n22857 = n4626 & ~n14452 ;
  assign n22858 = n22857 ^ n9317 ^ 1'b0 ;
  assign n22861 = n7244 ^ n6215 ^ 1'b0 ;
  assign n22862 = ~n2449 & n22861 ;
  assign n22863 = ~n2181 & n22862 ;
  assign n22864 = ~n5589 & n22863 ;
  assign n22859 = n2977 | n7208 ;
  assign n22860 = ~n10907 & n22859 ;
  assign n22865 = n22864 ^ n22860 ^ 1'b0 ;
  assign n22866 = ~n201 & n8234 ;
  assign n22867 = n12712 & n22866 ;
  assign n22868 = n13425 ^ n4756 ^ 1'b0 ;
  assign n22869 = n10900 & n22868 ;
  assign n22870 = n1024 & n3881 ;
  assign n22871 = n22869 | n22870 ;
  assign n22872 = n6193 & n16915 ;
  assign n22873 = ~n11920 & n22872 ;
  assign n22874 = n11443 & ~n12315 ;
  assign n22875 = ~n11955 & n22874 ;
  assign n22876 = n22875 ^ n18392 ^ 1'b0 ;
  assign n22883 = ( n7551 & n19220 ) | ( n7551 & n21813 ) | ( n19220 & n21813 ) ;
  assign n22877 = n18179 ^ n8456 ^ 1'b0 ;
  assign n22878 = n6265 & ~n22877 ;
  assign n22879 = n22878 ^ n19708 ^ 1'b0 ;
  assign n22880 = n436 & ~n22879 ;
  assign n22881 = n22880 ^ n18562 ^ 1'b0 ;
  assign n22882 = n8712 | n22881 ;
  assign n22884 = n22883 ^ n22882 ^ 1'b0 ;
  assign n22886 = n13253 ^ n10826 ^ 1'b0 ;
  assign n22885 = n14543 | n14658 ;
  assign n22887 = n22886 ^ n22885 ^ 1'b0 ;
  assign n22888 = ~n14124 & n15117 ;
  assign n22889 = ( ~n1308 & n5635 ) | ( ~n1308 & n22888 ) | ( n5635 & n22888 ) ;
  assign n22890 = n22889 ^ n21656 ^ 1'b0 ;
  assign n22891 = ( n5500 & n10540 ) | ( n5500 & n22180 ) | ( n10540 & n22180 ) ;
  assign n22892 = ( n2314 & n3569 ) | ( n2314 & n22891 ) | ( n3569 & n22891 ) ;
  assign n22893 = n10192 & ~n22892 ;
  assign n22894 = n8654 & ~n22893 ;
  assign n22895 = n3807 | n6389 ;
  assign n22896 = n14964 | n18486 ;
  assign n22897 = n22895 & ~n22896 ;
  assign n22898 = n800 & n5040 ;
  assign n22899 = n251 & n22898 ;
  assign n22900 = ( n1154 & n9524 ) | ( n1154 & n18465 ) | ( n9524 & n18465 ) ;
  assign n22901 = n20984 ^ n8584 ^ 1'b0 ;
  assign n22902 = n18553 & n22901 ;
  assign n22903 = n19562 ^ n4815 ^ n4703 ;
  assign n22904 = n5589 & ~n22903 ;
  assign n22905 = ~n5589 & n22904 ;
  assign n22906 = ~n4648 & n7289 ;
  assign n22907 = n15146 ^ n13011 ^ 1'b0 ;
  assign n22908 = n2886 | n22907 ;
  assign n22909 = n11052 & n13345 ;
  assign n22910 = n8319 & n14571 ;
  assign n22911 = n22910 ^ n13879 ^ 1'b0 ;
  assign n22913 = n7784 & n9792 ;
  assign n22912 = n14138 ^ n1320 ^ n709 ;
  assign n22914 = n22913 ^ n22912 ^ 1'b0 ;
  assign n22915 = ~n22911 & n22914 ;
  assign n22917 = n1883 ^ n493 ^ 1'b0 ;
  assign n22918 = ( n5809 & ~n14246 ) | ( n5809 & n22917 ) | ( ~n14246 & n22917 ) ;
  assign n22916 = n10368 ^ n8148 ^ 1'b0 ;
  assign n22919 = n22918 ^ n22916 ^ 1'b0 ;
  assign n22920 = ~n6240 & n22919 ;
  assign n22921 = n4998 ^ x3 ^ 1'b0 ;
  assign n22922 = n541 & n22921 ;
  assign n22923 = n14811 & n22922 ;
  assign n22924 = n2579 & ~n13067 ;
  assign n22925 = n10544 & ~n14507 ;
  assign n22926 = n22925 ^ n19173 ^ 1'b0 ;
  assign n22929 = n14852 | n19216 ;
  assign n22930 = ( n871 & ~n21332 ) | ( n871 & n22929 ) | ( ~n21332 & n22929 ) ;
  assign n22927 = ( n4113 & n4845 ) | ( n4113 & ~n11884 ) | ( n4845 & ~n11884 ) ;
  assign n22928 = n4422 & n22927 ;
  assign n22931 = n22930 ^ n22928 ^ 1'b0 ;
  assign n22932 = n10762 ^ n9603 ^ 1'b0 ;
  assign n22933 = n8603 | n22932 ;
  assign n22934 = n11575 | n22933 ;
  assign n22935 = n756 & ~n22934 ;
  assign n22936 = n12346 ^ n10333 ^ 1'b0 ;
  assign n22937 = ~n8478 & n22639 ;
  assign n22938 = ( n448 & ~n9273 ) | ( n448 & n22937 ) | ( ~n9273 & n22937 ) ;
  assign n22939 = n5834 & ~n13164 ;
  assign n22940 = n879 & ~n20369 ;
  assign n22941 = n1267 | n2706 ;
  assign n22942 = ( n5627 & ~n6717 ) | ( n5627 & n8341 ) | ( ~n6717 & n8341 ) ;
  assign n22943 = ~n237 & n1666 ;
  assign n22944 = n22943 ^ n3634 ^ 1'b0 ;
  assign n22945 = n22942 | n22944 ;
  assign n22946 = n22941 | n22945 ;
  assign n22947 = n10811 | n22946 ;
  assign n22948 = n17490 & ~n20970 ;
  assign n22949 = n16474 & n22948 ;
  assign n22950 = n22949 ^ n14623 ^ 1'b0 ;
  assign n22951 = n22950 ^ n18378 ^ n4944 ;
  assign n22952 = n4309 | n22951 ;
  assign n22953 = n2904 & n4856 ;
  assign n22954 = n22953 ^ n6860 ^ 1'b0 ;
  assign n22955 = n22954 ^ n10550 ^ 1'b0 ;
  assign n22956 = n20659 | n22955 ;
  assign n22957 = n12300 ^ n1078 ^ 1'b0 ;
  assign n22958 = ~n5456 & n22957 ;
  assign n22959 = ( ~n6297 & n7092 ) | ( ~n6297 & n14593 ) | ( n7092 & n14593 ) ;
  assign n22960 = n20203 ^ n9272 ^ 1'b0 ;
  assign n22961 = n22959 & ~n22960 ;
  assign n22962 = n57 & ~n22961 ;
  assign n22963 = ( n8846 & ~n9279 ) | ( n8846 & n20354 ) | ( ~n9279 & n20354 ) ;
  assign n22964 = n22963 ^ n22518 ^ 1'b0 ;
  assign n22965 = n696 & n8640 ;
  assign n22966 = n22965 ^ n9281 ^ 1'b0 ;
  assign n22970 = n7270 | n12502 ;
  assign n22967 = n630 ^ n604 ^ 1'b0 ;
  assign n22968 = n22967 ^ n9626 ^ n5145 ;
  assign n22969 = ~n5551 & n22968 ;
  assign n22971 = n22970 ^ n22969 ^ 1'b0 ;
  assign n22972 = n22966 & ~n22971 ;
  assign n22973 = ~n9982 & n19568 ;
  assign n22974 = ~n6406 & n22973 ;
  assign n22975 = n11983 ^ n6437 ^ 1'b0 ;
  assign n22978 = n2719 & ~n6230 ;
  assign n22979 = ~n5033 & n22978 ;
  assign n22976 = n15509 ^ n176 ^ 1'b0 ;
  assign n22977 = n16059 | n22976 ;
  assign n22980 = n22979 ^ n22977 ^ 1'b0 ;
  assign n22981 = n22980 ^ n16723 ^ 1'b0 ;
  assign n22982 = n22981 ^ n11877 ^ 1'b0 ;
  assign n22983 = n18931 | n22982 ;
  assign n22988 = n12877 ^ n153 ^ 1'b0 ;
  assign n22984 = n6870 ^ n6551 ^ 1'b0 ;
  assign n22985 = n14146 & ~n22984 ;
  assign n22986 = ~n14194 & n22985 ;
  assign n22987 = ~n8338 & n22986 ;
  assign n22989 = n22988 ^ n22987 ^ 1'b0 ;
  assign n22990 = ( n1210 & ~n4866 ) | ( n1210 & n13243 ) | ( ~n4866 & n13243 ) ;
  assign n22991 = n3406 & n7228 ;
  assign n22992 = n22990 & n22991 ;
  assign n22993 = n22992 ^ n9145 ^ 1'b0 ;
  assign n22994 = n16468 & ~n17466 ;
  assign n22995 = n22994 ^ n16220 ^ 1'b0 ;
  assign n22996 = n8753 & ~n11000 ;
  assign n22997 = ~n1502 & n19360 ;
  assign n22998 = ~n8287 & n22997 ;
  assign n22999 = ~n9013 & n12192 ;
  assign n23000 = n22999 ^ n5171 ^ 1'b0 ;
  assign n23001 = n8207 ^ n711 ^ 1'b0 ;
  assign n23002 = ~n5758 & n23001 ;
  assign n23003 = n23002 ^ n21151 ^ 1'b0 ;
  assign n23004 = n14995 ^ n10695 ^ n4944 ;
  assign n23005 = n350 & n23004 ;
  assign n23006 = n14695 ^ n2749 ^ 1'b0 ;
  assign n23007 = n23005 | n23006 ;
  assign n23011 = n8105 | n14620 ;
  assign n23012 = n23011 ^ n10816 ^ 1'b0 ;
  assign n23008 = n15631 ^ n10441 ^ n2104 ;
  assign n23009 = n16666 & ~n23008 ;
  assign n23010 = n5024 & ~n23009 ;
  assign n23013 = n23012 ^ n23010 ^ n10739 ;
  assign n23014 = n20288 ^ n14715 ^ n2110 ;
  assign n23015 = ( n2287 & n9397 ) | ( n2287 & ~n22612 ) | ( n9397 & ~n22612 ) ;
  assign n23018 = n20339 ^ n19775 ^ n4240 ;
  assign n23016 = ~n4757 & n12892 ;
  assign n23017 = n9495 & ~n23016 ;
  assign n23019 = n23018 ^ n23017 ^ 1'b0 ;
  assign n23020 = n17345 & n22094 ;
  assign n23021 = ~n2449 & n23020 ;
  assign n23022 = n10682 & n23021 ;
  assign n23023 = n5420 & ~n7265 ;
  assign n23025 = n2328 & n3398 ;
  assign n23024 = n6614 ^ n4078 ^ 1'b0 ;
  assign n23026 = n23025 ^ n23024 ^ n3710 ;
  assign n23027 = ( n89 & n5111 ) | ( n89 & n7046 ) | ( n5111 & n7046 ) ;
  assign n23028 = n10587 ^ n8907 ^ 1'b0 ;
  assign n23029 = n23028 ^ n7040 ^ 1'b0 ;
  assign n23030 = n21667 ^ n7541 ^ 1'b0 ;
  assign n23031 = n12423 ^ n9210 ^ 1'b0 ;
  assign n23032 = n8089 | n23031 ;
  assign n23033 = n14172 | n23032 ;
  assign n23037 = n3276 ^ n2913 ^ 1'b0 ;
  assign n23034 = n17166 & n22850 ;
  assign n23035 = n23034 ^ n18541 ^ 1'b0 ;
  assign n23036 = n12165 & ~n23035 ;
  assign n23038 = n23037 ^ n23036 ^ n3725 ;
  assign n23039 = n6616 & ~n10167 ;
  assign n23040 = ~n7935 & n23039 ;
  assign n23041 = n57 & n10835 ;
  assign n23042 = ~n12810 & n23041 ;
  assign n23043 = n2475 | n23042 ;
  assign n23044 = n23040 & ~n23043 ;
  assign n23045 = n18203 ^ n1015 ^ 1'b0 ;
  assign n23046 = ~n12036 & n23045 ;
  assign n23047 = n8526 ^ n2094 ^ 1'b0 ;
  assign n23048 = n11226 | n23047 ;
  assign n23049 = n4647 | n23048 ;
  assign n23050 = n8300 & n8787 ;
  assign n23051 = n12418 ^ n3061 ^ 1'b0 ;
  assign n23052 = n4345 | n23051 ;
  assign n23053 = n7827 | n19553 ;
  assign n23054 = n23053 ^ n7238 ^ 1'b0 ;
  assign n23055 = n23052 | n23054 ;
  assign n23056 = n5986 & n6527 ;
  assign n23057 = n23055 & n23056 ;
  assign n23058 = ~n18067 & n22536 ;
  assign n23059 = n12066 & n23058 ;
  assign n23060 = ~n3097 & n20087 ;
  assign n23061 = n22649 | n22743 ;
  assign n23062 = n23061 ^ n14554 ^ 1'b0 ;
  assign n23063 = n9115 ^ n6198 ^ 1'b0 ;
  assign n23064 = n11725 | n22427 ;
  assign n23065 = n11119 ^ n6896 ^ 1'b0 ;
  assign n23066 = n13546 ^ n360 ^ 1'b0 ;
  assign n23067 = n4647 & ~n16103 ;
  assign n23068 = n26 & n19216 ;
  assign n23069 = ~n2645 & n23068 ;
  assign n23070 = n23069 ^ n6111 ^ 1'b0 ;
  assign n23071 = n7856 & n23070 ;
  assign n23072 = n23071 ^ n14154 ^ 1'b0 ;
  assign n23073 = n23072 ^ n122 ^ 1'b0 ;
  assign n23074 = n22313 | n23073 ;
  assign n23075 = ( ~n1256 & n7383 ) | ( ~n1256 & n9667 ) | ( n7383 & n9667 ) ;
  assign n23076 = n23075 ^ n5311 ^ n1069 ;
  assign n23077 = n70 & n3500 ;
  assign n23078 = ~n2504 & n4622 ;
  assign n23079 = ~n3255 & n23078 ;
  assign n23080 = n23079 ^ n966 ^ 1'b0 ;
  assign n23081 = n23077 & ~n23080 ;
  assign n23082 = n10453 ^ n866 ^ 1'b0 ;
  assign n23083 = n226 | n23082 ;
  assign n23085 = ~n9820 & n12161 ;
  assign n23086 = n23085 ^ n10844 ^ 1'b0 ;
  assign n23084 = n4142 & n15953 ;
  assign n23087 = n23086 ^ n23084 ^ 1'b0 ;
  assign n23088 = n7146 | n10646 ;
  assign n23093 = n2579 & ~n19925 ;
  assign n23094 = n9619 & ~n23093 ;
  assign n23090 = n2964 ^ n2114 ^ n1435 ;
  assign n23089 = n978 ^ n842 ^ n532 ;
  assign n23091 = n23090 ^ n23089 ^ n4959 ;
  assign n23092 = n20781 & ~n23091 ;
  assign n23095 = n23094 ^ n23092 ^ 1'b0 ;
  assign n23096 = n23095 ^ n9643 ^ n523 ;
  assign n23097 = n2986 & n11223 ;
  assign n23098 = n3141 ^ n2106 ^ 1'b0 ;
  assign n23099 = n23097 & ~n23098 ;
  assign n23100 = ( ~n6578 & n10587 ) | ( ~n6578 & n23099 ) | ( n10587 & n23099 ) ;
  assign n23101 = n1918 & ~n9716 ;
  assign n23102 = n4113 & ~n9766 ;
  assign n23103 = n23102 ^ n6047 ^ 1'b0 ;
  assign n23104 = ( n5820 & n8093 ) | ( n5820 & ~n16922 ) | ( n8093 & ~n16922 ) ;
  assign n23105 = n23104 ^ n734 ^ 1'b0 ;
  assign n23106 = n3173 | n8171 ;
  assign n23107 = n7732 ^ n2837 ^ 1'b0 ;
  assign n23108 = n8159 | n23107 ;
  assign n23109 = n11383 ^ n7514 ^ 1'b0 ;
  assign n23110 = n23108 & ~n23109 ;
  assign n23111 = ( ~n2874 & n4704 ) | ( ~n2874 & n23110 ) | ( n4704 & n23110 ) ;
  assign n23112 = ( n19264 & ~n23106 ) | ( n19264 & n23111 ) | ( ~n23106 & n23111 ) ;
  assign n23113 = ~n4275 & n15005 ;
  assign n23114 = n5878 | n9753 ;
  assign n23115 = n8407 | n23114 ;
  assign n23116 = n12440 ^ n2605 ^ 1'b0 ;
  assign n23117 = n711 & n23116 ;
  assign n23118 = n23117 ^ n6576 ^ 1'b0 ;
  assign n23119 = n23115 & ~n23118 ;
  assign n23120 = ~n23113 & n23119 ;
  assign n23121 = n21494 ^ n2356 ^ 1'b0 ;
  assign n23122 = n15821 ^ n2070 ^ n398 ;
  assign n23123 = ~n4369 & n23122 ;
  assign n23124 = n23123 ^ n20834 ^ 1'b0 ;
  assign n23125 = n10946 ^ n588 ^ 1'b0 ;
  assign n23126 = n13081 & n23125 ;
  assign n23127 = ( n63 & ~n11383 ) | ( n63 & n12003 ) | ( ~n11383 & n12003 ) ;
  assign n23128 = ( n8515 & n15926 ) | ( n8515 & n23127 ) | ( n15926 & n23127 ) ;
  assign n23129 = n17850 & n23128 ;
  assign n23130 = ~n23126 & n23129 ;
  assign n23131 = n16414 ^ n12986 ^ 1'b0 ;
  assign n23132 = ( ~n3145 & n20066 ) | ( ~n3145 & n22979 ) | ( n20066 & n22979 ) ;
  assign n23133 = n10679 ^ n1459 ^ n702 ;
  assign n23134 = ~n14763 & n23133 ;
  assign n23135 = ~n23132 & n23134 ;
  assign n23136 = n1218 & n9360 ;
  assign n23137 = n20250 ^ n7479 ^ 1'b0 ;
  assign n23138 = n23137 ^ n22879 ^ n4864 ;
  assign n23139 = ( n1744 & n3350 ) | ( n1744 & n22084 ) | ( n3350 & n22084 ) ;
  assign n23140 = n23139 ^ n8019 ^ 1'b0 ;
  assign n23141 = n4900 | n23140 ;
  assign n23142 = n16738 | n23141 ;
  assign n23143 = n9685 & n13275 ;
  assign n23144 = n23143 ^ n22989 ^ 1'b0 ;
  assign n23145 = ( ~n6750 & n11134 ) | ( ~n6750 & n22267 ) | ( n11134 & n22267 ) ;
  assign n23146 = n14620 ^ n13651 ^ 1'b0 ;
  assign n23147 = ~n4863 & n23146 ;
  assign n23148 = n9042 ^ n6754 ^ 1'b0 ;
  assign n23149 = n5457 & ~n9580 ;
  assign n23150 = n14523 ^ n7768 ^ 1'b0 ;
  assign n23151 = n23150 ^ n2772 ^ n455 ;
  assign n23152 = ( n8447 & n13611 ) | ( n8447 & n16597 ) | ( n13611 & n16597 ) ;
  assign n23153 = n2374 & n19052 ;
  assign n23154 = n23153 ^ n5520 ^ 1'b0 ;
  assign n23155 = ~n23152 & n23154 ;
  assign n23156 = ( n6743 & n7543 ) | ( n6743 & n23155 ) | ( n7543 & n23155 ) ;
  assign n23157 = n15111 & ~n23156 ;
  assign n23158 = n18127 & n23157 ;
  assign n23159 = n9813 | n23158 ;
  assign n23160 = n5873 ^ n5366 ^ 1'b0 ;
  assign n23161 = ~n5891 & n23160 ;
  assign n23162 = n11973 ^ n11685 ^ n9298 ;
  assign n23163 = n20795 ^ n6415 ^ 1'b0 ;
  assign n23164 = n13749 | n23163 ;
  assign n23165 = n1562 | n10861 ;
  assign n23166 = n12003 ^ n5742 ^ 1'b0 ;
  assign n23167 = n10965 & ~n23166 ;
  assign n23168 = n1362 & n23167 ;
  assign n23169 = n3390 & n4599 ;
  assign n23170 = n15942 & n23169 ;
  assign n23171 = ~n23168 & n23170 ;
  assign n23172 = n13554 ^ n8947 ^ 1'b0 ;
  assign n23173 = n8257 & n23172 ;
  assign n23175 = n1691 | n10493 ;
  assign n23176 = n23175 ^ n10350 ^ 1'b0 ;
  assign n23174 = ( n440 & n4956 ) | ( n440 & n8889 ) | ( n4956 & n8889 ) ;
  assign n23177 = n23176 ^ n23174 ^ 1'b0 ;
  assign n23178 = n12918 ^ n2933 ^ 1'b0 ;
  assign n23179 = ( n787 & n18061 ) | ( n787 & n23178 ) | ( n18061 & n23178 ) ;
  assign n23180 = n15064 ^ n7169 ^ 1'b0 ;
  assign n23181 = n9748 & ~n23180 ;
  assign n23182 = n6954 | n12295 ;
  assign n23183 = n22812 | n23182 ;
  assign n23184 = n10842 | n13378 ;
  assign n23185 = n23183 | n23184 ;
  assign n23186 = ~n2271 & n3067 ;
  assign n23187 = n13942 & n23186 ;
  assign n23188 = ( n1931 & ~n12095 ) | ( n1931 & n13004 ) | ( ~n12095 & n13004 ) ;
  assign n23189 = n23188 ^ n4050 ^ 1'b0 ;
  assign n23190 = ~n7636 & n15824 ;
  assign n23191 = n16762 ^ n9417 ^ 1'b0 ;
  assign n23192 = n1969 & ~n6951 ;
  assign n23193 = ~n5406 & n23192 ;
  assign n23194 = n23193 ^ n8533 ^ n8077 ;
  assign n23195 = ( n17156 & n18739 ) | ( n17156 & n23194 ) | ( n18739 & n23194 ) ;
  assign n23196 = n6380 | n19468 ;
  assign n23197 = n23196 ^ n9402 ^ 1'b0 ;
  assign n23198 = n22599 ^ n4951 ^ 1'b0 ;
  assign n23199 = n612 & n23198 ;
  assign n23200 = ( n1917 & n11337 ) | ( n1917 & ~n19256 ) | ( n11337 & ~n19256 ) ;
  assign n23201 = n23199 & n23200 ;
  assign n23202 = ~n23197 & n23201 ;
  assign n23203 = ( n601 & ~n817 ) | ( n601 & n968 ) | ( ~n817 & n968 ) ;
  assign n23204 = n14583 & ~n23203 ;
  assign n23205 = n19714 ^ n15084 ^ 1'b0 ;
  assign n23207 = n9358 & n15229 ;
  assign n23206 = n91 & n10021 ;
  assign n23208 = n23207 ^ n23206 ^ 1'b0 ;
  assign n23209 = n7188 | n10708 ;
  assign n23210 = n23209 ^ n14445 ^ 1'b0 ;
  assign n23211 = n5231 & ~n6951 ;
  assign n23212 = n16189 & n20038 ;
  assign n23213 = n2622 | n5052 ;
  assign n23214 = n23213 ^ n1459 ^ 1'b0 ;
  assign n23215 = n8375 & n23214 ;
  assign n23216 = n4805 & ~n23215 ;
  assign n23217 = n1767 & n7505 ;
  assign n23219 = ~n1389 & n1854 ;
  assign n23220 = ~n1889 & n23219 ;
  assign n23221 = n2806 & ~n23220 ;
  assign n23218 = n1109 | n1287 ;
  assign n23222 = n23221 ^ n23218 ^ 1'b0 ;
  assign n23223 = n9683 | n15153 ;
  assign n23224 = n23223 ^ n4549 ^ 1'b0 ;
  assign n23225 = ( ~n1736 & n3634 ) | ( ~n1736 & n15889 ) | ( n3634 & n15889 ) ;
  assign n23230 = n976 | n4529 ;
  assign n23226 = n228 & n975 ;
  assign n23227 = n23226 ^ n1522 ^ 1'b0 ;
  assign n23228 = n8093 & n23227 ;
  assign n23229 = n23228 ^ n9081 ^ 1'b0 ;
  assign n23231 = n23230 ^ n23229 ^ 1'b0 ;
  assign n23232 = n22874 & n23231 ;
  assign n23233 = n1050 | n10709 ;
  assign n23234 = n23233 ^ n6292 ^ 1'b0 ;
  assign n23235 = n2677 & n18977 ;
  assign n23236 = n3789 | n16411 ;
  assign n23237 = ~n3870 & n23236 ;
  assign n23238 = n14781 ^ n7717 ^ 1'b0 ;
  assign n23239 = n1409 & ~n10677 ;
  assign n23240 = n14329 | n23239 ;
  assign n23241 = n4243 | n23240 ;
  assign n23242 = n23238 | n23241 ;
  assign n23243 = n2882 | n3435 ;
  assign n23244 = n2414 | n23243 ;
  assign n23245 = n23244 ^ n11363 ^ 1'b0 ;
  assign n23246 = n23245 ^ n3165 ^ 1'b0 ;
  assign n23247 = n434 & ~n23246 ;
  assign n23248 = n4671 ^ n3995 ^ 1'b0 ;
  assign n23249 = n23247 & n23248 ;
  assign n23250 = n23249 ^ n14047 ^ 1'b0 ;
  assign n23251 = n4427 ^ n890 ^ 1'b0 ;
  assign n23252 = ~n13473 & n23251 ;
  assign n23253 = n10070 & n11454 ;
  assign n23254 = ~n23252 & n23253 ;
  assign n23255 = n3953 ^ n361 ^ 1'b0 ;
  assign n23256 = ~n23254 & n23255 ;
  assign n23258 = n14185 ^ n6287 ^ n4835 ;
  assign n23257 = n5551 & ~n14229 ;
  assign n23259 = n23258 ^ n23257 ^ n5888 ;
  assign n23260 = n6481 | n18688 ;
  assign n23261 = n23260 ^ n8409 ^ 1'b0 ;
  assign n23262 = ( n17929 & n23200 ) | ( n17929 & n23261 ) | ( n23200 & n23261 ) ;
  assign n23263 = n6196 & ~n7056 ;
  assign n23264 = n23263 ^ n5469 ^ 1'b0 ;
  assign n23265 = n3530 & ~n23264 ;
  assign n23266 = ~n2695 & n23265 ;
  assign n23267 = n23266 ^ n15918 ^ 1'b0 ;
  assign n23268 = n20306 ^ n10183 ^ n349 ;
  assign n23269 = ( ~n6034 & n20070 ) | ( ~n6034 & n23268 ) | ( n20070 & n23268 ) ;
  assign n23270 = n6095 & ~n16551 ;
  assign n23271 = n23270 ^ n18570 ^ n15454 ;
  assign n23272 = ~n41 & n7633 ;
  assign n23273 = ~n7633 & n23272 ;
  assign n23274 = n991 & ~n23273 ;
  assign n23275 = n23273 & n23274 ;
  assign n23276 = n3608 ^ n1549 ^ 1'b0 ;
  assign n23277 = ~n954 & n23276 ;
  assign n23278 = n23277 ^ n18493 ^ 1'b0 ;
  assign n23279 = n1296 & ~n12181 ;
  assign n23280 = n3245 & ~n15153 ;
  assign n23281 = ~n169 & n23280 ;
  assign n23282 = n2725 & ~n3824 ;
  assign n23283 = n23282 ^ n6462 ^ n745 ;
  assign n23284 = n191 & ~n7468 ;
  assign n23285 = ~n20309 & n23284 ;
  assign n23286 = n23283 & ~n23285 ;
  assign n23287 = n23281 | n23286 ;
  assign n23288 = n7074 & ~n23287 ;
  assign n23289 = n1204 & n12056 ;
  assign n23290 = n23289 ^ n16823 ^ 1'b0 ;
  assign n23291 = n23290 ^ n12372 ^ 1'b0 ;
  assign n23292 = n15317 & ~n23291 ;
  assign n23294 = n15026 ^ n9694 ^ 1'b0 ;
  assign n23293 = n3949 & n18623 ;
  assign n23295 = n23294 ^ n23293 ^ 1'b0 ;
  assign n23296 = n5391 & ~n14316 ;
  assign n23297 = n14937 ^ n4345 ^ 1'b0 ;
  assign n23299 = ( n13945 & ~n19047 ) | ( n13945 & n20368 ) | ( ~n19047 & n20368 ) ;
  assign n23298 = ( ~n139 & n5873 ) | ( ~n139 & n6089 ) | ( n5873 & n6089 ) ;
  assign n23300 = n23299 ^ n23298 ^ n3076 ;
  assign n23301 = n188 & n2867 ;
  assign n23302 = ~n99 & n23301 ;
  assign n23303 = n13548 | n23302 ;
  assign n23304 = n23303 ^ n592 ^ 1'b0 ;
  assign n23305 = n13427 ^ n10705 ^ n10088 ;
  assign n23310 = n8665 & ~n10939 ;
  assign n23311 = n23310 ^ n4363 ^ 1'b0 ;
  assign n23309 = n1084 | n4962 ;
  assign n23312 = n23311 ^ n23309 ^ n6133 ;
  assign n23306 = n6783 | n10176 ;
  assign n23307 = n672 & n23306 ;
  assign n23308 = ~n760 & n23307 ;
  assign n23313 = n23312 ^ n23308 ^ n4536 ;
  assign n23314 = n14593 ^ n6181 ^ 1'b0 ;
  assign n23315 = ( x7 & n4346 ) | ( x7 & ~n7099 ) | ( n4346 & ~n7099 ) ;
  assign n23316 = n1443 & ~n23315 ;
  assign n23317 = n12339 ^ n4710 ^ 1'b0 ;
  assign n23318 = n23317 ^ n14136 ^ 1'b0 ;
  assign n23319 = n17841 ^ n16761 ^ 1'b0 ;
  assign n23320 = n4056 & ~n23319 ;
  assign n23321 = n7545 & ~n18234 ;
  assign n23322 = n955 & n23321 ;
  assign n23323 = n4565 & ~n23322 ;
  assign n23324 = ~n10966 & n23323 ;
  assign n23325 = n23324 ^ n6278 ^ 1'b0 ;
  assign n23326 = ~n9934 & n23325 ;
  assign n23327 = n11880 ^ n6668 ^ 1'b0 ;
  assign n23328 = n3784 & ~n23327 ;
  assign n23329 = n13427 ^ n10451 ^ n3168 ;
  assign n23330 = n15112 & n23329 ;
  assign n23333 = n4848 ^ n2230 ^ n1093 ;
  assign n23334 = n22161 ^ n15666 ^ 1'b0 ;
  assign n23335 = ~n23333 & n23334 ;
  assign n23331 = ~n2139 & n13382 ;
  assign n23332 = n20508 & n23331 ;
  assign n23336 = n23335 ^ n23332 ^ 1'b0 ;
  assign n23337 = n7402 & ~n23336 ;
  assign n23338 = n15349 ^ n4989 ^ n4841 ;
  assign n23339 = n7169 & n23338 ;
  assign n23340 = ~n580 & n23339 ;
  assign n23341 = n23340 ^ n13900 ^ 1'b0 ;
  assign n23342 = n21202 ^ n13644 ^ 1'b0 ;
  assign n23343 = n4986 | n13379 ;
  assign n23344 = n22966 ^ n18160 ^ 1'b0 ;
  assign n23345 = ~n3575 & n5693 ;
  assign n23346 = n12784 ^ n6995 ^ 1'b0 ;
  assign n23347 = n12808 & n23346 ;
  assign n23348 = n2735 | n17179 ;
  assign n23349 = n23348 ^ n19038 ^ 1'b0 ;
  assign n23355 = n8593 & ~n21508 ;
  assign n23353 = n6133 | n17226 ;
  assign n23354 = n23353 ^ n4944 ^ 1'b0 ;
  assign n23350 = ~n4896 & n8800 ;
  assign n23351 = n23350 ^ n21794 ^ 1'b0 ;
  assign n23352 = n4982 & ~n23351 ;
  assign n23356 = n23355 ^ n23354 ^ n23352 ;
  assign n23357 = ( ~n10397 & n14745 ) | ( ~n10397 & n15923 ) | ( n14745 & n15923 ) ;
  assign n23358 = n7802 & n9493 ;
  assign n23359 = n1353 & n23358 ;
  assign n23360 = n16356 & n20328 ;
  assign n23361 = ~n5612 & n23360 ;
  assign n23362 = n13516 ^ n1523 ^ 1'b0 ;
  assign n23364 = ( ~n263 & n4055 ) | ( ~n263 & n8700 ) | ( n4055 & n8700 ) ;
  assign n23363 = n5013 ^ n2225 ^ 1'b0 ;
  assign n23365 = n23364 ^ n23363 ^ 1'b0 ;
  assign n23366 = n8526 & n23365 ;
  assign n23367 = n5261 ^ n2030 ^ 1'b0 ;
  assign n23368 = n6286 & n23367 ;
  assign n23369 = ( n2790 & n12259 ) | ( n2790 & n23368 ) | ( n12259 & n23368 ) ;
  assign n23370 = n9060 & ~n21262 ;
  assign n23371 = n10433 & n23370 ;
  assign n23372 = n6399 | n8382 ;
  assign n23373 = n20805 | n23372 ;
  assign n23374 = n8254 & n23373 ;
  assign n23375 = n23374 ^ n20425 ^ 1'b0 ;
  assign n23376 = n350 & ~n8145 ;
  assign n23377 = n9734 & n11405 ;
  assign n23378 = n23376 & n23377 ;
  assign n23379 = n5683 & ~n6261 ;
  assign n23380 = n23379 ^ n11743 ^ 1'b0 ;
  assign n23381 = n3866 | n17411 ;
  assign n23382 = ~n1560 & n18555 ;
  assign n23383 = n18382 ^ n12191 ^ 1'b0 ;
  assign n23384 = n1189 & n5477 ;
  assign n23385 = n7543 & n15956 ;
  assign n23386 = n23385 ^ n15382 ^ 1'b0 ;
  assign n23387 = n22376 | n22681 ;
  assign n23388 = n4758 ^ n281 ^ 1'b0 ;
  assign n23389 = n2926 | n16635 ;
  assign n23390 = n23388 & ~n23389 ;
  assign n23391 = n4906 | n23390 ;
  assign n23392 = n12257 ^ n3029 ^ 1'b0 ;
  assign n23393 = n8520 | n8970 ;
  assign n23394 = n23392 & n23393 ;
  assign n23395 = n21471 ^ n20262 ^ 1'b0 ;
  assign n23396 = ~n4385 & n6238 ;
  assign n23397 = n23396 ^ n16389 ^ 1'b0 ;
  assign n23398 = n17940 | n23397 ;
  assign n23399 = n23047 ^ n12383 ^ n5162 ;
  assign n23400 = n23399 ^ n15631 ^ 1'b0 ;
  assign n23401 = n23400 ^ n11934 ^ n1131 ;
  assign n23402 = n23401 ^ n18048 ^ 1'b0 ;
  assign n23403 = n8539 ^ n3985 ^ 1'b0 ;
  assign n23404 = ~n14305 & n23403 ;
  assign n23405 = ~n2832 & n3786 ;
  assign n23406 = ~n17197 & n23405 ;
  assign n23407 = n9621 & ~n12002 ;
  assign n23408 = n4886 ^ n2587 ^ 1'b0 ;
  assign n23409 = n23407 & ~n23408 ;
  assign n23410 = n23409 ^ n63 ^ 1'b0 ;
  assign n23411 = n9204 ^ n953 ^ 1'b0 ;
  assign n23412 = n8127 | n18498 ;
  assign n23413 = ~n5032 & n23412 ;
  assign n23414 = n23413 ^ n12451 ^ 1'b0 ;
  assign n23415 = n12661 & ~n23414 ;
  assign n23416 = ~n18690 & n23415 ;
  assign n23418 = n6060 & ~n11711 ;
  assign n23417 = ~n1668 & n14907 ;
  assign n23419 = n23418 ^ n23417 ^ 1'b0 ;
  assign n23420 = n23419 ^ n13956 ^ 1'b0 ;
  assign n23422 = ~n8390 & n14282 ;
  assign n23423 = ~n12083 & n23422 ;
  assign n23421 = n3909 & n7575 ;
  assign n23424 = n23423 ^ n23421 ^ 1'b0 ;
  assign n23425 = n20848 & ~n23230 ;
  assign n23426 = n23425 ^ n11258 ^ 1'b0 ;
  assign n23428 = ~n1926 & n9935 ;
  assign n23427 = n578 & ~n18324 ;
  assign n23429 = n23428 ^ n23427 ^ 1'b0 ;
  assign n23430 = ~n23426 & n23429 ;
  assign n23431 = ( n6966 & n10189 ) | ( n6966 & ~n19282 ) | ( n10189 & ~n19282 ) ;
  assign n23432 = ( ~n9045 & n11170 ) | ( ~n9045 & n13266 ) | ( n11170 & n13266 ) ;
  assign n23433 = n23432 ^ n2405 ^ 1'b0 ;
  assign n23434 = n23433 ^ n5167 ^ 1'b0 ;
  assign n23435 = n6904 | n23434 ;
  assign n23436 = n8009 | n19092 ;
  assign n23437 = n12933 & ~n23436 ;
  assign n23438 = n7760 & ~n23437 ;
  assign n23439 = n23438 ^ n21773 ^ 1'b0 ;
  assign n23440 = ~n5546 & n7327 ;
  assign n23441 = n4930 & ~n9921 ;
  assign n23442 = n23440 & ~n23441 ;
  assign n23443 = ~n5667 & n17336 ;
  assign n23444 = ( n10347 & n20872 ) | ( n10347 & ~n23443 ) | ( n20872 & ~n23443 ) ;
  assign n23446 = n11587 ^ n8414 ^ n2880 ;
  assign n23447 = n12214 | n23446 ;
  assign n23445 = n1647 & n22040 ;
  assign n23448 = n23447 ^ n23445 ^ 1'b0 ;
  assign n23449 = n609 | n4830 ;
  assign n23450 = ~n21683 & n23449 ;
  assign n23451 = n23450 ^ n11245 ^ 1'b0 ;
  assign n23452 = n18106 | n18562 ;
  assign n23453 = n12460 | n23452 ;
  assign n23454 = n1316 | n23453 ;
  assign n23455 = ( n1864 & ~n5387 ) | ( n1864 & n6909 ) | ( ~n5387 & n6909 ) ;
  assign n23456 = n23455 ^ n4812 ^ 1'b0 ;
  assign n23457 = n12032 & ~n23456 ;
  assign n23458 = ~n4549 & n4943 ;
  assign n23459 = n6500 ^ n3000 ^ 1'b0 ;
  assign n23460 = ~n23458 & n23459 ;
  assign n23461 = ~n11719 & n23460 ;
  assign n23462 = n15770 | n23461 ;
  assign n23463 = n23462 ^ n5554 ^ 1'b0 ;
  assign n23464 = ~n2992 & n3362 ;
  assign n23465 = n23464 ^ n1676 ^ 1'b0 ;
  assign n23466 = n21387 & n23465 ;
  assign n23467 = n3898 & n23466 ;
  assign n23468 = n23467 ^ n14626 ^ 1'b0 ;
  assign n23469 = n16305 & n19367 ;
  assign n23470 = n2514 & n12321 ;
  assign n23471 = n9453 ^ n6064 ^ n4043 ;
  assign n23472 = n23470 & ~n23471 ;
  assign n23473 = n523 | n9813 ;
  assign n23474 = n23473 ^ n20648 ^ 1'b0 ;
  assign n23476 = ~n6776 & n10254 ;
  assign n23475 = n10657 & n15256 ;
  assign n23477 = n23476 ^ n23475 ^ 1'b0 ;
  assign n23478 = n8076 & n11873 ;
  assign n23479 = n23478 ^ n8342 ^ 1'b0 ;
  assign n23480 = n6756 ^ n4543 ^ 1'b0 ;
  assign n23481 = n15854 & n23480 ;
  assign n23482 = n12298 ^ n7240 ^ n1126 ;
  assign n23483 = n5806 & ~n23482 ;
  assign n23484 = n8301 | n8547 ;
  assign n23485 = n23484 ^ n2287 ^ 1'b0 ;
  assign n23486 = n2117 | n21679 ;
  assign n23487 = ( n3406 & n10815 ) | ( n3406 & n23486 ) | ( n10815 & n23486 ) ;
  assign n23488 = n13804 & ~n23487 ;
  assign n23489 = ~n2495 & n10095 ;
  assign n23490 = n46 & ~n11994 ;
  assign n23491 = n23490 ^ n9964 ^ 1'b0 ;
  assign n23492 = n23491 ^ n21202 ^ n11345 ;
  assign n23493 = n4195 ^ n3717 ^ 1'b0 ;
  assign n23494 = ~n23047 & n23493 ;
  assign n23495 = ~n23492 & n23494 ;
  assign n23496 = n19220 ^ n8486 ^ 1'b0 ;
  assign n23497 = n63 & n23496 ;
  assign n23498 = ~n10952 & n23497 ;
  assign n23499 = ~n9434 & n23498 ;
  assign n23500 = n9017 & ~n23499 ;
  assign n23501 = ( ~n4142 & n17046 ) | ( ~n4142 & n23500 ) | ( n17046 & n23500 ) ;
  assign n23502 = ~n5127 & n14074 ;
  assign n23503 = n23502 ^ n1600 ^ 1'b0 ;
  assign n23504 = n9376 ^ n5140 ^ 1'b0 ;
  assign n23505 = n23503 | n23504 ;
  assign n23506 = n997 & ~n23505 ;
  assign n23507 = n23506 ^ n11088 ^ 1'b0 ;
  assign n23508 = n1658 | n6582 ;
  assign n23509 = n18590 | n23508 ;
  assign n23510 = n23509 ^ n13004 ^ 1'b0 ;
  assign n23511 = n19823 ^ n14895 ^ 1'b0 ;
  assign n23512 = n23511 ^ n7925 ^ 1'b0 ;
  assign n23513 = n23510 | n23512 ;
  assign n23514 = n5891 ^ n1532 ^ 1'b0 ;
  assign n23515 = ~n6865 & n23514 ;
  assign n23516 = n5265 | n23515 ;
  assign n23517 = n9663 ^ n4752 ^ 1'b0 ;
  assign n23518 = n17665 & ~n21718 ;
  assign n23519 = n22834 & n23518 ;
  assign n23520 = n308 | n2203 ;
  assign n23521 = n4397 ^ n1374 ^ 1'b0 ;
  assign n23522 = n23520 | n23521 ;
  assign n23523 = n21955 ^ n41 ^ 1'b0 ;
  assign n23524 = ~n11632 & n23523 ;
  assign n23525 = n4136 & n7832 ;
  assign n23526 = n23525 ^ n15569 ^ 1'b0 ;
  assign n23527 = n23526 ^ n22290 ^ n1573 ;
  assign n23528 = n17335 ^ n4785 ^ 1'b0 ;
  assign n23529 = n3043 | n8143 ;
  assign n23530 = n23529 ^ n13689 ^ 1'b0 ;
  assign n23531 = n6275 & n11785 ;
  assign n23532 = n4427 ^ n331 ^ 1'b0 ;
  assign n23533 = n8551 & n10123 ;
  assign n23534 = n23533 ^ n6676 ^ 1'b0 ;
  assign n23535 = ~n23532 & n23534 ;
  assign n23536 = ~n16444 & n20363 ;
  assign n23545 = n1179 & ~n7319 ;
  assign n23546 = n23545 ^ n7126 ^ 1'b0 ;
  assign n23547 = n23546 ^ n1064 ^ 1'b0 ;
  assign n23548 = ~n9318 & n23547 ;
  assign n23549 = ~n498 & n11513 ;
  assign n23550 = n12490 & n23549 ;
  assign n23551 = ~n11634 & n23550 ;
  assign n23552 = n16489 & n23551 ;
  assign n23553 = n23548 & n23552 ;
  assign n23542 = n5080 | n17101 ;
  assign n23539 = x8 & ~n1704 ;
  assign n23538 = ~n4683 & n7272 ;
  assign n23537 = n12777 ^ n5675 ^ 1'b0 ;
  assign n23540 = n23539 ^ n23538 ^ n23537 ;
  assign n23541 = ~n15543 & n23540 ;
  assign n23543 = n23542 ^ n23541 ^ 1'b0 ;
  assign n23544 = ~n20357 & n23543 ;
  assign n23554 = n23553 ^ n23544 ^ 1'b0 ;
  assign n23555 = n5011 ^ n4578 ^ 1'b0 ;
  assign n23556 = n11915 | n23555 ;
  assign n23557 = n829 & ~n8542 ;
  assign n23558 = ~n601 & n23557 ;
  assign n23559 = n10793 ^ n9541 ^ 1'b0 ;
  assign n23560 = ~n3227 & n23559 ;
  assign n23561 = n17468 & n23560 ;
  assign n23562 = n23558 & n23561 ;
  assign n23563 = n208 | n6221 ;
  assign n23564 = n3094 | n23563 ;
  assign n23567 = n12327 & ~n14929 ;
  assign n23565 = n8421 & n16648 ;
  assign n23566 = ~n12289 & n23565 ;
  assign n23568 = n23567 ^ n23566 ^ 1'b0 ;
  assign n23569 = n10668 ^ n2550 ^ 1'b0 ;
  assign n23570 = n19726 ^ n18912 ^ 1'b0 ;
  assign n23571 = ~n3581 & n10438 ;
  assign n23572 = n1140 ^ n572 ^ 1'b0 ;
  assign n23573 = n23571 | n23572 ;
  assign n23574 = n23573 ^ n3326 ^ 1'b0 ;
  assign n23575 = ~n3274 & n5741 ;
  assign n23576 = ~n5051 & n23575 ;
  assign n23577 = n6704 ^ n2162 ^ 1'b0 ;
  assign n23578 = ~n7895 & n23577 ;
  assign n23579 = n23578 ^ n19210 ^ n5935 ;
  assign n23580 = n6556 | n18152 ;
  assign n23581 = n23580 ^ n6083 ^ 1'b0 ;
  assign n23582 = ( ~n1040 & n16802 ) | ( ~n1040 & n21482 ) | ( n16802 & n21482 ) ;
  assign n23583 = n3914 | n9805 ;
  assign n23584 = n6542 & n20644 ;
  assign n23585 = ~n23583 & n23584 ;
  assign n23587 = n119 & n624 ;
  assign n23588 = n23587 ^ n11225 ^ 1'b0 ;
  assign n23589 = n10722 | n23588 ;
  assign n23590 = n15632 & ~n23589 ;
  assign n23586 = n710 & ~n12006 ;
  assign n23591 = n23590 ^ n23586 ^ 1'b0 ;
  assign n23592 = n3560 & ~n17751 ;
  assign n23593 = n23592 ^ n15423 ^ n1182 ;
  assign n23594 = n23593 ^ n16359 ^ 1'b0 ;
  assign n23595 = n5815 | n23594 ;
  assign n23596 = ( n160 & ~n4222 ) | ( n160 & n4697 ) | ( ~n4222 & n4697 ) ;
  assign n23597 = n18928 & ~n20716 ;
  assign n23598 = ~n23596 & n23597 ;
  assign n23599 = n8888 | n21546 ;
  assign n23600 = n23599 ^ n11042 ^ 1'b0 ;
  assign n23601 = n21941 ^ n15693 ^ 1'b0 ;
  assign n23602 = n111 | n23601 ;
  assign n23603 = n14675 & ~n23602 ;
  assign n23604 = n21489 ^ n18894 ^ 1'b0 ;
  assign n23605 = ~n10523 & n23604 ;
  assign n23606 = ~n12272 & n17780 ;
  assign n23607 = n10503 | n23606 ;
  assign n23608 = n23607 ^ n13587 ^ 1'b0 ;
  assign n23609 = ~n3517 & n23608 ;
  assign n23619 = n6274 | n8157 ;
  assign n23610 = n4523 ^ n1902 ^ 1'b0 ;
  assign n23613 = n17389 ^ n1611 ^ 1'b0 ;
  assign n23614 = n12739 & ~n23613 ;
  assign n23611 = n15130 & n15402 ;
  assign n23612 = n1495 & ~n23611 ;
  assign n23615 = n23614 ^ n23612 ^ 1'b0 ;
  assign n23616 = n2199 & n23615 ;
  assign n23617 = n14688 & ~n23616 ;
  assign n23618 = ~n23610 & n23617 ;
  assign n23620 = n23619 ^ n23618 ^ 1'b0 ;
  assign n23621 = ~n4835 & n7507 ;
  assign n23622 = n23621 ^ n4303 ^ 1'b0 ;
  assign n23623 = n23622 ^ n16858 ^ n6845 ;
  assign n23624 = n5130 & ~n14930 ;
  assign n23625 = ~n113 & n23624 ;
  assign n23626 = n19785 | n23625 ;
  assign n23627 = n4149 & n4584 ;
  assign n23628 = n23627 ^ n10939 ^ 1'b0 ;
  assign n23629 = ( ~n8526 & n10662 ) | ( ~n8526 & n19529 ) | ( n10662 & n19529 ) ;
  assign n23630 = ~n11274 & n18074 ;
  assign n23631 = n23630 ^ n18193 ^ n12849 ;
  assign n23632 = n7471 & ~n17372 ;
  assign n23633 = n23632 ^ n15949 ^ 1'b0 ;
  assign n23634 = n3709 & n18157 ;
  assign n23635 = ~n13821 & n23634 ;
  assign n23636 = n6011 ^ n5353 ^ 1'b0 ;
  assign n23637 = n6149 ^ n4951 ^ 1'b0 ;
  assign n23638 = n23636 & ~n23637 ;
  assign n23639 = n21148 & n23486 ;
  assign n23640 = n16347 ^ n16070 ^ n5120 ;
  assign n23641 = n14923 | n16717 ;
  assign n23642 = n23641 ^ n6019 ^ 1'b0 ;
  assign n23643 = n1143 | n8603 ;
  assign n23644 = n23643 ^ n723 ^ 1'b0 ;
  assign n23645 = n21131 ^ n16948 ^ 1'b0 ;
  assign n23646 = n12915 & n14755 ;
  assign n23647 = n12845 | n23646 ;
  assign n23648 = n2561 & n15026 ;
  assign n23649 = n4858 ^ n3528 ^ 1'b0 ;
  assign n23650 = n5915 & ~n23649 ;
  assign n23651 = n23650 ^ n1988 ^ 1'b0 ;
  assign n23652 = n23648 & ~n23651 ;
  assign n23653 = n23652 ^ n2567 ^ 1'b0 ;
  assign n23654 = n8676 & ~n23653 ;
  assign n23655 = n13879 & n23654 ;
  assign n23656 = n23655 ^ n4710 ^ 1'b0 ;
  assign n23657 = n15552 & ~n23656 ;
  assign n23658 = n23657 ^ n17241 ^ 1'b0 ;
  assign n23659 = n13180 & ~n23658 ;
  assign n23660 = n11764 & n19580 ;
  assign n23661 = n4381 | n23660 ;
  assign n23662 = n172 & ~n8660 ;
  assign n23663 = n23662 ^ n145 ^ 1'b0 ;
  assign n23664 = n8857 | n23663 ;
  assign n23665 = n11606 | n23664 ;
  assign n23666 = ~n3959 & n4273 ;
  assign n23667 = n23666 ^ n263 ^ 1'b0 ;
  assign n23668 = n4214 ^ n2946 ^ 1'b0 ;
  assign n23669 = n19662 ^ n1533 ^ 1'b0 ;
  assign n23670 = n4875 & n7026 ;
  assign n23671 = n21198 ^ n2692 ^ 1'b0 ;
  assign n23672 = n23670 & n23671 ;
  assign n23673 = n3797 | n13866 ;
  assign n23674 = n23673 ^ n1545 ^ 1'b0 ;
  assign n23675 = ( n289 & n23672 ) | ( n289 & ~n23674 ) | ( n23672 & ~n23674 ) ;
  assign n23676 = n9109 | n23675 ;
  assign n23677 = n23676 ^ n6139 ^ 1'b0 ;
  assign n23678 = ~n5178 & n23677 ;
  assign n23679 = n10854 | n11219 ;
  assign n23680 = n2953 | n23679 ;
  assign n23681 = ~n22935 & n23664 ;
  assign n23682 = n7920 & ~n14951 ;
  assign n23683 = n23682 ^ n2729 ^ 1'b0 ;
  assign n23684 = n21336 ^ n10626 ^ n9145 ;
  assign n23685 = n23684 ^ n11667 ^ 1'b0 ;
  assign n23686 = n5867 ^ n4721 ^ 1'b0 ;
  assign n23687 = n23542 ^ n23137 ^ n20220 ;
  assign n23688 = n23687 ^ n13582 ^ 1'b0 ;
  assign n23689 = n23315 & ~n23688 ;
  assign n23690 = n2028 & ~n8807 ;
  assign n23691 = n23690 ^ n8660 ^ n4791 ;
  assign n23692 = n6000 ^ n2135 ^ 1'b0 ;
  assign n23693 = n11533 & n23692 ;
  assign n23694 = n17296 ^ n10353 ^ 1'b0 ;
  assign n23695 = n23693 & ~n23694 ;
  assign n23696 = ~n1603 & n7091 ;
  assign n23697 = n23696 ^ n620 ^ 1'b0 ;
  assign n23698 = n3140 & n23697 ;
  assign n23699 = n12451 & ~n12933 ;
  assign n23700 = n12933 & n23699 ;
  assign n23701 = n16098 | n23700 ;
  assign n23702 = n23700 & ~n23701 ;
  assign n23703 = n16415 & ~n17384 ;
  assign n23704 = n13729 & n23703 ;
  assign n23705 = ( n6487 & n17156 ) | ( n6487 & n23704 ) | ( n17156 & n23704 ) ;
  assign n23706 = n5813 & n7854 ;
  assign n23707 = ( ~n2853 & n19983 ) | ( ~n2853 & n23706 ) | ( n19983 & n23706 ) ;
  assign n23708 = n11943 ^ n6914 ^ 1'b0 ;
  assign n23709 = n2258 & n15849 ;
  assign n23710 = ~n1950 & n3749 ;
  assign n23711 = n1950 & n23710 ;
  assign n23712 = n3124 & ~n23711 ;
  assign n23713 = n23711 & n23712 ;
  assign n23714 = n23481 | n23713 ;
  assign n23715 = n23714 ^ n15608 ^ 1'b0 ;
  assign n23716 = n3505 | n5986 ;
  assign n23717 = n6011 ^ n2813 ^ 1'b0 ;
  assign n23718 = n1956 | n23717 ;
  assign n23719 = n23718 ^ n9732 ^ 1'b0 ;
  assign n23720 = ( ~n5279 & n6297 ) | ( ~n5279 & n16735 ) | ( n6297 & n16735 ) ;
  assign n23721 = ~n1609 & n12221 ;
  assign n23722 = n23721 ^ n16225 ^ 1'b0 ;
  assign n23723 = ( n21568 & n23720 ) | ( n21568 & n23722 ) | ( n23720 & n23722 ) ;
  assign n23724 = n98 & n10483 ;
  assign n23725 = n12289 ^ n10400 ^ 1'b0 ;
  assign n23726 = n893 & ~n23725 ;
  assign n23727 = n18919 ^ n1787 ^ 1'b0 ;
  assign n23728 = n4189 & n22698 ;
  assign n23729 = ~n5135 & n23728 ;
  assign n23730 = n3663 & ~n23729 ;
  assign n23733 = n6128 ^ n4627 ^ n1779 ;
  assign n23731 = n7838 ^ n5634 ^ n46 ;
  assign n23732 = n1493 | n23731 ;
  assign n23734 = n23733 ^ n23732 ^ 1'b0 ;
  assign n23735 = ~n6272 & n23734 ;
  assign n23736 = n4780 ^ n3581 ^ 1'b0 ;
  assign n23737 = n3765 | n8085 ;
  assign n23738 = n8733 & n20563 ;
  assign n23739 = ~n9072 & n11234 ;
  assign n23740 = n23738 & n23739 ;
  assign n23741 = n16168 ^ n6542 ^ 1'b0 ;
  assign n23742 = n14893 | n23741 ;
  assign n23744 = n5745 | n12103 ;
  assign n23743 = n6516 ^ n2846 ^ 1'b0 ;
  assign n23745 = n23744 ^ n23743 ^ 1'b0 ;
  assign n23746 = ~n23742 & n23745 ;
  assign n23747 = n23740 & n23746 ;
  assign n23748 = ( n2248 & ~n23737 ) | ( n2248 & n23747 ) | ( ~n23737 & n23747 ) ;
  assign n23749 = n21431 & ~n23748 ;
  assign n23750 = n23749 ^ n962 ^ 1'b0 ;
  assign n23751 = n9769 & n23750 ;
  assign n23752 = n21873 ^ n19424 ^ 1'b0 ;
  assign n23753 = n4113 | n21429 ;
  assign n23756 = n18863 ^ n4536 ^ 1'b0 ;
  assign n23754 = ~n870 & n21394 ;
  assign n23755 = n23754 ^ n9745 ^ 1'b0 ;
  assign n23757 = n23756 ^ n23755 ^ 1'b0 ;
  assign n23758 = n2249 & n3314 ;
  assign n23759 = n5380 | n23758 ;
  assign n23760 = n9416 ^ n7772 ^ n6762 ;
  assign n23761 = ( n5113 & n15323 ) | ( n5113 & ~n17082 ) | ( n15323 & ~n17082 ) ;
  assign n23762 = ( n2620 & n23760 ) | ( n2620 & ~n23761 ) | ( n23760 & ~n23761 ) ;
  assign n23763 = n23762 ^ n9283 ^ 1'b0 ;
  assign n23764 = n9935 & n19339 ;
  assign n23765 = n23764 ^ n11360 ^ 1'b0 ;
  assign n23766 = n3824 & n11947 ;
  assign n23767 = n23766 ^ n23286 ^ n3614 ;
  assign n23768 = n20571 ^ n18188 ^ 1'b0 ;
  assign n23769 = ~n1662 & n23768 ;
  assign n23770 = n15229 ^ n2633 ^ 1'b0 ;
  assign n23771 = ~n2787 & n23770 ;
  assign n23772 = n7134 & n16286 ;
  assign n23773 = n1437 & n23772 ;
  assign n23774 = n22670 ^ n19401 ^ n2298 ;
  assign n23775 = ( n1081 & n2050 ) | ( n1081 & ~n16728 ) | ( n2050 & ~n16728 ) ;
  assign n23776 = n13623 | n21906 ;
  assign n23777 = n9972 & n23776 ;
  assign n23778 = ~n18985 & n23777 ;
  assign n23779 = n23778 ^ n15675 ^ n1182 ;
  assign n23780 = n102 | n674 ;
  assign n23781 = n4729 ^ n3211 ^ n3207 ;
  assign n23782 = ~n23780 & n23781 ;
  assign n23783 = ~n940 & n23782 ;
  assign n23784 = ~n9765 & n10010 ;
  assign n23785 = ~n732 & n23784 ;
  assign n23787 = n16403 ^ n1832 ^ 1'b0 ;
  assign n23786 = n3198 | n7760 ;
  assign n23788 = n23787 ^ n23786 ^ 1'b0 ;
  assign n23796 = n8964 & n14293 ;
  assign n23797 = n2873 | n23796 ;
  assign n23789 = n6096 & n11608 ;
  assign n23790 = n14530 ^ x1 ^ 1'b0 ;
  assign n23791 = n1461 & n23790 ;
  assign n23792 = n6696 & ~n9149 ;
  assign n23793 = ~n23791 & n23792 ;
  assign n23794 = ( n1851 & n5016 ) | ( n1851 & ~n23793 ) | ( n5016 & ~n23793 ) ;
  assign n23795 = ( n1463 & ~n23789 ) | ( n1463 & n23794 ) | ( ~n23789 & n23794 ) ;
  assign n23798 = n23797 ^ n23795 ^ 1'b0 ;
  assign n23799 = ~n11612 & n22876 ;
  assign n23800 = n4505 & n23799 ;
  assign n23801 = ~n20188 & n21906 ;
  assign n23802 = n23801 ^ n9391 ^ 1'b0 ;
  assign n23803 = n644 | n23802 ;
  assign n23806 = n13422 ^ n403 ^ 1'b0 ;
  assign n23807 = ~n8692 & n23806 ;
  assign n23804 = ( n10962 & n11116 ) | ( n10962 & ~n21613 ) | ( n11116 & ~n21613 ) ;
  assign n23805 = n17825 & ~n23804 ;
  assign n23808 = n23807 ^ n23805 ^ 1'b0 ;
  assign n23809 = n149 & n1744 ;
  assign n23810 = n23809 ^ n12707 ^ 1'b0 ;
  assign n23811 = n23810 ^ n6039 ^ 1'b0 ;
  assign n23812 = n9774 & ~n23811 ;
  assign n23813 = n12571 | n23812 ;
  assign n23814 = n9379 ^ n369 ^ 1'b0 ;
  assign n23815 = n1260 & ~n13643 ;
  assign n23816 = ~n1260 & n23815 ;
  assign n23817 = n23816 ^ n281 ^ 1'b0 ;
  assign n23818 = n23817 ^ n23675 ^ n15978 ;
  assign n23819 = ( n6115 & n12273 ) | ( n6115 & n15085 ) | ( n12273 & n15085 ) ;
  assign n23820 = n9586 & n14319 ;
  assign n23821 = n23820 ^ n3755 ^ 1'b0 ;
  assign n23822 = ~n4298 & n23821 ;
  assign n23823 = n2296 & ~n4333 ;
  assign n23824 = n23823 ^ n6825 ^ 1'b0 ;
  assign n23825 = ~n8141 & n23824 ;
  assign n23826 = n23825 ^ n2586 ^ n1391 ;
  assign n23827 = n11262 ^ n2447 ^ 1'b0 ;
  assign n23828 = n23826 & n23827 ;
  assign n23829 = n2403 | n2836 ;
  assign n23830 = n23829 ^ n16776 ^ 1'b0 ;
  assign n23831 = n1454 & n12124 ;
  assign n23832 = n18252 ^ n7614 ^ 1'b0 ;
  assign n23833 = ( n11269 & n21564 ) | ( n11269 & n23832 ) | ( n21564 & n23832 ) ;
  assign n23835 = n8560 ^ n996 ^ 1'b0 ;
  assign n23836 = n10537 & n23835 ;
  assign n23834 = n15213 & n18716 ;
  assign n23837 = n23836 ^ n23834 ^ 1'b0 ;
  assign n23838 = n6088 & n23564 ;
  assign n23839 = n13478 ^ n6027 ^ 1'b0 ;
  assign n23840 = ~n1933 & n6131 ;
  assign n23841 = n23840 ^ n10685 ^ 1'b0 ;
  assign n23842 = ( ~n1416 & n13218 ) | ( ~n1416 & n23841 ) | ( n13218 & n23841 ) ;
  assign n23843 = n23842 ^ n17787 ^ 1'b0 ;
  assign n23844 = ~n23839 & n23843 ;
  assign n23845 = ~n20826 & n23844 ;
  assign n23846 = n5781 & n13917 ;
  assign n23847 = n21218 ^ n12939 ^ 1'b0 ;
  assign n23848 = n23847 ^ n1558 ^ 1'b0 ;
  assign n23849 = n10963 ^ n7398 ^ 1'b0 ;
  assign n23850 = n16612 & ~n16797 ;
  assign n23851 = n23850 ^ n6424 ^ 1'b0 ;
  assign n23852 = n2697 & ~n3284 ;
  assign n23853 = n21862 ^ n19080 ^ 1'b0 ;
  assign n23854 = ( n7167 & ~n23852 ) | ( n7167 & n23853 ) | ( ~n23852 & n23853 ) ;
  assign n23857 = n5135 ^ n1736 ^ 1'b0 ;
  assign n23858 = n7211 & n23857 ;
  assign n23855 = n4640 & ~n14893 ;
  assign n23856 = n23855 ^ n115 ^ 1'b0 ;
  assign n23859 = n23858 ^ n23856 ^ 1'b0 ;
  assign n23860 = n556 & n1945 ;
  assign n23861 = n23860 ^ n10569 ^ 1'b0 ;
  assign n23862 = n1974 & ~n23861 ;
  assign n23863 = n1868 ^ n78 ^ 1'b0 ;
  assign n23864 = n279 & n23863 ;
  assign n23865 = n14037 & ~n23571 ;
  assign n23866 = ~n23864 & n23865 ;
  assign n23867 = n18511 ^ n517 ^ 1'b0 ;
  assign n23869 = n13825 ^ n3191 ^ 1'b0 ;
  assign n23868 = n630 & n20940 ;
  assign n23870 = n23869 ^ n23868 ^ n12124 ;
  assign n23871 = n340 & n21303 ;
  assign n23872 = n23871 ^ n15037 ^ 1'b0 ;
  assign n23873 = n23872 ^ n10962 ^ 1'b0 ;
  assign n23874 = n8899 ^ n4887 ^ n2547 ;
  assign n23875 = n23874 ^ n18100 ^ n15375 ;
  assign n23876 = n9847 & ~n15065 ;
  assign n23877 = ( n4686 & n9904 ) | ( n4686 & ~n11258 ) | ( n9904 & ~n11258 ) ;
  assign n23878 = n23876 & n23877 ;
  assign n23879 = n23878 ^ n16460 ^ 1'b0 ;
  assign n23880 = n2041 & n13717 ;
  assign n23881 = n23880 ^ n3633 ^ 1'b0 ;
  assign n23882 = n10973 ^ n5029 ^ 1'b0 ;
  assign n23883 = n13962 & ~n23882 ;
  assign n23885 = ( n1397 & n3377 ) | ( n1397 & ~n18619 ) | ( n3377 & ~n18619 ) ;
  assign n23884 = ~n2604 & n5011 ;
  assign n23886 = n23885 ^ n23884 ^ 1'b0 ;
  assign n23887 = n23886 ^ n17656 ^ 1'b0 ;
  assign n23888 = n22318 & ~n23887 ;
  assign n23889 = n22142 ^ n16545 ^ n963 ;
  assign n23890 = ( n6914 & n10314 ) | ( n6914 & n22358 ) | ( n10314 & n22358 ) ;
  assign n23891 = n23890 ^ n15483 ^ 1'b0 ;
  assign n23892 = n2051 & n18981 ;
  assign n23893 = n18126 & n23892 ;
  assign n23894 = n23893 ^ n17347 ^ 1'b0 ;
  assign n23895 = ~n1189 & n9308 ;
  assign n23896 = ( n9645 & n15426 ) | ( n9645 & ~n23176 ) | ( n15426 & ~n23176 ) ;
  assign n23897 = n4290 & n23896 ;
  assign n23899 = ( ~n3962 & n8597 ) | ( ~n3962 & n15868 ) | ( n8597 & n15868 ) ;
  assign n23898 = n4549 | n16409 ;
  assign n23900 = n23899 ^ n23898 ^ 1'b0 ;
  assign n23901 = n6517 & n8672 ;
  assign n23902 = n22008 ^ n1655 ^ 1'b0 ;
  assign n23903 = ( n3599 & ~n5296 ) | ( n3599 & n6775 ) | ( ~n5296 & n6775 ) ;
  assign n23904 = n23903 ^ n17649 ^ 1'b0 ;
  assign n23905 = n12198 ^ n411 ^ 1'b0 ;
  assign n23906 = ~n908 & n17645 ;
  assign n23907 = ~n23905 & n23906 ;
  assign n23908 = ( n792 & n4683 ) | ( n792 & ~n12994 ) | ( n4683 & ~n12994 ) ;
  assign n23909 = n23908 ^ n12785 ^ 1'b0 ;
  assign n23910 = ( n2381 & n15136 ) | ( n2381 & ~n16440 ) | ( n15136 & ~n16440 ) ;
  assign n23911 = n7432 | n23910 ;
  assign n23912 = n2528 & ~n9504 ;
  assign n23913 = n22907 | n23912 ;
  assign n23914 = n15636 ^ n12481 ^ 1'b0 ;
  assign n23915 = n11108 ^ n9645 ^ 1'b0 ;
  assign n23916 = n1011 & n23915 ;
  assign n23917 = n23916 ^ n21886 ^ 1'b0 ;
  assign n23918 = n23917 ^ n12403 ^ 1'b0 ;
  assign n23919 = ( n4467 & ~n10265 ) | ( n4467 & n16485 ) | ( ~n10265 & n16485 ) ;
  assign n23921 = ~n1922 & n12771 ;
  assign n23922 = n23921 ^ n5813 ^ 1'b0 ;
  assign n23920 = ~n9519 & n17769 ;
  assign n23923 = n23922 ^ n23920 ^ n5786 ;
  assign n23924 = ~n3241 & n23923 ;
  assign n23925 = n23924 ^ n14582 ^ 1'b0 ;
  assign n23926 = ( n16981 & ~n23919 ) | ( n16981 & n23925 ) | ( ~n23919 & n23925 ) ;
  assign n23927 = n2130 & n2946 ;
  assign n23928 = n23927 ^ n1444 ^ 1'b0 ;
  assign n23929 = n20772 & n23928 ;
  assign n23930 = n15382 | n18073 ;
  assign n23931 = n17257 & n17993 ;
  assign n23932 = n5709 | n21210 ;
  assign n23933 = n23932 ^ n7418 ^ 1'b0 ;
  assign n23934 = n11680 ^ n4658 ^ 1'b0 ;
  assign n23935 = n18055 & n23934 ;
  assign n23936 = n15251 | n23935 ;
  assign n23937 = n23933 | n23936 ;
  assign n23938 = n2504 & n6324 ;
  assign n23939 = n5091 ^ n45 ^ 1'b0 ;
  assign n23940 = n15897 | n23939 ;
  assign n23948 = n12606 & ~n19091 ;
  assign n23949 = ( ~n4994 & n8245 ) | ( ~n4994 & n23948 ) | ( n8245 & n23948 ) ;
  assign n23941 = ( n4256 & n8720 ) | ( n4256 & ~n11636 ) | ( n8720 & ~n11636 ) ;
  assign n23942 = ( ~n3800 & n4842 ) | ( ~n3800 & n23941 ) | ( n4842 & n23941 ) ;
  assign n23943 = n8130 & ~n9625 ;
  assign n23944 = ( n5397 & n5438 ) | ( n5397 & ~n13952 ) | ( n5438 & ~n13952 ) ;
  assign n23945 = n23943 | n23944 ;
  assign n23946 = n14190 | n23945 ;
  assign n23947 = ~n23942 & n23946 ;
  assign n23950 = n23949 ^ n23947 ^ 1'b0 ;
  assign n23952 = n6625 ^ n1032 ^ 1'b0 ;
  assign n23953 = n11902 & n23952 ;
  assign n23951 = ~n3879 & n13239 ;
  assign n23954 = n23953 ^ n23951 ^ 1'b0 ;
  assign n23955 = n17057 ^ n22 ^ 1'b0 ;
  assign n23956 = n22362 ^ n16341 ^ n14125 ;
  assign n23957 = n963 & n6862 ;
  assign n23958 = ~n4819 & n23957 ;
  assign n23959 = n14872 & n23958 ;
  assign n23960 = n5495 | n21348 ;
  assign n23961 = ( n496 & n12058 ) | ( n496 & n23960 ) | ( n12058 & n23960 ) ;
  assign n23964 = n2901 & ~n3425 ;
  assign n23965 = ~n2510 & n23964 ;
  assign n23962 = n8061 ^ n4259 ^ 1'b0 ;
  assign n23963 = ( n6983 & n23221 ) | ( n6983 & ~n23962 ) | ( n23221 & ~n23962 ) ;
  assign n23966 = n23965 ^ n23963 ^ n7364 ;
  assign n23967 = n2627 & n5020 ;
  assign n23968 = n23967 ^ n19950 ^ n3997 ;
  assign n23969 = n23968 ^ n18412 ^ 1'b0 ;
  assign n23970 = n9362 & n23969 ;
  assign n23971 = ~n5210 & n10177 ;
  assign n23972 = ~n408 & n11400 ;
  assign n23973 = ~n5255 & n23972 ;
  assign n23974 = n23973 ^ n5224 ^ 1'b0 ;
  assign n23975 = n23974 ^ n17260 ^ 1'b0 ;
  assign n23976 = n7796 | n10744 ;
  assign n23977 = n11701 ^ n7492 ^ 1'b0 ;
  assign n23978 = n9868 | n23977 ;
  assign n23979 = n23976 & ~n23978 ;
  assign n23980 = n11823 ^ n8979 ^ n7574 ;
  assign n23981 = n6440 ^ n676 ^ 1'b0 ;
  assign n23982 = n738 & n23981 ;
  assign n23983 = n23980 & n23982 ;
  assign n23984 = n10199 | n23531 ;
  assign n23985 = n2256 | n4647 ;
  assign n23986 = ~n8690 & n23985 ;
  assign n23987 = n6572 & ~n23986 ;
  assign n23988 = ( n13002 & ~n23171 ) | ( n13002 & n23987 ) | ( ~n23171 & n23987 ) ;
  assign n23989 = n18510 ^ n11792 ^ 1'b0 ;
  assign n23990 = ( n5961 & n7807 ) | ( n5961 & n11582 ) | ( n7807 & n11582 ) ;
  assign n23991 = ~n772 & n23392 ;
  assign n23992 = ~n8539 & n23991 ;
  assign n23993 = n7300 ^ n2813 ^ 1'b0 ;
  assign n23994 = ~n23992 & n23993 ;
  assign n23995 = n17258 ^ n13287 ^ 1'b0 ;
  assign n23996 = n14850 & n23995 ;
  assign n23997 = n3187 & n5650 ;
  assign n23998 = n9354 & ~n22307 ;
  assign n23999 = n16777 & ~n23998 ;
  assign n24000 = n15605 & n16633 ;
  assign n24001 = n24000 ^ n12402 ^ n5880 ;
  assign n24002 = n7218 & n24001 ;
  assign n24003 = n24002 ^ n12405 ^ 1'b0 ;
  assign n24004 = n14236 ^ n3456 ^ n3043 ;
  assign n24005 = n18136 ^ n3346 ^ 1'b0 ;
  assign n24006 = ( n4743 & n9027 ) | ( n4743 & n10255 ) | ( n9027 & n10255 ) ;
  assign n24007 = ~n3361 & n24006 ;
  assign n24008 = ~n7860 & n14798 ;
  assign n24009 = n24008 ^ n5554 ^ 1'b0 ;
  assign n24010 = n24009 ^ n2928 ^ n2044 ;
  assign n24011 = n14134 | n15856 ;
  assign n24012 = n1641 & n2745 ;
  assign n24013 = n24012 ^ n16888 ^ 1'b0 ;
  assign n24014 = n6275 ^ n4540 ^ 1'b0 ;
  assign n24015 = n12830 ^ n4004 ^ 1'b0 ;
  assign n24016 = n2566 & n24015 ;
  assign n24017 = n20565 ^ n10294 ^ 1'b0 ;
  assign n24018 = n11204 ^ n7557 ^ 1'b0 ;
  assign n24019 = n24017 & ~n24018 ;
  assign n24020 = n2449 | n4605 ;
  assign n24021 = n10560 & ~n24020 ;
  assign n24022 = ~n3202 & n3454 ;
  assign n24023 = n24022 ^ n15498 ^ 1'b0 ;
  assign n24024 = n14247 & n24023 ;
  assign n24025 = ( ~n14443 & n24021 ) | ( ~n14443 & n24024 ) | ( n24021 & n24024 ) ;
  assign n24026 = n16207 ^ n10396 ^ 1'b0 ;
  assign n24027 = n4086 & n12578 ;
  assign n24028 = n245 & ~n7282 ;
  assign n24029 = ( n11253 & n20344 ) | ( n11253 & n24028 ) | ( n20344 & n24028 ) ;
  assign n24030 = n16264 ^ n10589 ^ n426 ;
  assign n24031 = n9815 & ~n10098 ;
  assign n24032 = n5736 & n24031 ;
  assign n24033 = n3864 ^ n741 ^ 1'b0 ;
  assign n24034 = n3997 & n24033 ;
  assign n24035 = n6882 | n13761 ;
  assign n24037 = n13330 ^ n6868 ^ 1'b0 ;
  assign n24038 = ~n8365 & n24037 ;
  assign n24039 = n5353 ^ n3729 ^ 1'b0 ;
  assign n24040 = n24038 & ~n24039 ;
  assign n24036 = n9910 ^ n9351 ^ 1'b0 ;
  assign n24041 = n24040 ^ n24036 ^ n9324 ;
  assign n24042 = n18771 ^ n6505 ^ 1'b0 ;
  assign n24043 = ~n24041 & n24042 ;
  assign n24044 = n735 & ~n9357 ;
  assign n24045 = n18061 & n24044 ;
  assign n24046 = n9701 & ~n16846 ;
  assign n24047 = n13920 ^ n711 ^ 1'b0 ;
  assign n24048 = n21339 ^ n1364 ^ 1'b0 ;
  assign n24049 = n976 & n24048 ;
  assign n24050 = n4318 & ~n5949 ;
  assign n24051 = n24050 ^ n10543 ^ 1'b0 ;
  assign n24052 = n450 & ~n20735 ;
  assign n24053 = n24052 ^ n11538 ^ 1'b0 ;
  assign n24054 = n11896 ^ n5425 ^ n3825 ;
  assign n24055 = n2505 | n13554 ;
  assign n24058 = n4835 | n23373 ;
  assign n24059 = n12590 & n24058 ;
  assign n24056 = n5797 & n12385 ;
  assign n24057 = n14890 & n24056 ;
  assign n24060 = n24059 ^ n24057 ^ n23215 ;
  assign n24061 = ( n2990 & ~n5073 ) | ( n2990 & n11329 ) | ( ~n5073 & n11329 ) ;
  assign n24062 = n15708 & ~n24061 ;
  assign n24065 = n8838 & ~n11915 ;
  assign n24066 = n17638 | n24065 ;
  assign n24067 = n24066 ^ n9821 ^ 1'b0 ;
  assign n24063 = ( n3912 & ~n5402 ) | ( n3912 & n8540 ) | ( ~n5402 & n8540 ) ;
  assign n24064 = n2541 & n24063 ;
  assign n24068 = n24067 ^ n24064 ^ 1'b0 ;
  assign n24069 = n24068 ^ n5455 ^ n61 ;
  assign n24071 = n7316 ^ n1668 ^ 1'b0 ;
  assign n24070 = n16561 ^ n855 ^ 1'b0 ;
  assign n24072 = n24071 ^ n24070 ^ 1'b0 ;
  assign n24073 = n24072 ^ n12558 ^ 1'b0 ;
  assign n24074 = ~n2727 & n6743 ;
  assign n24075 = ( n276 & n6001 ) | ( n276 & n24074 ) | ( n6001 & n24074 ) ;
  assign n24076 = n15360 ^ n10068 ^ 1'b0 ;
  assign n24077 = n24075 & n24076 ;
  assign n24078 = n18126 ^ n5639 ^ 1'b0 ;
  assign n24079 = n19755 & ~n24078 ;
  assign n24080 = n5106 & n24079 ;
  assign n24081 = n24080 ^ n14813 ^ 1'b0 ;
  assign n24082 = n15274 ^ n7323 ^ 1'b0 ;
  assign n24083 = n1384 ^ n865 ^ 1'b0 ;
  assign n24084 = ~n1859 & n24083 ;
  assign n24085 = n11794 ^ n2306 ^ 1'b0 ;
  assign n24086 = n24084 & ~n24085 ;
  assign n24087 = ( n14789 & n24082 ) | ( n14789 & ~n24086 ) | ( n24082 & ~n24086 ) ;
  assign n24088 = n15289 ^ n9328 ^ 1'b0 ;
  assign n24089 = n2736 & n24088 ;
  assign n24090 = ( n10897 & ~n13951 ) | ( n10897 & n24089 ) | ( ~n13951 & n24089 ) ;
  assign n24091 = n3460 ^ n1490 ^ 1'b0 ;
  assign n24092 = n3639 & ~n24091 ;
  assign n24093 = n3709 | n6987 ;
  assign n24094 = n24092 & ~n24093 ;
  assign n24095 = n24094 ^ n2102 ^ 1'b0 ;
  assign n24096 = n2030 | n18616 ;
  assign n24097 = n1177 & ~n12393 ;
  assign n24098 = n21294 ^ n19200 ^ 1'b0 ;
  assign n24099 = n24097 & n24098 ;
  assign n24100 = n73 | n22367 ;
  assign n24101 = n21387 ^ n4829 ^ 1'b0 ;
  assign n24102 = n9355 | n13449 ;
  assign n24103 = n24102 ^ n4576 ^ 1'b0 ;
  assign n24104 = ~n24101 & n24103 ;
  assign n24105 = ~n5800 & n14864 ;
  assign n24106 = n24105 ^ n362 ^ 1'b0 ;
  assign n24107 = n2823 & ~n13376 ;
  assign n24108 = n24107 ^ n4461 ^ 1'b0 ;
  assign n24109 = ~n14702 & n24108 ;
  assign n24115 = ~n2355 & n15009 ;
  assign n24110 = n8195 | n22101 ;
  assign n24111 = ( ~n4689 & n8630 ) | ( ~n4689 & n9946 ) | ( n8630 & n9946 ) ;
  assign n24112 = n24111 ^ n9599 ^ 1'b0 ;
  assign n24113 = n24110 | n24112 ;
  assign n24114 = n24113 ^ n3364 ^ 1'b0 ;
  assign n24116 = n24115 ^ n24114 ^ 1'b0 ;
  assign n24117 = n24116 ^ n13514 ^ 1'b0 ;
  assign n24118 = n7631 ^ n940 ^ 1'b0 ;
  assign n24119 = n24118 ^ n5417 ^ 1'b0 ;
  assign n24120 = n2170 ^ n283 ^ 1'b0 ;
  assign n24121 = n2503 | n24120 ;
  assign n24122 = n15472 ^ n3337 ^ 1'b0 ;
  assign n24123 = n7134 & ~n24122 ;
  assign n24124 = n24121 & n24123 ;
  assign n24125 = n9896 | n24124 ;
  assign n24126 = n24125 ^ n6147 ^ 1'b0 ;
  assign n24127 = n13740 ^ n119 ^ 1'b0 ;
  assign n24128 = ~n22210 & n24127 ;
  assign n24129 = n22893 ^ n6030 ^ 1'b0 ;
  assign n24130 = n296 | n24129 ;
  assign n24131 = n2849 | n4058 ;
  assign n24132 = n24131 ^ n11692 ^ 1'b0 ;
  assign n24133 = n9698 & n24132 ;
  assign n24134 = n24133 ^ n15898 ^ n7532 ;
  assign n24135 = n3007 ^ n1381 ^ 1'b0 ;
  assign n24136 = n24135 ^ n21038 ^ 1'b0 ;
  assign n24137 = n1069 & ~n17993 ;
  assign n24138 = n24137 ^ n9397 ^ 1'b0 ;
  assign n24139 = n15344 ^ n7545 ^ 1'b0 ;
  assign n24140 = n24138 & ~n24139 ;
  assign n24141 = n13379 ^ n9023 ^ 1'b0 ;
  assign n24142 = n6737 | n24141 ;
  assign n24143 = n3271 & ~n24142 ;
  assign n24144 = n24140 & ~n24143 ;
  assign n24145 = n24144 ^ n21409 ^ 1'b0 ;
  assign n24146 = n1982 | n22608 ;
  assign n24147 = n24146 ^ n886 ^ 1'b0 ;
  assign n24148 = n13467 | n21005 ;
  assign n24149 = n24148 ^ n21031 ^ 1'b0 ;
  assign n24150 = n99 & n9453 ;
  assign n24151 = n24149 & n24150 ;
  assign n24152 = n23756 ^ n12286 ^ n5310 ;
  assign n24153 = n3650 & ~n24152 ;
  assign n24160 = n16228 | n18770 ;
  assign n24161 = n3628 | n24160 ;
  assign n24162 = n24161 ^ n11599 ^ n1184 ;
  assign n24154 = n2280 & n2571 ;
  assign n24155 = n24154 ^ n209 ^ 1'b0 ;
  assign n24156 = n24155 ^ n1335 ^ 1'b0 ;
  assign n24157 = ~n10296 & n24156 ;
  assign n24158 = n24157 ^ n18478 ^ 1'b0 ;
  assign n24159 = n4319 & ~n24158 ;
  assign n24163 = n24162 ^ n24159 ^ 1'b0 ;
  assign n24165 = n4536 ^ n2645 ^ n2100 ;
  assign n24164 = n12402 ^ n1621 ^ 1'b0 ;
  assign n24166 = n24165 ^ n24164 ^ 1'b0 ;
  assign n24167 = n8176 & n24166 ;
  assign n24168 = n24167 ^ n5783 ^ 1'b0 ;
  assign n24169 = ( n581 & ~n2287 ) | ( n581 & n19658 ) | ( ~n2287 & n19658 ) ;
  assign n24170 = n7146 | n24169 ;
  assign n24171 = n24170 ^ n5352 ^ 1'b0 ;
  assign n24172 = ~n10926 & n14838 ;
  assign n24173 = ( n43 & ~n7065 ) | ( n43 & n9899 ) | ( ~n7065 & n9899 ) ;
  assign n24174 = n2857 | n4230 ;
  assign n24175 = n40 | n24174 ;
  assign n24176 = n24175 ^ n7323 ^ 1'b0 ;
  assign n24177 = n24173 & n24176 ;
  assign n24178 = ~n3386 & n4440 ;
  assign n24179 = ~n24177 & n24178 ;
  assign n24180 = n24172 & ~n24179 ;
  assign n24181 = n19047 ^ n8595 ^ n8037 ;
  assign n24182 = ~n10872 & n24181 ;
  assign n24183 = n11570 ^ n837 ^ 1'b0 ;
  assign n24184 = ~n20378 & n24183 ;
  assign n24185 = n24184 ^ n17325 ^ 1'b0 ;
  assign n24186 = ( ~n8523 & n13784 ) | ( ~n8523 & n16116 ) | ( n13784 & n16116 ) ;
  assign n24187 = n11603 ^ n3467 ^ n147 ;
  assign n24188 = n10682 & n24187 ;
  assign n24189 = n440 & n24188 ;
  assign n24190 = n24189 ^ n3628 ^ n3548 ;
  assign n24191 = n22161 ^ n17930 ^ 1'b0 ;
  assign n24192 = n24191 ^ n9452 ^ 1'b0 ;
  assign n24193 = n8242 ^ n1052 ^ n604 ;
  assign n24194 = n2089 | n24193 ;
  assign n24195 = ~n6636 & n10874 ;
  assign n24196 = ~n24194 & n24195 ;
  assign n24197 = n24196 ^ n6729 ^ 1'b0 ;
  assign n24198 = ~n801 & n5990 ;
  assign n24199 = n24198 ^ n177 ^ 1'b0 ;
  assign n24200 = n8577 | n11137 ;
  assign n24201 = n7601 & ~n9857 ;
  assign n24202 = ~n24200 & n24201 ;
  assign n24203 = n24202 ^ n574 ^ 1'b0 ;
  assign n24204 = n16963 | n24203 ;
  assign n24205 = n17359 ^ n12073 ^ n7330 ;
  assign n24206 = n24205 ^ n11097 ^ n7286 ;
  assign n24207 = ( n17399 & ~n17715 ) | ( n17399 & n24206 ) | ( ~n17715 & n24206 ) ;
  assign n24208 = n1558 & ~n20870 ;
  assign n24209 = n24208 ^ n1878 ^ 1'b0 ;
  assign n24210 = n24209 ^ n7954 ^ 1'b0 ;
  assign n24211 = n24210 ^ n14164 ^ 1'b0 ;
  assign n24212 = n1172 | n24211 ;
  assign n24217 = ~n3542 & n6743 ;
  assign n24214 = n2907 ^ n1503 ^ 1'b0 ;
  assign n24215 = n2345 & ~n24214 ;
  assign n24216 = n24215 ^ n4249 ^ 1'b0 ;
  assign n24218 = n24217 ^ n24216 ^ 1'b0 ;
  assign n24213 = ~n10189 & n23628 ;
  assign n24219 = n24218 ^ n24213 ^ 1'b0 ;
  assign n24220 = n10078 ^ n3161 ^ 1'b0 ;
  assign n24221 = n18126 ^ n833 ^ 1'b0 ;
  assign n24222 = n12493 & n24221 ;
  assign n24223 = n24222 ^ n4260 ^ 1'b0 ;
  assign n24224 = ~n24220 & n24223 ;
  assign n24228 = n1825 & ~n6366 ;
  assign n24229 = ~n20129 & n24228 ;
  assign n24225 = n9699 ^ n4216 ^ 1'b0 ;
  assign n24226 = n5706 & ~n24225 ;
  assign n24227 = n510 & ~n24226 ;
  assign n24230 = n24229 ^ n24227 ^ n20885 ;
  assign n24231 = n18389 ^ n3309 ^ 1'b0 ;
  assign n24232 = n4688 | n24231 ;
  assign n24233 = n24232 ^ n20245 ^ n2556 ;
  assign n24234 = n5877 & n19579 ;
  assign n24235 = n4976 ^ n3159 ^ 1'b0 ;
  assign n24236 = n24235 ^ n19580 ^ n8792 ;
  assign n24237 = n24236 ^ n15505 ^ n8014 ;
  assign n24238 = n24237 ^ n23298 ^ 1'b0 ;
  assign n24239 = n24234 & n24238 ;
  assign n24240 = n21190 ^ n2606 ^ 1'b0 ;
  assign n24241 = n2338 & ~n24240 ;
  assign n24242 = ~n6614 & n24241 ;
  assign n24243 = ( n134 & n6871 ) | ( n134 & ~n17505 ) | ( n6871 & ~n17505 ) ;
  assign n24244 = n23994 | n24243 ;
  assign n24245 = n15807 ^ n13513 ^ 1'b0 ;
  assign n24246 = n3586 & n24245 ;
  assign n24247 = n24246 ^ n1068 ^ n937 ;
  assign n24248 = n1940 & ~n18055 ;
  assign n24249 = n24248 ^ n9260 ^ 1'b0 ;
  assign n24250 = n1813 & n1990 ;
  assign n24251 = n2563 & n24250 ;
  assign n24252 = n24251 ^ n12225 ^ n11792 ;
  assign n24253 = n24252 ^ n15228 ^ 1'b0 ;
  assign n24254 = ~n24249 & n24253 ;
  assign n24255 = n10506 & n14280 ;
  assign n24256 = n9971 ^ n4638 ^ n1773 ;
  assign n24257 = n8595 ^ n7254 ^ 1'b0 ;
  assign n24258 = n22256 & ~n24257 ;
  assign n24259 = n24256 | n24258 ;
  assign n24260 = n24259 ^ n12765 ^ 1'b0 ;
  assign n24261 = n19946 ^ n19562 ^ n19210 ;
  assign n24262 = ( n2718 & n7270 ) | ( n2718 & n9138 ) | ( n7270 & n9138 ) ;
  assign n24263 = n4085 & ~n4120 ;
  assign n24264 = n24263 ^ n711 ^ 1'b0 ;
  assign n24265 = ( n17406 & n24262 ) | ( n17406 & ~n24264 ) | ( n24262 & ~n24264 ) ;
  assign n24266 = n5729 & n5778 ;
  assign n24267 = ~n2029 & n24266 ;
  assign n24268 = n10450 ^ n4629 ^ n2946 ;
  assign n24269 = n3932 & ~n24268 ;
  assign n24270 = n24269 ^ n8740 ^ 1'b0 ;
  assign n24271 = n24270 ^ n19399 ^ 1'b0 ;
  assign n24272 = n24271 ^ n19893 ^ 1'b0 ;
  assign n24273 = n24011 ^ n4004 ^ 1'b0 ;
  assign n24274 = n5968 & ~n17554 ;
  assign n24275 = n12194 ^ n7041 ^ n5249 ;
  assign n24278 = n2510 & ~n10674 ;
  assign n24276 = n4889 | n12115 ;
  assign n24277 = n18692 | n24276 ;
  assign n24279 = n24278 ^ n24277 ^ 1'b0 ;
  assign n24280 = n20401 & n24279 ;
  assign n24281 = ( n22527 & n24275 ) | ( n22527 & ~n24280 ) | ( n24275 & ~n24280 ) ;
  assign n24282 = n22722 ^ n13795 ^ n3730 ;
  assign n24283 = n619 & n24282 ;
  assign n24284 = n3277 ^ n455 ^ 1'b0 ;
  assign n24285 = ~n5796 & n24284 ;
  assign n24286 = n24285 ^ n8736 ^ 1'b0 ;
  assign n24287 = n614 & n20070 ;
  assign n24288 = n20368 ^ n14016 ^ n9006 ;
  assign n24289 = n24288 ^ n4721 ^ 1'b0 ;
  assign n24290 = n13157 ^ n11307 ^ n4570 ;
  assign n24291 = n2821 | n24290 ;
  assign n24292 = n5699 & ~n23962 ;
  assign n24293 = ~n797 & n8236 ;
  assign n24294 = n24293 ^ n23656 ^ 1'b0 ;
  assign n24295 = n6924 & ~n7099 ;
  assign n24296 = n24295 ^ n801 ^ 1'b0 ;
  assign n24297 = n24296 ^ n22464 ^ 1'b0 ;
  assign n24298 = n24294 & n24297 ;
  assign n24299 = n3819 & ~n14064 ;
  assign n24300 = n24299 ^ n17138 ^ 1'b0 ;
  assign n24301 = n1233 | n24300 ;
  assign n24302 = n24301 ^ n15276 ^ 1'b0 ;
  assign n24303 = n24302 ^ n21593 ^ 1'b0 ;
  assign n24304 = n4679 & n24303 ;
  assign n24305 = n63 & ~n1040 ;
  assign n24306 = n6535 | n24305 ;
  assign n24307 = n24306 ^ n5440 ^ 1'b0 ;
  assign n24308 = n24307 ^ n4976 ^ 1'b0 ;
  assign n24309 = n24308 ^ n12750 ^ 1'b0 ;
  assign n24310 = ~n9740 & n24309 ;
  assign n24311 = ( n6122 & n12540 ) | ( n6122 & ~n20177 ) | ( n12540 & ~n20177 ) ;
  assign n24312 = ( n10660 & n24310 ) | ( n10660 & ~n24311 ) | ( n24310 & ~n24311 ) ;
  assign n24313 = n17235 ^ n4805 ^ 1'b0 ;
  assign n24314 = ~n5209 & n24313 ;
  assign n24315 = n8187 & n24314 ;
  assign n24316 = n24315 ^ n23406 ^ 1'b0 ;
  assign n24317 = n19858 ^ n6382 ^ 1'b0 ;
  assign n24318 = n5861 & ~n24317 ;
  assign n24319 = ( n11470 & n18075 ) | ( n11470 & n20120 ) | ( n18075 & n20120 ) ;
  assign n24320 = ~n16303 & n24319 ;
  assign n24321 = n4536 & ~n24320 ;
  assign n24323 = ~n1628 & n6576 ;
  assign n24322 = n6251 ^ n3644 ^ 1'b0 ;
  assign n24324 = n24323 ^ n24322 ^ n14765 ;
  assign n24327 = ~n657 & n2946 ;
  assign n24325 = n2221 & n12856 ;
  assign n24326 = n10180 & n24325 ;
  assign n24328 = n24327 ^ n24326 ^ n3214 ;
  assign n24329 = ~n4660 & n7559 ;
  assign n24330 = n13113 | n24329 ;
  assign n24331 = n5217 | n9732 ;
  assign n24332 = n24331 ^ n18473 ^ 1'b0 ;
  assign n24333 = n24332 ^ n3264 ^ 1'b0 ;
  assign n24334 = n17450 & ~n24333 ;
  assign n24338 = ~n5127 & n13438 ;
  assign n24339 = n24338 ^ n3348 ^ 1'b0 ;
  assign n24335 = n4728 | n9737 ;
  assign n24336 = n24335 ^ n8534 ^ 1'b0 ;
  assign n24337 = n1681 | n24336 ;
  assign n24340 = n24339 ^ n24337 ^ n11635 ;
  assign n24341 = n11464 ^ n4290 ^ 1'b0 ;
  assign n24342 = n10769 | n24341 ;
  assign n24343 = n8502 | n24342 ;
  assign n24344 = n11944 & n14757 ;
  assign n24345 = ( n19210 & n20819 ) | ( n19210 & n24344 ) | ( n20819 & n24344 ) ;
  assign n24346 = n2937 & ~n21257 ;
  assign n24347 = n5699 | n8373 ;
  assign n24350 = n17751 | n20885 ;
  assign n24348 = n5053 | n9541 ;
  assign n24349 = n5589 & n24348 ;
  assign n24351 = n24350 ^ n24349 ^ 1'b0 ;
  assign n24352 = n4475 & ~n13090 ;
  assign n24353 = ~n15350 & n24352 ;
  assign n24354 = ( n9889 & n18499 ) | ( n9889 & n19191 ) | ( n18499 & n19191 ) ;
  assign n24355 = n24354 ^ n20319 ^ n1951 ;
  assign n24356 = ~n9072 & n19966 ;
  assign n24357 = n455 & ~n24356 ;
  assign n24358 = ( n2986 & n23882 ) | ( n2986 & n24357 ) | ( n23882 & n24357 ) ;
  assign n24359 = n12794 ^ n4861 ^ 1'b0 ;
  assign n24360 = n6261 ^ n3175 ^ 1'b0 ;
  assign n24361 = n8996 & ~n15826 ;
  assign n24362 = ~n6205 & n24361 ;
  assign n24363 = n24362 ^ n18528 ^ 1'b0 ;
  assign n24364 = n5796 | n24363 ;
  assign n24365 = n23406 ^ n17463 ^ n10652 ;
  assign n24366 = n8359 | n24365 ;
  assign n24367 = n42 | n2441 ;
  assign n24368 = n9929 ^ n566 ^ 1'b0 ;
  assign n24369 = n24368 ^ n10628 ^ 1'b0 ;
  assign n24370 = n23675 | n24369 ;
  assign n24371 = n14172 & n20919 ;
  assign n24372 = ~n4262 & n24371 ;
  assign n24373 = n9573 & n18928 ;
  assign n24374 = n17971 | n24373 ;
  assign n24375 = n13393 ^ n1097 ^ 1'b0 ;
  assign n24376 = ( ~n1826 & n24049 ) | ( ~n1826 & n24375 ) | ( n24049 & n24375 ) ;
  assign n24377 = n20681 ^ n12393 ^ 1'b0 ;
  assign n24378 = n7319 & ~n24377 ;
  assign n24379 = n15657 ^ n15432 ^ 1'b0 ;
  assign n24380 = n776 | n24379 ;
  assign n24381 = n2922 & ~n4750 ;
  assign n24382 = n24380 & n24381 ;
  assign n24383 = ( ~n125 & n6375 ) | ( ~n125 & n10124 ) | ( n6375 & n10124 ) ;
  assign n24384 = ~n19566 & n24383 ;
  assign n24385 = n15011 ^ n491 ^ 1'b0 ;
  assign n24386 = n16637 ^ n12477 ^ 1'b0 ;
  assign n24387 = n24386 ^ n22739 ^ 1'b0 ;
  assign n24388 = n5404 & n24387 ;
  assign n24389 = ( n6153 & n12901 ) | ( n6153 & ~n14612 ) | ( n12901 & ~n14612 ) ;
  assign n24390 = n4226 | n5725 ;
  assign n24391 = n24390 ^ n20535 ^ 1'b0 ;
  assign n24392 = ( n11080 & n23791 ) | ( n11080 & ~n24391 ) | ( n23791 & ~n24391 ) ;
  assign n24396 = n8584 ^ n6485 ^ 1'b0 ;
  assign n24397 = n5464 ^ n4373 ^ 1'b0 ;
  assign n24398 = n24397 ^ n922 ^ 1'b0 ;
  assign n24399 = n24396 & n24398 ;
  assign n24394 = n13078 ^ n9618 ^ n1515 ;
  assign n24393 = n3981 & ~n8147 ;
  assign n24395 = n24394 ^ n24393 ^ 1'b0 ;
  assign n24400 = n24399 ^ n24395 ^ 1'b0 ;
  assign n24401 = n32 & ~n12753 ;
  assign n24402 = n24401 ^ n4949 ^ 1'b0 ;
  assign n24403 = n4539 & ~n11113 ;
  assign n24404 = n24403 ^ n8912 ^ 1'b0 ;
  assign n24405 = n16672 ^ n12956 ^ 1'b0 ;
  assign n24406 = ( n4462 & n18620 ) | ( n4462 & n24405 ) | ( n18620 & n24405 ) ;
  assign n24407 = n20274 & n23998 ;
  assign n24408 = n12589 ^ n4388 ^ 1'b0 ;
  assign n24409 = n4189 | n24118 ;
  assign n24410 = n24408 | n24409 ;
  assign n24411 = n1904 & ~n18294 ;
  assign n24412 = n2650 | n24394 ;
  assign n24413 = n11462 | n13504 ;
  assign n24414 = n925 | n24413 ;
  assign n24415 = ( ~n24411 & n24412 ) | ( ~n24411 & n24414 ) | ( n24412 & n24414 ) ;
  assign n24418 = n7307 ^ n3329 ^ 1'b0 ;
  assign n24416 = n554 & ~n11568 ;
  assign n24417 = n24416 ^ n20369 ^ 1'b0 ;
  assign n24419 = n24418 ^ n24417 ^ 1'b0 ;
  assign n24420 = n20734 ^ n7823 ^ 1'b0 ;
  assign n24421 = n3059 | n24420 ;
  assign n24422 = n24421 ^ n8165 ^ 1'b0 ;
  assign n24423 = n3156 & ~n24422 ;
  assign n24424 = n24423 ^ n24333 ^ n18581 ;
  assign n24425 = n17122 & ~n21982 ;
  assign n24426 = n4199 | n9012 ;
  assign n24427 = n11578 | n24426 ;
  assign n24428 = n697 & n9146 ;
  assign n24429 = n24428 ^ n774 ^ 1'b0 ;
  assign n24430 = ( n7588 & ~n10079 ) | ( n7588 & n24429 ) | ( ~n10079 & n24429 ) ;
  assign n24431 = n2395 ^ n97 ^ 1'b0 ;
  assign n24432 = n19005 | n24431 ;
  assign n24433 = n10001 | n14333 ;
  assign n24434 = n12821 | n24433 ;
  assign n24435 = ~n24432 & n24434 ;
  assign n24436 = n20438 & n24435 ;
  assign n24437 = n4805 & n6455 ;
  assign n24438 = ~n2597 & n24437 ;
  assign n24439 = n11938 | n24438 ;
  assign n24440 = n2846 ^ n1460 ^ 1'b0 ;
  assign n24441 = ~n6895 & n24440 ;
  assign n24442 = ~n9079 & n24441 ;
  assign n24443 = n4352 ^ x3 ^ 1'b0 ;
  assign n24444 = n24443 ^ n9664 ^ n6533 ;
  assign n24445 = n7038 | n12456 ;
  assign n24446 = n16770 & ~n24445 ;
  assign n24447 = n4803 & ~n5769 ;
  assign n24448 = n24447 ^ n14533 ^ n556 ;
  assign n24449 = n8457 & ~n22837 ;
  assign n24450 = ~n22007 & n24449 ;
  assign n24451 = n23839 ^ n20689 ^ n1848 ;
  assign n24452 = n4992 ^ n876 ^ 1'b0 ;
  assign n24453 = ( ~n2603 & n3833 ) | ( ~n2603 & n24452 ) | ( n3833 & n24452 ) ;
  assign n24454 = n242 | n7784 ;
  assign n24455 = n194 & ~n4028 ;
  assign n24456 = n8351 & n24455 ;
  assign n24457 = n24456 ^ n6225 ^ 1'b0 ;
  assign n24458 = n4547 ^ n2427 ^ 1'b0 ;
  assign n24459 = n10794 & n13169 ;
  assign n24460 = ~n24458 & n24459 ;
  assign n24462 = n8372 ^ n3624 ^ 1'b0 ;
  assign n24461 = n8420 | n10178 ;
  assign n24463 = n24462 ^ n24461 ^ 1'b0 ;
  assign n24464 = n2701 | n24463 ;
  assign n24465 = n24464 ^ n19459 ^ 1'b0 ;
  assign n24466 = n17959 | n24465 ;
  assign n24467 = n24466 ^ n16539 ^ 1'b0 ;
  assign n24468 = n9553 ^ n2795 ^ 1'b0 ;
  assign n24469 = n5072 & n14427 ;
  assign n24470 = ~n24468 & n24469 ;
  assign n24471 = n21948 ^ n2277 ^ 1'b0 ;
  assign n24472 = n18948 | n24471 ;
  assign n24473 = n6150 & n24472 ;
  assign n24480 = n10799 ^ n709 ^ 1'b0 ;
  assign n24481 = ~n18239 & n24480 ;
  assign n24482 = n24481 ^ n18742 ^ 1'b0 ;
  assign n24474 = ( n2906 & n5044 ) | ( n2906 & ~n11429 ) | ( n5044 & ~n11429 ) ;
  assign n24475 = n3111 & n10917 ;
  assign n24476 = ~n14385 & n18290 ;
  assign n24477 = n24476 ^ n1290 ^ 1'b0 ;
  assign n24478 = ( ~n21820 & n24475 ) | ( ~n21820 & n24477 ) | ( n24475 & n24477 ) ;
  assign n24479 = ~n24474 & n24478 ;
  assign n24483 = n24482 ^ n24479 ^ 1'b0 ;
  assign n24484 = n4993 ^ n459 ^ 1'b0 ;
  assign n24485 = n11264 ^ n3473 ^ 1'b0 ;
  assign n24486 = n24485 ^ n5004 ^ 1'b0 ;
  assign n24487 = ~n3445 & n24486 ;
  assign n24488 = n23832 & n24487 ;
  assign n24489 = n18076 ^ n11988 ^ 1'b0 ;
  assign n24490 = n9981 ^ n4880 ^ 1'b0 ;
  assign n24492 = n14535 ^ n2044 ^ 1'b0 ;
  assign n24493 = ~n9991 & n24492 ;
  assign n24491 = n7207 | n7541 ;
  assign n24494 = n24493 ^ n24491 ^ 1'b0 ;
  assign n24495 = n10435 ^ n2719 ^ n1517 ;
  assign n24496 = n20535 ^ n5868 ^ 1'b0 ;
  assign n24497 = n12751 & ~n24496 ;
  assign n24498 = ~n2282 & n24497 ;
  assign n24499 = ~n16990 & n17556 ;
  assign n24500 = n15838 & n24499 ;
  assign n24501 = n24500 ^ n15516 ^ 1'b0 ;
  assign n24502 = n7626 ^ n1436 ^ 1'b0 ;
  assign n24503 = n9706 & ~n24502 ;
  assign n24504 = n19015 & n24503 ;
  assign n24505 = n18448 ^ n7011 ^ 1'b0 ;
  assign n24506 = n24505 ^ n6099 ^ 1'b0 ;
  assign n24507 = n993 & n24506 ;
  assign n24508 = n4969 & ~n12387 ;
  assign n24509 = n24508 ^ n2896 ^ 1'b0 ;
  assign n24510 = n10007 & n15776 ;
  assign n24511 = n11218 ^ n3413 ^ 1'b0 ;
  assign n24512 = ~n5053 & n13366 ;
  assign n24513 = n23646 ^ n4673 ^ n2828 ;
  assign n24514 = n1021 | n7807 ;
  assign n24515 = n24513 & ~n24514 ;
  assign n24516 = n14641 & ~n23426 ;
  assign n24517 = n3709 ^ n2535 ^ 1'b0 ;
  assign n24519 = ( ~n4723 & n13866 ) | ( ~n4723 & n18236 ) | ( n13866 & n18236 ) ;
  assign n24518 = ~n3680 & n4394 ;
  assign n24520 = n24519 ^ n24518 ^ n13444 ;
  assign n24521 = n17802 ^ n15026 ^ 1'b0 ;
  assign n24522 = ~n8697 & n24521 ;
  assign n24523 = ( ~n2100 & n5622 ) | ( ~n2100 & n13473 ) | ( n5622 & n13473 ) ;
  assign n24524 = ~n51 & n9169 ;
  assign n24525 = ~n24523 & n24524 ;
  assign n24526 = n11771 ^ n1836 ^ 1'b0 ;
  assign n24527 = n7870 & n24526 ;
  assign n24528 = n24527 ^ n2808 ^ 1'b0 ;
  assign n24529 = n24525 | n24528 ;
  assign n24530 = n24529 ^ n354 ^ 1'b0 ;
  assign n24531 = n1069 ^ n592 ^ n293 ;
  assign n24532 = n24531 ^ n4574 ^ n829 ;
  assign n24533 = n24532 ^ n24380 ^ 1'b0 ;
  assign n24534 = n21839 & ~n24533 ;
  assign n24535 = n5251 & n6155 ;
  assign n24536 = ~n1960 & n2990 ;
  assign n24537 = n1001 & n24536 ;
  assign n24538 = n3655 | n24537 ;
  assign n24539 = n9709 ^ n4663 ^ 1'b0 ;
  assign n24540 = n6549 & ~n24539 ;
  assign n24541 = n9919 & n24540 ;
  assign n24545 = ~n3663 & n13072 ;
  assign n24542 = n17303 ^ n6030 ^ 1'b0 ;
  assign n24543 = ~n13889 & n24542 ;
  assign n24544 = n12868 & n24543 ;
  assign n24546 = n24545 ^ n24544 ^ 1'b0 ;
  assign n24547 = n442 & ~n3568 ;
  assign n24548 = n1540 & ~n24547 ;
  assign n24549 = n24548 ^ n3868 ^ 1'b0 ;
  assign n24550 = n5944 & n16965 ;
  assign n24551 = n24550 ^ n448 ^ 1'b0 ;
  assign n24554 = n1262 & ~n12068 ;
  assign n24555 = ~n4342 & n24554 ;
  assign n24552 = n3508 & n12874 ;
  assign n24553 = n24552 ^ n2230 ^ 1'b0 ;
  assign n24556 = n24555 ^ n24553 ^ 1'b0 ;
  assign n24557 = ~n2577 & n15972 ;
  assign n24558 = n3241 ^ n2350 ^ 1'b0 ;
  assign n24559 = n710 & n24558 ;
  assign n24560 = n24559 ^ n5494 ^ 1'b0 ;
  assign n24561 = n20991 ^ n9084 ^ 1'b0 ;
  assign n24562 = n5068 ^ n2841 ^ 1'b0 ;
  assign n24563 = n24562 ^ n12491 ^ n6874 ;
  assign n24564 = n22003 ^ n16561 ^ 1'b0 ;
  assign n24565 = n13237 & ~n24564 ;
  assign n24566 = n9566 ^ n2879 ^ 1'b0 ;
  assign n24567 = n20172 & n24566 ;
  assign n24568 = ( n621 & ~n24565 ) | ( n621 & n24567 ) | ( ~n24565 & n24567 ) ;
  assign n24573 = ( n928 & n8060 ) | ( n928 & n8188 ) | ( n8060 & n8188 ) ;
  assign n24574 = n24573 ^ n923 ^ 1'b0 ;
  assign n24575 = ~n14125 & n24574 ;
  assign n24569 = n10915 ^ n1260 ^ 1'b0 ;
  assign n24570 = n24569 ^ n13526 ^ 1'b0 ;
  assign n24571 = n8740 & ~n24570 ;
  assign n24572 = ~n13139 & n24571 ;
  assign n24576 = n24575 ^ n24572 ^ 1'b0 ;
  assign n24577 = ( n2946 & ~n11829 ) | ( n2946 & n12321 ) | ( ~n11829 & n12321 ) ;
  assign n24578 = n5108 & ~n13819 ;
  assign n24579 = ~n20136 & n24578 ;
  assign n24580 = n13001 ^ n8265 ^ 1'b0 ;
  assign n24581 = n5740 ^ n3271 ^ 1'b0 ;
  assign n24582 = ~n24580 & n24581 ;
  assign n24583 = n15672 & n24582 ;
  assign n24584 = n24583 ^ n4297 ^ 1'b0 ;
  assign n24585 = n24579 | n24584 ;
  assign n24586 = n24585 ^ n12617 ^ 1'b0 ;
  assign n24587 = n24577 & ~n24586 ;
  assign n24588 = n11045 ^ n3636 ^ 1'b0 ;
  assign n24589 = n10391 | n24588 ;
  assign n24590 = n17168 ^ n3450 ^ 1'b0 ;
  assign n24591 = n22130 & n24590 ;
  assign n24592 = n9265 & ~n17637 ;
  assign n24593 = n2602 & n24592 ;
  assign n24594 = ~n8818 & n16594 ;
  assign n24595 = n24594 ^ n9246 ^ 1'b0 ;
  assign n24596 = n14179 ^ n2216 ^ 1'b0 ;
  assign n24597 = n18902 & ~n24596 ;
  assign n24598 = n12854 & n24597 ;
  assign n24599 = n7386 & ~n13632 ;
  assign n24600 = n14066 & n14119 ;
  assign n24601 = ( n1062 & n9795 ) | ( n1062 & n12468 ) | ( n9795 & n12468 ) ;
  assign n24602 = ( n4807 & n13804 ) | ( n4807 & ~n24601 ) | ( n13804 & ~n24601 ) ;
  assign n24603 = n24602 ^ n5815 ^ 1'b0 ;
  assign n24604 = ~n2418 & n24603 ;
  assign n24605 = n65 | n448 ;
  assign n24606 = n2050 ^ n1650 ^ 1'b0 ;
  assign n24607 = ~n13703 & n24606 ;
  assign n24608 = ~n13342 & n24607 ;
  assign n24609 = n24605 & n24608 ;
  assign n24610 = n15516 | n24609 ;
  assign n24611 = ( n5210 & n11100 ) | ( n5210 & ~n24610 ) | ( n11100 & ~n24610 ) ;
  assign n24612 = n12512 ^ n7000 ^ 1'b0 ;
  assign n24613 = ~n637 & n24612 ;
  assign n24614 = n24613 ^ n8470 ^ 1'b0 ;
  assign n24615 = ( n14350 & ~n19654 ) | ( n14350 & n24614 ) | ( ~n19654 & n24614 ) ;
  assign n24616 = n10453 ^ n4736 ^ 1'b0 ;
  assign n24617 = n16352 | n24616 ;
  assign n24618 = n3253 | n24617 ;
  assign n24619 = n11867 & n20509 ;
  assign n24620 = n16290 ^ n14849 ^ 1'b0 ;
  assign n24621 = n6374 & n24620 ;
  assign n24622 = n9805 ^ n5552 ^ 1'b0 ;
  assign n24623 = n24622 ^ n8378 ^ 1'b0 ;
  assign n24624 = n11359 ^ n8874 ^ 1'b0 ;
  assign n24625 = n24624 ^ n22453 ^ 1'b0 ;
  assign n24626 = n1654 | n3364 ;
  assign n24627 = n9783 | n24626 ;
  assign n24628 = ( n7558 & n17885 ) | ( n7558 & n24627 ) | ( n17885 & n24627 ) ;
  assign n24629 = n8130 ^ n4578 ^ 1'b0 ;
  assign n24630 = n13220 & n24629 ;
  assign n24631 = n2855 & n4350 ;
  assign n24632 = ~n3736 & n24631 ;
  assign n24633 = ~n24630 & n24632 ;
  assign n24634 = n24633 ^ n5725 ^ 1'b0 ;
  assign n24635 = ~n12206 & n24634 ;
  assign n24636 = n9977 & ~n24635 ;
  assign n24637 = n2020 & n3459 ;
  assign n24641 = ~n9377 & n10428 ;
  assign n24642 = n24641 ^ n4240 ^ 1'b0 ;
  assign n24643 = n14001 & n24642 ;
  assign n24644 = n12658 & n24643 ;
  assign n24638 = n19833 ^ n12221 ^ 1'b0 ;
  assign n24639 = n6215 | n24638 ;
  assign n24640 = n4640 & n24639 ;
  assign n24645 = n24644 ^ n24640 ^ 1'b0 ;
  assign n24646 = n3592 & ~n24645 ;
  assign n24647 = n10309 | n16979 ;
  assign n24648 = ~n6689 & n24647 ;
  assign n24649 = n1064 & n24648 ;
  assign n24650 = n22766 ^ n13829 ^ 1'b0 ;
  assign n24651 = n24649 | n24650 ;
  assign n24654 = n2082 | n22712 ;
  assign n24655 = n24654 ^ n4324 ^ 1'b0 ;
  assign n24656 = n24655 ^ n471 ^ n131 ;
  assign n24652 = n6793 ^ n5866 ^ n308 ;
  assign n24653 = n8353 & ~n24652 ;
  assign n24657 = n24656 ^ n24653 ^ 1'b0 ;
  assign n24658 = n4637 | n7659 ;
  assign n24659 = ~n12845 & n24658 ;
  assign n24660 = ( ~n4540 & n7975 ) | ( ~n4540 & n24659 ) | ( n7975 & n24659 ) ;
  assign n24661 = n8988 ^ n8395 ^ 1'b0 ;
  assign n24662 = n7304 & n24661 ;
  assign n24663 = n12959 ^ n10265 ^ n1312 ;
  assign n24664 = ( ~n1359 & n8166 ) | ( ~n1359 & n24663 ) | ( n8166 & n24663 ) ;
  assign n24665 = ~n15774 & n24664 ;
  assign n24666 = n19433 ^ n13138 ^ n10852 ;
  assign n24667 = n1036 & ~n24666 ;
  assign n24668 = n24665 & n24667 ;
  assign n24669 = n5118 ^ n2036 ^ 1'b0 ;
  assign n24670 = n132 | n24669 ;
  assign n24671 = n22673 ^ n12775 ^ n4318 ;
  assign n24672 = ( n1545 & n3508 ) | ( n1545 & ~n24671 ) | ( n3508 & ~n24671 ) ;
  assign n24673 = n6383 ^ n498 ^ 1'b0 ;
  assign n24674 = n1400 & n24673 ;
  assign n24675 = ( ~n176 & n3926 ) | ( ~n176 & n15320 ) | ( n3926 & n15320 ) ;
  assign n24676 = n2832 | n24675 ;
  assign n24677 = n24676 ^ n59 ^ 1'b0 ;
  assign n24678 = n24674 & n24677 ;
  assign n24679 = ( n3135 & n5316 ) | ( n3135 & n18835 ) | ( n5316 & n18835 ) ;
  assign n24680 = n15865 ^ n4913 ^ 1'b0 ;
  assign n24681 = n4516 | n24680 ;
  assign n24682 = n24681 ^ n665 ^ 1'b0 ;
  assign n24683 = ~n24679 & n24682 ;
  assign n24684 = n2565 | n11253 ;
  assign n24685 = n6064 | n22023 ;
  assign n24686 = n16025 | n24685 ;
  assign n24687 = n10548 ^ n6691 ^ n802 ;
  assign n24688 = n563 & n24380 ;
  assign n24689 = n24687 & n24688 ;
  assign n24690 = n20302 ^ n10957 ^ 1'b0 ;
  assign n24691 = ~n24689 & n24690 ;
  assign n24692 = n2207 | n24691 ;
  assign n24693 = ~n55 & n10088 ;
  assign n24694 = n24693 ^ n3305 ^ 1'b0 ;
  assign n24695 = ( ~n8751 & n12855 ) | ( ~n8751 & n24694 ) | ( n12855 & n24694 ) ;
  assign n24696 = n6493 | n9119 ;
  assign n24697 = n24696 ^ n18025 ^ 1'b0 ;
  assign n24698 = ( n3428 & n8411 ) | ( n3428 & n24697 ) | ( n8411 & n24697 ) ;
  assign n24699 = ~n9638 & n18161 ;
  assign n24700 = n24699 ^ n20602 ^ n14272 ;
  assign n24701 = n17836 ^ n16487 ^ 1'b0 ;
  assign n24702 = n17906 & n24701 ;
  assign n24704 = n5229 & ~n5515 ;
  assign n24705 = n24704 ^ n390 ^ 1'b0 ;
  assign n24703 = ~n10034 & n14386 ;
  assign n24706 = n24705 ^ n24703 ^ n6888 ;
  assign n24707 = ( ~n7759 & n9033 ) | ( ~n7759 & n14409 ) | ( n9033 & n14409 ) ;
  assign n24708 = n8297 | n24707 ;
  assign n24709 = n24708 ^ n698 ^ 1'b0 ;
  assign n24710 = n20362 ^ n11344 ^ 1'b0 ;
  assign n24711 = n22740 | n24710 ;
  assign n24712 = n37 & n2696 ;
  assign n24713 = n23097 ^ n20826 ^ n5179 ;
  assign n24714 = n7487 ^ n6696 ^ n6474 ;
  assign n24715 = n13276 | n24714 ;
  assign n24716 = n3606 ^ n3199 ^ 1'b0 ;
  assign n24717 = ( n7101 & n11386 ) | ( n7101 & n12289 ) | ( n11386 & n12289 ) ;
  assign n24718 = n24717 ^ n9263 ^ n1064 ;
  assign n24719 = ~n12059 & n24718 ;
  assign n24720 = ~n24716 & n24719 ;
  assign n24721 = n24251 & n24720 ;
  assign n24724 = n10219 ^ n8379 ^ n5092 ;
  assign n24722 = n2368 & n8746 ;
  assign n24723 = ~n13529 & n24722 ;
  assign n24725 = n24724 ^ n24723 ^ 1'b0 ;
  assign n24726 = ( n7976 & n15829 ) | ( n7976 & ~n24725 ) | ( n15829 & ~n24725 ) ;
  assign n24727 = ( n12808 & n14008 ) | ( n12808 & n16232 ) | ( n14008 & n16232 ) ;
  assign n24728 = ~n13153 & n24727 ;
  assign n24729 = ( ~n362 & n10282 ) | ( ~n362 & n20086 ) | ( n10282 & n20086 ) ;
  assign n24730 = n10583 & ~n15826 ;
  assign n24731 = n9683 & ~n24730 ;
  assign n24734 = n708 & ~n4920 ;
  assign n24735 = n2128 & n24734 ;
  assign n24732 = n4124 ^ n3789 ^ 1'b0 ;
  assign n24733 = n9899 & ~n24732 ;
  assign n24736 = n24735 ^ n24733 ^ 1'b0 ;
  assign n24737 = ( n4549 & n8833 ) | ( n4549 & n24736 ) | ( n8833 & n24736 ) ;
  assign n24738 = n9434 & n9529 ;
  assign n24739 = ~n601 & n24738 ;
  assign n24740 = n24737 & ~n24739 ;
  assign n24741 = n18773 ^ n2545 ^ 1'b0 ;
  assign n24742 = n2569 | n24741 ;
  assign n24743 = n6678 | n15250 ;
  assign n24744 = n9255 | n18074 ;
  assign n24745 = n14481 ^ n7977 ^ n217 ;
  assign n24746 = n24745 ^ n2319 ^ 1'b0 ;
  assign n24747 = n3837 ^ n1427 ^ 1'b0 ;
  assign n24748 = n7648 & ~n24747 ;
  assign n24749 = n8979 & ~n24748 ;
  assign n24750 = n24749 ^ n19917 ^ 1'b0 ;
  assign n24751 = n7516 & ~n24750 ;
  assign n24752 = n17376 ^ n3708 ^ 1'b0 ;
  assign n24753 = n2449 & n12845 ;
  assign n24754 = ~n3677 & n24753 ;
  assign n24755 = ( ~n2044 & n6511 ) | ( ~n2044 & n7102 ) | ( n6511 & n7102 ) ;
  assign n24756 = ~n909 & n24755 ;
  assign n24757 = n24756 ^ n8947 ^ 1'b0 ;
  assign n24758 = n16284 & ~n24757 ;
  assign n24759 = n24754 & n24758 ;
  assign n24760 = n12596 & n24759 ;
  assign n24761 = n4290 | n9141 ;
  assign n24762 = n10269 ^ n5430 ^ 1'b0 ;
  assign n24763 = ( ~n6758 & n24761 ) | ( ~n6758 & n24762 ) | ( n24761 & n24762 ) ;
  assign n24764 = n2257 ^ n352 ^ 1'b0 ;
  assign n24765 = n14450 & ~n18872 ;
  assign n24766 = ~n2722 & n19929 ;
  assign n24767 = ( ~n5197 & n8804 ) | ( ~n5197 & n9564 ) | ( n8804 & n9564 ) ;
  assign n24768 = n24766 & ~n24767 ;
  assign n24769 = n8424 ^ n4328 ^ 1'b0 ;
  assign n24770 = ~n16016 & n24769 ;
  assign n24771 = n24770 ^ n10751 ^ 1'b0 ;
  assign n24772 = n4334 | n9989 ;
  assign n24773 = ( n2606 & n18316 ) | ( n2606 & ~n24772 ) | ( n18316 & ~n24772 ) ;
  assign n24774 = n3707 | n22899 ;
  assign n24775 = n24774 ^ n1633 ^ 1'b0 ;
  assign n24776 = n23133 ^ n8560 ^ 1'b0 ;
  assign n24777 = n9216 ^ n5494 ^ 1'b0 ;
  assign n24778 = ~n20831 & n24777 ;
  assign n24779 = ~n14116 & n24778 ;
  assign n24780 = n24779 ^ n15182 ^ 1'b0 ;
  assign n24781 = ( n829 & ~n9796 ) | ( n829 & n24780 ) | ( ~n9796 & n24780 ) ;
  assign n24782 = n21146 ^ n11065 ^ 1'b0 ;
  assign n24785 = ( n220 & n2045 ) | ( n220 & ~n9202 ) | ( n2045 & ~n9202 ) ;
  assign n24783 = n7718 & ~n8713 ;
  assign n24784 = n836 & ~n24783 ;
  assign n24786 = n24785 ^ n24784 ^ 1'b0 ;
  assign n24787 = n24786 ^ n23320 ^ 1'b0 ;
  assign n24788 = n12285 | n12935 ;
  assign n24789 = ~n2297 & n8832 ;
  assign n24790 = n24788 & ~n24789 ;
  assign n24791 = n11833 | n24790 ;
  assign n24792 = n18556 & ~n24791 ;
  assign n24793 = n8975 & ~n11868 ;
  assign n24799 = n11942 & ~n22558 ;
  assign n24800 = n6460 | n24799 ;
  assign n24801 = n24800 ^ n10376 ^ 1'b0 ;
  assign n24794 = n3897 ^ n3305 ^ 1'b0 ;
  assign n24795 = n24794 ^ n19402 ^ 1'b0 ;
  assign n24796 = n21589 | n24795 ;
  assign n24797 = n24796 ^ n23177 ^ 1'b0 ;
  assign n24798 = n14845 & n24797 ;
  assign n24802 = n24801 ^ n24798 ^ 1'b0 ;
  assign n24803 = n16977 & ~n23911 ;
  assign n24804 = n13703 & n24803 ;
  assign n24807 = ~n5582 & n8693 ;
  assign n24805 = n1875 & ~n5008 ;
  assign n24806 = ~n5229 & n24805 ;
  assign n24808 = n24807 ^ n24806 ^ n19741 ;
  assign n24809 = ( n12754 & n18344 ) | ( n12754 & n18401 ) | ( n18344 & n18401 ) ;
  assign n24810 = n6193 | n24809 ;
  assign n24811 = n24810 ^ n16861 ^ 1'b0 ;
  assign n24812 = n1810 & ~n11023 ;
  assign n24813 = ~n13346 & n24812 ;
  assign n24814 = n8425 & n24813 ;
  assign n24815 = n6648 ^ n6239 ^ 1'b0 ;
  assign n24816 = ~n13362 & n13784 ;
  assign n24817 = n24816 ^ n24465 ^ 1'b0 ;
  assign n24818 = ( n17232 & n24815 ) | ( n17232 & n24817 ) | ( n24815 & n24817 ) ;
  assign n24819 = ~n20831 & n24818 ;
  assign n24820 = ~n3626 & n11554 ;
  assign n24821 = n24820 ^ n10178 ^ 1'b0 ;
  assign n24822 = n1556 ^ n1173 ^ 1'b0 ;
  assign n24823 = n209 & n11057 ;
  assign n24824 = n24823 ^ n11667 ^ 1'b0 ;
  assign n24825 = ( n19288 & n24822 ) | ( n19288 & n24824 ) | ( n24822 & n24824 ) ;
  assign n24826 = ~n9653 & n10352 ;
  assign n24827 = ~n18541 & n24826 ;
  assign n24828 = n3435 & ~n24827 ;
  assign n24829 = n24828 ^ n24805 ^ 1'b0 ;
  assign n24830 = n15437 ^ n2776 ^ 1'b0 ;
  assign n24831 = n11062 & n24830 ;
  assign n24832 = ~n18859 & n24831 ;
  assign n24833 = n3456 & ~n16042 ;
  assign n24834 = n24833 ^ n5305 ^ 1'b0 ;
  assign n24835 = n2561 & n5246 ;
  assign n24836 = ( n126 & ~n4164 ) | ( n126 & n24835 ) | ( ~n4164 & n24835 ) ;
  assign n24837 = n766 & n24836 ;
  assign n24838 = n7354 & ~n24837 ;
  assign n24839 = n19394 & n24838 ;
  assign n24840 = ~n3483 & n14282 ;
  assign n24841 = ( ~n644 & n5531 ) | ( ~n644 & n24840 ) | ( n5531 & n24840 ) ;
  assign n24842 = n24841 ^ n12779 ^ n2740 ;
  assign n24843 = n5129 ^ n1279 ^ 1'b0 ;
  assign n24844 = ~n24842 & n24843 ;
  assign n24845 = n3428 ^ n299 ^ 1'b0 ;
  assign n24846 = n24844 & ~n24845 ;
  assign n24847 = n24846 ^ n7932 ^ 1'b0 ;
  assign n24848 = ~n22620 & n24847 ;
  assign n24849 = n2537 | n13037 ;
  assign n24850 = n19807 & ~n24849 ;
  assign n24851 = n18786 ^ n9543 ^ 1'b0 ;
  assign n24852 = n4846 & n11105 ;
  assign n24853 = n15960 | n24852 ;
  assign n24854 = n24853 ^ n22588 ^ 1'b0 ;
  assign n24855 = n18522 ^ n14394 ^ 1'b0 ;
  assign n24856 = n7850 | n24855 ;
  assign n24857 = n6992 & ~n20426 ;
  assign n24858 = n24856 | n24857 ;
  assign n24859 = n1962 & ~n24858 ;
  assign n24860 = ( n492 & ~n1371 ) | ( n492 & n12080 ) | ( ~n1371 & n12080 ) ;
  assign n24861 = n24860 ^ n10564 ^ 1'b0 ;
  assign n24862 = n6287 | n24861 ;
  assign n24863 = n6274 & n12821 ;
  assign n24864 = n14187 & ~n18786 ;
  assign n24865 = n4733 & ~n5135 ;
  assign n24866 = ~n6101 & n24865 ;
  assign n24869 = n19172 ^ n12395 ^ 1'b0 ;
  assign n24867 = n2655 & n20281 ;
  assign n24868 = n21980 & n24867 ;
  assign n24870 = n24869 ^ n24868 ^ 1'b0 ;
  assign n24871 = ~n24866 & n24870 ;
  assign n24872 = n10382 ^ n8097 ^ 1'b0 ;
  assign n24873 = ~n2074 & n24872 ;
  assign n24874 = n24873 ^ n2205 ^ 1'b0 ;
  assign n24875 = ~n2131 & n24874 ;
  assign n24876 = n41 & n10876 ;
  assign n24877 = ( n5911 & n11567 ) | ( n5911 & ~n24876 ) | ( n11567 & ~n24876 ) ;
  assign n24878 = n10712 ^ n6678 ^ 1'b0 ;
  assign n24879 = n1069 & n24878 ;
  assign n24880 = n24879 ^ n2104 ^ 1'b0 ;
  assign n24881 = n24877 | n24880 ;
  assign n24882 = n4320 | n16495 ;
  assign n24883 = n14732 & ~n24882 ;
  assign n24884 = n11944 ^ n7469 ^ 1'b0 ;
  assign n24885 = ~n1805 & n24884 ;
  assign n24886 = ~n20064 & n24885 ;
  assign n24887 = n13882 & n24886 ;
  assign n24888 = ( n888 & n3708 ) | ( n888 & n18829 ) | ( n3708 & n18829 ) ;
  assign n24889 = n8854 ^ n5026 ^ 1'b0 ;
  assign n24891 = n7742 & n12184 ;
  assign n24890 = n17104 ^ n4685 ^ 1'b0 ;
  assign n24892 = n24891 ^ n24890 ^ 1'b0 ;
  assign n24893 = ~n11404 & n24892 ;
  assign n24894 = n17690 ^ n12073 ^ n11376 ;
  assign n24895 = n24893 & n24894 ;
  assign n24896 = ~n24889 & n24895 ;
  assign n24900 = ~n6449 & n20805 ;
  assign n24897 = n2818 ^ n2328 ^ 1'b0 ;
  assign n24898 = n24897 ^ n20062 ^ n12459 ;
  assign n24899 = n5477 | n24898 ;
  assign n24901 = n24900 ^ n24899 ^ 1'b0 ;
  assign n24902 = n6277 ^ n4656 ^ 1'b0 ;
  assign n24903 = n24902 ^ n9676 ^ n503 ;
  assign n24904 = n1853 & ~n24903 ;
  assign n24905 = n905 | n1201 ;
  assign n24906 = n9717 ^ n676 ^ 1'b0 ;
  assign n24907 = n10100 & ~n24906 ;
  assign n24908 = n24905 & n24907 ;
  assign n24909 = n19803 | n24908 ;
  assign n24910 = n15584 ^ n11249 ^ n7240 ;
  assign n24911 = n15809 ^ n7433 ^ 1'b0 ;
  assign n24912 = ( ~n194 & n17141 ) | ( ~n194 & n19665 ) | ( n17141 & n19665 ) ;
  assign n24913 = n24912 ^ n8201 ^ 1'b0 ;
  assign n24914 = ~n20720 & n24913 ;
  assign n24915 = n1198 | n3043 ;
  assign n24916 = n1298 & ~n24915 ;
  assign n24917 = n24916 ^ n5481 ^ 1'b0 ;
  assign n24918 = n13282 ^ n10226 ^ n105 ;
  assign n24920 = n1318 | n1926 ;
  assign n24921 = n1433 | n24920 ;
  assign n24919 = n411 | n7210 ;
  assign n24922 = n24921 ^ n24919 ^ 1'b0 ;
  assign n24923 = ( n3070 & n9299 ) | ( n3070 & ~n24922 ) | ( n9299 & ~n24922 ) ;
  assign n24924 = n24923 ^ n7255 ^ 1'b0 ;
  assign n24925 = n24918 & ~n24924 ;
  assign n24926 = n10905 & n24925 ;
  assign n24927 = ~n446 & n2314 ;
  assign n24928 = n7718 | n24927 ;
  assign n24929 = n24927 & ~n24928 ;
  assign n24930 = n6664 | n24929 ;
  assign n24931 = n24929 & ~n24930 ;
  assign n24932 = n6940 | n24931 ;
  assign n24933 = n6940 & ~n24932 ;
  assign n24934 = n17675 ^ n2770 ^ 1'b0 ;
  assign n24941 = n9610 & n16405 ;
  assign n24942 = n24941 ^ n15021 ^ 1'b0 ;
  assign n24935 = n10647 ^ n3688 ^ 1'b0 ;
  assign n24936 = n6380 | n24935 ;
  assign n24937 = n21316 ^ n6968 ^ 1'b0 ;
  assign n24938 = n649 & n24937 ;
  assign n24939 = ~n2983 & n24938 ;
  assign n24940 = ~n24936 & n24939 ;
  assign n24943 = n24942 ^ n24940 ^ 1'b0 ;
  assign n24945 = n11778 & n18575 ;
  assign n24946 = ~n11902 & n24945 ;
  assign n24944 = ~n10760 & n12727 ;
  assign n24947 = n24946 ^ n24944 ^ 1'b0 ;
  assign n24948 = n2909 & n4057 ;
  assign n24949 = n24948 ^ n15046 ^ 1'b0 ;
  assign n24950 = ( ~n20066 & n23001 ) | ( ~n20066 & n24949 ) | ( n23001 & n24949 ) ;
  assign n24951 = n13997 ^ n3240 ^ 1'b0 ;
  assign n24952 = ~n10537 & n11854 ;
  assign n24953 = n19038 | n21725 ;
  assign n24954 = ~n1134 & n22653 ;
  assign n24955 = n5567 & n24954 ;
  assign n24956 = n10040 ^ n4334 ^ 1'b0 ;
  assign n24957 = ( ~n15969 & n19280 ) | ( ~n15969 & n24956 ) | ( n19280 & n24956 ) ;
  assign n24958 = n14784 ^ n4383 ^ 1'b0 ;
  assign n24959 = n8508 ^ n3922 ^ n1744 ;
  assign n24960 = n24958 & ~n24959 ;
  assign n24961 = n21550 ^ n16127 ^ 1'b0 ;
  assign n24962 = n24961 ^ n2939 ^ 1'b0 ;
  assign n24963 = n24962 ^ n421 ^ 1'b0 ;
  assign n24964 = n8938 & n12339 ;
  assign n24965 = ~n3025 & n24964 ;
  assign n24966 = n16455 ^ n12698 ^ 1'b0 ;
  assign n24967 = n432 & ~n710 ;
  assign n24968 = n24967 ^ n11401 ^ 1'b0 ;
  assign n24970 = ( n5139 & n6155 ) | ( n5139 & n9583 ) | ( n6155 & n9583 ) ;
  assign n24971 = n10025 & n10793 ;
  assign n24972 = n24970 & n24971 ;
  assign n24969 = n2447 ^ n954 ^ 1'b0 ;
  assign n24973 = n24972 ^ n24969 ^ n16942 ;
  assign n24974 = n24973 ^ n14889 ^ 1'b0 ;
  assign n24975 = n18694 | n24974 ;
  assign n24976 = n14997 ^ n12867 ^ 1'b0 ;
  assign n24977 = n24976 ^ n4114 ^ 1'b0 ;
  assign n24978 = ~n8031 & n13133 ;
  assign n24979 = n4660 | n21419 ;
  assign n24980 = n24978 & ~n24979 ;
  assign n24981 = n14078 & ~n24980 ;
  assign n24982 = n24981 ^ n9884 ^ 1'b0 ;
  assign n24983 = n417 & n8110 ;
  assign n24984 = ~n436 & n24983 ;
  assign n24985 = n3931 | n24984 ;
  assign n24986 = n24982 & n24985 ;
  assign n24987 = n8738 ^ n4303 ^ 1'b0 ;
  assign n24988 = n9504 ^ n1768 ^ 1'b0 ;
  assign n24989 = n24837 ^ n15083 ^ 1'b0 ;
  assign n24990 = n7308 | n15879 ;
  assign n24991 = n24990 ^ n15217 ^ 1'b0 ;
  assign n24992 = n23378 | n24991 ;
  assign n24993 = n24992 ^ n99 ^ 1'b0 ;
  assign n24994 = n22766 ^ n1170 ^ 1'b0 ;
  assign n24995 = n614 | n24994 ;
  assign n24996 = ~n6320 & n7545 ;
  assign n24997 = n12961 | n24996 ;
  assign n24998 = n24997 ^ n51 ^ 1'b0 ;
  assign n24999 = n8076 & ~n24998 ;
  assign n25000 = ~n12928 & n24999 ;
  assign n25001 = n11927 | n25000 ;
  assign n25002 = n8130 & n15759 ;
  assign n25003 = n5402 | n8355 ;
  assign n25004 = n18353 | n25003 ;
  assign n25006 = ( ~n4775 & n9857 ) | ( ~n4775 & n15130 ) | ( n9857 & n15130 ) ;
  assign n25007 = n25006 ^ n19775 ^ 1'b0 ;
  assign n25008 = n5841 & ~n25007 ;
  assign n25005 = n10145 | n12150 ;
  assign n25009 = n25008 ^ n25005 ^ 1'b0 ;
  assign n25010 = n8594 ^ n4333 ^ 1'b0 ;
  assign n25011 = n15552 & ~n20959 ;
  assign n25012 = ~n12969 & n14846 ;
  assign n25013 = n25012 ^ n12632 ^ 1'b0 ;
  assign n25014 = n5706 ^ n5234 ^ 1'b0 ;
  assign n25015 = n1026 | n25014 ;
  assign n25016 = n22990 & ~n25015 ;
  assign n25017 = n4147 & ~n25016 ;
  assign n25018 = n25017 ^ n11082 ^ 1'b0 ;
  assign n25019 = n9884 ^ n5175 ^ 1'b0 ;
  assign n25020 = n9325 & n25019 ;
  assign n25021 = n2818 & n4704 ;
  assign n25022 = n25021 ^ n4225 ^ 1'b0 ;
  assign n25023 = n25022 ^ n8978 ^ 1'b0 ;
  assign n25024 = n7776 & ~n22954 ;
  assign n25025 = n11450 & n25024 ;
  assign n25026 = n23978 ^ n645 ^ 1'b0 ;
  assign n25028 = n14764 ^ n6213 ^ 1'b0 ;
  assign n25027 = n12026 & n20310 ;
  assign n25029 = n25028 ^ n25027 ^ 1'b0 ;
  assign n25032 = ~n4544 & n11225 ;
  assign n25030 = ( n7912 & ~n9623 ) | ( n7912 & n20943 ) | ( ~n9623 & n20943 ) ;
  assign n25031 = n25030 ^ n2463 ^ 1'b0 ;
  assign n25033 = n25032 ^ n25031 ^ 1'b0 ;
  assign n25034 = n4421 & n25033 ;
  assign n25035 = ~n14017 & n24202 ;
  assign n25036 = ( ~n532 & n10395 ) | ( ~n532 & n16301 ) | ( n10395 & n16301 ) ;
  assign n25038 = n15051 ^ n2864 ^ 1'b0 ;
  assign n25039 = n3144 | n25038 ;
  assign n25040 = n5321 | n25039 ;
  assign n25041 = n25040 ^ n1348 ^ 1'b0 ;
  assign n25037 = ~n3571 & n4712 ;
  assign n25042 = n25041 ^ n25037 ^ 1'b0 ;
  assign n25043 = n25042 ^ n23095 ^ 1'b0 ;
  assign n25044 = ~n13059 & n16765 ;
  assign n25045 = n24770 ^ n10878 ^ 1'b0 ;
  assign n25046 = n158 & ~n401 ;
  assign n25047 = n1399 & n25046 ;
  assign n25048 = n12707 | n25047 ;
  assign n25049 = n11403 ^ n7221 ^ 1'b0 ;
  assign n25050 = ~n12612 & n25049 ;
  assign n25051 = n15692 ^ n8465 ^ 1'b0 ;
  assign n25052 = n25050 & ~n25051 ;
  assign n25053 = ~n1768 & n4614 ;
  assign n25054 = n25053 ^ n10037 ^ 1'b0 ;
  assign n25055 = n10989 & ~n25054 ;
  assign n25056 = n25055 ^ n9143 ^ 1'b0 ;
  assign n25058 = n14343 ^ n12759 ^ 1'b0 ;
  assign n25057 = n15014 & ~n15503 ;
  assign n25059 = n25058 ^ n25057 ^ 1'b0 ;
  assign n25064 = n18111 ^ n10362 ^ n8906 ;
  assign n25062 = n1611 & ~n19346 ;
  assign n25063 = ~n40 & n25062 ;
  assign n25060 = n9295 ^ n1830 ^ 1'b0 ;
  assign n25061 = n5504 & n25060 ;
  assign n25065 = n25064 ^ n25063 ^ n25061 ;
  assign n25066 = n20011 ^ n15119 ^ 1'b0 ;
  assign n25067 = ~n12852 & n25066 ;
  assign n25068 = ~n9213 & n25067 ;
  assign n25069 = n25068 ^ n24902 ^ n6609 ;
  assign n25070 = n15653 ^ n205 ^ 1'b0 ;
  assign n25071 = n863 | n25070 ;
  assign n25072 = ( ~n879 & n4638 ) | ( ~n879 & n5001 ) | ( n4638 & n5001 ) ;
  assign n25073 = n5571 | n25072 ;
  assign n25074 = n3976 | n9973 ;
  assign n25075 = n916 & n25074 ;
  assign n25076 = n2208 & n25075 ;
  assign n25077 = n25076 ^ n523 ^ n294 ;
  assign n25078 = n5312 ^ n1789 ^ 1'b0 ;
  assign n25079 = n25077 & n25078 ;
  assign n25080 = n21707 & n25079 ;
  assign n25081 = ( n9760 & n17129 ) | ( n9760 & ~n25080 ) | ( n17129 & ~n25080 ) ;
  assign n25082 = ~n3514 & n25081 ;
  assign n25083 = n1108 & n5209 ;
  assign n25084 = n11132 | n14403 ;
  assign n25085 = n25084 ^ n9787 ^ 1'b0 ;
  assign n25086 = n25085 ^ n17424 ^ 1'b0 ;
  assign n25087 = n12694 ^ n8197 ^ 1'b0 ;
  assign n25088 = n25087 ^ n2791 ^ 1'b0 ;
  assign n25089 = n2583 & ~n25088 ;
  assign n25090 = n11339 | n25089 ;
  assign n25091 = ( ~n1345 & n2537 ) | ( ~n1345 & n11138 ) | ( n2537 & n11138 ) ;
  assign n25092 = n10734 ^ n9541 ^ 1'b0 ;
  assign n25093 = ~n25091 & n25092 ;
  assign n25094 = n18765 & n19785 ;
  assign n25095 = n16082 ^ n5554 ^ n1943 ;
  assign n25096 = n25095 ^ n20712 ^ 1'b0 ;
  assign n25097 = n10523 ^ n1505 ^ 1'b0 ;
  assign n25098 = n25097 ^ n17220 ^ 1'b0 ;
  assign n25099 = n20560 & n25098 ;
  assign n25100 = n2325 & ~n14827 ;
  assign n25101 = n6542 & ~n25100 ;
  assign n25102 = n11239 & n15617 ;
  assign n25103 = n25102 ^ n20815 ^ 1'b0 ;
  assign n25104 = n25103 ^ n21978 ^ 1'b0 ;
  assign n25105 = ~n25101 & n25104 ;
  assign n25107 = n16798 ^ n2977 ^ 1'b0 ;
  assign n25106 = ~n645 & n11135 ;
  assign n25108 = n25107 ^ n25106 ^ 1'b0 ;
  assign n25109 = n25108 ^ n7790 ^ 1'b0 ;
  assign n25110 = ~n954 & n25109 ;
  assign n25111 = n771 & n20062 ;
  assign n25112 = n10311 ^ n7572 ^ n3281 ;
  assign n25113 = n25112 ^ n16844 ^ n5554 ;
  assign n25114 = n1807 & n2979 ;
  assign n25115 = n25114 ^ n2787 ^ 1'b0 ;
  assign n25116 = n8909 | n25115 ;
  assign n25117 = n7287 ^ n882 ^ 1'b0 ;
  assign n25118 = n17441 ^ n902 ^ 1'b0 ;
  assign n25119 = n16567 & n25118 ;
  assign n25120 = n10743 & n25119 ;
  assign n25121 = n6553 ^ n2977 ^ 1'b0 ;
  assign n25122 = n2725 | n3770 ;
  assign n25123 = n25121 & ~n25122 ;
  assign n25124 = n15940 & ~n24135 ;
  assign n25125 = ~n8323 & n25124 ;
  assign n25126 = n25123 | n25125 ;
  assign n25127 = ~n13028 & n15542 ;
  assign n25128 = n25127 ^ n9666 ^ 1'b0 ;
  assign n25129 = ~n21619 & n25128 ;
  assign n25130 = n25126 & n25129 ;
  assign n25131 = n1003 & ~n11111 ;
  assign n25132 = ~n11396 & n15584 ;
  assign n25133 = n25132 ^ n18754 ^ 1'b0 ;
  assign n25134 = n865 | n25133 ;
  assign n25135 = n25131 | n25134 ;
  assign n25136 = ~n14784 & n25135 ;
  assign n25137 = n25136 ^ n22198 ^ 1'b0 ;
  assign n25142 = n5583 ^ n2051 ^ 1'b0 ;
  assign n25138 = n1625 | n2825 ;
  assign n25139 = n15395 & n25138 ;
  assign n25140 = n4480 & ~n25139 ;
  assign n25141 = n25140 ^ n7074 ^ 1'b0 ;
  assign n25143 = n25142 ^ n25141 ^ n22925 ;
  assign n25147 = n15493 ^ n12634 ^ 1'b0 ;
  assign n25148 = ( n5393 & ~n17226 ) | ( n5393 & n25147 ) | ( ~n17226 & n25147 ) ;
  assign n25149 = ( ~n7676 & n11095 ) | ( ~n7676 & n25148 ) | ( n11095 & n25148 ) ;
  assign n25144 = n7457 ^ n5372 ^ 1'b0 ;
  assign n25145 = n21906 & n25144 ;
  assign n25146 = n25145 ^ n1182 ^ 1'b0 ;
  assign n25150 = n25149 ^ n25146 ^ n9901 ;
  assign n25151 = ~n14752 & n25150 ;
  assign n25152 = n6157 & ~n14077 ;
  assign n25153 = n9263 ^ n7147 ^ 1'b0 ;
  assign n25154 = n4605 | n6682 ;
  assign n25158 = n1120 & ~n21041 ;
  assign n25159 = n25158 ^ n1160 ^ 1'b0 ;
  assign n25155 = n1265 & n12451 ;
  assign n25156 = n10147 & n25155 ;
  assign n25157 = n13493 & n25156 ;
  assign n25160 = n25159 ^ n25157 ^ 1'b0 ;
  assign n25161 = n200 | n1800 ;
  assign n25162 = n14170 ^ n9146 ^ 1'b0 ;
  assign n25163 = n12166 & ~n17603 ;
  assign n25164 = n1563 & ~n4719 ;
  assign n25165 = n7963 ^ n5446 ^ 1'b0 ;
  assign n25166 = n2935 & n25165 ;
  assign n25167 = n12383 ^ n864 ^ 1'b0 ;
  assign n25168 = n15742 | n25167 ;
  assign n25169 = n15991 & ~n25168 ;
  assign n25170 = n14495 & ~n25169 ;
  assign n25171 = n2612 & ~n6993 ;
  assign n25172 = ~n2821 & n4338 ;
  assign n25173 = n2821 & n25172 ;
  assign n25174 = n25173 ^ n10382 ^ 1'b0 ;
  assign n25175 = n5261 & n25174 ;
  assign n25176 = n25175 ^ n2674 ^ 1'b0 ;
  assign n25177 = n3409 & n3981 ;
  assign n25178 = n25177 ^ n12439 ^ n589 ;
  assign n25179 = n25178 ^ n18560 ^ 1'b0 ;
  assign n25180 = n5902 ^ n3379 ^ 1'b0 ;
  assign n25181 = ~n21169 & n25180 ;
  assign n25182 = n18330 ^ n9210 ^ n879 ;
  assign n25183 = n7122 ^ n1200 ^ 1'b0 ;
  assign n25184 = n25182 & n25183 ;
  assign n25185 = ( n12791 & n24177 ) | ( n12791 & n25184 ) | ( n24177 & n25184 ) ;
  assign n25186 = n11159 ^ n9732 ^ 1'b0 ;
  assign n25187 = n18201 & ~n25186 ;
  assign n25188 = n432 & ~n16412 ;
  assign n25189 = ~n25187 & n25188 ;
  assign n25190 = n13176 & n18470 ;
  assign n25191 = ~n16295 & n25190 ;
  assign n25192 = n11655 | n25191 ;
  assign n25193 = n11059 & ~n25192 ;
  assign n25194 = n17906 ^ n3774 ^ 1'b0 ;
  assign n25195 = n1343 & ~n19461 ;
  assign n25196 = n25195 ^ n10291 ^ n7481 ;
  assign n25197 = n25196 ^ n3973 ^ 1'b0 ;
  assign n25198 = n1848 & ~n8150 ;
  assign n25199 = n8882 & n25198 ;
  assign n25200 = n6369 ^ n4207 ^ 1'b0 ;
  assign n25201 = n15375 | n25200 ;
  assign n25202 = n25201 ^ n13165 ^ 1'b0 ;
  assign n25203 = ( n401 & ~n965 ) | ( n401 & n25202 ) | ( ~n965 & n25202 ) ;
  assign n25204 = ( n18882 & n25199 ) | ( n18882 & ~n25203 ) | ( n25199 & ~n25203 ) ;
  assign n25205 = n16298 ^ n10560 ^ 1'b0 ;
  assign n25206 = ~n7588 & n25205 ;
  assign n25207 = n3009 & n20458 ;
  assign n25208 = ~n25206 & n25207 ;
  assign n25209 = n25208 ^ n13038 ^ n1843 ;
  assign n25210 = n44 | n2343 ;
  assign n25211 = n12946 & n25210 ;
  assign n25212 = n25211 ^ n17013 ^ 1'b0 ;
  assign n25213 = n2930 & n24831 ;
  assign n25214 = n12976 & ~n13584 ;
  assign n25215 = n2345 & n25214 ;
  assign n25216 = n25215 ^ n9517 ^ 1'b0 ;
  assign n25217 = n7558 & ~n25216 ;
  assign n25218 = n23869 & n25217 ;
  assign n25219 = n25218 ^ n17214 ^ 1'b0 ;
  assign n25220 = n25219 ^ n18273 ^ n6251 ;
  assign n25221 = ~n3296 & n4039 ;
  assign n25222 = n6653 ^ n645 ^ 1'b0 ;
  assign n25223 = ~n24961 & n25222 ;
  assign n25224 = n2695 & ~n15674 ;
  assign n25225 = n8143 & n25224 ;
  assign n25226 = n2587 | n25225 ;
  assign n25227 = n25223 | n25226 ;
  assign n25228 = ( n15152 & n17893 ) | ( n15152 & ~n18454 ) | ( n17893 & ~n18454 ) ;
  assign n25229 = ~n16907 & n18353 ;
  assign n25230 = n25228 & n25229 ;
  assign n25231 = ~n11416 & n14175 ;
  assign n25232 = n25231 ^ n12005 ^ 1'b0 ;
  assign n25233 = n25232 ^ n12966 ^ 1'b0 ;
  assign n25234 = ( n811 & n3830 ) | ( n811 & n5016 ) | ( n3830 & n5016 ) ;
  assign n25235 = ~n7126 & n25234 ;
  assign n25236 = n25235 ^ n5822 ^ 1'b0 ;
  assign n25238 = n9884 ^ n978 ^ 1'b0 ;
  assign n25237 = ~n2304 & n3057 ;
  assign n25239 = n25238 ^ n25237 ^ 1'b0 ;
  assign n25240 = ~n2172 & n25239 ;
  assign n25241 = n22558 & n25240 ;
  assign n25242 = ~n8721 & n12551 ;
  assign n25243 = ~n16126 & n25242 ;
  assign n25244 = n24185 ^ n8509 ^ 1'b0 ;
  assign n25245 = n560 & n8456 ;
  assign n25246 = ~n9619 & n25245 ;
  assign n25247 = n25246 ^ n9041 ^ 1'b0 ;
  assign n25248 = n25247 ^ n19012 ^ n12611 ;
  assign n25249 = n5486 & n17798 ;
  assign n25250 = n25249 ^ n24976 ^ 1'b0 ;
  assign n25251 = n9467 ^ n4925 ^ 1'b0 ;
  assign n25252 = n18667 ^ n17371 ^ 1'b0 ;
  assign n25253 = n25251 & n25252 ;
  assign n25254 = n3263 | n8120 ;
  assign n25255 = n25254 ^ n10368 ^ 1'b0 ;
  assign n25256 = n7174 ^ n3876 ^ 1'b0 ;
  assign n25257 = n14046 & ~n25256 ;
  assign n25258 = n9345 & n23919 ;
  assign n25259 = n25257 & n25258 ;
  assign n25260 = n1095 & n2481 ;
  assign n25261 = n9055 ^ n2606 ^ 1'b0 ;
  assign n25262 = n8789 | n25261 ;
  assign n25263 = ( n1518 & n25260 ) | ( n1518 & ~n25262 ) | ( n25260 & ~n25262 ) ;
  assign n25264 = n1188 & n14125 ;
  assign n25265 = n25264 ^ n12861 ^ 1'b0 ;
  assign n25266 = n17525 ^ n4290 ^ 1'b0 ;
  assign n25267 = n6883 | n25266 ;
  assign n25268 = n25267 ^ n4280 ^ 1'b0 ;
  assign n25269 = n5484 & ~n13514 ;
  assign n25270 = ~n2534 & n25269 ;
  assign n25271 = ~n23345 & n25270 ;
  assign n25272 = n2765 ^ n2667 ^ 1'b0 ;
  assign n25273 = n19755 & ~n25272 ;
  assign n25274 = n180 & ~n17569 ;
  assign n25275 = ~n25273 & n25274 ;
  assign n25276 = n6739 ^ n1401 ^ 1'b0 ;
  assign n25277 = n22514 ^ n6743 ^ 1'b0 ;
  assign n25278 = n25276 & n25277 ;
  assign n25279 = ( ~n6720 & n11465 ) | ( ~n6720 & n15190 ) | ( n11465 & n15190 ) ;
  assign n25280 = n17736 | n25279 ;
  assign n25281 = n25280 ^ n3067 ^ 1'b0 ;
  assign n25282 = n9501 & ~n10803 ;
  assign n25283 = n1049 & ~n3856 ;
  assign n25284 = n25179 | n25283 ;
  assign n25285 = n25284 ^ n18707 ^ 1'b0 ;
  assign n25286 = ~n2871 & n5451 ;
  assign n25287 = n13057 & n25286 ;
  assign n25290 = n14755 ^ n11886 ^ 1'b0 ;
  assign n25288 = n8882 ^ n1751 ^ 1'b0 ;
  assign n25289 = n25288 ^ n1758 ^ 1'b0 ;
  assign n25291 = n25290 ^ n25289 ^ 1'b0 ;
  assign n25292 = n25291 ^ n16290 ^ n9408 ;
  assign n25293 = ~n10087 & n25292 ;
  assign n25294 = n24003 & ~n25293 ;
  assign n25295 = n11255 | n17183 ;
  assign n25296 = n13586 ^ n10122 ^ 1'b0 ;
  assign n25297 = n25295 | n25296 ;
  assign n25298 = ~n10084 & n25297 ;
  assign n25299 = n6466 & ~n7140 ;
  assign n25300 = n25299 ^ n12290 ^ 1'b0 ;
  assign n25301 = n13729 ^ n1026 ^ 1'b0 ;
  assign n25302 = ~n5074 & n5870 ;
  assign n25303 = n25302 ^ n17251 ^ 1'b0 ;
  assign n25304 = n25303 ^ n11695 ^ 1'b0 ;
  assign n25305 = n25301 | n25304 ;
  assign n25307 = n22716 ^ n21943 ^ 1'b0 ;
  assign n25306 = ~n1095 & n16255 ;
  assign n25308 = n25307 ^ n25306 ^ 1'b0 ;
  assign n25309 = n15960 ^ n12499 ^ 1'b0 ;
  assign n25310 = n20217 ^ n16745 ^ 1'b0 ;
  assign n25311 = n3199 & n16181 ;
  assign n25336 = n4673 | n11777 ;
  assign n25337 = n2113 | n25336 ;
  assign n25335 = n16836 ^ n6921 ^ 1'b0 ;
  assign n25312 = n661 | n1286 ;
  assign n25313 = n25312 ^ n20696 ^ 1'b0 ;
  assign n25315 = n2721 ^ n1602 ^ n142 ;
  assign n25318 = n1175 | n1492 ;
  assign n25316 = n3918 ^ n2101 ^ 1'b0 ;
  assign n25317 = n2245 | n25316 ;
  assign n25319 = n25318 ^ n25317 ^ 1'b0 ;
  assign n25320 = ~n25315 & n25319 ;
  assign n25314 = n1721 & n17768 ;
  assign n25321 = n25320 ^ n25314 ^ 1'b0 ;
  assign n25322 = n3786 & ~n20619 ;
  assign n25323 = n24927 & n25322 ;
  assign n25324 = ( n1442 & ~n5876 ) | ( n1442 & n25323 ) | ( ~n5876 & n25323 ) ;
  assign n25325 = ( n2992 & ~n4271 ) | ( n2992 & n25324 ) | ( ~n4271 & n25324 ) ;
  assign n25327 = n11450 & ~n13425 ;
  assign n25328 = n2422 & n25327 ;
  assign n25326 = n5261 ^ n2390 ^ 1'b0 ;
  assign n25329 = n25328 ^ n25326 ^ n1328 ;
  assign n25330 = n9583 & ~n18371 ;
  assign n25331 = n3483 & n25330 ;
  assign n25332 = n7707 & n25331 ;
  assign n25333 = ( n25325 & n25329 ) | ( n25325 & n25332 ) | ( n25329 & n25332 ) ;
  assign n25334 = ( n25313 & n25321 ) | ( n25313 & ~n25333 ) | ( n25321 & ~n25333 ) ;
  assign n25338 = n25337 ^ n25335 ^ n25334 ;
  assign n25339 = ~n9616 & n25222 ;
  assign n25340 = n25339 ^ n3361 ^ 1'b0 ;
  assign n25341 = n9808 & ~n13670 ;
  assign n25342 = n25341 ^ n23836 ^ n20356 ;
  assign n25343 = n10424 ^ n10227 ^ n10161 ;
  assign n25344 = n1093 | n12754 ;
  assign n25345 = n25344 ^ n11618 ^ 1'b0 ;
  assign n25346 = n25343 | n25345 ;
  assign n25347 = n18626 ^ n3734 ^ 1'b0 ;
  assign n25348 = n5022 & n25347 ;
  assign n25349 = n9167 ^ n2526 ^ 1'b0 ;
  assign n25350 = n1370 & ~n13523 ;
  assign n25351 = ~n4325 & n25350 ;
  assign n25352 = n25351 ^ n15789 ^ 1'b0 ;
  assign n25353 = ~n17057 & n20972 ;
  assign n25354 = n7842 ^ n2254 ^ 1'b0 ;
  assign n25355 = n23409 & ~n25354 ;
  assign n25356 = n12249 ^ n9533 ^ n7433 ;
  assign n25357 = n25356 ^ n21719 ^ n10919 ;
  assign n25358 = n1261 & ~n6504 ;
  assign n25363 = n5026 ^ n3997 ^ 1'b0 ;
  assign n25364 = ~n1928 & n25363 ;
  assign n25365 = n14796 | n25364 ;
  assign n25361 = n434 & n4287 ;
  assign n25359 = n937 | n3048 ;
  assign n25360 = n25359 ^ n22797 ^ 1'b0 ;
  assign n25362 = n25361 ^ n25360 ^ n19026 ;
  assign n25366 = n25365 ^ n25362 ^ n7011 ;
  assign n25367 = n21600 | n25366 ;
  assign n25368 = n25367 ^ n21269 ^ 1'b0 ;
  assign n25369 = n4434 ^ n4226 ^ 1'b0 ;
  assign n25370 = n3710 & ~n25369 ;
  assign n25371 = ( n8616 & n10511 ) | ( n8616 & n25370 ) | ( n10511 & n25370 ) ;
  assign n25372 = n7506 | n25371 ;
  assign n25373 = n20931 ^ n1762 ^ n111 ;
  assign n25374 = n7884 & ~n10272 ;
  assign n25375 = n3085 | n25374 ;
  assign n25376 = n3824 & n5393 ;
  assign n25377 = n25376 ^ n19664 ^ 1'b0 ;
  assign n25378 = ( n1276 & n9770 ) | ( n1276 & n25377 ) | ( n9770 & n25377 ) ;
  assign n25379 = n12983 | n17915 ;
  assign n25380 = n9180 | n25379 ;
  assign n25382 = ( n2213 & n6357 ) | ( n2213 & ~n13949 ) | ( n6357 & ~n13949 ) ;
  assign n25381 = n2139 & ~n5678 ;
  assign n25383 = n25382 ^ n25381 ^ 1'b0 ;
  assign n25389 = n7383 ^ n2276 ^ 1'b0 ;
  assign n25384 = n12840 ^ n1710 ^ 1'b0 ;
  assign n25385 = n3478 | n25384 ;
  assign n25386 = n24627 ^ n11686 ^ 1'b0 ;
  assign n25387 = n25385 | n25386 ;
  assign n25388 = n25387 ^ n5251 ^ 1'b0 ;
  assign n25390 = n25389 ^ n25388 ^ n3581 ;
  assign n25391 = n16405 ^ n6556 ^ 1'b0 ;
  assign n25392 = n25391 ^ n6435 ^ 1'b0 ;
  assign n25393 = ~n19045 & n20242 ;
  assign n25394 = ~n475 & n14945 ;
  assign n25395 = n3660 & n22862 ;
  assign n25396 = n25395 ^ n13155 ^ 1'b0 ;
  assign n25397 = ( ~n1802 & n5906 ) | ( ~n1802 & n6022 ) | ( n5906 & n6022 ) ;
  assign n25398 = n17788 | n25397 ;
  assign n25399 = n25398 ^ n17608 ^ 1'b0 ;
  assign n25400 = n25396 & ~n25399 ;
  assign n25401 = n19988 ^ n4230 ^ 1'b0 ;
  assign n25402 = n25400 | n25401 ;
  assign n25403 = n10526 | n25402 ;
  assign n25404 = ~n3541 & n3893 ;
  assign n25405 = ( n2135 & n12135 ) | ( n2135 & n25404 ) | ( n12135 & n25404 ) ;
  assign n25408 = ~n1532 & n2523 ;
  assign n25409 = n10108 & n25408 ;
  assign n25406 = n11614 ^ n5244 ^ n2242 ;
  assign n25407 = n25406 ^ n21873 ^ 1'b0 ;
  assign n25410 = n25409 ^ n25407 ^ n12971 ;
  assign n25411 = n15053 ^ n7032 ^ 1'b0 ;
  assign n25412 = ~n5656 & n25411 ;
  assign n25413 = n25412 ^ n1605 ^ 1'b0 ;
  assign n25414 = ~n3170 & n11696 ;
  assign n25415 = n15953 & n25414 ;
  assign n25416 = n7918 & ~n25415 ;
  assign n25417 = n11488 ^ n3176 ^ 1'b0 ;
  assign n25418 = n3025 & ~n4945 ;
  assign n25419 = ~n25417 & n25418 ;
  assign n25420 = n25419 ^ n18034 ^ n4543 ;
  assign n25421 = n25420 ^ n17259 ^ n1512 ;
  assign n25422 = n25421 ^ n2823 ^ 1'b0 ;
  assign n25423 = n2431 & ~n25422 ;
  assign n25424 = n17849 & ~n19147 ;
  assign n25425 = ~n6646 & n25424 ;
  assign n25426 = n19892 | n20574 ;
  assign n25427 = n25426 ^ n17572 ^ 1'b0 ;
  assign n25428 = n25230 ^ n9541 ^ 1'b0 ;
  assign n25430 = n16691 ^ n8824 ^ 1'b0 ;
  assign n25431 = ~n5509 & n25430 ;
  assign n25429 = n6647 ^ n2657 ^ 1'b0 ;
  assign n25432 = n25431 ^ n25429 ^ 1'b0 ;
  assign n25433 = n2797 & n6985 ;
  assign n25434 = n5836 ^ n1131 ^ 1'b0 ;
  assign n25435 = n11736 | n25434 ;
  assign n25436 = n10435 ^ n7585 ^ 1'b0 ;
  assign n25438 = n14951 ^ n12456 ^ 1'b0 ;
  assign n25439 = ~n1848 & n25438 ;
  assign n25437 = n7252 ^ n6953 ^ 1'b0 ;
  assign n25440 = n25439 ^ n25437 ^ 1'b0 ;
  assign n25441 = n3433 & ~n25440 ;
  assign n25442 = n9667 ^ n1360 ^ 1'b0 ;
  assign n25443 = ( n861 & n8894 ) | ( n861 & n16914 ) | ( n8894 & n16914 ) ;
  assign n25444 = n18127 & ~n22895 ;
  assign n25445 = n2889 ^ n490 ^ 1'b0 ;
  assign n25446 = n25445 ^ n21345 ^ 1'b0 ;
  assign n25447 = n23089 & ~n25446 ;
  assign n25448 = n4217 & ~n11998 ;
  assign n25449 = n2885 & n25448 ;
  assign n25450 = ~n891 & n14580 ;
  assign n25451 = n9450 & ~n16914 ;
  assign n25453 = ~n7686 & n19501 ;
  assign n25452 = n24187 ^ n19971 ^ n13272 ;
  assign n25454 = n25453 ^ n25452 ^ 1'b0 ;
  assign n25455 = n14049 | n25454 ;
  assign n25456 = n25455 ^ n17133 ^ 1'b0 ;
  assign n25457 = ~n12869 & n14485 ;
  assign n25458 = n8337 & n21587 ;
  assign n25459 = ~n3732 & n25458 ;
  assign n25460 = n2228 | n25459 ;
  assign n25461 = n8470 | n20155 ;
  assign n25462 = ~n18021 & n25461 ;
  assign n25463 = ~n17902 & n25462 ;
  assign n25464 = n2359 & n25463 ;
  assign n25465 = n12514 & ~n16556 ;
  assign n25466 = n25464 & n25465 ;
  assign n25469 = n11220 & n11247 ;
  assign n25467 = n8275 | n10316 ;
  assign n25468 = n5992 | n25467 ;
  assign n25470 = n25469 ^ n25468 ^ 1'b0 ;
  assign n25471 = n9303 ^ n1439 ^ 1'b0 ;
  assign n25472 = n18522 & ~n25471 ;
  assign n25473 = n25194 & ~n25472 ;
  assign n25474 = n6365 & ~n20044 ;
  assign n25475 = n7795 & n25474 ;
  assign n25476 = n17659 | n25475 ;
  assign n25477 = n16159 ^ n15643 ^ n13371 ;
  assign n25478 = n25477 ^ n16173 ^ n8558 ;
  assign n25479 = n18242 & n19455 ;
  assign n25480 = n18819 ^ n11701 ^ 1'b0 ;
  assign n25481 = n25480 ^ n6743 ^ 1'b0 ;
  assign n25482 = n25479 & n25481 ;
  assign n25483 = n13069 & ~n25482 ;
  assign n25484 = n25483 ^ n18467 ^ 1'b0 ;
  assign n25485 = n6866 | n10313 ;
  assign n25486 = n25485 ^ n5640 ^ 1'b0 ;
  assign n25487 = ~n21469 & n25486 ;
  assign n25488 = n1023 ^ n884 ^ 1'b0 ;
  assign n25489 = ~n5037 & n25488 ;
  assign n25490 = ~n2686 & n7580 ;
  assign n25491 = ( n13760 & n14914 ) | ( n13760 & ~n23126 ) | ( n14914 & ~n23126 ) ;
  assign n25492 = n7219 | n13062 ;
  assign n25493 = ~n7440 & n10243 ;
  assign n25494 = ~n13907 & n25493 ;
  assign n25495 = n9753 | n23744 ;
  assign n25496 = n1944 & ~n25495 ;
  assign n25497 = n15926 ^ n2174 ^ 1'b0 ;
  assign n25498 = n21242 & ~n25497 ;
  assign n25499 = ( n1419 & n5399 ) | ( n1419 & n18063 ) | ( n5399 & n18063 ) ;
  assign n25500 = ~n10378 & n25499 ;
  assign n25501 = n8590 & n19689 ;
  assign n25502 = n8177 ^ n4104 ^ 1'b0 ;
  assign n25503 = n25502 ^ n15932 ^ 1'b0 ;
  assign n25504 = n17831 ^ n612 ^ 1'b0 ;
  assign n25505 = ( n1848 & n2732 ) | ( n1848 & n25504 ) | ( n2732 & n25504 ) ;
  assign n25506 = n5716 & ~n12805 ;
  assign n25509 = n2698 | n8172 ;
  assign n25507 = n6716 ^ n4945 ^ 1'b0 ;
  assign n25508 = n4154 | n25507 ;
  assign n25510 = n25509 ^ n25508 ^ 1'b0 ;
  assign n25511 = n12834 ^ n4892 ^ 1'b0 ;
  assign n25512 = ~n2566 & n21780 ;
  assign n25513 = n25511 & n25512 ;
  assign n25514 = n1866 & n2357 ;
  assign n25515 = ~n4631 & n25514 ;
  assign n25516 = n8972 | n24917 ;
  assign n25517 = n25516 ^ n15360 ^ 1'b0 ;
  assign n25518 = n601 & n14656 ;
  assign n25519 = n18813 | n25518 ;
  assign n25521 = n1382 & n10993 ;
  assign n25520 = ~n4193 & n16094 ;
  assign n25522 = n25521 ^ n25520 ^ 1'b0 ;
  assign n25523 = n25522 ^ n16295 ^ n10502 ;
  assign n25524 = ~n25519 & n25523 ;
  assign n25525 = n6916 | n18707 ;
  assign n25526 = n13391 & ~n14873 ;
  assign n25527 = ~n10830 & n25526 ;
  assign n25528 = n21935 & n25527 ;
  assign n25530 = n7705 & ~n17888 ;
  assign n25531 = n25530 ^ n18008 ^ 1'b0 ;
  assign n25529 = n2528 & ~n3093 ;
  assign n25532 = n25531 ^ n25529 ^ 1'b0 ;
  assign n25533 = ~n276 & n25532 ;
  assign n25534 = ( ~n2094 & n9275 ) | ( ~n2094 & n17531 ) | ( n9275 & n17531 ) ;
  assign n25535 = n25318 ^ n1885 ^ 1'b0 ;
  assign n25536 = ~n9635 & n24755 ;
  assign n25537 = n25536 ^ n8292 ^ 1'b0 ;
  assign n25538 = ~n22441 & n22608 ;
  assign n25539 = n7361 ^ n4311 ^ 1'b0 ;
  assign n25540 = n25539 ^ n19092 ^ n6462 ;
  assign n25541 = n25540 ^ n24951 ^ 1'b0 ;
  assign n25542 = n24615 | n25541 ;
  assign n25543 = n3688 ^ n2541 ^ 1'b0 ;
  assign n25544 = n25543 ^ n9321 ^ 1'b0 ;
  assign n25545 = n15666 ^ n9539 ^ 1'b0 ;
  assign n25546 = n25545 ^ n11415 ^ 1'b0 ;
  assign n25547 = ( n1402 & n4204 ) | ( n1402 & n18150 ) | ( n4204 & n18150 ) ;
  assign n25548 = n25547 ^ n20053 ^ 1'b0 ;
  assign n25549 = n9000 & n9939 ;
  assign n25550 = n1017 & ~n25549 ;
  assign n25551 = ( n306 & n20487 ) | ( n306 & n25550 ) | ( n20487 & n25550 ) ;
  assign n25552 = n1825 & ~n25551 ;
  assign n25553 = n8323 ^ n8097 ^ n5796 ;
  assign n25554 = n25553 ^ n6820 ^ 1'b0 ;
  assign n25555 = n12306 & ~n24215 ;
  assign n25556 = ~n2557 & n25555 ;
  assign n25557 = n10372 | n14981 ;
  assign n25558 = n8296 | n25557 ;
  assign n25559 = n4928 ^ n1160 ^ n656 ;
  assign n25560 = n25559 ^ n9258 ^ n6440 ;
  assign n25561 = n1471 & n25560 ;
  assign n25562 = n13726 & n25561 ;
  assign n25563 = n25562 ^ n23217 ^ n19994 ;
  assign n25564 = n6309 | n11266 ;
  assign n25565 = n6968 | n25564 ;
  assign n25566 = n19761 & n25565 ;
  assign n25567 = n17224 ^ n5218 ^ 1'b0 ;
  assign n25568 = n17383 & n25567 ;
  assign n25569 = n12898 & n25568 ;
  assign n25570 = ( n2662 & n6051 ) | ( n2662 & ~n21816 ) | ( n6051 & ~n21816 ) ;
  assign n25571 = n8271 ^ n4624 ^ 1'b0 ;
  assign n25572 = n22862 & ~n25571 ;
  assign n25573 = ( n119 & n9802 ) | ( n119 & ~n25572 ) | ( n9802 & ~n25572 ) ;
  assign n25574 = n22569 ^ n18435 ^ 1'b0 ;
  assign n25575 = n8740 & n25574 ;
  assign n25576 = n17919 ^ n10631 ^ 1'b0 ;
  assign n25577 = n20456 ^ n19810 ^ n10905 ;
  assign n25578 = n25577 ^ n12076 ^ 1'b0 ;
  assign n25579 = n25578 ^ n24502 ^ n9935 ;
  assign n25580 = ~n1556 & n7472 ;
  assign n25581 = n25580 ^ n12090 ^ n9186 ;
  assign n25582 = n7929 & n25581 ;
  assign n25583 = n1153 & ~n19559 ;
  assign n25584 = n25583 ^ n15697 ^ 1'b0 ;
  assign n25585 = n1172 & ~n5102 ;
  assign n25586 = n17432 & n19081 ;
  assign n25587 = n25017 ^ n3404 ^ 1'b0 ;
  assign n25588 = n18133 & ~n25587 ;
  assign n25589 = n8506 & n12575 ;
  assign n25590 = ~n11598 & n25589 ;
  assign n25591 = ( n461 & n5536 ) | ( n461 & ~n12761 ) | ( n5536 & ~n12761 ) ;
  assign n25592 = ( n2999 & n9382 ) | ( n2999 & n25591 ) | ( n9382 & n25591 ) ;
  assign n25593 = n25592 ^ n17110 ^ 1'b0 ;
  assign n25594 = n25590 | n25593 ;
  assign n25595 = ~n18889 & n25594 ;
  assign n25596 = n18252 ^ n5324 ^ n1677 ;
  assign n25597 = ~n1069 & n25596 ;
  assign n25598 = ~n11429 & n25597 ;
  assign n25599 = n5315 & ~n11832 ;
  assign n25600 = n25599 ^ n16305 ^ 1'b0 ;
  assign n25601 = n14255 ^ n11184 ^ 1'b0 ;
  assign n25602 = n2387 | n8117 ;
  assign n25603 = n1543 | n25602 ;
  assign n25604 = ( n8864 & n14586 ) | ( n8864 & n25603 ) | ( n14586 & n25603 ) ;
  assign n25605 = ~n8751 & n24375 ;
  assign n25606 = ~n25604 & n25605 ;
  assign n25607 = n25601 | n25606 ;
  assign n25608 = n25607 ^ n139 ^ 1'b0 ;
  assign n25609 = ( ~n112 & n6036 ) | ( ~n112 & n12771 ) | ( n6036 & n12771 ) ;
  assign n25610 = n14997 ^ n14678 ^ n4708 ;
  assign n25611 = n25610 ^ n20666 ^ n18583 ;
  assign n25612 = n9961 ^ n9589 ^ 1'b0 ;
  assign n25613 = n287 | n25612 ;
  assign n25614 = n25611 & ~n25613 ;
  assign n25615 = n25614 ^ n17450 ^ n4318 ;
  assign n25616 = n8146 & n14441 ;
  assign n25617 = n25616 ^ n809 ^ 1'b0 ;
  assign n25618 = ~n3648 & n25617 ;
  assign n25619 = ~n102 & n11841 ;
  assign n25620 = n25619 ^ n12896 ^ 1'b0 ;
  assign n25621 = n25620 ^ n6739 ^ 1'b0 ;
  assign n25622 = n11796 & n22959 ;
  assign n25623 = n7002 ^ n5898 ^ 1'b0 ;
  assign n25624 = n714 | n17813 ;
  assign n25625 = ~n6784 & n25624 ;
  assign n25626 = n7041 & n25625 ;
  assign n25627 = n25623 & n25626 ;
  assign n25628 = n24869 | n25627 ;
  assign n25629 = n25622 | n25628 ;
  assign n25632 = n7675 ^ n2020 ^ 1'b0 ;
  assign n25633 = n1888 & n25632 ;
  assign n25634 = n25633 ^ n7267 ^ 1'b0 ;
  assign n25635 = n12631 & n25634 ;
  assign n25630 = n18977 ^ n676 ^ 1'b0 ;
  assign n25631 = n25630 ^ n10830 ^ 1'b0 ;
  assign n25636 = n25635 ^ n25631 ^ 1'b0 ;
  assign n25637 = n22377 & n25636 ;
  assign n25638 = n25637 ^ n23295 ^ n2339 ;
  assign n25639 = ( n826 & ~n10110 ) | ( n826 & n17439 ) | ( ~n10110 & n17439 ) ;
  assign n25640 = ~n8325 & n18546 ;
  assign n25641 = ( n1848 & n10424 ) | ( n1848 & ~n25640 ) | ( n10424 & ~n25640 ) ;
  assign n25642 = n7884 ^ n2599 ^ 1'b0 ;
  assign n25643 = n8204 & n25642 ;
  assign n25644 = n2231 | n16882 ;
  assign n25645 = n25644 ^ n19146 ^ 1'b0 ;
  assign n25646 = n25643 & ~n25645 ;
  assign n25647 = n9191 ^ n7303 ^ 1'b0 ;
  assign n25648 = n1623 & n25647 ;
  assign n25649 = n25648 ^ n9823 ^ 1'b0 ;
  assign n25650 = n22813 & n25649 ;
  assign n25651 = ( ~n2470 & n11103 ) | ( ~n2470 & n23767 ) | ( n11103 & n23767 ) ;
  assign n25654 = n1942 | n8824 ;
  assign n25655 = n25654 ^ n14573 ^ 1'b0 ;
  assign n25653 = n19894 ^ n969 ^ 1'b0 ;
  assign n25652 = n5873 & ~n15095 ;
  assign n25656 = n25655 ^ n25653 ^ n25652 ;
  assign n25657 = n1373 & n5040 ;
  assign n25658 = n25657 ^ n10808 ^ 1'b0 ;
  assign n25659 = ( n6217 & n16712 ) | ( n6217 & n25658 ) | ( n16712 & n25658 ) ;
  assign n25660 = ~n6076 & n18973 ;
  assign n25661 = n7985 ^ n3043 ^ 1'b0 ;
  assign n25662 = n7326 ^ n6819 ^ 1'b0 ;
  assign n25663 = ~n4223 & n25662 ;
  assign n25664 = n451 & n25663 ;
  assign n25665 = n18828 ^ n13827 ^ 1'b0 ;
  assign n25666 = ~n25664 & n25665 ;
  assign n25667 = n21119 ^ n10848 ^ 1'b0 ;
  assign n25668 = n20343 | n25667 ;
  assign n25669 = n25668 ^ n24952 ^ 1'b0 ;
  assign n25670 = n6263 | n12554 ;
  assign n25671 = n2606 & n8163 ;
  assign n25672 = n25671 ^ n25413 ^ n8015 ;
  assign n25673 = n5428 & ~n16426 ;
  assign n25674 = n17468 ^ n11740 ^ n1566 ;
  assign n25675 = n25674 ^ n8074 ^ 1'b0 ;
  assign n25676 = n6745 & ~n25675 ;
  assign n25677 = ~n3309 & n4520 ;
  assign n25680 = n1406 & n3654 ;
  assign n25681 = ~n7949 & n25680 ;
  assign n25678 = n10897 & n11172 ;
  assign n25679 = n19756 & n25678 ;
  assign n25682 = n25681 ^ n25679 ^ 1'b0 ;
  assign n25683 = n4549 ^ n283 ^ 1'b0 ;
  assign n25684 = n23369 & ~n25683 ;
  assign n25685 = n1518 | n11218 ;
  assign n25686 = n22477 & ~n25685 ;
  assign n25687 = n25686 ^ n7906 ^ 1'b0 ;
  assign n25688 = ( n1848 & ~n8058 ) | ( n1848 & n14282 ) | ( ~n8058 & n14282 ) ;
  assign n25689 = n25688 ^ n2729 ^ 1'b0 ;
  assign n25690 = n17308 & n25689 ;
  assign n25691 = n2549 & n25690 ;
  assign n25692 = ~n11349 & n14462 ;
  assign n25693 = n22502 | n25496 ;
  assign n25694 = n10141 | n25693 ;
  assign n25695 = ~n1421 & n2135 ;
  assign n25696 = ~n3223 & n25695 ;
  assign n25697 = n22850 ^ n14507 ^ n8849 ;
  assign n25698 = n12641 | n15420 ;
  assign n25699 = n16644 ^ n3987 ^ 1'b0 ;
  assign n25700 = n25698 & ~n25699 ;
  assign n25701 = n22869 ^ n3973 ^ 1'b0 ;
  assign n25702 = n6243 & ~n25701 ;
  assign n25707 = n10391 ^ n4691 ^ 1'b0 ;
  assign n25703 = ~n829 & n17671 ;
  assign n25704 = n25703 ^ n7627 ^ 1'b0 ;
  assign n25705 = n25704 ^ n2917 ^ 1'b0 ;
  assign n25706 = n2868 & n25705 ;
  assign n25708 = n25707 ^ n25706 ^ 1'b0 ;
  assign n25709 = n22104 | n25708 ;
  assign n25710 = n22646 ^ n17355 ^ 1'b0 ;
  assign n25711 = n23676 ^ n5550 ^ 1'b0 ;
  assign n25712 = n15563 ^ n2764 ^ 1'b0 ;
  assign n25713 = n13209 & n25712 ;
  assign n25714 = n25529 ^ n12093 ^ 1'b0 ;
  assign n25715 = n1658 | n13301 ;
  assign n25716 = n12257 | n25715 ;
  assign n25717 = n3918 & n25716 ;
  assign n25718 = n25717 ^ n9479 ^ 1'b0 ;
  assign n25719 = n6600 & ~n22461 ;
  assign n25720 = n25719 ^ x10 ^ 1'b0 ;
  assign n25721 = n6837 ^ n6801 ^ n4526 ;
  assign n25722 = ~n14603 & n25721 ;
  assign n25723 = ~n472 & n12373 ;
  assign n25724 = n2741 & n25723 ;
  assign n25725 = ~n5860 & n13940 ;
  assign n25726 = ~n25724 & n25725 ;
  assign n25727 = ~n7129 & n16922 ;
  assign n25728 = n24936 ^ n11638 ^ n688 ;
  assign n25729 = n3582 | n25728 ;
  assign n25730 = n25727 & ~n25729 ;
  assign n25731 = n9911 & n10743 ;
  assign n25732 = ~n21593 & n25731 ;
  assign n25733 = n25732 ^ n4848 ^ 1'b0 ;
  assign n25735 = n24096 ^ n5552 ^ 1'b0 ;
  assign n25736 = n1956 | n25735 ;
  assign n25734 = n11433 & n15610 ;
  assign n25737 = n25736 ^ n25734 ^ 1'b0 ;
  assign n25738 = n13314 ^ n13067 ^ n3008 ;
  assign n25740 = n458 | n14057 ;
  assign n25741 = ( n574 & ~n8618 ) | ( n574 & n25740 ) | ( ~n8618 & n25740 ) ;
  assign n25739 = n3455 & ~n8426 ;
  assign n25742 = n25741 ^ n25739 ^ 1'b0 ;
  assign n25743 = n8145 & ~n25742 ;
  assign n25744 = n2712 & ~n22809 ;
  assign n25745 = ~n4792 & n15879 ;
  assign n25746 = n3871 | n23780 ;
  assign n25747 = n6093 & ~n25746 ;
  assign n25748 = n25747 ^ n17743 ^ 1'b0 ;
  assign n25749 = ~n5790 & n25748 ;
  assign n25750 = n19986 & n25749 ;
  assign n25751 = n25750 ^ n11724 ^ n5315 ;
  assign n25752 = n22604 ^ n1927 ^ 1'b0 ;
  assign n25753 = n12101 ^ n7193 ^ 1'b0 ;
  assign n25754 = n1999 | n25753 ;
  assign n25755 = n6062 ^ n3162 ^ 1'b0 ;
  assign n25756 = n25755 ^ n4180 ^ 1'b0 ;
  assign n25757 = n12439 | n25756 ;
  assign n25759 = n6643 ^ n1201 ^ 1'b0 ;
  assign n25760 = n5920 & n25759 ;
  assign n25758 = n1766 | n7071 ;
  assign n25761 = n25760 ^ n25758 ^ 1'b0 ;
  assign n25762 = n25761 ^ n20666 ^ n18601 ;
  assign n25763 = n5652 ^ n5631 ^ 1'b0 ;
  assign n25764 = n11668 & ~n25763 ;
  assign n25765 = n7219 ^ n6877 ^ 1'b0 ;
  assign n25766 = ~n10423 & n25765 ;
  assign n25767 = n22558 ^ n645 ^ 1'b0 ;
  assign n25768 = n25767 ^ n13947 ^ n10626 ;
  assign n25769 = n7243 ^ n3620 ^ 1'b0 ;
  assign n25770 = n25769 ^ n4462 ^ 1'b0 ;
  assign n25771 = ~n3658 & n25770 ;
  assign n25772 = ( ~n23982 & n25768 ) | ( ~n23982 & n25771 ) | ( n25768 & n25771 ) ;
  assign n25773 = n2535 | n2579 ;
  assign n25774 = n15579 | n18739 ;
  assign n25775 = ~n4259 & n16178 ;
  assign n25776 = n11356 ^ n7813 ^ 1'b0 ;
  assign n25777 = n25775 | n25776 ;
  assign n25778 = ~n24707 & n25777 ;
  assign n25779 = n11234 | n11906 ;
  assign n25780 = n25779 ^ n4285 ^ 1'b0 ;
  assign n25781 = ~n2627 & n25780 ;
  assign n25782 = ~n2137 & n9454 ;
  assign n25783 = n25782 ^ n8907 ^ 1'b0 ;
  assign n25784 = n21840 | n22651 ;
  assign n25785 = n25784 ^ n5162 ^ 1'b0 ;
  assign n25786 = ( ~n17128 & n25783 ) | ( ~n17128 & n25785 ) | ( n25783 & n25785 ) ;
  assign n25787 = n1540 | n4214 ;
  assign n25788 = ~n1381 & n1948 ;
  assign n25789 = n25788 ^ n13172 ^ 1'b0 ;
  assign n25790 = n25787 | n25789 ;
  assign n25791 = n4450 | n25790 ;
  assign n25792 = n25791 ^ n10122 ^ n4514 ;
  assign n25793 = ( n7104 & n11542 ) | ( n7104 & ~n25792 ) | ( n11542 & ~n25792 ) ;
  assign n25794 = n5456 & n18417 ;
  assign n25795 = ( n3148 & n6835 ) | ( n3148 & n20310 ) | ( n6835 & n20310 ) ;
  assign n25796 = ~n5965 & n25795 ;
  assign n25797 = n25796 ^ n17640 ^ n11042 ;
  assign n25798 = n22151 ^ n12992 ^ 1'b0 ;
  assign n25799 = n2471 & n21132 ;
  assign n25800 = ~n1403 & n25799 ;
  assign n25801 = n25800 ^ n15257 ^ 1'b0 ;
  assign n25802 = n25801 ^ n19360 ^ 1'b0 ;
  assign n25803 = n6774 | n25802 ;
  assign n25804 = n13749 ^ n4260 ^ 1'b0 ;
  assign n25805 = n17085 & n25804 ;
  assign n25806 = ~n19091 & n25805 ;
  assign n25807 = n3224 ^ n2523 ^ 1'b0 ;
  assign n25808 = ~n16116 & n25807 ;
  assign n25809 = n4412 | n17849 ;
  assign n25810 = n25809 ^ n760 ^ 1'b0 ;
  assign n25813 = n14493 | n15759 ;
  assign n25814 = n25813 ^ n14125 ^ n2720 ;
  assign n25811 = n13008 ^ n3495 ^ 1'b0 ;
  assign n25812 = ( n1672 & n3700 ) | ( n1672 & n25811 ) | ( n3700 & n25811 ) ;
  assign n25815 = n25814 ^ n25812 ^ n19355 ;
  assign n25816 = ~n8131 & n19840 ;
  assign n25817 = n25816 ^ n13009 ^ 1'b0 ;
  assign n25818 = n6491 ^ n2805 ^ 1'b0 ;
  assign n25819 = n6027 & n15490 ;
  assign n25820 = ( n10260 & n25818 ) | ( n10260 & n25819 ) | ( n25818 & n25819 ) ;
  assign n25821 = n4396 ^ n149 ^ 1'b0 ;
  assign n25822 = n1569 | n25821 ;
  assign n25823 = n2623 & ~n14462 ;
  assign n25824 = n25822 & n25823 ;
  assign n25825 = n25824 ^ n12852 ^ 1'b0 ;
  assign n25826 = ~n11219 & n25825 ;
  assign n25827 = n9496 & n13225 ;
  assign n25828 = n25827 ^ n3394 ^ 1'b0 ;
  assign n25829 = n4132 | n25828 ;
  assign n25830 = n17162 ^ n5270 ^ 1'b0 ;
  assign n25831 = n25829 | n25830 ;
  assign n25832 = n13991 ^ n7788 ^ 1'b0 ;
  assign n25833 = n2335 ^ n1234 ^ 1'b0 ;
  assign n25834 = ( ~n9851 & n21119 ) | ( ~n9851 & n25833 ) | ( n21119 & n25833 ) ;
  assign n25835 = n447 & ~n718 ;
  assign n25836 = n2696 | n13143 ;
  assign n25837 = n25836 ^ n5022 ^ 1'b0 ;
  assign n25838 = n57 & ~n5538 ;
  assign n25839 = n25838 ^ n2425 ^ 1'b0 ;
  assign n25840 = n18686 & ~n25839 ;
  assign n25841 = n25837 & n25840 ;
  assign n25842 = n5735 & n10369 ;
  assign n25843 = n6462 & n11462 ;
  assign n25844 = n25 | n117 ;
  assign n25845 = n25 & ~n25844 ;
  assign n25846 = n236 & ~n25845 ;
  assign n25847 = n25845 & n25846 ;
  assign n25848 = n107 & ~n1073 ;
  assign n25849 = ~n107 & n25848 ;
  assign n25850 = n1004 & ~n25849 ;
  assign n25851 = n25849 & n25850 ;
  assign n25852 = n20 | n143 ;
  assign n25853 = n20 & ~n25852 ;
  assign n25854 = n25853 ^ n451 ^ 1'b0 ;
  assign n25855 = ~n25851 & n25854 ;
  assign n25856 = ~n13124 & n25855 ;
  assign n25857 = n25847 & n25856 ;
  assign n25858 = n25857 ^ n24891 ^ 1'b0 ;
  assign n25868 = ~n5099 & n6829 ;
  assign n25869 = ~n6829 & n25868 ;
  assign n25870 = n10108 | n25869 ;
  assign n25871 = n25869 & ~n25870 ;
  assign n25859 = n440 | n1936 ;
  assign n25860 = n1936 & ~n25859 ;
  assign n25861 = n237 & ~n25860 ;
  assign n25862 = n25860 & n25861 ;
  assign n25863 = x3 & n254 ;
  assign n25864 = ~x3 & n25863 ;
  assign n25865 = n25862 & ~n25864 ;
  assign n25866 = n4461 & n25865 ;
  assign n25867 = n25866 ^ n14715 ^ 1'b0 ;
  assign n25872 = n25871 ^ n25867 ^ 1'b0 ;
  assign n25873 = n25858 & ~n25872 ;
  assign n25874 = n6053 & ~n6168 ;
  assign n25875 = n6168 & n25874 ;
  assign n25876 = ~n1979 & n25875 ;
  assign n25877 = ( n4918 & ~n5359 ) | ( n4918 & n7774 ) | ( ~n5359 & n7774 ) ;
  assign n25878 = ~n1045 & n25877 ;
  assign n25879 = n25878 ^ n10380 ^ n7343 ;
  assign n25880 = n2405 & ~n18486 ;
  assign n25881 = n8421 ^ n7598 ^ n1628 ;
  assign n25882 = n25881 ^ n17452 ^ n984 ;
  assign n25889 = n11188 ^ n6948 ^ n448 ;
  assign n25888 = ( n4292 & n12311 ) | ( n4292 & ~n19397 ) | ( n12311 & ~n19397 ) ;
  assign n25890 = n25889 ^ n25888 ^ 1'b0 ;
  assign n25883 = n1868 | n13476 ;
  assign n25884 = n25883 ^ n6246 ^ 1'b0 ;
  assign n25885 = n25884 ^ n9376 ^ 1'b0 ;
  assign n25886 = n25885 ^ n16265 ^ n12143 ;
  assign n25887 = ( n4697 & n10952 ) | ( n4697 & n25886 ) | ( n10952 & n25886 ) ;
  assign n25891 = n25890 ^ n25887 ^ n8039 ;
  assign n25893 = n25315 ^ n7969 ^ 1'b0 ;
  assign n25892 = n4835 | n16504 ;
  assign n25894 = n25893 ^ n25892 ^ 1'b0 ;
  assign n25895 = n4271 | n23074 ;
  assign n25896 = n24952 | n25895 ;
  assign n25897 = ~n11260 & n21837 ;
  assign n25898 = n21526 | n25897 ;
  assign n25899 = ~n33 & n24487 ;
  assign n25900 = n5104 & n25899 ;
  assign n25901 = n25900 ^ n6457 ^ 1'b0 ;
  assign n25902 = n23001 & n25901 ;
  assign n25903 = n10321 ^ n8027 ^ 1'b0 ;
  assign n25904 = ( ~n5878 & n9492 ) | ( ~n5878 & n25903 ) | ( n9492 & n25903 ) ;
  assign n25905 = n25904 ^ n3114 ^ 1'b0 ;
  assign n25906 = n4163 & n12165 ;
  assign n25907 = ~n3153 & n25906 ;
  assign n25908 = n25907 ^ n8105 ^ n2432 ;
  assign n25909 = n25908 ^ n17168 ^ 1'b0 ;
  assign n25910 = n386 & n14664 ;
  assign n25911 = n5866 ^ n686 ^ 1'b0 ;
  assign n25912 = n25910 & n25911 ;
  assign n25913 = n25912 ^ n17825 ^ 1'b0 ;
  assign n25914 = n25913 ^ n5327 ^ 1'b0 ;
  assign n25915 = n8746 & ~n11013 ;
  assign n25916 = n25915 ^ n10066 ^ 1'b0 ;
  assign n25917 = n25916 ^ n10930 ^ 1'b0 ;
  assign n25918 = ~n11353 & n25917 ;
  assign n25919 = ~n1930 & n18996 ;
  assign n25921 = n3923 ^ n3471 ^ 1'b0 ;
  assign n25920 = ~n5831 & n9779 ;
  assign n25922 = n25921 ^ n25920 ^ 1'b0 ;
  assign n25923 = ~n25919 & n25922 ;
  assign n25924 = n23294 ^ n9546 ^ 1'b0 ;
  assign n25925 = n18733 ^ n15371 ^ 1'b0 ;
  assign n25926 = n12659 | n25925 ;
  assign n25927 = n9052 ^ n7627 ^ n6222 ;
  assign n25928 = n328 & n25927 ;
  assign n25929 = ~n4948 & n25928 ;
  assign n25930 = n3237 & n19903 ;
  assign n25931 = n13391 ^ n12139 ^ 1'b0 ;
  assign n25932 = n5380 ^ n4663 ^ 1'b0 ;
  assign n25933 = n1815 | n25932 ;
  assign n25934 = ( n607 & ~n873 ) | ( n607 & n2605 ) | ( ~n873 & n2605 ) ;
  assign n25935 = ( n63 & n5537 ) | ( n63 & ~n10095 ) | ( n5537 & ~n10095 ) ;
  assign n25936 = n15405 ^ n6261 ^ 1'b0 ;
  assign n25937 = n25935 & n25936 ;
  assign n25938 = ~n25934 & n25937 ;
  assign n25939 = ~n18639 & n25938 ;
  assign n25940 = n12234 ^ n12034 ^ 1'b0 ;
  assign n25941 = ( n3491 & ~n5495 ) | ( n3491 & n17681 ) | ( ~n5495 & n17681 ) ;
  assign n25942 = n25941 ^ n220 ^ 1'b0 ;
  assign n25943 = n13393 & ~n25942 ;
  assign n25945 = n8463 ^ n4638 ^ 1'b0 ;
  assign n25946 = ~n13354 & n25945 ;
  assign n25944 = n113 & n15142 ;
  assign n25947 = n25946 ^ n25944 ^ 1'b0 ;
  assign n25948 = n17637 ^ n3541 ^ 1'b0 ;
  assign n25949 = n6360 & n25948 ;
  assign n25950 = n18745 ^ n15433 ^ 1'b0 ;
  assign n25951 = n25949 & n25950 ;
  assign n25952 = n17155 & n25951 ;
  assign n25953 = n5732 & ~n10316 ;
  assign n25954 = n4004 & n6142 ;
  assign n25955 = ~n592 & n1600 ;
  assign n25956 = n25955 ^ n6902 ^ n6689 ;
  assign n25957 = ~n9923 & n25956 ;
  assign n25958 = ~n3635 & n7443 ;
  assign n25959 = n25958 ^ n7021 ^ 1'b0 ;
  assign n25960 = ~n11589 & n25959 ;
  assign n25961 = ~n8416 & n25960 ;
  assign n25962 = ~n3869 & n25961 ;
  assign n25963 = n129 & n5088 ;
  assign n25964 = ~n4614 & n25963 ;
  assign n25965 = n25964 ^ n1237 ^ 1'b0 ;
  assign n25966 = n17622 | n24011 ;
  assign n25967 = n13689 | n15014 ;
  assign n25968 = n19503 ^ n5137 ^ 1'b0 ;
  assign n25969 = n25968 ^ n6790 ^ 1'b0 ;
  assign n25970 = n3899 & ~n11430 ;
  assign n25971 = n25970 ^ n8294 ^ n3922 ;
  assign n25972 = n1192 & n25971 ;
  assign n25973 = n1926 & n22862 ;
  assign n25974 = n25973 ^ n11497 ^ 1'b0 ;
  assign n25975 = n22176 | n25974 ;
  assign n25976 = n1650 ^ n1411 ^ n32 ;
  assign n25977 = n13569 ^ n12271 ^ 1'b0 ;
  assign n25978 = n25976 | n25977 ;
  assign n25979 = n19787 ^ n12681 ^ 1'b0 ;
  assign n25980 = n22020 | n25979 ;
  assign n25981 = n21604 | n25980 ;
  assign n25982 = n17496 & n25981 ;
  assign n25983 = ~n6428 & n25982 ;
  assign n25984 = n21182 | n25983 ;
  assign n25985 = ~n3784 & n25984 ;
  assign n25986 = n7774 & n13479 ;
  assign n25987 = n2278 & n25986 ;
  assign n25988 = n25987 ^ n6682 ^ 1'b0 ;
  assign n25995 = n312 & ~n1176 ;
  assign n25989 = ~n1503 & n12135 ;
  assign n25990 = ~n24418 & n25989 ;
  assign n25991 = n14375 & ~n25990 ;
  assign n25992 = n25991 ^ n22814 ^ 1'b0 ;
  assign n25993 = n25992 ^ n11644 ^ 1'b0 ;
  assign n25994 = n7120 & n25993 ;
  assign n25996 = n25995 ^ n25994 ^ 1'b0 ;
  assign n25997 = n20647 & n25996 ;
  assign n25998 = n7118 & n20413 ;
  assign n25999 = n25998 ^ n4948 ^ 1'b0 ;
  assign n26001 = n20805 ^ n8226 ^ n4915 ;
  assign n26000 = n6433 & ~n18294 ;
  assign n26002 = n26001 ^ n26000 ^ 1'b0 ;
  assign n26003 = ~n40 & n1138 ;
  assign n26004 = ~n12169 & n26003 ;
  assign n26005 = n2298 | n2750 ;
  assign n26006 = n26004 & ~n26005 ;
  assign n26007 = n7319 & n18245 ;
  assign n26008 = ~n14462 & n26007 ;
  assign n26009 = ( n10773 & n15687 ) | ( n10773 & n26008 ) | ( n15687 & n26008 ) ;
  assign n26010 = n10053 ^ n2326 ^ n195 ;
  assign n26011 = n2177 & ~n26010 ;
  assign n26012 = n26011 ^ n2433 ^ 1'b0 ;
  assign n26013 = ~n176 & n26012 ;
  assign n26014 = n8584 & ~n14665 ;
  assign n26015 = n26014 ^ n13172 ^ 1'b0 ;
  assign n26016 = n4104 & ~n4689 ;
  assign n26017 = ~n26015 & n26016 ;
  assign n26018 = n26013 & ~n26017 ;
  assign n26019 = ~n5305 & n26018 ;
  assign n26020 = n16797 | n19991 ;
  assign n26021 = n18196 & ~n26020 ;
  assign n26022 = n16922 ^ n5916 ^ 1'b0 ;
  assign n26023 = n14719 | n26022 ;
  assign n26024 = n26023 ^ n6723 ^ 1'b0 ;
  assign n26025 = ~n24417 & n26024 ;
  assign n26026 = n9003 | n17619 ;
  assign n26027 = ( n6771 & n18994 ) | ( n6771 & n26026 ) | ( n18994 & n26026 ) ;
  assign n26028 = n162 | n9827 ;
  assign n26029 = n26028 ^ n2722 ^ 1'b0 ;
  assign n26030 = n18619 ^ n4802 ^ 1'b0 ;
  assign n26031 = ~n15729 & n26030 ;
  assign n26032 = ~n5159 & n23113 ;
  assign n26034 = n16557 ^ n2011 ^ 1'b0 ;
  assign n26033 = n2857 | n7464 ;
  assign n26035 = n26034 ^ n26033 ^ 1'b0 ;
  assign n26036 = ~n25724 & n26035 ;
  assign n26037 = ~n1387 & n22454 ;
  assign n26038 = n26037 ^ n10352 ^ 1'b0 ;
  assign n26039 = n8134 | n26038 ;
  assign n26042 = n523 ^ n166 ^ 1'b0 ;
  assign n26043 = n2022 & n26042 ;
  assign n26044 = n310 & n26043 ;
  assign n26045 = ~n13692 & n26044 ;
  assign n26040 = n5612 & ~n18733 ;
  assign n26041 = n26040 ^ n12830 ^ 1'b0 ;
  assign n26046 = n26045 ^ n26041 ^ 1'b0 ;
  assign n26047 = n14146 & ~n26046 ;
  assign n26048 = n12975 ^ n6704 ^ n481 ;
  assign n26049 = n26048 ^ n14503 ^ 1'b0 ;
  assign n26050 = n7006 & n26049 ;
  assign n26051 = ( n1175 & n2095 ) | ( n1175 & n22085 ) | ( n2095 & n22085 ) ;
  assign n26052 = n2890 & ~n26051 ;
  assign n26053 = n26052 ^ n884 ^ 1'b0 ;
  assign n26054 = n598 | n13199 ;
  assign n26055 = n26053 & ~n26054 ;
  assign n26056 = n18280 & ~n26055 ;
  assign n26057 = n26056 ^ n14290 ^ 1'b0 ;
  assign n26058 = n21853 ^ n11345 ^ 1'b0 ;
  assign n26059 = n533 & ~n26058 ;
  assign n26060 = ( n5935 & ~n6040 ) | ( n5935 & n19886 ) | ( ~n6040 & n19886 ) ;
  assign n26061 = n15382 ^ n12990 ^ 1'b0 ;
  assign n26063 = n344 & ~n771 ;
  assign n26064 = ( n299 & n4620 ) | ( n299 & n20044 ) | ( n4620 & n20044 ) ;
  assign n26065 = n7059 ^ n1471 ^ 1'b0 ;
  assign n26066 = n26064 & n26065 ;
  assign n26067 = ~n26063 & n26066 ;
  assign n26062 = n3119 & n16506 ;
  assign n26068 = n26067 ^ n26062 ^ 1'b0 ;
  assign n26069 = n25232 ^ n21870 ^ n4971 ;
  assign n26070 = ~n12279 & n25093 ;
  assign n26071 = n26070 ^ n17841 ^ 1'b0 ;
  assign n26072 = n802 | n18490 ;
  assign n26073 = n13004 & ~n26072 ;
  assign n26074 = n26073 ^ n2505 ^ 1'b0 ;
  assign n26075 = ~n6490 & n18669 ;
  assign n26077 = ( n1315 & ~n18389 ) | ( n1315 & n20272 ) | ( ~n18389 & n20272 ) ;
  assign n26076 = n4913 | n8376 ;
  assign n26078 = n26077 ^ n26076 ^ 1'b0 ;
  assign n26079 = n4345 & n8640 ;
  assign n26080 = ~n17774 & n26079 ;
  assign n26081 = ~n1853 & n26080 ;
  assign n26082 = ~n2628 & n8203 ;
  assign n26083 = n26082 ^ n17567 ^ 1'b0 ;
  assign n26084 = n2230 & ~n9098 ;
  assign n26085 = n965 & n26084 ;
  assign n26086 = n26085 ^ n14635 ^ n5511 ;
  assign n26087 = n2080 & n13410 ;
  assign n26088 = ~n8054 & n13097 ;
  assign n26089 = n13003 ^ n619 ^ 1'b0 ;
  assign n26090 = n5968 & ~n26089 ;
  assign n26091 = n26088 | n26090 ;
  assign n26092 = n14532 ^ n8471 ^ 1'b0 ;
  assign n26093 = n18286 ^ n18036 ^ 1'b0 ;
  assign n26095 = ~n2795 & n14134 ;
  assign n26096 = ~n4425 & n26095 ;
  assign n26094 = n6919 & ~n14112 ;
  assign n26097 = n26096 ^ n26094 ^ 1'b0 ;
  assign n26098 = ~n26093 & n26097 ;
  assign n26099 = n23443 ^ n21335 ^ n3422 ;
  assign n26100 = ~n7485 & n26099 ;
  assign n26101 = n2488 & n24441 ;
  assign n26102 = n6662 & ~n6819 ;
  assign n26103 = ~n4183 & n26102 ;
  assign n26104 = n21880 ^ n11492 ^ 1'b0 ;
  assign n26105 = n26103 & n26104 ;
  assign n26106 = n25704 | n25922 ;
  assign n26107 = n1378 | n2787 ;
  assign n26108 = n26107 ^ n10477 ^ 1'b0 ;
  assign n26109 = n25182 & ~n26108 ;
  assign n26110 = n26109 ^ n13845 ^ 1'b0 ;
  assign n26111 = n8228 | n26110 ;
  assign n26112 = n19608 ^ n8166 ^ 1'b0 ;
  assign n26113 = n7265 & ~n26112 ;
  assign n26114 = n26113 ^ n7441 ^ 1'b0 ;
  assign n26115 = n20693 ^ n15411 ^ 1'b0 ;
  assign n26116 = n11846 & n19961 ;
  assign n26117 = n2816 & n11222 ;
  assign n26118 = n26117 ^ n19147 ^ 1'b0 ;
  assign n26119 = ~n473 & n1490 ;
  assign n26120 = n18399 & n26119 ;
  assign n26121 = n7935 & ~n22851 ;
  assign n26122 = ~n9504 & n26121 ;
  assign n26123 = n10784 ^ n2382 ^ 1'b0 ;
  assign n26124 = n20436 ^ n3699 ^ 1'b0 ;
  assign n26125 = n9159 & ~n14920 ;
  assign n26126 = n14321 ^ n5051 ^ 1'b0 ;
  assign n26127 = ~n12456 & n26126 ;
  assign n26128 = n26127 ^ n8220 ^ n1463 ;
  assign n26129 = ( n8844 & n11671 ) | ( n8844 & ~n23798 ) | ( n11671 & ~n23798 ) ;
  assign n26134 = n221 & ~n20149 ;
  assign n26135 = ~n23440 & n26134 ;
  assign n26130 = n24441 ^ n7164 ^ n6275 ;
  assign n26131 = n5182 & ~n26130 ;
  assign n26132 = n24927 & n26131 ;
  assign n26133 = n13646 & ~n26132 ;
  assign n26136 = n26135 ^ n26133 ^ 1'b0 ;
  assign n26137 = n2615 & n20671 ;
  assign n26138 = n26137 ^ n23719 ^ 1'b0 ;
  assign n26139 = n25843 ^ n4992 ^ n2297 ;
  assign n26140 = n601 & ~n9374 ;
  assign n26141 = n26140 ^ n12872 ^ 1'b0 ;
  assign n26142 = n5484 & n26141 ;
  assign n26143 = n26142 ^ n20255 ^ 1'b0 ;
  assign n26144 = ( n2030 & n4514 ) | ( n2030 & n11611 ) | ( n4514 & n11611 ) ;
  assign n26145 = n26144 ^ n3832 ^ 1'b0 ;
  assign n26146 = ( ~n3824 & n8149 ) | ( ~n3824 & n26145 ) | ( n8149 & n26145 ) ;
  assign n26147 = n11243 & n13844 ;
  assign n26148 = n26147 ^ n24835 ^ 1'b0 ;
  assign n26149 = n14152 ^ n3016 ^ 1'b0 ;
  assign n26150 = n37 & ~n13199 ;
  assign n26151 = n26149 & n26150 ;
  assign n26152 = ( n2004 & n11132 ) | ( n2004 & n15065 ) | ( n11132 & n15065 ) ;
  assign n26153 = n26151 | n26152 ;
  assign n26154 = n26153 ^ n14426 ^ 1'b0 ;
  assign n26155 = n501 & ~n26154 ;
  assign n26156 = n9075 & ~n22839 ;
  assign n26157 = n23723 ^ n20869 ^ 1'b0 ;
  assign n26158 = n14626 ^ n4114 ^ 1'b0 ;
  assign n26159 = n21482 ^ n3467 ^ 1'b0 ;
  assign n26160 = ~n5617 & n17761 ;
  assign n26161 = ( n12995 & ~n26159 ) | ( n12995 & n26160 ) | ( ~n26159 & n26160 ) ;
  assign n26164 = n4097 ^ n2802 ^ n850 ;
  assign n26163 = n2416 & ~n4318 ;
  assign n26165 = n26164 ^ n26163 ^ 1'b0 ;
  assign n26162 = ( n3387 & n6005 ) | ( n3387 & ~n6430 ) | ( n6005 & ~n6430 ) ;
  assign n26166 = n26165 ^ n26162 ^ 1'b0 ;
  assign n26167 = n24065 ^ n318 ^ 1'b0 ;
  assign n26168 = n23858 ^ n9971 ^ 1'b0 ;
  assign n26169 = ~n778 & n26168 ;
  assign n26170 = n21146 & n26161 ;
  assign n26171 = ( n8185 & ~n12644 ) | ( n8185 & n20061 ) | ( ~n12644 & n20061 ) ;
  assign n26172 = n26171 ^ n24770 ^ n24010 ;
  assign n26173 = n5725 & n17287 ;
  assign n26174 = n9750 & ~n14926 ;
  assign n26175 = n101 & n26174 ;
  assign n26176 = n21679 & ~n26175 ;
  assign n26177 = n26176 ^ n23841 ^ 1'b0 ;
  assign n26178 = n7352 | n26177 ;
  assign n26179 = n8157 & ~n25260 ;
  assign n26180 = ( ~n1866 & n6168 ) | ( ~n1866 & n26179 ) | ( n6168 & n26179 ) ;
  assign n26181 = ( n369 & n11209 ) | ( n369 & ~n11614 ) | ( n11209 & ~n11614 ) ;
  assign n26182 = n205 | n6292 ;
  assign n26183 = n6069 | n26182 ;
  assign n26184 = n4702 | n26183 ;
  assign n26185 = n483 & n4199 ;
  assign n26186 = n4340 & ~n26185 ;
  assign n26187 = ( ~n6785 & n11271 ) | ( ~n6785 & n16620 ) | ( n11271 & n16620 ) ;
  assign n26188 = n2605 & ~n26187 ;
  assign n26189 = n17459 ^ n13689 ^ 1'b0 ;
  assign n26190 = n26189 ^ n19991 ^ 1'b0 ;
  assign n26191 = n6687 ^ n835 ^ 1'b0 ;
  assign n26192 = n25445 | n26191 ;
  assign n26193 = n26192 ^ n24168 ^ n13594 ;
  assign n26194 = n11440 ^ n1006 ^ 1'b0 ;
  assign n26195 = n17149 & ~n26194 ;
  assign n26196 = n26195 ^ n4072 ^ n1071 ;
  assign n26197 = ~n6255 & n21837 ;
  assign n26198 = ~n6273 & n26197 ;
  assign n26199 = ~n8607 & n12135 ;
  assign n26200 = n26199 ^ n2677 ^ 1'b0 ;
  assign n26201 = n10659 ^ n3353 ^ 1'b0 ;
  assign n26204 = n2617 & ~n11204 ;
  assign n26202 = n3883 & ~n5571 ;
  assign n26203 = n26202 ^ n4932 ^ 1'b0 ;
  assign n26205 = n26204 ^ n26203 ^ n5473 ;
  assign n26206 = n26205 ^ n5099 ^ 1'b0 ;
  assign n26207 = n25494 | n26206 ;
  assign n26208 = n26207 ^ n4410 ^ 1'b0 ;
  assign n26209 = n4454 | n8591 ;
  assign n26210 = n10420 & n19275 ;
  assign n26211 = n10408 ^ n2664 ^ 1'b0 ;
  assign n26212 = n26210 & n26211 ;
  assign n26213 = n22290 ^ n14813 ^ 1'b0 ;
  assign n26214 = n22080 ^ n2211 ^ 1'b0 ;
  assign n26215 = ~n945 & n1826 ;
  assign n26216 = n26215 ^ n874 ^ 1'b0 ;
  assign n26217 = n26216 ^ n15674 ^ 1'b0 ;
  assign n26218 = n4220 ^ n1312 ^ 1'b0 ;
  assign n26219 = ( n6454 & n7225 ) | ( n6454 & ~n26218 ) | ( n7225 & ~n26218 ) ;
  assign n26221 = n2083 ^ n1172 ^ 1'b0 ;
  assign n26220 = n12567 ^ n2403 ^ 1'b0 ;
  assign n26222 = n26221 ^ n26220 ^ 1'b0 ;
  assign n26223 = n26219 | n26222 ;
  assign n26231 = n12680 ^ n5673 ^ 1'b0 ;
  assign n26232 = ~n8638 & n18498 ;
  assign n26233 = ~n16641 & n26232 ;
  assign n26234 = n26233 ^ n19755 ^ 1'b0 ;
  assign n26235 = n26231 & ~n26234 ;
  assign n26229 = n20044 ^ n10798 ^ 1'b0 ;
  assign n26226 = ( n12131 & ~n15145 ) | ( n12131 & n17784 ) | ( ~n15145 & n17784 ) ;
  assign n26224 = n3082 & n5070 ;
  assign n26225 = n11247 | n26224 ;
  assign n26227 = n26226 ^ n26225 ^ 1'b0 ;
  assign n26228 = n26227 ^ n21473 ^ 1'b0 ;
  assign n26230 = n26229 ^ n26228 ^ 1'b0 ;
  assign n26236 = n26235 ^ n26230 ^ 1'b0 ;
  assign n26237 = n7655 | n26236 ;
  assign n26238 = n3193 & ~n12995 ;
  assign n26239 = n21543 & n26238 ;
  assign n26240 = n3181 & n6868 ;
  assign n26241 = ~n1616 & n26240 ;
  assign n26242 = n6488 ^ n4683 ^ 1'b0 ;
  assign n26243 = n19620 & ~n26242 ;
  assign n26244 = ~n1591 & n26243 ;
  assign n26245 = n9020 & n26244 ;
  assign n26246 = ( n3912 & ~n14470 ) | ( n3912 & n26245 ) | ( ~n14470 & n26245 ) ;
  assign n26247 = n24866 & n26246 ;
  assign n26248 = ( n19193 & n26241 ) | ( n19193 & ~n26247 ) | ( n26241 & ~n26247 ) ;
  assign n26249 = ~n5832 & n14646 ;
  assign n26250 = n26249 ^ n6337 ^ 1'b0 ;
  assign n26251 = ( n7089 & ~n23893 ) | ( n7089 & n24024 ) | ( ~n23893 & n24024 ) ;
  assign n26252 = n16897 ^ n10549 ^ 1'b0 ;
  assign n26253 = n10668 & ~n26252 ;
  assign n26254 = n18210 & ~n26253 ;
  assign n26255 = ~n26251 & n26254 ;
  assign n26256 = n16556 ^ n14646 ^ 1'b0 ;
  assign n26257 = n19458 | n26256 ;
  assign n26258 = n16156 & n26257 ;
  assign n26259 = ( ~n6049 & n7215 ) | ( ~n6049 & n17381 ) | ( n7215 & n17381 ) ;
  assign n26260 = n204 | n26259 ;
  assign n26261 = n5504 | n26260 ;
  assign n26262 = n19270 | n26261 ;
  assign n26263 = n26262 ^ n7125 ^ 1'b0 ;
  assign n26264 = n5830 | n26263 ;
  assign n26265 = n6107 & n7125 ;
  assign n26266 = n26265 ^ n11924 ^ 1'b0 ;
  assign n26267 = n3564 | n26266 ;
  assign n26268 = n15687 | n26267 ;
  assign n26269 = ~n12138 & n26268 ;
  assign n26270 = ~n15919 & n17680 ;
  assign n26271 = n26270 ^ n777 ^ 1'b0 ;
  assign n26272 = n26271 ^ n6147 ^ 1'b0 ;
  assign n26273 = n13559 & ~n26272 ;
  assign n26274 = n21213 ^ n19146 ^ 1'b0 ;
  assign n26275 = ~n6091 & n26274 ;
  assign n26276 = n15906 & n17530 ;
  assign n26277 = n13561 & ~n26276 ;
  assign n26278 = n5732 ^ n4990 ^ 1'b0 ;
  assign n26279 = ( n2653 & n26277 ) | ( n2653 & n26278 ) | ( n26277 & n26278 ) ;
  assign n26280 = n26279 ^ n886 ^ 1'b0 ;
  assign n26281 = n12763 & n26280 ;
  assign n26282 = n11445 & n22988 ;
  assign n26283 = n10973 & n26282 ;
  assign n26284 = n536 ^ n85 ^ 1'b0 ;
  assign n26285 = ~n15276 & n26284 ;
  assign n26286 = n8886 ^ n8616 ^ n8226 ;
  assign n26287 = n6867 ^ n6128 ^ 1'b0 ;
  assign n26288 = n26287 ^ n15772 ^ n8595 ;
  assign n26289 = n26288 ^ n20960 ^ n9161 ;
  assign n26290 = ( n4405 & ~n26286 ) | ( n4405 & n26289 ) | ( ~n26286 & n26289 ) ;
  assign n26291 = n22669 ^ n558 ^ 1'b0 ;
  assign n26292 = ~n5420 & n26291 ;
  assign n26293 = n19525 ^ n3824 ^ 1'b0 ;
  assign n26294 = ( n18270 & ~n19090 ) | ( n18270 & n23662 ) | ( ~n19090 & n23662 ) ;
  assign n26295 = n26 | n26294 ;
  assign n26296 = n7915 ^ n6951 ^ 1'b0 ;
  assign n26297 = n1553 & n26296 ;
  assign n26298 = n3976 & n8610 ;
  assign n26299 = n26298 ^ n6911 ^ 1'b0 ;
  assign n26300 = ~n26297 & n26299 ;
  assign n26301 = n26300 ^ n17185 ^ n4188 ;
  assign n26302 = n4559 ^ n1243 ^ 1'b0 ;
  assign n26303 = ~n21076 & n26302 ;
  assign n26304 = ~n6775 & n26303 ;
  assign n26305 = n12219 & ~n23363 ;
  assign n26306 = n21652 ^ n10479 ^ 1'b0 ;
  assign n26307 = n4258 & n26306 ;
  assign n26308 = n26305 & n26307 ;
  assign n26309 = n9659 & n16588 ;
  assign n26310 = ( n777 & ~n4804 ) | ( n777 & n15420 ) | ( ~n4804 & n15420 ) ;
  assign n26311 = ~n4298 & n8389 ;
  assign n26312 = n4298 & n26311 ;
  assign n26313 = n26310 | n26312 ;
  assign n26314 = ~n20715 & n26313 ;
  assign n26315 = n26314 ^ n12169 ^ 1'b0 ;
  assign n26316 = n6602 ^ n4743 ^ n2805 ;
  assign n26317 = n4508 & n26316 ;
  assign n26318 = n25135 & ~n26317 ;
  assign n26319 = n6005 ^ n4127 ^ 1'b0 ;
  assign n26320 = n26319 ^ n3175 ^ 1'b0 ;
  assign n26321 = n18027 ^ n3059 ^ 1'b0 ;
  assign n26322 = n4239 & ~n26321 ;
  assign n26323 = n21073 & n22422 ;
  assign n26324 = n26323 ^ n3408 ^ 1'b0 ;
  assign n26325 = ~n18290 & n18880 ;
  assign n26326 = n22317 ^ n11880 ^ 1'b0 ;
  assign n26327 = n14507 ^ n8801 ^ 1'b0 ;
  assign n26328 = ~n4289 & n26327 ;
  assign n26329 = n26328 ^ n18601 ^ 1'b0 ;
  assign n26330 = n1264 | n26329 ;
  assign n26331 = ( ~n2731 & n18093 ) | ( ~n2731 & n20125 ) | ( n18093 & n20125 ) ;
  assign n26332 = n5272 & ~n16522 ;
  assign n26333 = n23860 ^ n19135 ^ n2568 ;
  assign n26334 = n17734 ^ n10372 ^ 1'b0 ;
  assign n26335 = n9598 | n26334 ;
  assign n26336 = n77 & ~n26335 ;
  assign n26337 = n2144 & ~n19258 ;
  assign n26338 = n26337 ^ n3945 ^ 1'b0 ;
  assign n26339 = n12920 ^ n4330 ^ 1'b0 ;
  assign n26340 = n18164 & n26339 ;
  assign n26341 = n4852 | n6441 ;
  assign n26342 = n356 & n1064 ;
  assign n26343 = ~n4207 & n26342 ;
  assign n26344 = n7417 ^ n3009 ^ 1'b0 ;
  assign n26345 = ~n8211 & n26344 ;
  assign n26346 = n26345 ^ n15563 ^ 1'b0 ;
  assign n26347 = n11288 | n26346 ;
  assign n26348 = n7502 | n26347 ;
  assign n26349 = n3109 | n10587 ;
  assign n26350 = n16058 ^ n3959 ^ n882 ;
  assign n26351 = ( ~n3469 & n25897 ) | ( ~n3469 & n26350 ) | ( n25897 & n26350 ) ;
  assign n26352 = n498 | n6316 ;
  assign n26353 = n26352 ^ n17369 ^ 1'b0 ;
  assign n26354 = n26029 ^ n11615 ^ 1'b0 ;
  assign n26355 = ~n1175 & n26354 ;
  assign n26356 = n13903 ^ n7898 ^ 1'b0 ;
  assign n26357 = n1244 ^ n592 ^ 1'b0 ;
  assign n26358 = n19518 | n26357 ;
  assign n26359 = n26356 | n26358 ;
  assign n26360 = ~n4141 & n13524 ;
  assign n26361 = ~n10820 & n26360 ;
  assign n26362 = ~n21810 & n26361 ;
  assign n26364 = n5953 & ~n13493 ;
  assign n26365 = n1613 & n26364 ;
  assign n26366 = n2627 & ~n11786 ;
  assign n26367 = ( ~n342 & n2131 ) | ( ~n342 & n26366 ) | ( n2131 & n26366 ) ;
  assign n26368 = n26367 ^ n12249 ^ 1'b0 ;
  assign n26369 = ~n26365 & n26368 ;
  assign n26363 = n23483 ^ n134 ^ 1'b0 ;
  assign n26370 = n26369 ^ n26363 ^ n14386 ;
  assign n26371 = n4009 ^ n756 ^ 1'b0 ;
  assign n26372 = n20740 ^ n6731 ^ 1'b0 ;
  assign n26373 = n9324 | n26372 ;
  assign n26374 = n5987 | n26373 ;
  assign n26375 = n26374 ^ n9108 ^ 1'b0 ;
  assign n26376 = ~n26371 & n26375 ;
  assign n26377 = ( n13071 & n13758 ) | ( n13071 & ~n26376 ) | ( n13758 & ~n26376 ) ;
  assign n26378 = n14961 ^ n1992 ^ 1'b0 ;
  assign n26379 = n26378 ^ n5904 ^ 1'b0 ;
  assign n26380 = n3222 | n26379 ;
  assign n26381 = n24736 ^ n4226 ^ 1'b0 ;
  assign n26382 = n25706 ^ n7150 ^ 1'b0 ;
  assign n26383 = n11772 & n26382 ;
  assign n26384 = n13069 ^ n7001 ^ 1'b0 ;
  assign n26385 = n6579 & n26384 ;
  assign n26386 = n10094 & n19405 ;
  assign n26387 = n26386 ^ n9933 ^ 1'b0 ;
  assign n26388 = n1412 | n22864 ;
  assign n26389 = n7249 ^ n5303 ^ n3353 ;
  assign n26390 = n11288 ^ n8294 ^ 1'b0 ;
  assign n26391 = n5791 | n26390 ;
  assign n26392 = ( n11859 & n26389 ) | ( n11859 & n26391 ) | ( n26389 & n26391 ) ;
  assign n26393 = ~n7505 & n26392 ;
  assign n26394 = n26393 ^ n2230 ^ n717 ;
  assign n26395 = n12548 ^ n953 ^ 1'b0 ;
  assign n26396 = n26395 ^ n14999 ^ 1'b0 ;
  assign n26397 = ~n1654 & n8341 ;
  assign n26398 = n10679 & n26397 ;
  assign n26399 = n4675 & n9583 ;
  assign n26400 = n10360 | n16116 ;
  assign n26401 = ~n23729 & n26400 ;
  assign n26402 = ~n11988 & n19273 ;
  assign n26403 = n24063 ^ n6131 ^ 1'b0 ;
  assign n26404 = n14267 & ~n26403 ;
  assign n26405 = n4251 & ~n26404 ;
  assign n26406 = n11927 ^ n6067 ^ 1'b0 ;
  assign n26407 = n13963 & n26406 ;
  assign n26408 = n6039 & n11021 ;
  assign n26409 = n5845 ^ n3943 ^ n350 ;
  assign n26410 = n26409 ^ n22970 ^ 1'b0 ;
  assign n26411 = n4629 & ~n15259 ;
  assign n26412 = ~n26410 & n26411 ;
  assign n26413 = n26408 | n26412 ;
  assign n26414 = n26407 | n26413 ;
  assign n26415 = n9436 ^ n9149 ^ n1775 ;
  assign n26416 = n5855 | n11239 ;
  assign n26417 = ~n1625 & n25254 ;
  assign n26418 = n26417 ^ n11107 ^ 1'b0 ;
  assign n26419 = n9027 ^ n541 ^ 1'b0 ;
  assign n26420 = n22008 & n23005 ;
  assign n26421 = n40 | n121 ;
  assign n26422 = n3805 & n7653 ;
  assign n26423 = n26421 & n26422 ;
  assign n26424 = n8029 & n16059 ;
  assign n26425 = n6205 | n15702 ;
  assign n26426 = n26425 ^ n9479 ^ 1'b0 ;
  assign n26427 = n11134 ^ n423 ^ 1'b0 ;
  assign n26428 = ~n26426 & n26427 ;
  assign n26429 = n26428 ^ n764 ^ 1'b0 ;
  assign n26430 = n26424 & ~n26429 ;
  assign n26431 = n17343 & ~n20720 ;
  assign n26432 = n17576 & n26431 ;
  assign n26433 = n3423 & n15338 ;
  assign n26434 = n26433 ^ n1391 ^ 1'b0 ;
  assign n26435 = n10263 & ~n26434 ;
  assign n26436 = n26435 ^ n12213 ^ 1'b0 ;
  assign n26437 = ( n6249 & n12164 ) | ( n6249 & ~n14508 ) | ( n12164 & ~n14508 ) ;
  assign n26438 = n26437 ^ n13755 ^ 1'b0 ;
  assign n26439 = ( n11072 & n20073 ) | ( n11072 & ~n26438 ) | ( n20073 & ~n26438 ) ;
  assign n26440 = ( n7069 & n7641 ) | ( n7069 & ~n14392 ) | ( n7641 & ~n14392 ) ;
  assign n26441 = ( n361 & n6259 ) | ( n361 & n26440 ) | ( n6259 & n26440 ) ;
  assign n26442 = n26441 ^ n20021 ^ 1'b0 ;
  assign n26443 = n23335 ^ n15784 ^ 1'b0 ;
  assign n26444 = n3989 & ~n26443 ;
  assign n26445 = ~n1050 & n5223 ;
  assign n26450 = n13037 ^ n5022 ^ 1'b0 ;
  assign n26446 = n5298 | n7644 ;
  assign n26447 = n5083 ^ n4291 ^ 1'b0 ;
  assign n26448 = n2019 | n26447 ;
  assign n26449 = n26446 & ~n26448 ;
  assign n26451 = n26450 ^ n26449 ^ 1'b0 ;
  assign n26452 = ( ~n40 & n12916 ) | ( ~n40 & n26451 ) | ( n12916 & n26451 ) ;
  assign n26453 = n2511 | n10564 ;
  assign n26454 = n192 & n19229 ;
  assign n26455 = ~n26453 & n26454 ;
  assign n26457 = n10465 ^ n3167 ^ n345 ;
  assign n26456 = n110 & n8621 ;
  assign n26458 = n26457 ^ n26456 ^ 1'b0 ;
  assign n26459 = n19698 & ~n26458 ;
  assign n26460 = n7896 | n19322 ;
  assign n26461 = n21081 ^ n4366 ^ n2925 ;
  assign n26462 = ~n3060 & n26461 ;
  assign n26463 = n1359 & ~n13567 ;
  assign n26464 = n26463 ^ n1068 ^ 1'b0 ;
  assign n26465 = ( n16787 & n18679 ) | ( n16787 & n22097 ) | ( n18679 & n22097 ) ;
  assign n26466 = n18386 ^ n5061 ^ 1'b0 ;
  assign n26467 = ~n3554 & n26466 ;
  assign n26468 = n26465 & ~n26467 ;
  assign n26469 = n510 & n7365 ;
  assign n26470 = n26469 ^ n20970 ^ 1'b0 ;
  assign n26471 = n17731 ^ n13561 ^ 1'b0 ;
  assign n26475 = n5840 ^ n2640 ^ 1'b0 ;
  assign n26476 = n5774 & n26475 ;
  assign n26472 = ~n665 & n899 ;
  assign n26473 = n7543 & n26472 ;
  assign n26474 = n26473 ^ n19348 ^ n6278 ;
  assign n26477 = n26476 ^ n26474 ^ 1'b0 ;
  assign n26478 = n17574 & ~n26477 ;
  assign n26479 = n2694 & n25289 ;
  assign n26480 = ~n25953 & n26479 ;
  assign n26481 = n9687 ^ n7903 ^ 1'b0 ;
  assign n26482 = n14290 & n21316 ;
  assign n26483 = n6983 & n22684 ;
  assign n26484 = n11671 & n26483 ;
  assign n26485 = n26482 | n26484 ;
  assign n26486 = n1156 | n26485 ;
  assign n26487 = n15157 & n15607 ;
  assign n26488 = ~n20353 & n26487 ;
  assign n26489 = n1293 & n16337 ;
  assign n26490 = n26489 ^ n791 ^ 1'b0 ;
  assign n26491 = n5264 & ~n26490 ;
  assign n26492 = n1900 & n2021 ;
  assign n26493 = n26492 ^ n6574 ^ 1'b0 ;
  assign n26495 = n2797 & ~n24696 ;
  assign n26494 = ~n4602 & n23529 ;
  assign n26496 = n26495 ^ n26494 ^ 1'b0 ;
  assign n26497 = n10127 | n26496 ;
  assign n26498 = n14523 & ~n26497 ;
  assign n26499 = n5212 ^ n4427 ^ 1'b0 ;
  assign n26500 = n19778 ^ n13270 ^ n5657 ;
  assign n26501 = ( n5550 & n8154 ) | ( n5550 & n25738 ) | ( n8154 & n25738 ) ;
  assign n26502 = n13865 | n17306 ;
  assign n26503 = n9060 ^ n711 ^ 1'b0 ;
  assign n26504 = n13112 ^ n12303 ^ n2606 ;
  assign n26505 = n6664 | n26504 ;
  assign n26506 = n9736 & n14008 ;
  assign n26507 = n26505 & n26506 ;
  assign n26508 = ~n5384 & n23200 ;
  assign n26509 = ~n23200 & n26508 ;
  assign n26510 = n13758 ^ n9336 ^ 1'b0 ;
  assign n26511 = n26510 ^ n26132 ^ n18319 ;
  assign n26512 = n7298 & n10910 ;
  assign n26513 = n26512 ^ n8884 ^ 1'b0 ;
  assign n26514 = n8903 | n26513 ;
  assign n26515 = n19727 & ~n26514 ;
  assign n26516 = n20471 ^ n2460 ^ 1'b0 ;
  assign n26517 = n20598 ^ n5712 ^ 1'b0 ;
  assign n26518 = ~n7596 & n26517 ;
  assign n26519 = n7308 | n26518 ;
  assign n26520 = n250 | n25677 ;
  assign n26521 = n16539 | n26520 ;
  assign n26522 = n3309 & ~n8122 ;
  assign n26523 = ~n17755 & n26522 ;
  assign n26524 = ~n51 & n7378 ;
  assign n26525 = ~n7378 & n26524 ;
  assign n26526 = ~n3951 & n10676 ;
  assign n26527 = ~n686 & n26526 ;
  assign n26528 = n26525 & n26527 ;
  assign n26529 = n15964 & n26528 ;
  assign n26530 = n14445 | n19602 ;
  assign n26531 = n8476 | n26530 ;
  assign n26532 = x7 & ~n879 ;
  assign n26533 = n4222 & n26532 ;
  assign n26534 = n26533 ^ n23152 ^ n1000 ;
  assign n26535 = n686 | n26106 ;
  assign n26536 = n26535 ^ n5867 ^ 1'b0 ;
  assign n26537 = n4886 ^ n1147 ^ 1'b0 ;
  assign n26538 = n848 & n26537 ;
  assign n26539 = n26538 ^ n22123 ^ 1'b0 ;
  assign n26540 = n8912 & ~n20792 ;
  assign n26541 = n26540 ^ n1182 ^ 1'b0 ;
  assign n26542 = ~n100 & n8341 ;
  assign n26543 = n26542 ^ n809 ^ 1'b0 ;
  assign n26544 = n14893 ^ n990 ^ 1'b0 ;
  assign n26545 = n491 & n7776 ;
  assign n26546 = n26545 ^ n2230 ^ 1'b0 ;
  assign n26547 = n15969 ^ n10684 ^ 1'b0 ;
  assign n26548 = ~n6415 & n26547 ;
  assign n26549 = ( n2933 & n5212 ) | ( n2933 & ~n26548 ) | ( n5212 & ~n26548 ) ;
  assign n26550 = n18519 ^ n9656 ^ 1'b0 ;
  assign n26553 = n12433 ^ n5838 ^ 1'b0 ;
  assign n26551 = n13467 | n15865 ;
  assign n26552 = n532 | n26551 ;
  assign n26554 = n26553 ^ n26552 ^ 1'b0 ;
  assign n26555 = n9309 ^ n6337 ^ 1'b0 ;
  assign n26556 = ~n3229 & n26555 ;
  assign n26557 = ~n15932 & n22876 ;
  assign n26558 = ~n2827 & n18061 ;
  assign n26559 = n1875 & n26558 ;
  assign n26560 = n12220 ^ n11680 ^ n3120 ;
  assign n26561 = n10885 | n15320 ;
  assign n26562 = n26561 ^ n3066 ^ 1'b0 ;
  assign n26563 = ( ~n1751 & n4102 ) | ( ~n1751 & n12540 ) | ( n4102 & n12540 ) ;
  assign n26564 = n2943 ^ n263 ^ 1'b0 ;
  assign n26565 = ~n26563 & n26564 ;
  assign n26566 = n11155 ^ n8067 ^ n1940 ;
  assign n26567 = n23747 & n26566 ;
  assign n26568 = n10756 ^ n8418 ^ 1'b0 ;
  assign n26569 = n5908 & ~n26568 ;
  assign n26570 = n26569 ^ n2606 ^ 1'b0 ;
  assign n26571 = n9809 & ~n16556 ;
  assign n26572 = n3792 | n26571 ;
  assign n26573 = n1599 & ~n1681 ;
  assign n26574 = ( ~n5394 & n18221 ) | ( ~n5394 & n26573 ) | ( n18221 & n26573 ) ;
  assign n26575 = n3870 | n17505 ;
  assign n26584 = n2725 | n7400 ;
  assign n26585 = n20092 & n26584 ;
  assign n26586 = ~n20448 & n26585 ;
  assign n26583 = n25620 ^ n3717 ^ 1'b0 ;
  assign n26580 = n8338 ^ n3582 ^ 1'b0 ;
  assign n26581 = n18406 & ~n26580 ;
  assign n26577 = ~n19201 & n24307 ;
  assign n26578 = n26577 ^ n6471 ^ 1'b0 ;
  assign n26576 = n24485 ^ n18709 ^ n13643 ;
  assign n26579 = n26578 ^ n26576 ^ 1'b0 ;
  assign n26582 = n26581 ^ n26579 ^ n21381 ;
  assign n26587 = n26586 ^ n26583 ^ n26582 ;
  assign n26588 = n26211 ^ n22314 ^ n18804 ;
  assign n26589 = n14729 & ~n26588 ;
  assign n26590 = n26589 ^ n8158 ^ 1'b0 ;
  assign n26591 = n5227 & n9093 ;
  assign n26592 = ~n3049 & n26591 ;
  assign n26593 = ~n181 & n19687 ;
  assign n26594 = ~n3473 & n4262 ;
  assign n26595 = n26594 ^ n225 ^ 1'b0 ;
  assign n26596 = n24380 ^ n3818 ^ 1'b0 ;
  assign n26597 = ( n45 & ~n26595 ) | ( n45 & n26596 ) | ( ~n26595 & n26596 ) ;
  assign n26598 = n15089 | n15346 ;
  assign n26599 = n9014 & ~n26598 ;
  assign n26600 = ( n2421 & n19081 ) | ( n2421 & n26599 ) | ( n19081 & n26599 ) ;
  assign n26601 = n16357 ^ n2526 ^ 1'b0 ;
  assign n26602 = ( n15772 & ~n26600 ) | ( n15772 & n26601 ) | ( ~n26600 & n26601 ) ;
  assign n26603 = n1339 & n15903 ;
  assign n26604 = n17266 | n26603 ;
  assign n26605 = n26604 ^ n14771 ^ 1'b0 ;
  assign n26606 = ~n10625 & n20137 ;
  assign n26607 = n26606 ^ n20417 ^ 1'b0 ;
  assign n26608 = n9715 ^ n2945 ^ 1'b0 ;
  assign n26609 = ~n10516 & n26608 ;
  assign n26610 = n26609 ^ n19867 ^ 1'b0 ;
  assign n26611 = n2145 & ~n3179 ;
  assign n26612 = n442 | n4782 ;
  assign n26613 = n26612 ^ n19209 ^ 1'b0 ;
  assign n26614 = ~n26611 & n26613 ;
  assign n26615 = ~n7342 & n26614 ;
  assign n26616 = ~n12963 & n26615 ;
  assign n26617 = n6458 & ~n9811 ;
  assign n26618 = n26617 ^ n849 ^ 1'b0 ;
  assign n26619 = n26618 ^ n25047 ^ n7937 ;
  assign n26620 = n21503 | n26619 ;
  assign n26621 = n4490 ^ n1942 ^ 1'b0 ;
  assign n26622 = n26621 ^ n25325 ^ 1'b0 ;
  assign n26623 = n26620 | n26622 ;
  assign n26624 = n3406 ^ n3241 ^ 1'b0 ;
  assign n26625 = n26624 ^ n20672 ^ 1'b0 ;
  assign n26626 = n19450 & n26625 ;
  assign n26627 = n23861 ^ n19705 ^ n181 ;
  assign n26628 = n7516 & n13684 ;
  assign n26630 = n750 & ~n8519 ;
  assign n26629 = n2682 & n7932 ;
  assign n26631 = n26630 ^ n26629 ^ 1'b0 ;
  assign n26632 = n14508 & n26631 ;
  assign n26633 = n26632 ^ n11938 ^ 1'b0 ;
  assign n26634 = ~n26628 & n26633 ;
  assign n26635 = n5768 ^ n1953 ^ 1'b0 ;
  assign n26636 = n26635 ^ n9086 ^ n1409 ;
  assign n26637 = n9360 & ~n17162 ;
  assign n26638 = n10684 & n26637 ;
  assign n26639 = ~n1213 & n26638 ;
  assign n26640 = n9385 & ~n26220 ;
  assign n26641 = ~n11502 & n23270 ;
  assign n26642 = n21549 ^ n9124 ^ 1'b0 ;
  assign n26643 = n26642 ^ n13876 ^ n6143 ;
  assign n26644 = n26641 & n26643 ;
  assign n26645 = n13595 ^ n12591 ^ 1'b0 ;
  assign n26647 = n9511 ^ n7788 ^ 1'b0 ;
  assign n26648 = n2065 | n26647 ;
  assign n26646 = ~n9076 & n19791 ;
  assign n26649 = n26648 ^ n26646 ^ 1'b0 ;
  assign n26650 = n20819 ^ n3918 ^ n1155 ;
  assign n26651 = n1650 & ~n13351 ;
  assign n26652 = n24934 & n26651 ;
  assign n26653 = n26652 ^ n15919 ^ 1'b0 ;
  assign n26654 = n7707 ^ n4156 ^ n2180 ;
  assign n26655 = n4330 & n26654 ;
  assign n26656 = n8411 ^ n945 ^ 1'b0 ;
  assign n26657 = n23882 ^ n2418 ^ 1'b0 ;
  assign n26658 = n13943 | n19322 ;
  assign n26659 = n26657 & ~n26658 ;
  assign n26660 = n10218 ^ n7864 ^ 1'b0 ;
  assign n26661 = n11134 ^ n10785 ^ 1'b0 ;
  assign n26662 = n16549 & ~n26661 ;
  assign n26663 = ( n10689 & n26049 ) | ( n10689 & ~n26662 ) | ( n26049 & ~n26662 ) ;
  assign n26674 = n7377 ^ n3537 ^ 1'b0 ;
  assign n26669 = n21552 ^ n115 ^ 1'b0 ;
  assign n26670 = n25363 ^ n6821 ^ 1'b0 ;
  assign n26671 = n26669 & n26670 ;
  assign n26672 = n26671 ^ n11140 ^ n4331 ;
  assign n26668 = n21190 ^ n11274 ^ 1'b0 ;
  assign n26673 = n26672 ^ n26668 ^ n16963 ;
  assign n26664 = n1332 | n1516 ;
  assign n26665 = n11429 & ~n18875 ;
  assign n26666 = n15274 | n26665 ;
  assign n26667 = n26664 & ~n26666 ;
  assign n26675 = n26674 ^ n26673 ^ n26667 ;
  assign n26676 = n10180 ^ n780 ^ 1'b0 ;
  assign n26677 = n8480 & ~n26676 ;
  assign n26678 = n16274 ^ n15796 ^ 1'b0 ;
  assign n26679 = n26677 & ~n26678 ;
  assign n26680 = n5673 ^ n3114 ^ 1'b0 ;
  assign n26681 = n26680 ^ n18841 ^ 1'b0 ;
  assign n26682 = ~n1052 & n5781 ;
  assign n26683 = n26682 ^ n19826 ^ 1'b0 ;
  assign n26684 = n16166 & ~n26683 ;
  assign n26685 = n26684 ^ n2628 ^ 1'b0 ;
  assign n26686 = ~n23802 & n26685 ;
  assign n26687 = n26686 ^ n3202 ^ 1'b0 ;
  assign n26688 = n14730 & ~n25312 ;
  assign n26689 = n2494 ^ n1529 ^ 1'b0 ;
  assign n26690 = n26688 | n26689 ;
  assign n26691 = n26251 & n26690 ;
  assign n26692 = ( n2544 & ~n7485 ) | ( n2544 & n12589 ) | ( ~n7485 & n12589 ) ;
  assign n26694 = x2 & ~n22227 ;
  assign n26693 = n15345 ^ n13735 ^ 1'b0 ;
  assign n26695 = n26694 ^ n26693 ^ n7326 ;
  assign n26696 = n401 & n6049 ;
  assign n26697 = n26696 ^ n16190 ^ 1'b0 ;
  assign n26698 = n9147 & n14151 ;
  assign n26699 = n4454 & n26698 ;
  assign n26700 = n25624 ^ n2534 ^ 1'b0 ;
  assign n26701 = n15373 ^ n4387 ^ 1'b0 ;
  assign n26702 = n32 | n26701 ;
  assign n26703 = n23021 ^ n879 ^ 1'b0 ;
  assign n26704 = n23946 & n26703 ;
  assign n26705 = ( ~n2926 & n7572 ) | ( ~n2926 & n16678 ) | ( n7572 & n16678 ) ;
  assign n26706 = n2056 | n4937 ;
  assign n26707 = n26705 & ~n26706 ;
  assign n26719 = ~n7753 & n12780 ;
  assign n26720 = n16342 & ~n26719 ;
  assign n26721 = n9634 | n26720 ;
  assign n26722 = n18048 & ~n26721 ;
  assign n26708 = n3298 ^ n744 ^ 1'b0 ;
  assign n26709 = ( ~n9905 & n17793 ) | ( ~n9905 & n26708 ) | ( n17793 & n26708 ) ;
  assign n26715 = n9951 & n14512 ;
  assign n26710 = n4903 & n11725 ;
  assign n26711 = ( ~n2966 & n11194 ) | ( ~n2966 & n12880 ) | ( n11194 & n12880 ) ;
  assign n26712 = n8009 ^ n2466 ^ 1'b0 ;
  assign n26713 = n26711 & n26712 ;
  assign n26714 = ~n26710 & n26713 ;
  assign n26716 = n26715 ^ n26714 ^ 1'b0 ;
  assign n26717 = n26709 & ~n26716 ;
  assign n26718 = ~n10574 & n26717 ;
  assign n26723 = n26722 ^ n26718 ^ 1'b0 ;
  assign n26726 = ~n7221 & n21563 ;
  assign n26727 = n26726 ^ n1875 ^ 1'b0 ;
  assign n26724 = n7736 ^ n7483 ^ n1610 ;
  assign n26725 = n14593 & ~n26724 ;
  assign n26728 = n26727 ^ n26725 ^ 1'b0 ;
  assign n26729 = n926 ^ n115 ^ 1'b0 ;
  assign n26730 = n26729 ^ n4632 ^ 1'b0 ;
  assign n26731 = n17605 ^ n11402 ^ 1'b0 ;
  assign n26732 = n4093 & ~n26731 ;
  assign n26733 = n24110 & n26732 ;
  assign n26734 = n18664 & ~n26733 ;
  assign n26735 = n26734 ^ n18245 ^ 1'b0 ;
  assign n26736 = n7672 & ~n22514 ;
  assign n26737 = n1897 & n12046 ;
  assign n26739 = n15213 ^ n2650 ^ 1'b0 ;
  assign n26740 = n5848 & ~n26739 ;
  assign n26738 = n15119 & n23650 ;
  assign n26741 = n26740 ^ n26738 ^ 1'b0 ;
  assign n26742 = n26741 ^ n16882 ^ 1'b0 ;
  assign n26743 = ~n26737 & n26742 ;
  assign n26744 = n18330 ^ n9014 ^ 1'b0 ;
  assign n26745 = n26744 ^ n12642 ^ 1'b0 ;
  assign n26746 = ~n7154 & n22433 ;
  assign n26747 = n1553 & n26746 ;
  assign n26748 = n3786 & n5679 ;
  assign n26749 = ~n3786 & n26748 ;
  assign n26750 = n26749 ^ n26694 ^ 1'b0 ;
  assign n26751 = n10417 & n26750 ;
  assign n26752 = n26751 ^ n17407 ^ 1'b0 ;
  assign n26753 = n6491 ^ n43 ^ 1'b0 ;
  assign n26754 = n8755 | n26753 ;
  assign n26755 = n26754 ^ n9879 ^ n4717 ;
  assign n26756 = n20462 ^ n6638 ^ 1'b0 ;
  assign n26757 = n19731 & n26756 ;
  assign n26758 = n8681 | n23217 ;
  assign n26759 = n9036 ^ n6720 ^ n249 ;
  assign n26760 = n8086 & n10388 ;
  assign n26761 = ~n26759 & n26760 ;
  assign n26762 = n2953 & n10077 ;
  assign n26763 = n26762 ^ n16210 ^ 1'b0 ;
  assign n26764 = n26679 ^ n11697 ^ 1'b0 ;
  assign n26765 = n16187 ^ n12142 ^ n6470 ;
  assign n26766 = n9487 | n13932 ;
  assign n26767 = n6743 ^ n2928 ^ 1'b0 ;
  assign n26768 = n877 & ~n26767 ;
  assign n26769 = ~n26766 & n26768 ;
  assign n26770 = n24565 ^ n22839 ^ n16932 ;
  assign n26771 = n15595 & n18674 ;
  assign n26772 = ( n16156 & n23005 ) | ( n16156 & n26771 ) | ( n23005 & n26771 ) ;
  assign n26773 = n5042 ^ n3221 ^ 1'b0 ;
  assign n26774 = ~n19973 & n26773 ;
  assign n26775 = n1080 ^ n1040 ^ 1'b0 ;
  assign n26776 = n26775 ^ n20475 ^ n4273 ;
  assign n26777 = ~n7356 & n26776 ;
  assign n26778 = n7114 & n26777 ;
  assign n26779 = ( n2130 & ~n3964 ) | ( n2130 & n22657 ) | ( ~n3964 & n22657 ) ;
  assign n26780 = n26778 | n26779 ;
  assign n26782 = n13941 & n17736 ;
  assign n26783 = ~n15654 & n26782 ;
  assign n26781 = n62 | n801 ;
  assign n26784 = n26783 ^ n26781 ^ 1'b0 ;
  assign n26785 = ~n2697 & n6766 ;
  assign n26786 = n16829 & n26785 ;
  assign n26787 = n7790 | n26786 ;
  assign n26788 = n14158 & ~n26787 ;
  assign n26789 = ( n4207 & n15534 ) | ( n4207 & n16025 ) | ( n15534 & n16025 ) ;
  assign n26790 = n230 & ~n2339 ;
  assign n26791 = ( ~n1551 & n26789 ) | ( ~n1551 & n26790 ) | ( n26789 & n26790 ) ;
  assign n26792 = n1228 & n3307 ;
  assign n26793 = n26792 ^ n18594 ^ 1'b0 ;
  assign n26794 = ( n20921 & n21323 ) | ( n20921 & ~n26144 ) | ( n21323 & ~n26144 ) ;
  assign n26795 = ~n6014 & n14866 ;
  assign n26796 = n25163 & ~n26795 ;
  assign n26797 = n7554 | n13860 ;
  assign n26798 = n26797 ^ n434 ^ 1'b0 ;
  assign n26799 = n26798 ^ n15720 ^ 1'b0 ;
  assign n26800 = n13784 ^ n5809 ^ 1'b0 ;
  assign n26802 = n11555 & n22597 ;
  assign n26801 = ~n1064 & n21050 ;
  assign n26803 = n26802 ^ n26801 ^ 1'b0 ;
  assign n26804 = n1088 & n19224 ;
  assign n26805 = ~n2216 & n26804 ;
  assign n26806 = n26805 ^ n6581 ^ 1'b0 ;
  assign n26807 = ( n1143 & ~n2327 ) | ( n1143 & n16944 ) | ( ~n2327 & n16944 ) ;
  assign n26809 = ~n816 & n9036 ;
  assign n26810 = n8604 & ~n26809 ;
  assign n26811 = n350 | n3855 ;
  assign n26812 = n26810 & ~n26811 ;
  assign n26808 = n1082 & ~n3772 ;
  assign n26813 = n26812 ^ n26808 ^ 1'b0 ;
  assign n26814 = n10958 ^ n10018 ^ 1'b0 ;
  assign n26815 = n12095 | n26814 ;
  assign n26816 = n19520 & n20552 ;
  assign n26817 = n26815 & n26816 ;
  assign n26818 = ~n3096 & n8414 ;
  assign n26822 = n192 & n6871 ;
  assign n26820 = n9869 ^ n5702 ^ 1'b0 ;
  assign n26819 = ~n1223 & n16870 ;
  assign n26821 = n26820 ^ n26819 ^ 1'b0 ;
  assign n26823 = n26822 ^ n26821 ^ n23956 ;
  assign n26824 = n26823 ^ n25726 ^ 1'b0 ;
  assign n26826 = n2999 ^ n2192 ^ 1'b0 ;
  assign n26827 = n7195 | n26826 ;
  assign n26828 = n26827 ^ n17630 ^ n8442 ;
  assign n26825 = ~n6556 & n6759 ;
  assign n26829 = n26828 ^ n26825 ^ 1'b0 ;
  assign n26830 = n1840 | n2337 ;
  assign n26831 = n26830 ^ n8753 ^ 1'b0 ;
  assign n26832 = n26831 ^ n6632 ^ 1'b0 ;
  assign n26833 = n5684 & ~n6505 ;
  assign n26834 = n26833 ^ n10788 ^ 1'b0 ;
  assign n26835 = n6590 & ~n13151 ;
  assign n26836 = n26835 ^ n14848 ^ 1'b0 ;
  assign n26837 = n26836 ^ n10266 ^ n10252 ;
  assign n26838 = n7168 ^ n1105 ^ 1'b0 ;
  assign n26839 = n26837 | n26838 ;
  assign n26840 = n4165 & ~n23220 ;
  assign n26841 = n9995 & n26840 ;
  assign n26842 = n5919 & n25010 ;
  assign n26843 = n26841 & n26842 ;
  assign n26844 = ~n9667 & n14397 ;
  assign n26845 = n6727 & n26844 ;
  assign n26846 = n205 | n26845 ;
  assign n26847 = n26846 ^ n5867 ^ 1'b0 ;
  assign n26848 = n5197 ^ n3679 ^ 1'b0 ;
  assign n26849 = n11934 & n26848 ;
  assign n26851 = n1460 & ~n5965 ;
  assign n26852 = n26851 ^ n6644 ^ 1'b0 ;
  assign n26853 = n26852 ^ n10826 ^ n7240 ;
  assign n26850 = n14338 & ~n19189 ;
  assign n26854 = n26853 ^ n26850 ^ n14914 ;
  assign n26855 = n26849 & n26854 ;
  assign n26857 = ( n13769 & n16989 ) | ( n13769 & ~n25289 ) | ( n16989 & ~n25289 ) ;
  assign n26856 = n4681 & n6376 ;
  assign n26858 = n26857 ^ n26856 ^ 1'b0 ;
  assign n26859 = n16910 ^ n5817 ^ 1'b0 ;
  assign n26860 = n26859 ^ n6104 ^ n1457 ;
  assign n26861 = n12590 | n14150 ;
  assign n26862 = n26860 & ~n26861 ;
  assign n26863 = n7586 | n19638 ;
  assign n26864 = n26863 ^ n19787 ^ 1'b0 ;
  assign n26865 = n26864 ^ n25678 ^ n1818 ;
  assign n26866 = n11320 ^ n9145 ^ n2657 ;
  assign n26867 = n4733 & ~n23836 ;
  assign n26868 = n26867 ^ n22292 ^ 1'b0 ;
  assign n26869 = n21892 & ~n26868 ;
  assign n26870 = n26869 ^ n5982 ^ 1'b0 ;
  assign n26871 = n8395 & n19569 ;
  assign n26872 = n10897 ^ n3189 ^ 1'b0 ;
  assign n26873 = n14470 & ~n26872 ;
  assign n26874 = n25879 ^ n8127 ^ 1'b0 ;
  assign n26875 = n1951 | n2266 ;
  assign n26876 = ( n6199 & ~n15315 ) | ( n6199 & n26875 ) | ( ~n15315 & n26875 ) ;
  assign n26877 = n15103 ^ n1081 ^ 1'b0 ;
  assign n26881 = n14076 | n26094 ;
  assign n26882 = n26881 ^ n12168 ^ 1'b0 ;
  assign n26878 = n2631 | n8039 ;
  assign n26879 = n26878 ^ n22040 ^ 1'b0 ;
  assign n26880 = n20417 | n26879 ;
  assign n26883 = n26882 ^ n26880 ^ 1'b0 ;
  assign n26884 = n12893 ^ n6384 ^ 1'b0 ;
  assign n26885 = ( n20772 & n23837 ) | ( n20772 & n26884 ) | ( n23837 & n26884 ) ;
  assign n26886 = n26754 ^ n11064 ^ 1'b0 ;
  assign n26887 = n26886 ^ n25741 ^ n17897 ;
  assign n26888 = n24329 ^ n18695 ^ n5948 ;
  assign n26889 = n26888 ^ n8895 ^ 1'b0 ;
  assign n26890 = n5053 | n8612 ;
  assign n26891 = n8612 & ~n26890 ;
  assign n26892 = n15009 & ~n26891 ;
  assign n26896 = n4570 & n5818 ;
  assign n26897 = ~n4570 & n26896 ;
  assign n26898 = n8302 & ~n26897 ;
  assign n26899 = n26897 & n26898 ;
  assign n26900 = n2130 & ~n26899 ;
  assign n26901 = ~n2130 & n26900 ;
  assign n26902 = n1408 & n7977 ;
  assign n26903 = ~n1408 & n26902 ;
  assign n26904 = ~n19891 & n26903 ;
  assign n26905 = n26901 | n26904 ;
  assign n26893 = n3285 | n26088 ;
  assign n26894 = n26088 & ~n26893 ;
  assign n26895 = n6745 & ~n26894 ;
  assign n26906 = n26905 ^ n26895 ^ 1'b0 ;
  assign n26907 = n26892 & ~n26906 ;
  assign n26908 = x1 & n17956 ;
  assign n26909 = n25239 ^ n18835 ^ 1'b0 ;
  assign n26910 = n20031 ^ n7697 ^ 1'b0 ;
  assign n26911 = n1050 & ~n26910 ;
  assign n26912 = n26911 ^ n7011 ^ 1'b0 ;
  assign n26913 = n26912 ^ n3268 ^ 1'b0 ;
  assign n26914 = n26913 ^ n4434 ^ 1'b0 ;
  assign n26915 = ~n26909 & n26914 ;
  assign n26916 = ~n4549 & n9511 ;
  assign n26917 = n24028 & n26916 ;
  assign n26918 = ( n10424 & ~n23680 ) | ( n10424 & n26917 ) | ( ~n23680 & n26917 ) ;
  assign n26919 = ( n1380 & ~n6895 ) | ( n1380 & n18938 ) | ( ~n6895 & n18938 ) ;
  assign n26920 = ~n15604 & n22101 ;
  assign n26921 = n6191 & n26920 ;
  assign n26922 = ~n10390 & n26921 ;
  assign n26923 = n481 | n4846 ;
  assign n26924 = n26923 ^ n18622 ^ n498 ;
  assign n26925 = ( n4247 & n21848 ) | ( n4247 & ~n26924 ) | ( n21848 & ~n26924 ) ;
  assign n26926 = n16522 ^ n14052 ^ 1'b0 ;
  assign n26927 = n26926 ^ n21654 ^ 1'b0 ;
  assign n26928 = n3309 | n4446 ;
  assign n26929 = n13771 ^ n1311 ^ 1'b0 ;
  assign n26930 = n26929 ^ n1484 ^ 1'b0 ;
  assign n26931 = n26930 ^ n23426 ^ 1'b0 ;
  assign n26932 = n10654 | n16510 ;
  assign n26933 = n26932 ^ n25637 ^ 1'b0 ;
  assign n26934 = n36 | n5554 ;
  assign n26935 = n22942 & ~n26934 ;
  assign n26936 = ( n6302 & n8633 ) | ( n6302 & ~n14067 ) | ( n8633 & ~n14067 ) ;
  assign n26937 = n8392 ^ n5597 ^ 1'b0 ;
  assign n26938 = n12046 ^ n9027 ^ 1'b0 ;
  assign n26939 = ~n6660 & n16589 ;
  assign n26940 = ~n9013 & n10329 ;
  assign n26941 = ( n1979 & n9751 ) | ( n1979 & ~n26940 ) | ( n9751 & ~n26940 ) ;
  assign n26942 = n26941 ^ n1545 ^ 1'b0 ;
  assign n26943 = n8247 & ~n26942 ;
  assign n26944 = n2751 & n4153 ;
  assign n26945 = n18548 | n26944 ;
  assign n26946 = n26945 ^ n11921 ^ 1'b0 ;
  assign n26947 = n8480 | n26946 ;
  assign n26948 = n11896 & ~n26947 ;
  assign n26949 = n15486 | n24907 ;
  assign n26950 = n5461 ^ n4878 ^ 1'b0 ;
  assign n26951 = n1138 | n26950 ;
  assign n26952 = n9517 | n26951 ;
  assign n26953 = n13769 ^ n3245 ^ 1'b0 ;
  assign n26954 = n1694 & n26953 ;
  assign n26955 = n14188 ^ n11249 ^ n4667 ;
  assign n26956 = n18074 | n18876 ;
  assign n26957 = n25785 ^ n6754 ^ 1'b0 ;
  assign n26958 = ~n26956 & n26957 ;
  assign n26959 = n3877 | n14880 ;
  assign n26960 = n26959 ^ n11700 ^ 1'b0 ;
  assign n26961 = n1439 & ~n19721 ;
  assign n26962 = n26961 ^ n19928 ^ 1'b0 ;
  assign n26963 = n3906 & n15878 ;
  assign n26964 = n26963 ^ n22230 ^ 1'b0 ;
  assign n26965 = n2044 & n9494 ;
  assign n26966 = n9795 & ~n9904 ;
  assign n26967 = n7251 | n26966 ;
  assign n26968 = n8404 & ~n26967 ;
  assign n26969 = n26336 ^ n7408 ^ 1'b0 ;
  assign n26970 = ~n2192 & n2677 ;
  assign n26971 = n22394 ^ n8165 ^ 1'b0 ;
  assign n26972 = n26971 ^ n24585 ^ n11575 ;
  assign n26973 = n4927 & ~n20995 ;
  assign n26974 = n26972 & n26973 ;
  assign n26981 = n4533 & n21321 ;
  assign n26982 = n26981 ^ n26391 ^ 1'b0 ;
  assign n26975 = n1395 & n7272 ;
  assign n26976 = n4205 & ~n14475 ;
  assign n26977 = n20781 ^ n2254 ^ 1'b0 ;
  assign n26978 = ( n26266 & n26976 ) | ( n26266 & ~n26977 ) | ( n26976 & ~n26977 ) ;
  assign n26979 = n26975 | n26978 ;
  assign n26980 = n11490 & ~n26979 ;
  assign n26983 = n26982 ^ n26980 ^ 1'b0 ;
  assign n26984 = n16182 & n19185 ;
  assign n26985 = n26983 & n26984 ;
  assign n26986 = ~n12606 & n21138 ;
  assign n26987 = n26986 ^ n1433 ^ 1'b0 ;
  assign n26988 = n21914 ^ n19920 ^ 1'b0 ;
  assign n26989 = n8073 ^ n3696 ^ 1'b0 ;
  assign n26990 = n4638 & ~n26989 ;
  assign n26991 = n26990 ^ n21849 ^ 1'b0 ;
  assign n26992 = n8644 | n16601 ;
  assign n26993 = ( n21163 & n24624 ) | ( n21163 & ~n26992 ) | ( n24624 & ~n26992 ) ;
  assign n26994 = n1664 & ~n12304 ;
  assign n26995 = ~n10990 & n26994 ;
  assign n26996 = n17661 & n26995 ;
  assign n26997 = n26996 ^ n4551 ^ n1248 ;
  assign n26999 = x2 & n6893 ;
  assign n27000 = ~n328 & n26999 ;
  assign n26998 = ~n2114 & n17290 ;
  assign n27001 = n27000 ^ n26998 ^ 1'b0 ;
  assign n27002 = n8799 & n27001 ;
  assign n27003 = n27002 ^ n15024 ^ 1'b0 ;
  assign n27004 = n27003 ^ n15876 ^ 1'b0 ;
  assign n27005 = n26997 | n27004 ;
  assign n27006 = n22511 & ~n27005 ;
  assign n27007 = ~n1841 & n2589 ;
  assign n27008 = n27007 ^ n12701 ^ 1'b0 ;
  assign n27009 = n766 & n27008 ;
  assign n27010 = ( ~n3919 & n4897 ) | ( ~n3919 & n25455 ) | ( n4897 & n25455 ) ;
  assign n27011 = n12551 ^ n9524 ^ n6189 ;
  assign n27012 = n27011 ^ n7657 ^ 1'b0 ;
  assign n27013 = n80 | n1114 ;
  assign n27014 = n22929 & ~n26720 ;
  assign n27015 = n27014 ^ n11988 ^ 1'b0 ;
  assign n27016 = n9732 | n25076 ;
  assign n27017 = n25076 & ~n27016 ;
  assign n27018 = n27017 ^ n16274 ^ 1'b0 ;
  assign n27019 = n3739 & ~n8397 ;
  assign n27020 = ~n26618 & n27019 ;
  assign n27021 = n27020 ^ n16816 ^ 1'b0 ;
  assign n27022 = n22507 | n27021 ;
  assign n27023 = n7860 | n11736 ;
  assign n27024 = n27022 & ~n27023 ;
  assign n27025 = n27024 ^ n18433 ^ 1'b0 ;
  assign n27026 = n27018 & n27025 ;
  assign n27027 = n25366 ^ n11393 ^ 1'b0 ;
  assign n27028 = n4700 & ~n23088 ;
  assign n27029 = n5353 | n6019 ;
  assign n27030 = n17687 & ~n27029 ;
  assign n27031 = n21740 & n27030 ;
  assign n27032 = n8593 ^ n77 ^ 1'b0 ;
  assign n27033 = n22698 ^ n9211 ^ 1'b0 ;
  assign n27034 = ( ~n8470 & n25790 ) | ( ~n8470 & n27033 ) | ( n25790 & n27033 ) ;
  assign n27035 = n20735 ^ n543 ^ 1'b0 ;
  assign n27036 = n27035 ^ n11872 ^ n8470 ;
  assign n27037 = n20106 ^ n3159 ^ 1'b0 ;
  assign n27038 = n10883 & ~n27037 ;
  assign n27046 = n1575 ^ n1125 ^ n879 ;
  assign n27047 = n9758 & n27046 ;
  assign n27048 = n27047 ^ n13796 ^ 1'b0 ;
  assign n27049 = n8183 & n27048 ;
  assign n27050 = n2549 & n27049 ;
  assign n27040 = ~n1986 & n19580 ;
  assign n27039 = n4526 | n14273 ;
  assign n27041 = n27040 ^ n27039 ^ 1'b0 ;
  assign n27042 = n11249 ^ n4635 ^ 1'b0 ;
  assign n27043 = n27041 & n27042 ;
  assign n27044 = n27043 ^ n11633 ^ n4804 ;
  assign n27045 = ~n1235 & n27044 ;
  assign n27051 = n27050 ^ n27045 ^ 1'b0 ;
  assign n27052 = n20756 ^ n6220 ^ 1'b0 ;
  assign n27053 = n21048 & ~n27052 ;
  assign n27054 = n14172 & n26470 ;
  assign n27055 = n27054 ^ n18254 ^ 1'b0 ;
  assign n27056 = n9213 & n13025 ;
  assign n27057 = n27056 ^ n18324 ^ n3840 ;
  assign n27058 = ( n5068 & ~n15850 ) | ( n5068 & n24191 ) | ( ~n15850 & n24191 ) ;
  assign n27065 = n136 & n780 ;
  assign n27066 = n27065 ^ n2196 ^ 1'b0 ;
  assign n27067 = n27066 ^ n5581 ^ 1'b0 ;
  assign n27068 = ~n7151 & n27067 ;
  assign n27062 = ~n711 & n5724 ;
  assign n27063 = n4595 & n27062 ;
  assign n27064 = ~n8789 & n27063 ;
  assign n27059 = n12678 ^ n1129 ^ 1'b0 ;
  assign n27060 = n27059 ^ n4307 ^ 1'b0 ;
  assign n27061 = ~n13965 & n27060 ;
  assign n27069 = n27068 ^ n27064 ^ n27061 ;
  assign n27070 = n27069 ^ n19004 ^ 1'b0 ;
  assign n27077 = n13972 ^ n6925 ^ 1'b0 ;
  assign n27078 = n2509 & n27077 ;
  assign n27071 = n3205 & n12327 ;
  assign n27072 = n4617 & n27071 ;
  assign n27073 = n1664 & ~n27072 ;
  assign n27074 = n6272 & n27073 ;
  assign n27075 = n27074 ^ n3868 ^ 1'b0 ;
  assign n27076 = n7873 | n27075 ;
  assign n27079 = n27078 ^ n27076 ^ n1389 ;
  assign n27080 = n9206 ^ n3909 ^ 1'b0 ;
  assign n27081 = n27079 | n27080 ;
  assign n27082 = n10125 & n27081 ;
  assign n27083 = n9755 & ~n10592 ;
  assign n27084 = n27083 ^ n9634 ^ 1'b0 ;
  assign n27085 = n16935 ^ n16452 ^ n3888 ;
  assign n27086 = n361 | n8373 ;
  assign n27087 = n27085 | n27086 ;
  assign n27088 = ( n23654 & n26805 ) | ( n23654 & ~n27087 ) | ( n26805 & ~n27087 ) ;
  assign n27089 = n652 & n10204 ;
  assign n27090 = n20693 ^ n14860 ^ 1'b0 ;
  assign n27091 = n20205 ^ n7435 ^ 1'b0 ;
  assign n27092 = n11053 | n12937 ;
  assign n27093 = ~n6768 & n27092 ;
  assign n27094 = n27093 ^ n9983 ^ 1'b0 ;
  assign n27095 = n26077 ^ n3753 ^ 1'b0 ;
  assign n27096 = ( ~n1526 & n2021 ) | ( ~n1526 & n7584 ) | ( n2021 & n7584 ) ;
  assign n27097 = n7080 & n27096 ;
  assign n27098 = n4258 & ~n27097 ;
  assign n27099 = ~n5392 & n27098 ;
  assign n27100 = n7084 ^ n4548 ^ 1'b0 ;
  assign n27101 = ( n12153 & n25549 ) | ( n12153 & n27100 ) | ( n25549 & n27100 ) ;
  assign n27102 = n27101 ^ n17394 ^ 1'b0 ;
  assign n27110 = n3070 ^ n2142 ^ 1'b0 ;
  assign n27111 = n1577 & n27110 ;
  assign n27112 = ( n126 & ~n11968 ) | ( n126 & n27111 ) | ( ~n11968 & n27111 ) ;
  assign n27103 = n6940 ^ n6925 ^ 1'b0 ;
  assign n27105 = n5750 & ~n9839 ;
  assign n27104 = n5725 & ~n21424 ;
  assign n27106 = n27105 ^ n27104 ^ 1'b0 ;
  assign n27107 = n27103 | n27106 ;
  assign n27108 = n15228 ^ n10267 ^ 1'b0 ;
  assign n27109 = ~n27107 & n27108 ;
  assign n27113 = n27112 ^ n27109 ^ 1'b0 ;
  assign n27114 = n11443 & ~n16400 ;
  assign n27115 = n27114 ^ n23016 ^ 1'b0 ;
  assign n27124 = n2360 & ~n5987 ;
  assign n27125 = n7796 & n27124 ;
  assign n27121 = n7322 & n20413 ;
  assign n27122 = ~n4622 & n27121 ;
  assign n27117 = n8678 ^ n3810 ^ n2802 ;
  assign n27118 = n1940 & ~n27117 ;
  assign n27119 = ~n4413 & n27118 ;
  assign n27116 = n4717 & ~n5517 ;
  assign n27120 = n27119 ^ n27116 ^ 1'b0 ;
  assign n27123 = n27122 ^ n27120 ^ 1'b0 ;
  assign n27126 = n27125 ^ n27123 ^ 1'b0 ;
  assign n27128 = n4296 | n9279 ;
  assign n27127 = ~n9704 & n12810 ;
  assign n27129 = n27128 ^ n27127 ^ 1'b0 ;
  assign n27130 = n21550 ^ n2622 ^ 1'b0 ;
  assign n27131 = n16527 | n27130 ;
  assign n27132 = ( ~n2281 & n11120 ) | ( ~n2281 & n11914 ) | ( n11120 & n11914 ) ;
  assign n27133 = n11642 ^ n654 ^ 1'b0 ;
  assign n27134 = n8500 ^ n6647 ^ 1'b0 ;
  assign n27135 = n24361 & ~n27134 ;
  assign n27136 = ~n5954 & n6471 ;
  assign n27137 = n1207 | n27136 ;
  assign n27138 = n27135 | n27137 ;
  assign n27139 = n647 & n27138 ;
  assign n27140 = ~n5240 & n27139 ;
  assign n27141 = n5678 | n22087 ;
  assign n27142 = n24268 & ~n27141 ;
  assign n27143 = n12823 & n27142 ;
  assign n27144 = ~n17698 & n27143 ;
  assign n27145 = n5997 ^ n4328 ^ 1'b0 ;
  assign n27146 = n5897 | n27145 ;
  assign n27147 = n9829 & ~n18403 ;
  assign n27148 = n7288 | n27147 ;
  assign n27149 = n1766 & n2039 ;
  assign n27150 = n5361 & n15889 ;
  assign n27151 = ~n27149 & n27150 ;
  assign n27152 = n8638 & n10507 ;
  assign n27153 = n1048 | n21373 ;
  assign n27154 = n7927 | n27153 ;
  assign n27155 = n15850 & n21240 ;
  assign n27156 = n27155 ^ n26566 ^ 1'b0 ;
  assign n27157 = n21131 & ~n27156 ;
  assign n27158 = n10745 & n27157 ;
  assign n27159 = n6557 ^ n5348 ^ 1'b0 ;
  assign n27160 = ~n18378 & n27159 ;
  assign n27161 = n22130 ^ n15430 ^ 1'b0 ;
  assign n27162 = n27161 ^ n20658 ^ n5554 ;
  assign n27163 = n22362 ^ n10264 ^ 1'b0 ;
  assign n27164 = ( n1800 & n5729 ) | ( n1800 & n27163 ) | ( n5729 & n27163 ) ;
  assign n27166 = n12486 & n13682 ;
  assign n27167 = n27166 ^ n395 ^ 1'b0 ;
  assign n27168 = ( n7508 & n21471 ) | ( n7508 & ~n27167 ) | ( n21471 & ~n27167 ) ;
  assign n27165 = n11387 | n21178 ;
  assign n27169 = n27168 ^ n27165 ^ 1'b0 ;
  assign n27170 = n9251 ^ n3381 ^ 1'b0 ;
  assign n27171 = n586 & ~n27170 ;
  assign n27172 = n27171 ^ n4269 ^ 1'b0 ;
  assign n27173 = n9049 | n27172 ;
  assign n27174 = ~n11134 & n17559 ;
  assign n27175 = ~n478 & n27174 ;
  assign n27176 = n78 | n18505 ;
  assign n27177 = n9583 | n27176 ;
  assign n27178 = n1540 | n2909 ;
  assign n27179 = n18831 & n27178 ;
  assign n27180 = ~n6939 & n27179 ;
  assign n27181 = n1974 & ~n27180 ;
  assign n27182 = n27181 ^ n16379 ^ 1'b0 ;
  assign n27183 = ~n27177 & n27182 ;
  assign n27184 = n27183 ^ n18501 ^ n16094 ;
  assign n27185 = n8208 & n26553 ;
  assign n27186 = ( n8696 & ~n25976 ) | ( n8696 & n27185 ) | ( ~n25976 & n27185 ) ;
  assign n27187 = n5026 | n17020 ;
  assign n27188 = n27187 ^ n4624 ^ 1'b0 ;
  assign n27189 = n27186 & n27188 ;
  assign n27191 = n7900 ^ n1895 ^ 1'b0 ;
  assign n27190 = ~n1766 & n6683 ;
  assign n27192 = n27191 ^ n27190 ^ 1'b0 ;
  assign n27193 = n16286 ^ n919 ^ 1'b0 ;
  assign n27194 = n26051 | n27193 ;
  assign n27195 = ~n19968 & n21371 ;
  assign n27196 = n3081 & n27195 ;
  assign n27197 = n381 & ~n437 ;
  assign n27198 = n27197 ^ n269 ^ 1'b0 ;
  assign n27199 = ~n9791 & n14683 ;
  assign n27200 = n6168 & n27199 ;
  assign n27201 = ( n1206 & n3412 ) | ( n1206 & ~n27200 ) | ( n3412 & ~n27200 ) ;
  assign n27202 = n17310 ^ n2712 ^ 1'b0 ;
  assign n27203 = n12499 & ~n14724 ;
  assign n27204 = n27203 ^ n9005 ^ 1'b0 ;
  assign n27205 = n6771 | n27204 ;
  assign n27206 = ( ~n7860 & n17666 ) | ( ~n7860 & n27205 ) | ( n17666 & n27205 ) ;
  assign n27207 = n2752 | n11811 ;
  assign n27208 = n27207 ^ n4937 ^ 1'b0 ;
  assign n27209 = n14765 & ~n15749 ;
  assign n27210 = n16177 & ~n27209 ;
  assign n27211 = ( ~n18000 & n27208 ) | ( ~n18000 & n27210 ) | ( n27208 & n27210 ) ;
  assign n27212 = n7523 | n13591 ;
  assign n27213 = n3790 & ~n27212 ;
  assign n27214 = ~n251 & n7428 ;
  assign n27215 = n2421 & ~n7830 ;
  assign n27216 = n27215 ^ n3187 ^ 1'b0 ;
  assign n27217 = n7482 ^ n6774 ^ 1'b0 ;
  assign n27218 = n27217 ^ n867 ^ 1'b0 ;
  assign n27219 = ~n27216 & n27218 ;
  assign n27220 = n19727 ^ n16286 ^ 1'b0 ;
  assign n27221 = n20216 & n27220 ;
  assign n27222 = n19150 & n24038 ;
  assign n27223 = n5404 & ~n19108 ;
  assign n27224 = ~n7142 & n27223 ;
  assign n27225 = n878 & ~n27224 ;
  assign n27226 = n27225 ^ n14533 ^ 1'b0 ;
  assign n27227 = n27222 & n27226 ;
  assign n27228 = ~n27221 & n27227 ;
  assign n27229 = n24092 ^ n6699 ^ 1'b0 ;
  assign n27230 = n3027 | n27229 ;
  assign n27231 = ( ~n1962 & n16882 ) | ( ~n1962 & n27230 ) | ( n16882 & n27230 ) ;
  assign n27232 = n22903 ^ n966 ^ 1'b0 ;
  assign n27233 = n4352 & ~n4792 ;
  assign n27234 = n10934 & n27233 ;
  assign n27235 = ~n37 & n27234 ;
  assign n27236 = n15124 & n18963 ;
  assign n27237 = n27236 ^ n9226 ^ 1'b0 ;
  assign n27238 = ~n5967 & n27237 ;
  assign n27239 = n27238 ^ n22524 ^ 1'b0 ;
  assign n27240 = n686 | n21953 ;
  assign n27241 = n27240 ^ n205 ^ 1'b0 ;
  assign n27242 = n27241 ^ n14960 ^ n9528 ;
  assign n27243 = ( n510 & n1370 ) | ( n510 & n24189 ) | ( n1370 & n24189 ) ;
  assign n27244 = n5036 & n19509 ;
  assign n27245 = n3481 & ~n19665 ;
  assign n27246 = n27245 ^ n7137 ^ 1'b0 ;
  assign n27247 = n19172 ^ n16341 ^ n16234 ;
  assign n27248 = n27247 ^ n536 ^ 1'b0 ;
  assign n27249 = n26227 & n27248 ;
  assign n27250 = n9626 | n19212 ;
  assign n27251 = ( ~n5250 & n12106 ) | ( ~n5250 & n27250 ) | ( n12106 & n27250 ) ;
  assign n27252 = n24804 ^ n19058 ^ n8985 ;
  assign n27253 = ~n2391 & n15670 ;
  assign n27254 = n12480 ^ n2845 ^ 1'b0 ;
  assign n27255 = n27253 & ~n27254 ;
  assign n27256 = n27255 ^ n20861 ^ 1'b0 ;
  assign n27257 = n18457 ^ n9108 ^ 1'b0 ;
  assign n27258 = n17147 ^ n13233 ^ n6770 ;
  assign n27259 = n7053 ^ n3054 ^ 1'b0 ;
  assign n27260 = n21862 ^ n21752 ^ 1'b0 ;
  assign n27261 = n10516 ^ n7462 ^ 1'b0 ;
  assign n27262 = ~n14497 & n27261 ;
  assign n27263 = n27262 ^ n2907 ^ 1'b0 ;
  assign n27264 = ~n27260 & n27263 ;
  assign n27266 = n3729 & ~n14476 ;
  assign n27265 = ~n5623 & n18692 ;
  assign n27267 = n27266 ^ n27265 ^ 1'b0 ;
  assign n27268 = n27267 ^ n26392 ^ 1'b0 ;
  assign n27269 = n12155 | n27268 ;
  assign n27272 = n18553 & n23646 ;
  assign n27270 = ( n4068 & n14452 ) | ( n4068 & ~n15005 ) | ( n14452 & ~n15005 ) ;
  assign n27271 = n15776 & ~n27270 ;
  assign n27273 = n27272 ^ n27271 ^ 1'b0 ;
  assign n27274 = n20751 ^ n5259 ^ 1'b0 ;
  assign n27275 = n27273 & n27274 ;
  assign n27276 = n10825 ^ n4141 ^ 1'b0 ;
  assign n27277 = n27276 ^ n1970 ^ n319 ;
  assign n27278 = ( ~n2173 & n23672 ) | ( ~n2173 & n27277 ) | ( n23672 & n27277 ) ;
  assign n27279 = n27278 ^ n18252 ^ 1'b0 ;
  assign n27280 = n16971 ^ n8979 ^ 1'b0 ;
  assign n27281 = n12877 ^ n12770 ^ n2403 ;
  assign n27282 = n27280 | n27281 ;
  assign n27283 = n3595 & ~n18048 ;
  assign n27284 = ~n7271 & n17625 ;
  assign n27285 = n4558 & n27284 ;
  assign n27286 = n24264 ^ n797 ^ 1'b0 ;
  assign n27287 = n11062 ^ n8408 ^ 1'b0 ;
  assign n27288 = n13498 & n27117 ;
  assign n27289 = ( x10 & ~n10792 ) | ( x10 & n27288 ) | ( ~n10792 & n27288 ) ;
  assign n27290 = n1858 & ~n27289 ;
  assign n27291 = n19497 ^ n14229 ^ 1'b0 ;
  assign n27292 = ~n2806 & n27291 ;
  assign n27293 = n23352 ^ n6227 ^ 1'b0 ;
  assign n27294 = ( n8128 & ~n27292 ) | ( n8128 & n27293 ) | ( ~n27292 & n27293 ) ;
  assign n27295 = n27063 ^ n9954 ^ 1'b0 ;
  assign n27296 = n4019 & ~n20648 ;
  assign n27297 = n27296 ^ n8740 ^ 1'b0 ;
  assign n27298 = ( ~n26699 & n27295 ) | ( ~n26699 & n27297 ) | ( n27295 & n27297 ) ;
  assign n27299 = n13567 ^ n8639 ^ n8058 ;
  assign n27300 = n21810 ^ n6866 ^ 1'b0 ;
  assign n27301 = n143 | n27300 ;
  assign n27302 = ~n5435 & n21943 ;
  assign n27303 = n11233 ^ n5234 ^ 1'b0 ;
  assign n27304 = n14674 | n27303 ;
  assign n27305 = n1124 | n27304 ;
  assign n27306 = n27305 ^ n14035 ^ 1'b0 ;
  assign n27307 = n1888 & ~n27306 ;
  assign n27308 = ~n6353 & n27307 ;
  assign n27311 = n2379 & ~n15876 ;
  assign n27312 = n27311 ^ n3382 ^ 1'b0 ;
  assign n27309 = n6383 ^ n3075 ^ 1'b0 ;
  assign n27310 = n9769 & n27309 ;
  assign n27313 = n27312 ^ n27310 ^ 1'b0 ;
  assign n27314 = n22996 ^ n17700 ^ 1'b0 ;
  assign n27315 = n1761 | n10971 ;
  assign n27316 = n21001 | n26185 ;
  assign n27317 = n18986 ^ n5563 ^ 1'b0 ;
  assign n27318 = n27317 ^ n25916 ^ n22729 ;
  assign n27319 = n4721 & ~n20426 ;
  assign n27326 = n8873 & n13426 ;
  assign n27327 = ~n13426 & n27326 ;
  assign n27323 = n5904 & ~n16755 ;
  assign n27324 = n16755 & n27323 ;
  assign n27325 = n5933 | n27324 ;
  assign n27328 = n27327 ^ n27325 ^ 1'b0 ;
  assign n27321 = n1506 & ~n23214 ;
  assign n27320 = n3909 & ~n9866 ;
  assign n27322 = n27321 ^ n27320 ^ 1'b0 ;
  assign n27329 = n27328 ^ n27322 ^ 1'b0 ;
  assign n27330 = n22723 & ~n27329 ;
  assign n27333 = n9935 ^ n7103 ^ 1'b0 ;
  assign n27334 = n8453 | n27333 ;
  assign n27335 = n27334 ^ n24984 ^ n6298 ;
  assign n27336 = n27335 ^ n15126 ^ 1'b0 ;
  assign n27331 = n16517 ^ n11819 ^ n6138 ;
  assign n27332 = n15990 & n27331 ;
  assign n27337 = n27336 ^ n27332 ^ 1'b0 ;
  assign n27338 = n2828 | n25562 ;
  assign n27344 = n5773 ^ n5628 ^ n1143 ;
  assign n27339 = ~n5831 & n8090 ;
  assign n27340 = n3904 ^ n2820 ^ 1'b0 ;
  assign n27341 = n17319 | n27340 ;
  assign n27342 = ( n9618 & n12799 ) | ( n9618 & ~n27341 ) | ( n12799 & ~n27341 ) ;
  assign n27343 = n27339 | n27342 ;
  assign n27345 = n27344 ^ n27343 ^ 1'b0 ;
  assign n27346 = n1134 | n1913 ;
  assign n27347 = n1894 & ~n27346 ;
  assign n27348 = n11605 & ~n12177 ;
  assign n27349 = n13006 | n27348 ;
  assign n27350 = n27347 & ~n27349 ;
  assign n27351 = ~n59 & n3595 ;
  assign n27352 = n4113 & ~n15160 ;
  assign n27353 = n27352 ^ n7183 ^ 1'b0 ;
  assign n27354 = n27351 & n27353 ;
  assign n27355 = n5464 & n7836 ;
  assign n27356 = n1000 & n8782 ;
  assign n27357 = n27356 ^ n4411 ^ 1'b0 ;
  assign n27358 = ~n13378 & n24534 ;
  assign n27359 = n17994 & n20188 ;
  assign n27360 = ~n26146 & n27359 ;
  assign n27361 = n27360 ^ n10780 ^ 1'b0 ;
  assign n27362 = n14347 & n17946 ;
  assign n27363 = n27362 ^ n26288 ^ 1'b0 ;
  assign n27364 = ( n7617 & ~n10296 ) | ( n7617 & n11475 ) | ( ~n10296 & n11475 ) ;
  assign n27365 = n19677 & ~n27364 ;
  assign n27366 = n27365 ^ n795 ^ 1'b0 ;
  assign n27367 = n27363 | n27366 ;
  assign n27368 = n20850 & ~n25089 ;
  assign n27369 = n6062 & n27368 ;
  assign n27370 = n6426 | n11603 ;
  assign n27371 = n9830 | n27370 ;
  assign n27372 = n7297 & n10797 ;
  assign n27373 = n3109 | n15928 ;
  assign n27374 = n6362 & ~n27373 ;
  assign n27375 = n12946 & ~n14977 ;
  assign n27376 = n2651 & n27375 ;
  assign n27377 = ( n27372 & n27374 ) | ( n27372 & ~n27376 ) | ( n27374 & ~n27376 ) ;
  assign n27378 = n21627 ^ n21344 ^ 1'b0 ;
  assign n27379 = n27377 & n27378 ;
  assign n27380 = n17222 & n27379 ;
  assign n27381 = n4445 | n27380 ;
  assign n27382 = ( n3508 & n7917 ) | ( n3508 & ~n22315 ) | ( n7917 & ~n22315 ) ;
  assign n27383 = n7665 & n27382 ;
  assign n27384 = ~n20811 & n27383 ;
  assign n27385 = n12159 | n25121 ;
  assign n27389 = n15543 ^ n1569 ^ 1'b0 ;
  assign n27390 = ~n3491 & n27389 ;
  assign n27386 = n2068 | n8424 ;
  assign n27387 = n1258 | n27386 ;
  assign n27388 = n6506 & n27387 ;
  assign n27391 = n27390 ^ n27388 ^ 1'b0 ;
  assign n27392 = ~n27385 & n27391 ;
  assign n27393 = n13111 ^ n12800 ^ n9146 ;
  assign n27394 = n14106 & ~n27393 ;
  assign n27395 = n4275 & n27394 ;
  assign n27396 = n14619 | n20872 ;
  assign n27397 = n27396 ^ n13477 ^ 1'b0 ;
  assign n27398 = n2377 & n6050 ;
  assign n27399 = n4088 & n27398 ;
  assign n27400 = n11768 | n24942 ;
  assign n27410 = n11572 & n22716 ;
  assign n27401 = ~n36 & n8524 ;
  assign n27402 = n27401 ^ n11059 ^ 1'b0 ;
  assign n27403 = ~n10987 & n20817 ;
  assign n27404 = n6890 ^ n250 ^ 1'b0 ;
  assign n27405 = ~n2650 & n27404 ;
  assign n27406 = n550 & n27405 ;
  assign n27407 = n13374 & n27406 ;
  assign n27408 = n27407 ^ n20332 ^ 1'b0 ;
  assign n27409 = ( n27402 & n27403 ) | ( n27402 & n27408 ) | ( n27403 & n27408 ) ;
  assign n27411 = n27410 ^ n27409 ^ n12555 ;
  assign n27412 = n1100 | n15053 ;
  assign n27413 = n8467 | n27412 ;
  assign n27414 = n5420 & ~n20848 ;
  assign n27415 = n1154 ^ n776 ^ 1'b0 ;
  assign n27416 = n13196 ^ n12853 ^ n7702 ;
  assign n27417 = n27415 | n27416 ;
  assign n27418 = n23193 ^ n2731 ^ 1'b0 ;
  assign n27419 = ~n5099 & n27418 ;
  assign n27420 = n18193 | n27419 ;
  assign n27421 = n18099 & ~n27420 ;
  assign n27422 = n5741 & ~n8150 ;
  assign n27423 = n27422 ^ n21116 ^ 1'b0 ;
  assign n27424 = n12010 ^ n1818 ^ 1'b0 ;
  assign n27425 = n184 & ~n624 ;
  assign n27426 = n22312 ^ n18882 ^ 1'b0 ;
  assign n27427 = ~n7665 & n13396 ;
  assign n27428 = n27427 ^ n13243 ^ 1'b0 ;
  assign n27429 = n21408 ^ n13123 ^ 1'b0 ;
  assign n27430 = n17445 & n24646 ;
  assign n27431 = n27429 & n27430 ;
  assign n27432 = n17535 ^ n9555 ^ 1'b0 ;
  assign n27433 = n3195 & ~n27432 ;
  assign n27434 = n19959 ^ n16812 ^ 1'b0 ;
  assign n27435 = n11722 | n27434 ;
  assign n27436 = n19793 ^ n13712 ^ 1'b0 ;
  assign n27437 = n20041 & ~n27436 ;
  assign n27438 = ~n18266 & n27437 ;
  assign n27439 = n5980 ^ n4318 ^ 1'b0 ;
  assign n27440 = n27439 ^ n19347 ^ n2922 ;
  assign n27441 = n27440 ^ n5175 ^ 1'b0 ;
  assign n27442 = n8018 ^ n40 ^ 1'b0 ;
  assign n27443 = ( ~n5262 & n22052 ) | ( ~n5262 & n25708 ) | ( n22052 & n25708 ) ;
  assign n27444 = n22521 ^ n10517 ^ n4683 ;
  assign n27445 = ( n929 & n9997 ) | ( n929 & n27444 ) | ( n9997 & n27444 ) ;
  assign n27446 = n8652 & ~n11260 ;
  assign n27447 = n17258 & n27446 ;
  assign n27448 = n24660 ^ n18192 ^ 1'b0 ;
  assign n27449 = n18716 ^ n2922 ^ 1'b0 ;
  assign n27450 = ~n11241 & n21062 ;
  assign n27451 = ( n11245 & ~n27449 ) | ( n11245 & n27450 ) | ( ~n27449 & n27450 ) ;
  assign n27453 = ~n2759 & n3975 ;
  assign n27454 = n7282 & n27453 ;
  assign n27452 = ( n5790 & n8774 ) | ( n5790 & ~n17247 ) | ( n8774 & ~n17247 ) ;
  assign n27455 = n27454 ^ n27452 ^ 1'b0 ;
  assign n27456 = ~n12401 & n27455 ;
  assign n27457 = n21667 ^ n4334 ^ 1'b0 ;
  assign n27458 = n5109 & n27457 ;
  assign n27459 = n7707 & ~n15962 ;
  assign n27460 = n12389 ^ n615 ^ 1'b0 ;
  assign n27461 = n2695 | n6093 ;
  assign n27462 = n6059 & n13546 ;
  assign n27463 = ~n18692 & n27462 ;
  assign n27464 = n6652 | n7118 ;
  assign n27465 = n27464 ^ n2411 ^ 1'b0 ;
  assign n27466 = n27465 ^ n8318 ^ 1'b0 ;
  assign n27467 = n5346 & n27466 ;
  assign n27477 = n2367 & n14879 ;
  assign n27472 = ( n945 & n4758 ) | ( n945 & n8232 ) | ( n4758 & n8232 ) ;
  assign n27473 = ~n15095 & n27472 ;
  assign n27474 = n27473 ^ n6282 ^ 1'b0 ;
  assign n27468 = n33 | n4930 ;
  assign n27469 = n7052 & ~n27468 ;
  assign n27470 = n7860 ^ n51 ^ 1'b0 ;
  assign n27471 = ~n27469 & n27470 ;
  assign n27475 = n27474 ^ n27471 ^ n15934 ;
  assign n27476 = ~n14332 & n27475 ;
  assign n27478 = n27477 ^ n27476 ^ 1'b0 ;
  assign n27479 = n20368 ^ n5720 ^ n3401 ;
  assign n27480 = n10171 & ~n27479 ;
  assign n27481 = n23225 & n27480 ;
  assign n27482 = n1109 | n18401 ;
  assign n27483 = n27482 ^ n4670 ^ 1'b0 ;
  assign n27484 = ( n26104 & n27104 ) | ( n26104 & n27483 ) | ( n27104 & n27483 ) ;
  assign n27485 = n22023 ^ n20650 ^ 1'b0 ;
  assign n27486 = n4736 & ~n27485 ;
  assign n27487 = n11335 | n21195 ;
  assign n27488 = n10843 & ~n27487 ;
  assign n27489 = n6460 & n19936 ;
  assign n27490 = n5175 ^ n2135 ^ 1'b0 ;
  assign n27491 = n7551 & n27490 ;
  assign n27492 = n10430 | n26421 ;
  assign n27493 = n27492 ^ n13455 ^ 1'b0 ;
  assign n27494 = ( ~n10178 & n12823 ) | ( ~n10178 & n27493 ) | ( n12823 & n27493 ) ;
  assign n27495 = n9351 & n16974 ;
  assign n27496 = ~n27494 & n27495 ;
  assign n27497 = n7704 & n11219 ;
  assign n27498 = ~n4290 & n6251 ;
  assign n27501 = n26418 ^ n7620 ^ 1'b0 ;
  assign n27502 = n12032 & ~n27501 ;
  assign n27499 = n8440 & ~n9507 ;
  assign n27500 = ~n9968 & n27499 ;
  assign n27503 = n27502 ^ n27500 ^ 1'b0 ;
  assign n27504 = n4421 & ~n6407 ;
  assign n27505 = n27504 ^ n3691 ^ 1'b0 ;
  assign n27506 = ~n2023 & n27505 ;
  assign n27507 = n10098 & n27506 ;
  assign n27508 = n27507 ^ n3776 ^ 1'b0 ;
  assign n27509 = n8424 | n21339 ;
  assign n27510 = n20052 & ~n24644 ;
  assign n27511 = ~n9332 & n27510 ;
  assign n27512 = n27511 ^ n1368 ^ 1'b0 ;
  assign n27513 = n21075 ^ n1220 ^ 1'b0 ;
  assign n27514 = n4993 | n27513 ;
  assign n27515 = ( n4803 & n9935 ) | ( n4803 & ~n27514 ) | ( n9935 & ~n27514 ) ;
  assign n27516 = ( n4452 & n18184 ) | ( n4452 & n27515 ) | ( n18184 & n27515 ) ;
  assign n27517 = n27516 ^ n17136 ^ n4072 ;
  assign n27518 = ~n1248 & n18076 ;
  assign n27519 = n6403 & ~n27518 ;
  assign n27520 = ~n718 & n1029 ;
  assign n27521 = n27520 ^ n4974 ^ 1'b0 ;
  assign n27522 = n27521 ^ n26664 ^ n20343 ;
  assign n27523 = n27522 ^ n15987 ^ 1'b0 ;
  assign n27526 = n5749 & ~n9615 ;
  assign n27524 = n3503 | n11633 ;
  assign n27525 = n27524 ^ n1393 ^ 1'b0 ;
  assign n27527 = n27526 ^ n27525 ^ 1'b0 ;
  assign n27528 = n3370 & ~n9238 ;
  assign n27529 = n27527 & n27528 ;
  assign n27530 = n8556 & ~n10802 ;
  assign n27531 = n6107 ^ n6094 ^ n1319 ;
  assign n27532 = n6628 & n27531 ;
  assign n27533 = n15982 ^ n13275 ^ n5722 ;
  assign n27534 = ( ~n14220 & n24601 ) | ( ~n14220 & n27533 ) | ( n24601 & n27533 ) ;
  assign n27535 = n9318 & n9560 ;
  assign n27536 = n8085 & n27535 ;
  assign n27537 = ~n5475 & n7823 ;
  assign n27538 = ~n27536 & n27537 ;
  assign n27539 = n3198 ^ n1532 ^ 1'b0 ;
  assign n27540 = ~n1353 & n27539 ;
  assign n27541 = n18716 & n27540 ;
  assign n27542 = n27541 ^ n20614 ^ 1'b0 ;
  assign n27543 = n4275 | n4964 ;
  assign n27544 = n1368 & n21878 ;
  assign n27545 = n27543 & n27544 ;
  assign n27546 = n6919 | n27545 ;
  assign n27547 = n19868 & ~n27546 ;
  assign n27548 = n11830 ^ n3637 ^ n1138 ;
  assign n27549 = ( n3387 & n21914 ) | ( n3387 & n27548 ) | ( n21914 & n27548 ) ;
  assign n27550 = n3784 | n9918 ;
  assign n27551 = n8103 | n24109 ;
  assign n27552 = n1535 ^ n865 ^ 1'b0 ;
  assign n27553 = n4691 & n27552 ;
  assign n27554 = n13340 ^ n5483 ^ 1'b0 ;
  assign n27555 = ~n27553 & n27554 ;
  assign n27556 = n2377 & ~n2791 ;
  assign n27557 = n11888 ^ n435 ^ 1'b0 ;
  assign n27558 = n16450 & n27557 ;
  assign n27559 = n4567 & n27558 ;
  assign n27560 = n17035 ^ n6852 ^ n6020 ;
  assign n27561 = n194 & ~n2664 ;
  assign n27562 = ~n9372 & n27561 ;
  assign n27563 = n2304 | n27562 ;
  assign n27564 = n3112 & ~n27515 ;
  assign n27565 = n27564 ^ n18082 ^ 1'b0 ;
  assign n27566 = ~n27563 & n27565 ;
  assign n27567 = x10 & n27566 ;
  assign n27568 = ~n27560 & n27567 ;
  assign n27569 = n818 & ~n7916 ;
  assign n27570 = n27569 ^ n12053 ^ 1'b0 ;
  assign n27571 = n191 & n7605 ;
  assign n27572 = n11275 & n27571 ;
  assign n27573 = n24732 ^ n4207 ^ 1'b0 ;
  assign n27574 = n20859 & n27573 ;
  assign n27575 = ~n13467 & n27574 ;
  assign n27576 = ~n10874 & n27575 ;
  assign n27577 = ( n443 & ~n14100 ) | ( n443 & n27576 ) | ( ~n14100 & n27576 ) ;
  assign n27578 = ( n12077 & n23308 ) | ( n12077 & n27577 ) | ( n23308 & n27577 ) ;
  assign n27579 = n4506 | n16343 ;
  assign n27580 = n15385 | n27579 ;
  assign n27581 = ~n9669 & n14700 ;
  assign n27582 = n27581 ^ n3817 ^ 1'b0 ;
  assign n27583 = n24485 & n27582 ;
  assign n27584 = n1262 ^ n87 ^ 1'b0 ;
  assign n27585 = n27584 ^ n5372 ^ 1'b0 ;
  assign n27586 = n22394 | n27585 ;
  assign n27587 = n8071 ^ n6050 ^ 1'b0 ;
  assign n27588 = n2775 & ~n27587 ;
  assign n27589 = n18394 ^ n572 ^ 1'b0 ;
  assign n27590 = n23306 & ~n27589 ;
  assign n27591 = n20399 ^ n617 ^ 1'b0 ;
  assign n27592 = n13658 ^ n11429 ^ 1'b0 ;
  assign n27593 = n27592 ^ n23492 ^ n14551 ;
  assign n27594 = n6847 & ~n11748 ;
  assign n27595 = n5157 & ~n27594 ;
  assign n27596 = ~n20858 & n27595 ;
  assign n27597 = n4388 ^ n3784 ^ 1'b0 ;
  assign n27598 = n27596 & ~n27597 ;
  assign n27599 = n3916 & n8183 ;
  assign n27600 = n15013 & n27599 ;
  assign n27601 = n14214 ^ n6451 ^ 1'b0 ;
  assign n27602 = n23729 ^ n4330 ^ 1'b0 ;
  assign n27603 = n2422 | n12267 ;
  assign n27604 = n5773 & ~n27603 ;
  assign n27605 = n7976 ^ n6683 ^ 1'b0 ;
  assign n27606 = n3460 | n27605 ;
  assign n27607 = n4493 & ~n6666 ;
  assign n27608 = n22662 & n27607 ;
  assign n27609 = ~n12322 & n27608 ;
  assign n27610 = n27609 ^ n22988 ^ 1'b0 ;
  assign n27611 = n2209 ^ n63 ^ 1'b0 ;
  assign n27612 = n1625 | n27611 ;
  assign n27613 = n16213 & n27612 ;
  assign n27614 = n23081 ^ n16556 ^ 1'b0 ;
  assign n27615 = n18955 | n27614 ;
  assign n27616 = n10861 | n21414 ;
  assign n27617 = n2456 | n27616 ;
  assign n27618 = n19792 | n22239 ;
  assign n27619 = n3506 ^ n3408 ^ 1'b0 ;
  assign n27620 = ~n1993 & n27619 ;
  assign n27621 = n5311 | n6536 ;
  assign n27622 = n27621 ^ n8141 ^ 1'b0 ;
  assign n27623 = n27622 ^ n21076 ^ n5137 ;
  assign n27624 = n23128 ^ n16234 ^ 1'b0 ;
  assign n27625 = n23505 | n27624 ;
  assign n27626 = n21110 ^ n2230 ^ 1'b0 ;
  assign n27627 = n4965 & n27626 ;
  assign n27628 = n27627 ^ n3303 ^ 1'b0 ;
  assign n27629 = n19135 & n27628 ;
  assign n27630 = ~n18001 & n27629 ;
  assign n27631 = ~n2005 & n16974 ;
  assign n27632 = n27631 ^ n6131 ^ n2917 ;
  assign n27634 = ( n4724 & n12138 ) | ( n4724 & n19014 ) | ( n12138 & n19014 ) ;
  assign n27635 = n27634 ^ n27582 ^ 1'b0 ;
  assign n27633 = n18496 & n27234 ;
  assign n27636 = n27635 ^ n27633 ^ n14089 ;
  assign n27637 = n18775 ^ n6801 ^ n4694 ;
  assign n27638 = ( n1003 & n9211 ) | ( n1003 & n25553 ) | ( n9211 & n25553 ) ;
  assign n27639 = ~n10208 & n17649 ;
  assign n27640 = ~n27638 & n27639 ;
  assign n27641 = n16727 & ~n25291 ;
  assign n27642 = n5486 & ~n12788 ;
  assign n27643 = n27642 ^ n18177 ^ n18157 ;
  assign n27644 = n27641 | n27643 ;
  assign n27646 = n3079 & ~n19865 ;
  assign n27647 = ~n4041 & n27646 ;
  assign n27645 = ( n7638 & ~n21029 ) | ( n7638 & n21382 ) | ( ~n21029 & n21382 ) ;
  assign n27648 = n27647 ^ n27645 ^ 1'b0 ;
  assign n27649 = ~n692 & n9352 ;
  assign n27650 = n2904 & n10953 ;
  assign n27651 = n10579 & n27650 ;
  assign n27652 = ( n1386 & n27649 ) | ( n1386 & n27651 ) | ( n27649 & n27651 ) ;
  assign n27653 = ( n25893 & n26873 ) | ( n25893 & n27652 ) | ( n26873 & n27652 ) ;
  assign n27654 = n6087 ^ n3134 ^ 1'b0 ;
  assign n27655 = n7969 ^ n682 ^ 1'b0 ;
  assign n27656 = ~n3263 & n4992 ;
  assign n27657 = n17736 & n25839 ;
  assign n27661 = ( ~n113 & n1255 ) | ( ~n113 & n5935 ) | ( n1255 & n5935 ) ;
  assign n27658 = ~n209 & n780 ;
  assign n27659 = n9070 | n10433 ;
  assign n27660 = n27658 & ~n27659 ;
  assign n27662 = n27661 ^ n27660 ^ n11898 ;
  assign n27663 = n2369 & ~n16593 ;
  assign n27664 = n27663 ^ n9530 ^ 1'b0 ;
  assign n27665 = n21996 ^ n12932 ^ 1'b0 ;
  assign n27666 = n13438 & ~n27665 ;
  assign n27667 = n27666 ^ n6376 ^ 1'b0 ;
  assign n27668 = n9275 & n27667 ;
  assign n27669 = n4382 | n4531 ;
  assign n27670 = n27669 ^ n1558 ^ 1'b0 ;
  assign n27671 = ~n4345 & n27670 ;
  assign n27672 = n1303 ^ n762 ^ 1'b0 ;
  assign n27673 = ~n884 & n27672 ;
  assign n27674 = n26963 ^ n2849 ^ 1'b0 ;
  assign n27675 = ~n17384 & n27674 ;
  assign n27676 = n27673 & n27675 ;
  assign n27677 = n27671 & n27676 ;
  assign n27678 = n6437 ^ n3819 ^ 1'b0 ;
  assign n27679 = n17922 | n21809 ;
  assign n27680 = n23001 ^ n12135 ^ 1'b0 ;
  assign n27681 = n6650 | n8455 ;
  assign n27682 = n20943 ^ n17959 ^ 1'b0 ;
  assign n27683 = n6810 ^ n794 ^ 1'b0 ;
  assign n27684 = ( n2104 & ~n22677 ) | ( n2104 & n26226 ) | ( ~n22677 & n26226 ) ;
  assign n27685 = n609 & ~n1176 ;
  assign n27686 = ~n5596 & n27685 ;
  assign n27687 = n27686 ^ n605 ^ 1'b0 ;
  assign n27688 = n17299 | n27687 ;
  assign n27689 = n15349 ^ n1088 ^ 1'b0 ;
  assign n27690 = n7215 & n27689 ;
  assign n27691 = n27690 ^ n4536 ^ 1'b0 ;
  assign n27692 = n1906 | n8109 ;
  assign n27693 = n27692 ^ n4923 ^ 1'b0 ;
  assign n27694 = ~n21005 & n27693 ;
  assign n27695 = ( n27688 & ~n27691 ) | ( n27688 & n27694 ) | ( ~n27691 & n27694 ) ;
  assign n27696 = n1647 & ~n5907 ;
  assign n27697 = n27696 ^ n2314 ^ 1'b0 ;
  assign n27698 = n3635 & n24411 ;
  assign n27699 = n27698 ^ n14761 ^ 1'b0 ;
  assign n27700 = n27699 ^ n13224 ^ 1'b0 ;
  assign n27701 = n27700 ^ n11941 ^ 1'b0 ;
  assign n27705 = n744 | n19961 ;
  assign n27706 = n744 & ~n27705 ;
  assign n27702 = n2658 | n3892 ;
  assign n27703 = n3892 & ~n27702 ;
  assign n27704 = n4657 | n27703 ;
  assign n27707 = n27706 ^ n27704 ^ 1'b0 ;
  assign n27708 = ~n4246 & n4458 ;
  assign n27709 = n4246 & n27708 ;
  assign n27710 = n2249 & ~n27709 ;
  assign n27711 = ~n2249 & n27710 ;
  assign n27712 = n27707 | n27711 ;
  assign n27713 = n27707 & ~n27712 ;
  assign n27714 = x10 | n11066 ;
  assign n27715 = n11066 & ~n27714 ;
  assign n27716 = n27715 ^ n18768 ^ 1'b0 ;
  assign n27717 = ~n27713 & n27716 ;
  assign n27718 = n27713 & n27717 ;
  assign n27719 = n1654 ^ n1481 ^ 1'b0 ;
  assign n27720 = ~n126 & n27719 ;
  assign n27721 = n27720 ^ n24344 ^ n1115 ;
  assign n27722 = n27718 & n27721 ;
  assign n27723 = ~n10108 & n10540 ;
  assign n27724 = n27723 ^ n24483 ^ 1'b0 ;
  assign n27725 = n10833 ^ n5965 ^ 1'b0 ;
  assign n27726 = n17746 & n27725 ;
  assign n27727 = n27726 ^ n16323 ^ n2339 ;
  assign n27728 = n19645 ^ n13567 ^ 1'b0 ;
  assign n27729 = n8546 & ~n27728 ;
  assign n27730 = n27729 ^ n21931 ^ n8291 ;
  assign n27731 = n5509 ^ n5400 ^ 1'b0 ;
  assign n27732 = n4614 & n27731 ;
  assign n27733 = ~n17468 & n27732 ;
  assign n27734 = n13905 ^ n10581 ^ 1'b0 ;
  assign n27735 = n10393 & ~n27734 ;
  assign n27736 = n7071 | n10180 ;
  assign n27737 = n27736 ^ n6045 ^ 1'b0 ;
  assign n27738 = n27737 ^ n19887 ^ 1'b0 ;
  assign n27739 = ~n3926 & n8977 ;
  assign n27740 = ~n1681 & n27739 ;
  assign n27741 = n6142 & n21506 ;
  assign n27742 = n27741 ^ n1543 ^ 1'b0 ;
  assign n27743 = n4402 & ~n27742 ;
  assign n27744 = n27743 ^ n12692 ^ 1'b0 ;
  assign n27745 = n17526 ^ n8888 ^ 1'b0 ;
  assign n27746 = n12678 ^ n2105 ^ 1'b0 ;
  assign n27747 = ( ~n503 & n2126 ) | ( ~n503 & n16771 ) | ( n2126 & n16771 ) ;
  assign n27748 = n5769 | n6225 ;
  assign n27749 = n296 & ~n16812 ;
  assign n27750 = n14748 & ~n22077 ;
  assign n27751 = n27749 & n27750 ;
  assign n27754 = n442 & ~n18501 ;
  assign n27755 = n16499 & n27754 ;
  assign n27752 = n3383 & ~n5587 ;
  assign n27753 = n27752 ^ n8872 ^ n2338 ;
  assign n27756 = n27755 ^ n27753 ^ 1'b0 ;
  assign n27757 = n23005 ^ n21463 ^ 1'b0 ;
  assign n27758 = ( n1088 & n4457 ) | ( n1088 & ~n27757 ) | ( n4457 & ~n27757 ) ;
  assign n27759 = ~n10962 & n13263 ;
  assign n27760 = n6805 & n27759 ;
  assign n27761 = ~n27758 & n27760 ;
  assign n27762 = n213 & n9027 ;
  assign n27763 = n12697 & ~n22945 ;
  assign n27764 = n27763 ^ n7526 ^ 1'b0 ;
  assign n27765 = n8730 & n25482 ;
  assign n27766 = n27765 ^ n1550 ^ 1'b0 ;
  assign n27767 = n24689 & ~n27766 ;
  assign n27768 = n27767 ^ n18272 ^ 1'b0 ;
  assign n27769 = n7046 ^ n100 ^ 1'b0 ;
  assign n27770 = n22377 & n27769 ;
  assign n27771 = ~n1777 & n2122 ;
  assign n27772 = n27770 & n27771 ;
  assign n27773 = n3551 & ~n9130 ;
  assign n27774 = n10057 & n27773 ;
  assign n27775 = n10993 & ~n12461 ;
  assign n27776 = n25687 ^ n10102 ^ 1'b0 ;
  assign n27777 = n24786 ^ n7197 ^ 1'b0 ;
  assign n27778 = n20705 ^ n19544 ^ n11749 ;
  assign n27779 = n25436 ^ n18193 ^ 1'b0 ;
  assign n27780 = n13441 & ~n27779 ;
  assign n27781 = ( ~n5599 & n9946 ) | ( ~n5599 & n10038 ) | ( n9946 & n10038 ) ;
  assign n27782 = n17513 | n27781 ;
  assign n27783 = n27782 ^ n893 ^ 1'b0 ;
  assign n27784 = n661 & ~n27783 ;
  assign n27785 = n27784 ^ n401 ^ 1'b0 ;
  assign n27786 = ~n423 & n13937 ;
  assign n27787 = n27786 ^ n4652 ^ 1'b0 ;
  assign n27788 = n8692 | n27787 ;
  assign n27789 = n27788 ^ n13865 ^ 1'b0 ;
  assign n27790 = n27789 ^ n6896 ^ 1'b0 ;
  assign n27791 = n3797 | n27790 ;
  assign n27792 = ( ~n3541 & n10650 ) | ( ~n3541 & n27791 ) | ( n10650 & n27791 ) ;
  assign n27793 = n27792 ^ n13572 ^ 1'b0 ;
  assign n27794 = ( n7631 & n11302 ) | ( n7631 & n27793 ) | ( n11302 & n27793 ) ;
  assign n27796 = n20811 ^ n947 ^ 1'b0 ;
  assign n27797 = n506 & ~n27796 ;
  assign n27795 = n1344 & ~n5160 ;
  assign n27798 = n27797 ^ n27795 ^ 1'b0 ;
  assign n27799 = n8841 & ~n19041 ;
  assign n27800 = n3500 | n27799 ;
  assign n27801 = n7496 & ~n27800 ;
  assign n27802 = n22516 & ~n25475 ;
  assign n27803 = n10339 & n27802 ;
  assign n27804 = ~n9385 & n24481 ;
  assign n27805 = ~n15781 & n27804 ;
  assign n27806 = n27805 ^ n5174 ^ n4160 ;
  assign n27807 = ~n471 & n27806 ;
  assign n27808 = n7334 & ~n8021 ;
  assign n27809 = ~n21264 & n27808 ;
  assign n27810 = ~n1856 & n27809 ;
  assign n27811 = n27810 ^ n7478 ^ n7071 ;
  assign n27812 = ( n1619 & ~n27807 ) | ( n1619 & n27811 ) | ( ~n27807 & n27811 ) ;
  assign n27813 = n23505 ^ n10446 ^ 1'b0 ;
  assign n27814 = ~n5751 & n8603 ;
  assign n27815 = n1025 & n1470 ;
  assign n27816 = n10004 & n27815 ;
  assign n27817 = n27816 ^ n26810 ^ 1'b0 ;
  assign n27818 = ~n27814 & n27817 ;
  assign n27819 = n3665 ^ n947 ^ 1'b0 ;
  assign n27820 = n27818 & ~n27819 ;
  assign n27821 = n25637 ^ n19973 ^ 1'b0 ;
  assign n27822 = n19188 & ~n25328 ;
  assign n27823 = n16282 ^ n1731 ^ 1'b0 ;
  assign n27824 = ~n8209 & n15325 ;
  assign n27825 = n27824 ^ n3313 ^ 1'b0 ;
  assign n27826 = ( n3120 & ~n17424 ) | ( n3120 & n27825 ) | ( ~n17424 & n27825 ) ;
  assign n27827 = n27826 ^ n25998 ^ 1'b0 ;
  assign n27828 = n27823 & n27827 ;
  assign n27829 = ~n694 & n4520 ;
  assign n27830 = n11262 & n27829 ;
  assign n27831 = ~n23329 & n27830 ;
  assign n27832 = ~n23511 & n26679 ;
  assign n27833 = ~n16731 & n27832 ;
  assign n27834 = n2759 | n15373 ;
  assign n27835 = n27834 ^ n705 ^ 1'b0 ;
  assign n27836 = ( n9094 & n25930 ) | ( n9094 & ~n27835 ) | ( n25930 & ~n27835 ) ;
  assign n27839 = ~n686 & n8943 ;
  assign n27840 = ~n20622 & n27839 ;
  assign n27837 = ~n4308 & n20956 ;
  assign n27838 = n27837 ^ n18387 ^ 1'b0 ;
  assign n27841 = n27840 ^ n27838 ^ 1'b0 ;
  assign n27842 = n15938 & ~n27841 ;
  assign n27843 = n27842 ^ n22512 ^ n8251 ;
  assign n27844 = n7680 & ~n23362 ;
  assign n27845 = n20089 ^ n8355 ^ n1015 ;
  assign n27846 = n27845 ^ n26029 ^ n3491 ;
  assign n27847 = n27846 ^ n24234 ^ 1'b0 ;
  assign n27848 = n448 | n1233 ;
  assign n27849 = n27848 ^ n22823 ^ 1'b0 ;
  assign n27850 = n2072 | n11829 ;
  assign n27851 = n1826 | n27850 ;
  assign n27852 = ~n8265 & n27851 ;
  assign n27853 = n27852 ^ n12214 ^ 1'b0 ;
  assign n27854 = ~n17180 & n27853 ;
  assign n27855 = n7512 ^ n6528 ^ n1587 ;
  assign n27856 = ~n381 & n27855 ;
  assign n27857 = n27856 ^ n6560 ^ 1'b0 ;
  assign n27858 = n14842 ^ n12151 ^ n3248 ;
  assign n27859 = n603 & n1771 ;
  assign n27860 = ~n9283 & n15385 ;
  assign n27861 = n25528 ^ n4102 ^ 1'b0 ;
  assign n27862 = n27860 & n27861 ;
  assign n27863 = n9509 ^ n4685 ^ 1'b0 ;
  assign n27864 = n7798 & ~n21021 ;
  assign n27865 = n27864 ^ n15340 ^ 1'b0 ;
  assign n27866 = n27865 ^ n26664 ^ 1'b0 ;
  assign n27868 = n15815 ^ n7675 ^ 1'b0 ;
  assign n27867 = ( ~x4 & n8729 ) | ( ~x4 & n17915 ) | ( n8729 & n17915 ) ;
  assign n27869 = n27868 ^ n27867 ^ 1'b0 ;
  assign n27870 = n3077 & n5712 ;
  assign n27871 = ~n9959 & n27870 ;
  assign n27872 = n23411 & ~n27871 ;
  assign n27873 = n27872 ^ n2328 ^ 1'b0 ;
  assign n27874 = n5948 ^ n4487 ^ 1'b0 ;
  assign n27875 = n13754 & ~n27874 ;
  assign n27876 = n1079 & n27875 ;
  assign n27877 = n3413 ^ n1921 ^ 1'b0 ;
  assign n27878 = n4525 & n27877 ;
  assign n27879 = n19947 ^ n11221 ^ 1'b0 ;
  assign n27880 = n1650 & n27879 ;
  assign n27881 = n4249 & n27880 ;
  assign n27882 = ~n27878 & n27881 ;
  assign n27884 = ( n6814 & n11182 ) | ( n6814 & ~n16351 ) | ( n11182 & ~n16351 ) ;
  assign n27883 = n17748 ^ n624 ^ 1'b0 ;
  assign n27885 = n27884 ^ n27883 ^ 1'b0 ;
  assign n27886 = n27885 ^ n23258 ^ 1'b0 ;
  assign n27887 = n10129 & n23455 ;
  assign n27888 = ~n17277 & n27887 ;
  assign n27889 = n16468 ^ n16082 ^ 1'b0 ;
  assign n27890 = ~n27888 & n27889 ;
  assign n27891 = n20142 ^ n6681 ^ 1'b0 ;
  assign n27892 = ~n2408 & n23950 ;
  assign n27893 = n7312 & ~n9837 ;
  assign n27894 = n21396 ^ n7577 ^ n6738 ;
  assign n27895 = n195 & n16838 ;
  assign n27896 = n27895 ^ n9496 ^ 1'b0 ;
  assign n27897 = n10634 ^ n3031 ^ 1'b0 ;
  assign n27898 = n27897 ^ n22424 ^ 1'b0 ;
  assign n27899 = n12999 | n27898 ;
  assign n27900 = ( x11 & n27896 ) | ( x11 & ~n27899 ) | ( n27896 & ~n27899 ) ;
  assign n27901 = n11785 & n19056 ;
  assign n27902 = ~n11166 & n27901 ;
  assign n27903 = n27902 ^ n7240 ^ 1'b0 ;
  assign n27904 = n27903 ^ n723 ^ 1'b0 ;
  assign n27905 = n27904 ^ n5794 ^ 1'b0 ;
  assign n27906 = n6746 & n27905 ;
  assign n27907 = n18010 ^ n7617 ^ 1'b0 ;
  assign n27908 = ~n14972 & n18669 ;
  assign n27909 = n15212 ^ n7553 ^ 1'b0 ;
  assign n27910 = n18203 ^ n12866 ^ 1'b0 ;
  assign n27911 = n4970 & n10934 ;
  assign n27912 = ~n6129 & n27911 ;
  assign n27913 = n27494 & ~n27912 ;
  assign n27914 = n27913 ^ n13477 ^ n8414 ;
  assign n27916 = ( n539 & ~n881 ) | ( n539 & n4136 ) | ( ~n881 & n4136 ) ;
  assign n27915 = n5811 ^ n15 ^ 1'b0 ;
  assign n27917 = n27916 ^ n27915 ^ n4858 ;
  assign n27918 = n27917 ^ n8163 ^ 1'b0 ;
  assign n27920 = n12918 ^ n3153 ^ n312 ;
  assign n27919 = n4829 ^ n690 ^ 1'b0 ;
  assign n27921 = n27920 ^ n27919 ^ 1'b0 ;
  assign n27922 = n17825 ^ n5043 ^ 1'b0 ;
  assign n27924 = n25445 ^ n984 ^ 1'b0 ;
  assign n27923 = n2221 & ~n6169 ;
  assign n27925 = n27924 ^ n27923 ^ 1'b0 ;
  assign n27926 = ~n5396 & n16625 ;
  assign n27927 = ( n465 & n4285 ) | ( n465 & n4661 ) | ( n4285 & n4661 ) ;
  assign n27928 = n16155 | n27927 ;
  assign n27929 = n3981 & n12708 ;
  assign n27930 = n27929 ^ n1402 ^ 1'b0 ;
  assign n27931 = n27930 ^ n2985 ^ 1'b0 ;
  assign n27932 = n10953 & n27931 ;
  assign n27933 = n8318 | n27932 ;
  assign n27934 = ~n11829 & n24115 ;
  assign n27935 = n27934 ^ n1145 ^ 1'b0 ;
  assign n27936 = n915 | n15013 ;
  assign n27937 = n3329 | n5975 ;
  assign n27938 = ( ~n27935 & n27936 ) | ( ~n27935 & n27937 ) | ( n27936 & n27937 ) ;
  assign n27939 = n11808 ^ n11655 ^ 1'b0 ;
  assign n27940 = ~n14251 & n27939 ;
  assign n27944 = n25112 ^ n5129 ^ 1'b0 ;
  assign n27945 = n605 & ~n27944 ;
  assign n27943 = n1443 & n4989 ;
  assign n27946 = n27945 ^ n27943 ^ 1'b0 ;
  assign n27941 = n12088 & ~n14475 ;
  assign n27942 = n2070 & ~n27941 ;
  assign n27947 = n27946 ^ n27942 ^ 1'b0 ;
  assign n27948 = n18771 | n27947 ;
  assign n27949 = n1930 | n2321 ;
  assign n27950 = n27949 ^ n1933 ^ 1'b0 ;
  assign n27951 = n27950 ^ n4570 ^ n1223 ;
  assign n27952 = ( n17785 & n24011 ) | ( n17785 & n27951 ) | ( n24011 & n27951 ) ;
  assign n27953 = ~n313 & n27952 ;
  assign n27954 = n24193 & n27953 ;
  assign n27955 = n27954 ^ n26106 ^ 1'b0 ;
  assign n27956 = n23687 & n27955 ;
  assign n27957 = n9733 & ~n13072 ;
  assign n27958 = n19364 & n27957 ;
  assign n27959 = n10239 ^ n6954 ^ 1'b0 ;
  assign n27960 = n11250 | n27959 ;
  assign n27961 = n14454 ^ n12684 ^ 1'b0 ;
  assign n27962 = n984 & ~n27961 ;
  assign n27963 = n8590 ^ n7776 ^ 1'b0 ;
  assign n27964 = n2808 & n9250 ;
  assign n27965 = n17795 ^ n7383 ^ 1'b0 ;
  assign n27966 = n27964 & n27965 ;
  assign n27967 = n12817 ^ n6763 ^ 1'b0 ;
  assign n27968 = n19817 ^ n6977 ^ n438 ;
  assign n27969 = n27968 ^ n9309 ^ n1039 ;
  assign n27970 = ( ~n22791 & n27967 ) | ( ~n22791 & n27969 ) | ( n27967 & n27969 ) ;
  assign n27971 = n14530 ^ n5348 ^ 1'b0 ;
  assign n27972 = n27971 ^ n18975 ^ n16096 ;
  assign n27973 = n27972 ^ n15349 ^ 1'b0 ;
  assign n27974 = n7392 | n27973 ;
  assign n27975 = n984 | n15826 ;
  assign n27976 = n6285 & n27975 ;
  assign n27977 = n27976 ^ n3446 ^ 1'b0 ;
  assign n27978 = n13951 ^ n4438 ^ n1937 ;
  assign n27981 = n481 | n2422 ;
  assign n27982 = n6040 | n27981 ;
  assign n27983 = ~n5053 & n8733 ;
  assign n27984 = n10079 & n27983 ;
  assign n27985 = ( n7366 & ~n27982 ) | ( n7366 & n27984 ) | ( ~n27982 & n27984 ) ;
  assign n27979 = n5226 ^ n430 ^ 1'b0 ;
  assign n27980 = n25487 & n27979 ;
  assign n27986 = n27985 ^ n27980 ^ 1'b0 ;
  assign n27987 = n14646 ^ n923 ^ 1'b0 ;
  assign n27993 = ~n18954 & n26013 ;
  assign n27994 = ~n16679 & n27993 ;
  assign n27988 = ~n7779 & n14102 ;
  assign n27989 = n27988 ^ n5069 ^ 1'b0 ;
  assign n27990 = n14417 & ~n27989 ;
  assign n27991 = ~n6115 & n27990 ;
  assign n27992 = ( n3934 & ~n11718 ) | ( n3934 & n27991 ) | ( ~n11718 & n27991 ) ;
  assign n27995 = n27994 ^ n27992 ^ 1'b0 ;
  assign n27996 = n8203 ^ n6711 ^ 1'b0 ;
  assign n27997 = n18893 | n27996 ;
  assign n28002 = n16858 ^ n16203 ^ 1'b0 ;
  assign n28003 = n28002 ^ n6109 ^ 1'b0 ;
  assign n27998 = n6759 ^ n4688 ^ n2664 ;
  assign n27999 = n14332 | n27998 ;
  assign n28000 = n4140 | n27999 ;
  assign n28001 = ~n496 & n28000 ;
  assign n28004 = n28003 ^ n28001 ^ 1'b0 ;
  assign n28005 = ~n3593 & n20230 ;
  assign n28006 = n28005 ^ n747 ^ 1'b0 ;
  assign n28007 = ~n18472 & n28006 ;
  assign n28008 = n25635 ^ n13783 ^ 1'b0 ;
  assign n28009 = ~n12936 & n28008 ;
  assign n28010 = n16343 ^ n11365 ^ n4500 ;
  assign n28011 = n19289 ^ n5866 ^ 1'b0 ;
  assign n28012 = n24984 | n28011 ;
  assign n28013 = n22329 ^ n4056 ^ 1'b0 ;
  assign n28014 = ~n9759 & n12661 ;
  assign n28015 = n10347 & ~n28014 ;
  assign n28016 = ~n6384 & n28015 ;
  assign n28017 = n5914 & n12351 ;
  assign n28018 = ( ~n20078 & n21352 ) | ( ~n20078 & n28017 ) | ( n21352 & n28017 ) ;
  assign n28023 = ~n2387 & n25610 ;
  assign n28024 = n28023 ^ n7801 ^ n4584 ;
  assign n28020 = n5424 & ~n12664 ;
  assign n28019 = ~n7342 & n14247 ;
  assign n28021 = n28020 ^ n28019 ^ n3590 ;
  assign n28022 = ~n8262 & n28021 ;
  assign n28025 = n28024 ^ n28022 ^ 1'b0 ;
  assign n28026 = n7752 ^ n4541 ^ 1'b0 ;
  assign n28027 = n28026 ^ n14446 ^ 1'b0 ;
  assign n28028 = n28025 & n28027 ;
  assign n28029 = ( n1553 & ~n10922 ) | ( n1553 & n27159 ) | ( ~n10922 & n27159 ) ;
  assign n28030 = n3362 | n28029 ;
  assign n28031 = ~n22890 & n23579 ;
  assign n28032 = n21471 ^ n6157 ^ 1'b0 ;
  assign n28033 = n28031 & ~n28032 ;
  assign n28034 = n28033 ^ n2368 ^ 1'b0 ;
  assign n28037 = ( n1728 & n11751 ) | ( n1728 & n19886 ) | ( n11751 & n19886 ) ;
  assign n28038 = n28037 ^ n10564 ^ 1'b0 ;
  assign n28039 = n16781 | n28038 ;
  assign n28035 = n1952 & n8748 ;
  assign n28036 = ~n996 & n28035 ;
  assign n28040 = n28039 ^ n28036 ^ 1'b0 ;
  assign n28041 = n15366 ^ n3177 ^ 1'b0 ;
  assign n28042 = n8020 & n28041 ;
  assign n28043 = ~n17919 & n28042 ;
  assign n28044 = n28043 ^ n667 ^ 1'b0 ;
  assign n28045 = n28044 ^ n1972 ^ 1'b0 ;
  assign n28046 = n8808 & ~n28045 ;
  assign n28047 = n1150 & ~n2124 ;
  assign n28048 = n28047 ^ n3770 ^ 1'b0 ;
  assign n28049 = n27004 | n28048 ;
  assign n28050 = n19472 | n28049 ;
  assign n28051 = n23596 | n28050 ;
  assign n28052 = ( n125 & ~n10950 ) | ( n125 & n14418 ) | ( ~n10950 & n14418 ) ;
  assign n28053 = n28052 ^ n23538 ^ n19092 ;
  assign n28054 = n11372 & ~n27759 ;
  assign n28055 = n6222 & n13136 ;
  assign n28056 = n2451 & n28055 ;
  assign n28057 = n6460 ^ n494 ^ 1'b0 ;
  assign n28058 = n3826 & n28057 ;
  assign n28059 = n28058 ^ n19985 ^ 1'b0 ;
  assign n28060 = ~n8070 & n22223 ;
  assign n28062 = n21504 ^ n3162 ^ 1'b0 ;
  assign n28063 = n28062 ^ n20339 ^ n6383 ;
  assign n28061 = ~n10054 & n13907 ;
  assign n28064 = n28063 ^ n28061 ^ 1'b0 ;
  assign n28065 = ~n15441 & n15746 ;
  assign n28067 = n9085 ^ n7974 ^ 1'b0 ;
  assign n28068 = n6304 & ~n28067 ;
  assign n28069 = n11762 & n28068 ;
  assign n28070 = n28069 ^ n14646 ^ 1'b0 ;
  assign n28071 = n28070 ^ n13397 ^ 1'b0 ;
  assign n28066 = n19280 ^ n11923 ^ n11652 ;
  assign n28072 = n28071 ^ n28066 ^ n16158 ;
  assign n28073 = n6776 ^ n741 ^ 1'b0 ;
  assign n28074 = n4104 & n14886 ;
  assign n28075 = ~n25624 & n28074 ;
  assign n28077 = n1078 & n21453 ;
  assign n28076 = ~n7425 & n14392 ;
  assign n28078 = n28077 ^ n28076 ^ 1'b0 ;
  assign n28079 = n4941 & n14164 ;
  assign n28080 = ( n14678 & n28078 ) | ( n14678 & ~n28079 ) | ( n28078 & ~n28079 ) ;
  assign n28083 = n8681 | n21193 ;
  assign n28084 = ~n4469 & n9676 ;
  assign n28085 = n8259 | n12945 ;
  assign n28086 = ( n11558 & n25738 ) | ( n11558 & n28085 ) | ( n25738 & n28085 ) ;
  assign n28087 = ( n11480 & ~n28084 ) | ( n11480 & n28086 ) | ( ~n28084 & n28086 ) ;
  assign n28088 = n28083 & n28087 ;
  assign n28081 = n7140 & n11084 ;
  assign n28082 = n28081 ^ n23721 ^ n6389 ;
  assign n28089 = n28088 ^ n28082 ^ 1'b0 ;
  assign n28090 = n9279 & n17669 ;
  assign n28091 = n28090 ^ n21146 ^ n2911 ;
  assign n28092 = n10734 ^ n4249 ^ 1'b0 ;
  assign n28093 = ~n5458 & n28092 ;
  assign n28094 = ~n28091 & n28093 ;
  assign n28095 = n829 & n28094 ;
  assign n28096 = ( ~n2284 & n3979 ) | ( ~n2284 & n4115 ) | ( n3979 & n4115 ) ;
  assign n28097 = n28096 ^ n14247 ^ n8733 ;
  assign n28098 = ( n432 & ~n7320 ) | ( n432 & n28097 ) | ( ~n7320 & n28097 ) ;
  assign n28099 = n1450 & n11260 ;
  assign n28100 = n126 | n7377 ;
  assign n28101 = ( ~n473 & n2216 ) | ( ~n473 & n28100 ) | ( n2216 & n28100 ) ;
  assign n28102 = n2541 & n8474 ;
  assign n28103 = n11000 & n28102 ;
  assign n28104 = n22110 ^ n21776 ^ 1'b0 ;
  assign n28105 = ~n13298 & n28104 ;
  assign n28106 = ~n654 & n9805 ;
  assign n28107 = n8039 & n28106 ;
  assign n28108 = n12046 & ~n28107 ;
  assign n28109 = n28108 ^ n20289 ^ 1'b0 ;
  assign n28110 = n9135 & n11120 ;
  assign n28111 = ~n5094 & n28110 ;
  assign n28112 = n5042 | n28111 ;
  assign n28113 = n5127 ^ n4799 ^ 1'b0 ;
  assign n28114 = n20050 & n28113 ;
  assign n28115 = n12080 ^ n11273 ^ 1'b0 ;
  assign n28116 = n28114 & n28115 ;
  assign n28117 = n5844 & n13670 ;
  assign n28118 = ( n143 & ~n8659 ) | ( n143 & n19097 ) | ( ~n8659 & n19097 ) ;
  assign n28119 = n28118 ^ n15184 ^ 1'b0 ;
  assign n28120 = n1031 | n14026 ;
  assign n28121 = n3925 & n28120 ;
  assign n28122 = ~n1630 & n5102 ;
  assign n28123 = n22658 ^ n11435 ^ 1'b0 ;
  assign n28124 = n13449 ^ n4240 ^ 1'b0 ;
  assign n28125 = n28123 & n28124 ;
  assign n28126 = n2987 | n12589 ;
  assign n28127 = n962 | n23079 ;
  assign n28128 = n28127 ^ n5479 ^ 1'b0 ;
  assign n28129 = n28128 ^ n563 ^ 1'b0 ;
  assign n28130 = ~n24615 & n28129 ;
  assign n28131 = n28130 ^ n9474 ^ n5570 ;
  assign n28132 = n6569 ^ n1083 ^ 1'b0 ;
  assign n28133 = ( ~n2797 & n20383 ) | ( ~n2797 & n28132 ) | ( n20383 & n28132 ) ;
  assign n28134 = ~n17402 & n18566 ;
  assign n28135 = n28134 ^ n27267 ^ 1'b0 ;
  assign n28136 = ( ~n5930 & n19294 ) | ( ~n5930 & n26694 ) | ( n19294 & n26694 ) ;
  assign n28137 = ~n3308 & n14190 ;
  assign n28138 = n28137 ^ n1102 ^ 1'b0 ;
  assign n28139 = n28138 ^ n24605 ^ 1'b0 ;
  assign n28140 = n13240 ^ n1552 ^ 1'b0 ;
  assign n28141 = ( n2397 & ~n28139 ) | ( n2397 & n28140 ) | ( ~n28139 & n28140 ) ;
  assign n28142 = n7704 & n8165 ;
  assign n28143 = n28142 ^ n22622 ^ n11225 ;
  assign n28144 = n27843 | n28143 ;
  assign n28145 = n14386 | n28144 ;
  assign n28146 = n676 | n11036 ;
  assign n28149 = n19616 ^ n17614 ^ n8467 ;
  assign n28147 = n18562 ^ n18109 ^ n17079 ;
  assign n28148 = ~n27040 & n28147 ;
  assign n28150 = n28149 ^ n28148 ^ 1'b0 ;
  assign n28151 = ( ~n3090 & n13078 ) | ( ~n3090 & n19909 ) | ( n13078 & n19909 ) ;
  assign n28152 = n5716 & ~n11602 ;
  assign n28153 = n15910 & n28152 ;
  assign n28154 = n28153 ^ n27596 ^ n16981 ;
  assign n28155 = n12404 ^ n3773 ^ n903 ;
  assign n28156 = n28155 ^ n26310 ^ n12556 ;
  assign n28157 = n16605 ^ n9804 ^ 1'b0 ;
  assign n28158 = n20394 ^ n101 ^ 1'b0 ;
  assign n28159 = n28158 ^ n10586 ^ 1'b0 ;
  assign n28160 = n2416 ^ n381 ^ 1'b0 ;
  assign n28161 = n28160 ^ n11341 ^ 1'b0 ;
  assign n28162 = n14158 | n28161 ;
  assign n28163 = n10446 ^ n4858 ^ 1'b0 ;
  assign n28164 = n28162 | n28163 ;
  assign n28165 = n10408 & ~n28164 ;
  assign n28166 = n7629 & n19159 ;
  assign n28167 = n28166 ^ n28014 ^ 1'b0 ;
  assign n28168 = n28167 ^ n863 ^ 1'b0 ;
  assign n28169 = n28168 ^ n14854 ^ 1'b0 ;
  assign n28170 = n1965 | n6301 ;
  assign n28171 = n826 & n998 ;
  assign n28172 = ~n2672 & n2922 ;
  assign n28173 = n9898 & n28172 ;
  assign n28174 = n28173 ^ n15332 ^ n7650 ;
  assign n28175 = n28174 ^ n23571 ^ n18017 ;
  assign n28176 = n8684 & ~n19613 ;
  assign n28177 = n22176 ^ n9852 ^ 1'b0 ;
  assign n28178 = n28177 ^ n4892 ^ n3310 ;
  assign n28179 = n5675 ^ n1122 ^ 1'b0 ;
  assign n28180 = n19529 | n28179 ;
  assign n28181 = ( n1980 & ~n3807 ) | ( n1980 & n10950 ) | ( ~n3807 & n10950 ) ;
  assign n28182 = n28181 ^ n5885 ^ 1'b0 ;
  assign n28183 = n28182 ^ n8755 ^ 1'b0 ;
  assign n28184 = ~n2122 & n11091 ;
  assign n28185 = n28184 ^ n3985 ^ 1'b0 ;
  assign n28186 = ~n10240 & n28185 ;
  assign n28187 = n8051 & n28186 ;
  assign n28188 = ~n2082 & n18889 ;
  assign n28189 = ~n4298 & n28188 ;
  assign n28190 = n28189 ^ n6445 ^ 1'b0 ;
  assign n28191 = n14136 ^ n4004 ^ n1143 ;
  assign n28192 = n28191 ^ n7250 ^ 1'b0 ;
  assign n28193 = ~n26728 & n28192 ;
  assign n28194 = n4068 | n11946 ;
  assign n28195 = n28194 ^ n465 ^ 1'b0 ;
  assign n28196 = n6593 & ~n28195 ;
  assign n28197 = n20582 & n28196 ;
  assign n28198 = n12021 & n19751 ;
  assign n28199 = n28198 ^ n14980 ^ 1'b0 ;
  assign n28200 = n28199 ^ n20235 ^ n2951 ;
  assign n28201 = ~n10035 & n28200 ;
  assign n28202 = n16355 & n28201 ;
  assign n28203 = n21749 ^ n11844 ^ n5353 ;
  assign n28204 = ( n20130 & n25160 ) | ( n20130 & ~n28203 ) | ( n25160 & ~n28203 ) ;
  assign n28205 = n381 & ~n8017 ;
  assign n28206 = ~n7943 & n28205 ;
  assign n28207 = n28206 ^ n24924 ^ 1'b0 ;
  assign n28208 = n3778 & n28207 ;
  assign n28209 = n3567 | n3760 ;
  assign n28210 = n28209 ^ n6713 ^ 1'b0 ;
  assign n28211 = n16620 & ~n28210 ;
  assign n28215 = n11839 & n22394 ;
  assign n28212 = n8168 ^ n6059 ^ n578 ;
  assign n28213 = n4212 | n16129 ;
  assign n28214 = n28212 & n28213 ;
  assign n28216 = n28215 ^ n28214 ^ 1'b0 ;
  assign n28217 = n2969 & n11184 ;
  assign n28218 = n3326 ^ n2268 ^ 1'b0 ;
  assign n28219 = n21713 & n28218 ;
  assign n28220 = n17390 ^ n10450 ^ 1'b0 ;
  assign n28221 = ~n12779 & n28220 ;
  assign n28222 = n5639 & ~n10695 ;
  assign n28223 = n28222 ^ n6414 ^ 1'b0 ;
  assign n28224 = n3269 | n28223 ;
  assign n28225 = n8041 | n28224 ;
  assign n28226 = n19493 ^ n12180 ^ 1'b0 ;
  assign n28227 = n8028 & n28226 ;
  assign n28228 = ~n4187 & n5393 ;
  assign n28229 = n804 & n28228 ;
  assign n28230 = n17761 ^ n7046 ^ n4188 ;
  assign n28231 = n9794 & ~n28230 ;
  assign n28232 = n13717 & ~n28231 ;
  assign n28233 = n28229 & n28232 ;
  assign n28234 = n3869 ^ n2728 ^ 1'b0 ;
  assign n28235 = n14965 ^ n6003 ^ 1'b0 ;
  assign n28236 = ( n23376 & n27875 ) | ( n23376 & n28235 ) | ( n27875 & n28235 ) ;
  assign n28237 = ( n14465 & n15671 ) | ( n14465 & n28236 ) | ( n15671 & n28236 ) ;
  assign n28238 = n28237 ^ n18239 ^ 1'b0 ;
  assign n28239 = n19185 & n27293 ;
  assign n28240 = n9573 & n28239 ;
  assign n28241 = n10230 ^ n5791 ^ n2118 ;
  assign n28242 = n11832 ^ n7621 ^ 1'b0 ;
  assign n28243 = n3385 & ~n28242 ;
  assign n28244 = n28243 ^ n3128 ^ 1'b0 ;
  assign n28245 = n4066 | n26840 ;
  assign n28246 = ~n4096 & n18911 ;
  assign n28247 = n2951 & n8832 ;
  assign n28248 = n7572 ^ n3730 ^ 1'b0 ;
  assign n28249 = n7599 & n27171 ;
  assign n28250 = n9936 & n28249 ;
  assign n28251 = n17473 | n28250 ;
  assign n28252 = n17096 ^ n10971 ^ 1'b0 ;
  assign n28253 = ( n2436 & n17378 ) | ( n2436 & n28252 ) | ( n17378 & n28252 ) ;
  assign n28254 = n17986 ^ n8923 ^ 1'b0 ;
  assign n28256 = ~n10744 & n19234 ;
  assign n28257 = n28256 ^ n11980 ^ 1'b0 ;
  assign n28255 = n5771 ^ n3755 ^ 1'b0 ;
  assign n28258 = n28257 ^ n28255 ^ 1'b0 ;
  assign n28259 = n28254 | n28258 ;
  assign n28260 = n8654 ^ n4368 ^ 1'b0 ;
  assign n28261 = n7621 & n28260 ;
  assign n28262 = n4404 | n26220 ;
  assign n28263 = n23976 ^ n14156 ^ 1'b0 ;
  assign n28264 = ~n172 & n4994 ;
  assign n28265 = n28263 & n28264 ;
  assign n28266 = ~n16096 & n18063 ;
  assign n28267 = n28266 ^ n13857 ^ 1'b0 ;
  assign n28268 = n1929 & ~n8480 ;
  assign n28269 = n28268 ^ n2569 ^ 1'b0 ;
  assign n28271 = n5994 & ~n28230 ;
  assign n28272 = ~n9103 & n28271 ;
  assign n28273 = n28174 & n28272 ;
  assign n28270 = n22448 ^ n3495 ^ 1'b0 ;
  assign n28274 = n28273 ^ n28270 ^ 1'b0 ;
  assign n28275 = n26916 | n28274 ;
  assign n28276 = n18687 & ~n27294 ;
  assign n28277 = ~n7489 & n28276 ;
  assign n28278 = n7407 & ~n20934 ;
  assign n28279 = n6441 ^ n4402 ^ 1'b0 ;
  assign n28280 = n1945 | n28279 ;
  assign n28281 = n28280 ^ n23650 ^ 1'b0 ;
  assign n28282 = n28281 ^ n14967 ^ 1'b0 ;
  assign n28283 = n2898 | n9049 ;
  assign n28284 = n28283 ^ n11595 ^ 1'b0 ;
  assign n28285 = n28282 & ~n28284 ;
  assign n28286 = ~n706 & n16329 ;
  assign n28287 = ~n2740 & n9463 ;
  assign n28288 = n10062 & n28287 ;
  assign n28289 = n10989 & ~n15176 ;
  assign n28290 = ~n14013 & n28289 ;
  assign n28291 = n8429 & ~n28290 ;
  assign n28292 = n739 | n4237 ;
  assign n28293 = n28292 ^ n6753 ^ 1'b0 ;
  assign n28294 = n28291 & ~n28293 ;
  assign n28295 = n16094 & ~n17843 ;
  assign n28296 = n11802 | n18583 ;
  assign n28297 = n28296 ^ n11153 ^ 1'b0 ;
  assign n28298 = n20173 | n28297 ;
  assign n28299 = n15472 | n28298 ;
  assign n28300 = n9739 ^ n2760 ^ 1'b0 ;
  assign n28301 = ~n17518 & n28300 ;
  assign n28302 = ~n23186 & n28301 ;
  assign n28303 = n4712 & n18002 ;
  assign n28304 = ~n14452 & n28303 ;
  assign n28310 = n12075 ^ n1506 ^ 1'b0 ;
  assign n28311 = n8824 & ~n28310 ;
  assign n28307 = n9220 ^ n3119 ^ 1'b0 ;
  assign n28305 = n13418 ^ n9192 ^ 1'b0 ;
  assign n28306 = ~n3286 & n28305 ;
  assign n28308 = n28307 ^ n28306 ^ 1'b0 ;
  assign n28309 = n6901 & n28308 ;
  assign n28312 = n28311 ^ n28309 ^ 1'b0 ;
  assign n28313 = n15046 ^ n6674 ^ 1'b0 ;
  assign n28314 = n16060 & n28313 ;
  assign n28315 = n4717 & ~n22781 ;
  assign n28316 = n13056 & n28315 ;
  assign n28317 = n5068 ^ n4275 ^ 1'b0 ;
  assign n28318 = ~n28316 & n28317 ;
  assign n28319 = n46 & n1523 ;
  assign n28320 = ( n3632 & n7778 ) | ( n3632 & ~n25658 ) | ( n7778 & ~n25658 ) ;
  assign n28321 = ( ~n776 & n2427 ) | ( ~n776 & n3135 ) | ( n2427 & n3135 ) ;
  assign n28322 = n8149 & ~n20911 ;
  assign n28323 = n6322 & n28322 ;
  assign n28324 = n28323 ^ n11254 ^ 1'b0 ;
  assign n28325 = ( n6598 & n28321 ) | ( n6598 & n28324 ) | ( n28321 & n28324 ) ;
  assign n28326 = n10737 ^ n6858 ^ 1'b0 ;
  assign n28327 = n8555 | n10430 ;
  assign n28328 = n28327 ^ n5127 ^ 1'b0 ;
  assign n28329 = n9107 & ~n28328 ;
  assign n28331 = ~n14658 & n19904 ;
  assign n28330 = n15056 & n27903 ;
  assign n28332 = n28331 ^ n28330 ^ 1'b0 ;
  assign n28333 = ( n6096 & n8105 ) | ( n6096 & ~n13695 ) | ( n8105 & ~n13695 ) ;
  assign n28334 = n28333 ^ n16546 ^ 1'b0 ;
  assign n28335 = ( n14763 & n27297 ) | ( n14763 & n28334 ) | ( n27297 & n28334 ) ;
  assign n28336 = n14744 & ~n21363 ;
  assign n28337 = n19350 & ~n26297 ;
  assign n28338 = n4637 ^ n1674 ^ 1'b0 ;
  assign n28339 = ~n8119 & n28338 ;
  assign n28340 = n28339 ^ n13325 ^ 1'b0 ;
  assign n28341 = n518 | n28340 ;
  assign n28342 = n25087 ^ n21723 ^ 1'b0 ;
  assign n28343 = n21836 ^ n1401 ^ 1'b0 ;
  assign n28344 = n28342 & n28343 ;
  assign n28345 = n10282 ^ n2358 ^ 1'b0 ;
  assign n28346 = ~n4222 & n28345 ;
  assign n28347 = n28346 ^ n9313 ^ 1'b0 ;
  assign n28348 = ( n8640 & n16207 ) | ( n8640 & n28347 ) | ( n16207 & n28347 ) ;
  assign n28349 = n17608 ^ n1592 ^ n813 ;
  assign n28350 = n4177 & n28349 ;
  assign n28351 = n9397 ^ n1000 ^ 1'b0 ;
  assign n28352 = n12925 & n28351 ;
  assign n28353 = n8980 ^ n5483 ^ 1'b0 ;
  assign n28354 = n28352 & ~n28353 ;
  assign n28355 = n5494 ^ n4052 ^ 1'b0 ;
  assign n28356 = ( n13020 & ~n15976 ) | ( n13020 & n28355 ) | ( ~n15976 & n28355 ) ;
  assign n28357 = n28356 ^ n17199 ^ 1'b0 ;
  assign n28358 = n11864 ^ n6452 ^ 1'b0 ;
  assign n28362 = n5168 ^ n842 ^ 1'b0 ;
  assign n28363 = n7975 & ~n28362 ;
  assign n28364 = ~n9941 & n28363 ;
  assign n28360 = n14975 ^ n11567 ^ 1'b0 ;
  assign n28361 = n11964 & ~n28360 ;
  assign n28365 = n28364 ^ n28361 ^ 1'b0 ;
  assign n28359 = n7017 & ~n18234 ;
  assign n28366 = n28365 ^ n28359 ^ n4315 ;
  assign n28367 = n21506 ^ n179 ^ 1'b0 ;
  assign n28368 = n22705 & ~n28367 ;
  assign n28369 = n28063 & n28368 ;
  assign n28370 = n28369 ^ n12826 ^ 1'b0 ;
  assign n28371 = n22883 ^ n19893 ^ n7710 ;
  assign n28372 = n8607 ^ n5269 ^ 1'b0 ;
  assign n28373 = n250 | n28372 ;
  assign n28374 = n28373 ^ n24727 ^ n1264 ;
  assign n28375 = n3003 & n7389 ;
  assign n28376 = n17580 & n28375 ;
  assign n28377 = n21156 & n25479 ;
  assign n28378 = n466 & n28377 ;
  assign n28379 = n19292 & ~n23796 ;
  assign n28380 = n28379 ^ n6320 ^ 1'b0 ;
  assign n28381 = n6183 & n17719 ;
  assign n28382 = n3157 & ~n18835 ;
  assign n28383 = ~n7008 & n7613 ;
  assign n28384 = n28383 ^ n710 ^ 1'b0 ;
  assign n28385 = ( n24236 & n26146 ) | ( n24236 & ~n28384 ) | ( n26146 & ~n28384 ) ;
  assign n28386 = n9550 ^ n5552 ^ 1'b0 ;
  assign n28387 = n7322 & n23532 ;
  assign n28388 = n28387 ^ n24996 ^ 1'b0 ;
  assign n28389 = n9984 ^ n3725 ^ 1'b0 ;
  assign n28390 = n20534 & ~n28389 ;
  assign n28391 = n28390 ^ n15903 ^ 1'b0 ;
  assign n28392 = n17900 ^ n2117 ^ 1'b0 ;
  assign n28393 = n2911 & n11161 ;
  assign n28394 = n27064 ^ n6576 ^ 1'b0 ;
  assign n28395 = ~n6510 & n15830 ;
  assign n28396 = n28394 & n28395 ;
  assign n28397 = n28393 & ~n28396 ;
  assign n28398 = n2747 & n12754 ;
  assign n28399 = ( n11644 & n28397 ) | ( n11644 & ~n28398 ) | ( n28397 & ~n28398 ) ;
  assign n28400 = n5279 ^ n1308 ^ 1'b0 ;
  assign n28401 = n9173 & ~n28400 ;
  assign n28402 = ~n16084 & n28401 ;
  assign n28403 = n23686 ^ n14222 ^ 1'b0 ;
  assign n28404 = n23225 & ~n28403 ;
  assign n28405 = ~n11751 & n28404 ;
  assign n28406 = n12586 ^ n9036 ^ 1'b0 ;
  assign n28407 = n16575 & n28406 ;
  assign n28408 = n8931 ^ n5656 ^ 1'b0 ;
  assign n28409 = n3819 & n15632 ;
  assign n28410 = n2190 & n28409 ;
  assign n28411 = ~n19004 & n23252 ;
  assign n28412 = n28411 ^ n10519 ^ 1'b0 ;
  assign n28414 = ~n15134 & n16047 ;
  assign n28415 = n27187 | n28414 ;
  assign n28416 = n28415 ^ n1630 ^ 1'b0 ;
  assign n28413 = n22038 | n23860 ;
  assign n28417 = n28416 ^ n28413 ^ 1'b0 ;
  assign n28418 = ~n5627 & n12578 ;
  assign n28419 = n28418 ^ n5783 ^ 1'b0 ;
  assign n28420 = n19205 ^ n3573 ^ 1'b0 ;
  assign n28421 = n10430 | n28420 ;
  assign n28422 = n28421 ^ n806 ^ 1'b0 ;
  assign n28423 = n28419 & ~n28422 ;
  assign n28424 = n18579 & n22580 ;
  assign n28425 = n9694 ^ n1507 ^ n688 ;
  assign n28426 = n18518 & n21212 ;
  assign n28427 = n28425 & n28426 ;
  assign n28428 = n777 & ~n15046 ;
  assign n28429 = ~n13346 & n17923 ;
  assign n28430 = n28428 & n28429 ;
  assign n28431 = ~n28427 & n28430 ;
  assign n28432 = n20216 ^ n13849 ^ n12093 ;
  assign n28433 = ( ~n7810 & n17675 ) | ( ~n7810 & n28432 ) | ( n17675 & n28432 ) ;
  assign n28435 = n95 | n545 ;
  assign n28434 = n2504 & ~n5870 ;
  assign n28436 = n28435 ^ n28434 ^ 1'b0 ;
  assign n28437 = n1446 & ~n28436 ;
  assign n28438 = n28437 ^ n18680 ^ 1'b0 ;
  assign n28439 = n10243 & ~n28438 ;
  assign n28440 = n28439 ^ n2425 ^ 1'b0 ;
  assign n28441 = ~n6535 & n15145 ;
  assign n28442 = n11059 ^ n3196 ^ 1'b0 ;
  assign n28443 = n20136 & n28442 ;
  assign n28444 = n28443 ^ n19189 ^ 1'b0 ;
  assign n28445 = n15190 & n15341 ;
  assign n28446 = n28445 ^ n2414 ^ 1'b0 ;
  assign n28447 = n5250 | n28446 ;
  assign n28448 = n21781 ^ n20815 ^ 1'b0 ;
  assign n28449 = ~n22488 & n28448 ;
  assign n28450 = ~n10785 & n28449 ;
  assign n28451 = n15850 ^ n7216 ^ 1'b0 ;
  assign n28453 = ~n5051 & n8725 ;
  assign n28452 = n14086 | n16190 ;
  assign n28454 = n28453 ^ n28452 ^ 1'b0 ;
  assign n28455 = n28454 ^ n16236 ^ 1'b0 ;
  assign n28456 = ( n7711 & ~n11250 ) | ( n7711 & n17608 ) | ( ~n11250 & n17608 ) ;
  assign n28457 = ( n4769 & ~n11788 ) | ( n4769 & n11955 ) | ( ~n11788 & n11955 ) ;
  assign n28458 = ( n13007 & ~n28456 ) | ( n13007 & n28457 ) | ( ~n28456 & n28457 ) ;
  assign n28459 = n12298 & ~n19775 ;
  assign n28460 = n5716 & ~n28459 ;
  assign n28461 = n8413 & n26570 ;
  assign n28462 = n12460 & n28461 ;
  assign n28463 = ~n3580 & n5484 ;
  assign n28464 = n28463 ^ n6032 ^ 1'b0 ;
  assign n28465 = n28464 ^ n8750 ^ 1'b0 ;
  assign n28466 = n3517 & n10356 ;
  assign n28467 = n28466 ^ n17760 ^ 1'b0 ;
  assign n28471 = n15730 ^ n4487 ^ n2955 ;
  assign n28468 = n7970 ^ n7433 ^ n3574 ;
  assign n28469 = n7828 & ~n28468 ;
  assign n28470 = ~n27011 & n28469 ;
  assign n28472 = n28471 ^ n28470 ^ n27975 ;
  assign n28473 = ~n14658 & n28472 ;
  assign n28474 = n24819 ^ n7091 ^ 1'b0 ;
  assign n28475 = n1612 & n28474 ;
  assign n28476 = n19829 ^ n1812 ^ 1'b0 ;
  assign n28477 = n8558 ^ n4477 ^ 1'b0 ;
  assign n28478 = n777 & ~n28477 ;
  assign n28479 = n4488 | n16910 ;
  assign n28480 = n3060 | n28479 ;
  assign n28481 = ~n28478 & n28480 ;
  assign n28482 = n24124 ^ n22271 ^ 1'b0 ;
  assign n28483 = n25824 ^ n17589 ^ 1'b0 ;
  assign n28485 = n2775 & n15756 ;
  assign n28486 = ~n22309 & n28485 ;
  assign n28484 = n9230 & n12028 ;
  assign n28487 = n28486 ^ n28484 ^ 1'b0 ;
  assign n28488 = n26069 ^ n8456 ^ 1'b0 ;
  assign n28489 = n12641 | n28488 ;
  assign n28490 = n9057 ^ n8848 ^ 1'b0 ;
  assign n28491 = n8885 & ~n28490 ;
  assign n28492 = n19238 ^ n10118 ^ n7468 ;
  assign n28493 = n28492 ^ n835 ^ 1'b0 ;
  assign n28494 = n27371 & n28493 ;
  assign n28495 = n3750 & n14879 ;
  assign n28496 = n28495 ^ n16394 ^ n3630 ;
  assign n28497 = n8356 | n24553 ;
  assign n28498 = n28497 ^ n1490 ^ 1'b0 ;
  assign n28499 = ( n6122 & ~n10999 ) | ( n6122 & n28498 ) | ( ~n10999 & n28498 ) ;
  assign n28500 = n15172 ^ n4994 ^ 1'b0 ;
  assign n28502 = n2589 & n19979 ;
  assign n28503 = ~n4093 & n28502 ;
  assign n28501 = ( n4131 & n10688 ) | ( n4131 & n16925 ) | ( n10688 & n16925 ) ;
  assign n28504 = n28503 ^ n28501 ^ 1'b0 ;
  assign n28505 = n28500 & ~n28504 ;
  assign n28506 = n2313 & ~n10724 ;
  assign n28507 = ( ~n18053 & n20118 ) | ( ~n18053 & n20911 ) | ( n20118 & n20911 ) ;
  assign n28508 = ( n5651 & ~n16694 ) | ( n5651 & n28507 ) | ( ~n16694 & n28507 ) ;
  assign n28509 = n5768 & ~n11453 ;
  assign n28510 = n1448 & n28509 ;
  assign n28511 = n28510 ^ n9680 ^ n4918 ;
  assign n28512 = ( n4848 & n27149 ) | ( n4848 & n28511 ) | ( n27149 & n28511 ) ;
  assign n28513 = n8119 ^ n5596 ^ 1'b0 ;
  assign n28514 = n28512 & ~n28513 ;
  assign n28515 = n28448 ^ n18832 ^ n7585 ;
  assign n28516 = n21262 ^ n18857 ^ 1'b0 ;
  assign n28517 = ~n7270 & n28516 ;
  assign n28518 = n11306 & n24772 ;
  assign n28519 = n12113 ^ n10311 ^ 1'b0 ;
  assign n28520 = n4471 | n28519 ;
  assign n28525 = n7196 & ~n9613 ;
  assign n28521 = n17966 ^ n1089 ^ 1'b0 ;
  assign n28522 = n6415 & n28521 ;
  assign n28523 = n28522 ^ n6743 ^ 1'b0 ;
  assign n28524 = ~n4275 & n28523 ;
  assign n28526 = n28525 ^ n28524 ^ n742 ;
  assign n28527 = n28526 ^ n18779 ^ n5645 ;
  assign n28528 = n11860 ^ n10010 ^ 1'b0 ;
  assign n28529 = ~n78 & n28528 ;
  assign n28530 = ~n28527 & n28529 ;
  assign n28531 = n28530 ^ n10062 ^ 1'b0 ;
  assign n28532 = n1133 ^ n811 ^ 1'b0 ;
  assign n28533 = ~n17542 & n28532 ;
  assign n28534 = n13708 ^ n11254 ^ n351 ;
  assign n28535 = n28534 ^ n2849 ^ 1'b0 ;
  assign n28536 = n27033 ^ n17488 ^ 1'b0 ;
  assign n28537 = n11083 | n26473 ;
  assign n28538 = n11250 & ~n28537 ;
  assign n28539 = n28536 & n28538 ;
  assign n28540 = ~n563 & n15161 ;
  assign n28541 = n27138 ^ n1666 ^ 1'b0 ;
  assign n28542 = n6128 | n10164 ;
  assign n28543 = n28542 ^ n1446 ^ 1'b0 ;
  assign n28544 = n28543 ^ n13842 ^ 1'b0 ;
  assign n28545 = ~n21724 & n28544 ;
  assign n28546 = ~n6933 & n28545 ;
  assign n28547 = n28546 ^ n13063 ^ 1'b0 ;
  assign n28548 = n14616 ^ n10543 ^ n5298 ;
  assign n28549 = n28548 ^ n17999 ^ 1'b0 ;
  assign n28550 = ~n10339 & n28549 ;
  assign n28552 = ~n3375 & n9388 ;
  assign n28553 = ~n9388 & n28552 ;
  assign n28551 = n8206 & ~n8764 ;
  assign n28554 = n28553 ^ n28551 ^ 1'b0 ;
  assign n28555 = n2054 | n2676 ;
  assign n28556 = n2054 & ~n28555 ;
  assign n28557 = ~n640 & n28556 ;
  assign n28558 = ~n20830 & n28557 ;
  assign n28559 = ( n26978 & n28554 ) | ( n26978 & n28558 ) | ( n28554 & n28558 ) ;
  assign n28560 = n3768 & n8972 ;
  assign n28561 = n7078 & n8874 ;
  assign n28562 = n6872 | n23734 ;
  assign n28563 = n28562 ^ n25279 ^ 1'b0 ;
  assign n28564 = ~n6720 & n10382 ;
  assign n28565 = n5818 & ~n28564 ;
  assign n28566 = n6568 ^ n3293 ^ 1'b0 ;
  assign n28567 = n24531 & ~n28566 ;
  assign n28568 = n28567 ^ n26770 ^ 1'b0 ;
  assign n28569 = n14413 & n22722 ;
  assign n28570 = ~n2958 & n28569 ;
  assign n28571 = ( n16666 & ~n24217 ) | ( n16666 & n26799 ) | ( ~n24217 & n26799 ) ;
  assign n28572 = n2550 | n13825 ;
  assign n28573 = n6020 & ~n28572 ;
  assign n28574 = n14600 & n28573 ;
  assign n28575 = n526 & ~n2603 ;
  assign n28576 = ~n17075 & n28575 ;
  assign n28577 = n6122 | n28576 ;
  assign n28578 = n28577 ^ n27426 ^ 1'b0 ;
  assign n28579 = n25646 ^ n7272 ^ 1'b0 ;
  assign n28580 = n8672 | n28579 ;
  assign n28581 = ~n2231 & n12247 ;
  assign n28582 = ~n12156 & n28581 ;
  assign n28583 = n19081 | n28582 ;
  assign n28584 = n25698 ^ n15197 ^ 1'b0 ;
  assign n28585 = n8967 ^ n2977 ^ 1'b0 ;
  assign n28586 = n28584 & ~n28585 ;
  assign n28588 = n2885 & ~n22736 ;
  assign n28589 = n28588 ^ n19234 ^ 1'b0 ;
  assign n28587 = n11782 | n16746 ;
  assign n28590 = n28589 ^ n28587 ^ 1'b0 ;
  assign n28591 = n7644 ^ n1805 ^ 1'b0 ;
  assign n28592 = n4053 & ~n28591 ;
  assign n28593 = n4817 & n28592 ;
  assign n28594 = n113 & ~n16684 ;
  assign n28595 = n18162 | n19718 ;
  assign n28596 = n28595 ^ n10985 ^ 1'b0 ;
  assign n28597 = n28596 ^ n23242 ^ 1'b0 ;
  assign n28598 = n24013 & n28597 ;
  assign n28600 = n2899 & n17153 ;
  assign n28599 = n13960 | n14297 ;
  assign n28601 = n28600 ^ n28599 ^ 1'b0 ;
  assign n28602 = n12894 ^ n8262 ^ 1'b0 ;
  assign n28607 = n3851 ^ n2876 ^ 1'b0 ;
  assign n28603 = n4228 ^ n176 ^ 1'b0 ;
  assign n28604 = n12604 & ~n28603 ;
  assign n28605 = ~n5725 & n7540 ;
  assign n28606 = ~n28604 & n28605 ;
  assign n28608 = n28607 ^ n28606 ^ 1'b0 ;
  assign n28609 = ~n24268 & n28608 ;
  assign n28610 = n7886 & ~n15662 ;
  assign n28611 = n944 & ~n15775 ;
  assign n28612 = n6684 & n28611 ;
  assign n28613 = ~n15973 & n23765 ;
  assign n28614 = n10448 | n28613 ;
  assign n28615 = n287 & ~n28614 ;
  assign n28616 = n4864 & n7144 ;
  assign n28617 = ( n117 & ~n17964 ) | ( n117 & n21110 ) | ( ~n17964 & n21110 ) ;
  assign n28620 = n1256 & n6914 ;
  assign n28621 = n17885 ^ n9673 ^ 1'b0 ;
  assign n28622 = ~n28620 & n28621 ;
  assign n28618 = n13895 | n16236 ;
  assign n28619 = n28618 ^ n22891 ^ 1'b0 ;
  assign n28623 = n28622 ^ n28619 ^ n2020 ;
  assign n28624 = n24252 | n27941 ;
  assign n28625 = n4411 | n5175 ;
  assign n28626 = ~n251 & n697 ;
  assign n28627 = n2346 & n28626 ;
  assign n28628 = n10263 & ~n28627 ;
  assign n28629 = n15424 & n28628 ;
  assign n28630 = n3450 ^ n59 ^ 1'b0 ;
  assign n28631 = n5570 & n28630 ;
  assign n28632 = n28631 ^ n8639 ^ 1'b0 ;
  assign n28633 = n27055 | n28632 ;
  assign n28634 = n22441 ^ n4112 ^ 1'b0 ;
  assign n28635 = n4364 & ~n15118 ;
  assign n28636 = ( n12088 & ~n12185 ) | ( n12088 & n28635 ) | ( ~n12185 & n28635 ) ;
  assign n28637 = n28636 ^ n20856 ^ 1'b0 ;
  assign n28638 = ( n8962 & ~n28634 ) | ( n8962 & n28637 ) | ( ~n28634 & n28637 ) ;
  assign n28641 = ~n9066 & n12497 ;
  assign n28639 = n3870 & n4784 ;
  assign n28640 = n28639 ^ n24579 ^ n5803 ;
  assign n28642 = n28641 ^ n28640 ^ n19032 ;
  assign n28643 = n7255 | n9281 ;
  assign n28644 = n28643 ^ n23344 ^ 1'b0 ;
  assign n28645 = n11344 ^ n2169 ^ 1'b0 ;
  assign n28646 = n809 | n8543 ;
  assign n28647 = n28646 ^ n23833 ^ 1'b0 ;
  assign n28648 = n28645 | n28647 ;
  assign n28649 = ~n9643 & n10357 ;
  assign n28650 = ( n3973 & ~n4090 ) | ( n3973 & n28649 ) | ( ~n4090 & n28649 ) ;
  assign n28652 = ~n14936 & n20108 ;
  assign n28651 = n8190 & n22115 ;
  assign n28653 = n28652 ^ n28651 ^ 1'b0 ;
  assign n28654 = n1036 & ~n1720 ;
  assign n28655 = ~n20793 & n28654 ;
  assign n28656 = n21565 ^ n3212 ^ 1'b0 ;
  assign n28657 = n28655 | n28656 ;
  assign n28658 = n3825 & ~n26860 ;
  assign n28659 = n3512 | n16973 ;
  assign n28660 = n28659 ^ n11668 ^ 1'b0 ;
  assign n28661 = n9450 | n12288 ;
  assign n28662 = n28661 ^ n19710 ^ 1'b0 ;
  assign n28663 = n2759 | n3461 ;
  assign n28664 = n28663 ^ n5601 ^ 1'b0 ;
  assign n28665 = n20118 | n28664 ;
  assign n28666 = n18611 & ~n28665 ;
  assign n28667 = n837 | n24748 ;
  assign n28668 = ~n20645 & n28667 ;
  assign n28669 = n28668 ^ n28203 ^ 1'b0 ;
  assign n28670 = ( n874 & n11480 ) | ( n874 & n15550 ) | ( n11480 & n15550 ) ;
  assign n28671 = n1341 & ~n28670 ;
  assign n28672 = n28669 & n28671 ;
  assign n28677 = ~n9745 & n15347 ;
  assign n28678 = ~n5388 & n28677 ;
  assign n28679 = n398 | n28678 ;
  assign n28680 = n3060 | n28679 ;
  assign n28681 = ( n4847 & n6402 ) | ( n4847 & n28680 ) | ( n6402 & n28680 ) ;
  assign n28673 = ~n5781 & n24714 ;
  assign n28674 = n3867 & n28673 ;
  assign n28675 = ( n3855 & n13899 ) | ( n3855 & ~n28674 ) | ( n13899 & ~n28674 ) ;
  assign n28676 = n25718 & ~n28675 ;
  assign n28682 = n28681 ^ n28676 ^ 1'b0 ;
  assign n28683 = ( n2857 & ~n7244 ) | ( n2857 & n11147 ) | ( ~n7244 & n11147 ) ;
  assign n28684 = n8728 & ~n28683 ;
  assign n28685 = n5559 ^ n1475 ^ 1'b0 ;
  assign n28686 = n7567 | n10546 ;
  assign n28687 = n28686 ^ n4752 ^ 1'b0 ;
  assign n28688 = n14821 & ~n28687 ;
  assign n28689 = ~n12330 & n28688 ;
  assign n28690 = n14292 ^ n8209 ^ 1'b0 ;
  assign n28691 = ~n20068 & n28690 ;
  assign n28692 = ~n13561 & n28691 ;
  assign n28693 = n6208 & n12123 ;
  assign n28694 = n11379 & ~n27142 ;
  assign n28695 = ~n28693 & n28694 ;
  assign n28696 = n3894 | n26109 ;
  assign n28697 = n4590 | n8479 ;
  assign n28698 = ( n3456 & n5688 ) | ( n3456 & ~n28697 ) | ( n5688 & ~n28697 ) ;
  assign n28699 = n5651 & ~n10200 ;
  assign n28700 = ~n22628 & n28699 ;
  assign n28701 = n28700 ^ n7008 ^ 1'b0 ;
  assign n28702 = n24485 | n27097 ;
  assign n28703 = n16419 ^ n1085 ^ 1'b0 ;
  assign n28704 = n1134 & ~n28703 ;
  assign n28705 = ~n2997 & n11507 ;
  assign n28706 = n20614 ^ n2603 ^ 1'b0 ;
  assign n28707 = n4204 | n5290 ;
  assign n28708 = n20193 ^ n6725 ^ 1'b0 ;
  assign n28709 = n22483 ^ n6546 ^ 1'b0 ;
  assign n28710 = n10111 | n28709 ;
  assign n28711 = n22937 | n28710 ;
  assign n28712 = n24881 ^ n7233 ^ 1'b0 ;
  assign n28713 = n6445 | n27521 ;
  assign n28714 = n9851 ^ n6181 ^ 1'b0 ;
  assign n28715 = n28714 ^ n19443 ^ n3460 ;
  assign n28716 = ( n13023 & n17301 ) | ( n13023 & n22078 ) | ( n17301 & n22078 ) ;
  assign n28717 = ~n23346 & n28716 ;
  assign n28718 = n28717 ^ n14719 ^ 1'b0 ;
  assign n28719 = n28718 ^ n2588 ^ 1'b0 ;
  assign n28720 = n1188 & ~n2621 ;
  assign n28721 = ~n962 & n28720 ;
  assign n28722 = n960 | n28721 ;
  assign n28723 = n371 & ~n17024 ;
  assign n28724 = ~n17031 & n24013 ;
  assign n28725 = ~n1512 & n11959 ;
  assign n28726 = n28725 ^ n5352 ^ 1'b0 ;
  assign n28727 = ( ~n70 & n3322 ) | ( ~n70 & n28726 ) | ( n3322 & n28726 ) ;
  assign n28728 = n373 & ~n28727 ;
  assign n28729 = n28728 ^ n11485 ^ 1'b0 ;
  assign n28730 = n6851 & n28729 ;
  assign n28731 = ~n15308 & n28730 ;
  assign n28732 = n27069 ^ n9930 ^ 1'b0 ;
  assign n28733 = n22202 & ~n28732 ;
  assign n28734 = n390 | n5790 ;
  assign n28735 = n14077 | n28734 ;
  assign n28736 = n28735 ^ n5837 ^ 1'b0 ;
  assign n28737 = ~n4894 & n9218 ;
  assign n28738 = n115 | n4177 ;
  assign n28739 = n17676 ^ n14913 ^ n13425 ;
  assign n28740 = ~n14553 & n28739 ;
  assign n28741 = n19727 ^ n3469 ^ 1'b0 ;
  assign n28742 = n4483 | n28741 ;
  assign n28743 = n28742 ^ n12687 ^ 1'b0 ;
  assign n28744 = ~n9131 & n28743 ;
  assign n28745 = n20705 ^ n10516 ^ 1'b0 ;
  assign n28747 = n14308 ^ n6703 ^ n6157 ;
  assign n28746 = n27147 ^ n14849 ^ 1'b0 ;
  assign n28748 = n28747 ^ n28746 ^ 1'b0 ;
  assign n28749 = n24165 ^ n16861 ^ 1'b0 ;
  assign n28750 = n20736 & n24865 ;
  assign n28751 = ~n28749 & n28750 ;
  assign n28752 = ~n8269 & n24283 ;
  assign n28753 = ~n2989 & n4212 ;
  assign n28754 = n22160 ^ n1929 ^ 1'b0 ;
  assign n28755 = n19729 | n28754 ;
  assign n28756 = n14649 ^ n6541 ^ 1'b0 ;
  assign n28757 = ~n5554 & n28756 ;
  assign n28758 = ~n27684 & n28757 ;
  assign n28759 = n11258 & ~n11961 ;
  assign n28760 = n19672 & n28759 ;
  assign n28761 = n28760 ^ n9152 ^ 1'b0 ;
  assign n28762 = ~n23928 & n28761 ;
  assign n28763 = n16349 & n28762 ;
  assign n28764 = ( n6845 & n14895 ) | ( n6845 & n28763 ) | ( n14895 & n28763 ) ;
  assign n28765 = n12188 & n15063 ;
  assign n28767 = ~n6700 & n11123 ;
  assign n28766 = n10385 & n17744 ;
  assign n28768 = n28767 ^ n28766 ^ 1'b0 ;
  assign n28769 = n15900 ^ n13041 ^ 1'b0 ;
  assign n28770 = n28769 ^ n8763 ^ 1'b0 ;
  assign n28771 = n694 | n28770 ;
  assign n28772 = n2281 & ~n25680 ;
  assign n28773 = n354 & n28772 ;
  assign n28774 = n28773 ^ n12990 ^ 1'b0 ;
  assign n28775 = n14526 ^ n2650 ^ 1'b0 ;
  assign n28776 = ~n10677 & n17900 ;
  assign n28777 = n28776 ^ n411 ^ 1'b0 ;
  assign n28778 = n17650 ^ n6879 ^ 1'b0 ;
  assign n28779 = n3987 & n28778 ;
  assign n28780 = n6753 & ~n12335 ;
  assign n28781 = n1505 | n8563 ;
  assign n28782 = n441 | n28781 ;
  assign n28783 = n28782 ^ n14559 ^ 1'b0 ;
  assign n28784 = n2344 & n28783 ;
  assign n28785 = n2741 & n24714 ;
  assign n28786 = ~n18912 & n28785 ;
  assign n28787 = ( n28780 & n28784 ) | ( n28780 & n28786 ) | ( n28784 & n28786 ) ;
  assign n28788 = n19052 ^ n11535 ^ 1'b0 ;
  assign n28789 = ~n7268 & n8382 ;
  assign n28790 = n17210 & n27607 ;
  assign n28791 = n1959 & n28790 ;
  assign n28792 = n28791 ^ n11511 ^ 1'b0 ;
  assign n28794 = n5135 ^ n1856 ^ 1'b0 ;
  assign n28795 = n9109 & ~n28794 ;
  assign n28793 = n959 & ~n9073 ;
  assign n28796 = n28795 ^ n28793 ^ 1'b0 ;
  assign n28797 = ~n1426 & n16262 ;
  assign n28798 = n7916 & n28797 ;
  assign n28799 = n28798 ^ n10723 ^ 1'b0 ;
  assign n28800 = n10279 & ~n13693 ;
  assign n28801 = n26929 ^ n10073 ^ n1825 ;
  assign n28802 = n16794 & n28801 ;
  assign n28803 = n28802 ^ n27579 ^ 1'b0 ;
  assign n28804 = n1984 ^ n1296 ^ 1'b0 ;
  assign n28805 = n17878 & ~n28804 ;
  assign n28806 = n28805 ^ n6030 ^ n5149 ;
  assign n28807 = n439 | n13700 ;
  assign n28808 = n28807 ^ n2553 ^ 1'b0 ;
  assign n28809 = n7253 | n9192 ;
  assign n28810 = n6608 & ~n28809 ;
  assign n28811 = n28810 ^ n28360 ^ 1'b0 ;
  assign n28812 = n1317 | n28811 ;
  assign n28813 = n28808 & ~n28812 ;
  assign n28814 = n28813 ^ n12146 ^ n3038 ;
  assign n28815 = n19198 & n20991 ;
  assign n28816 = n4471 & n28815 ;
  assign n28817 = ~n2597 & n6537 ;
  assign n28818 = n11736 ^ n9601 ^ 1'b0 ;
  assign n28819 = n6443 & ~n10209 ;
  assign n28820 = n2889 | n28819 ;
  assign n28821 = n28820 ^ n181 ^ 1'b0 ;
  assign n28828 = n19925 ^ n9564 ^ 1'b0 ;
  assign n28827 = n10897 ^ n9939 ^ 1'b0 ;
  assign n28822 = n5896 & n9439 ;
  assign n28823 = n28822 ^ n27521 ^ 1'b0 ;
  assign n28824 = n4572 & ~n10512 ;
  assign n28825 = ~n13631 & n28824 ;
  assign n28826 = n28823 & ~n28825 ;
  assign n28829 = n28828 ^ n28827 ^ n28826 ;
  assign n28830 = n1704 & n4330 ;
  assign n28831 = n3541 & ~n6498 ;
  assign n28832 = n3385 & ~n3489 ;
  assign n28833 = ~n2999 & n28832 ;
  assign n28834 = n9600 & ~n10494 ;
  assign n28835 = ~n15514 & n28834 ;
  assign n28836 = n28835 ^ n18022 ^ 1'b0 ;
  assign n28837 = ~n28833 & n28836 ;
  assign n28838 = n28837 ^ n26462 ^ n2934 ;
  assign n28839 = n10448 | n15464 ;
  assign n28840 = ~n22674 & n25609 ;
  assign n28841 = n2729 & ~n6583 ;
  assign n28842 = n2509 & n28841 ;
  assign n28843 = ~n10905 & n28842 ;
  assign n28844 = n4239 | n5502 ;
  assign n28845 = n2899 | n28844 ;
  assign n28846 = n28845 ^ n12127 ^ 1'b0 ;
  assign n28847 = n19691 & ~n28846 ;
  assign n28848 = ( n3446 & n28843 ) | ( n3446 & n28847 ) | ( n28843 & n28847 ) ;
  assign n28849 = n16876 ^ n15217 ^ 1'b0 ;
  assign n28850 = n10305 ^ n7718 ^ 1'b0 ;
  assign n28851 = ~n3059 & n28850 ;
  assign n28852 = n11411 & n28851 ;
  assign n28853 = n28852 ^ n16966 ^ 1'b0 ;
  assign n28854 = n27171 ^ n15569 ^ 1'b0 ;
  assign n28855 = n293 | n28854 ;
  assign n28856 = n6144 | n28855 ;
  assign n28857 = n28856 ^ n15910 ^ 1'b0 ;
  assign n28858 = n12165 & ~n28857 ;
  assign n28859 = ~n8931 & n15056 ;
  assign n28860 = n28859 ^ n19743 ^ 1'b0 ;
  assign n28863 = n4490 & n15682 ;
  assign n28861 = n598 & n14164 ;
  assign n28862 = ~n14370 & n28861 ;
  assign n28864 = n28863 ^ n28862 ^ 1'b0 ;
  assign n28868 = n4048 ^ n1400 ^ 1'b0 ;
  assign n28865 = n18909 ^ n13359 ^ 1'b0 ;
  assign n28866 = n4330 & n28865 ;
  assign n28867 = n16578 | n28866 ;
  assign n28869 = n28868 ^ n28867 ^ n19635 ;
  assign n28870 = n28869 ^ n26308 ^ n2523 ;
  assign n28873 = ~n2485 & n5806 ;
  assign n28871 = n27875 ^ n12071 ^ 1'b0 ;
  assign n28872 = n4750 | n28871 ;
  assign n28874 = n28873 ^ n28872 ^ 1'b0 ;
  assign n28875 = n3591 | n19236 ;
  assign n28876 = n28875 ^ n4859 ^ 1'b0 ;
  assign n28877 = ~n12548 & n16118 ;
  assign n28878 = ~n28876 & n28877 ;
  assign n28879 = n28878 ^ n15150 ^ 1'b0 ;
  assign n28880 = n28301 ^ n12629 ^ 1'b0 ;
  assign n28883 = ( n1995 & n4121 ) | ( n1995 & ~n4869 ) | ( n4121 & ~n4869 ) ;
  assign n28884 = n28883 ^ n9955 ^ 1'b0 ;
  assign n28885 = n5197 | n28884 ;
  assign n28881 = n22290 ^ n7772 ^ 1'b0 ;
  assign n28882 = n14252 | n28881 ;
  assign n28886 = n28885 ^ n28882 ^ n17667 ;
  assign n28887 = n10646 & ~n28886 ;
  assign n28888 = n11078 & ~n23861 ;
  assign n28889 = n2928 & n28888 ;
  assign n28890 = n1118 & n28368 ;
  assign n28894 = n4743 & n13717 ;
  assign n28895 = n28894 ^ n2884 ^ 1'b0 ;
  assign n28891 = ~n13585 & n18455 ;
  assign n28892 = ( ~n11544 & n19869 ) | ( ~n11544 & n28891 ) | ( n19869 & n28891 ) ;
  assign n28893 = n283 & n28892 ;
  assign n28896 = n28895 ^ n28893 ^ 1'b0 ;
  assign n28897 = n28153 & n28896 ;
  assign n28898 = n7554 ^ n5501 ^ 1'b0 ;
  assign n28899 = n28898 ^ n3584 ^ 1'b0 ;
  assign n28900 = n8421 | n9314 ;
  assign n28901 = n10647 | n28900 ;
  assign n28902 = n28901 ^ n17824 ^ 1'b0 ;
  assign n28903 = ~n14738 & n27068 ;
  assign n28904 = n25885 ^ n2563 ^ 1'b0 ;
  assign n28905 = n28903 | n28904 ;
  assign n28906 = n17226 & ~n28905 ;
  assign n28907 = n21649 ^ n5589 ^ 1'b0 ;
  assign n28908 = ~n25437 & n28907 ;
  assign n28909 = n21562 ^ n5796 ^ 1'b0 ;
  assign n28910 = n24028 & ~n28909 ;
  assign n28911 = n28910 ^ n26188 ^ 1'b0 ;
  assign n28912 = n16570 & ~n28146 ;
  assign n28913 = ~n28911 & n28912 ;
  assign n28914 = n17175 & n18907 ;
  assign n28915 = n28914 ^ n1636 ^ 1'b0 ;
  assign n28916 = n6457 ^ n2556 ^ 1'b0 ;
  assign n28917 = n11611 | n28916 ;
  assign n28918 = ~n5399 & n22120 ;
  assign n28919 = n28918 ^ n5175 ^ 1'b0 ;
  assign n28920 = n17232 ^ n636 ^ 1'b0 ;
  assign n28921 = n20514 | n28618 ;
  assign n28922 = n8516 | n28921 ;
  assign n28923 = n12119 & n28922 ;
  assign n28929 = ( ~n230 & n4859 ) | ( ~n230 & n14617 ) | ( n4859 & n14617 ) ;
  assign n28924 = ~n5581 & n22712 ;
  assign n28925 = n5957 & ~n17243 ;
  assign n28926 = n28925 ^ n1535 ^ 1'b0 ;
  assign n28927 = ~n28924 & n28926 ;
  assign n28928 = ~n18741 & n28927 ;
  assign n28930 = n28929 ^ n28928 ^ n249 ;
  assign n28931 = n19497 ^ n13572 ^ 1'b0 ;
  assign n28932 = ~n28930 & n28931 ;
  assign n28933 = n1803 ^ n813 ^ n26 ;
  assign n28934 = n28933 ^ n3245 ^ n1563 ;
  assign n28935 = n10348 & ~n11876 ;
  assign n28936 = ~n7208 & n28935 ;
  assign n28937 = n12747 ^ n6511 ^ 1'b0 ;
  assign n28938 = n22844 ^ n16010 ^ 1'b0 ;
  assign n28939 = n2131 | n10376 ;
  assign n28940 = n28939 ^ n8660 ^ 1'b0 ;
  assign n28941 = n28688 | n28940 ;
  assign n28942 = n1647 & ~n8117 ;
  assign n28943 = n12758 & n28942 ;
  assign n28944 = n13772 ^ n9118 ^ n7196 ;
  assign n28945 = ( n14299 & ~n15725 ) | ( n14299 & n28944 ) | ( ~n15725 & n28944 ) ;
  assign n28946 = n27385 ^ n835 ^ 1'b0 ;
  assign n28947 = n7778 & ~n28946 ;
  assign n28948 = n16567 & ~n22407 ;
  assign n28949 = ~n28947 & n28948 ;
  assign n28951 = ~n4230 & n13258 ;
  assign n28950 = n2124 & n6305 ;
  assign n28952 = n28951 ^ n28950 ^ 1'b0 ;
  assign n28953 = ~n8397 & n28952 ;
  assign n28954 = ~n3608 & n26130 ;
  assign n28955 = n8552 ^ n2525 ^ n1185 ;
  assign n28956 = n17445 & ~n28955 ;
  assign n28957 = ~n24266 & n28956 ;
  assign n28958 = n28957 ^ n3805 ^ 1'b0 ;
  assign n28959 = ~n13815 & n16060 ;
  assign n28960 = n28959 ^ n1932 ^ 1'b0 ;
  assign n28961 = ~n2232 & n9815 ;
  assign n28962 = n28961 ^ n25792 ^ n22688 ;
  assign n28963 = n5169 | n7588 ;
  assign n28964 = n28963 ^ n4827 ^ 1'b0 ;
  assign n28965 = n10983 | n28964 ;
  assign n28966 = n28965 ^ n11029 ^ 1'b0 ;
  assign n28967 = n6053 & ~n8008 ;
  assign n28968 = n8450 & n28967 ;
  assign n28969 = n4732 & ~n7014 ;
  assign n28970 = n19304 ^ n1164 ^ 1'b0 ;
  assign n28971 = ~n10080 & n28970 ;
  assign n28972 = n28971 ^ n12869 ^ 1'b0 ;
  assign n28973 = n6521 & n28972 ;
  assign n28974 = n6097 & ~n17207 ;
  assign n28975 = n3153 & ~n28974 ;
  assign n28976 = n23446 ^ n3395 ^ 1'b0 ;
  assign n28978 = n21409 ^ n15618 ^ 1'b0 ;
  assign n28979 = n28978 ^ n14287 ^ 1'b0 ;
  assign n28977 = ~n25184 & n28545 ;
  assign n28980 = n28979 ^ n28977 ^ 1'b0 ;
  assign n28981 = n15573 ^ n1940 ^ 1'b0 ;
  assign n28982 = n13726 ^ n6302 ^ 1'b0 ;
  assign n28983 = n1307 & n7864 ;
  assign n28984 = ( n1851 & n3971 ) | ( n1851 & n5066 ) | ( n3971 & n5066 ) ;
  assign n28985 = ~n115 & n6101 ;
  assign n28986 = n28984 & n28985 ;
  assign n28987 = n4195 & ~n28986 ;
  assign n28988 = n28983 & n28987 ;
  assign n28989 = n2758 | n28988 ;
  assign n28990 = ( n4004 & n7768 ) | ( n4004 & ~n11777 ) | ( n7768 & ~n11777 ) ;
  assign n28991 = n25688 ^ n11161 ^ 1'b0 ;
  assign n28992 = n28991 ^ n5941 ^ 1'b0 ;
  assign n28993 = n7129 ^ n342 ^ 1'b0 ;
  assign n28994 = n676 | n12866 ;
  assign n28995 = n28993 | n28994 ;
  assign n28996 = n21849 ^ n3035 ^ 1'b0 ;
  assign n28997 = ~n21868 & n22081 ;
  assign n28998 = n2451 | n12898 ;
  assign n28999 = n1537 & ~n28998 ;
  assign n29000 = ~n3803 & n16755 ;
  assign n29001 = ~n13565 & n29000 ;
  assign n29002 = n29001 ^ n2584 ^ 1'b0 ;
  assign n29003 = n2587 & n24655 ;
  assign n29004 = ~n20951 & n29003 ;
  assign n29005 = n29004 ^ n2011 ^ 1'b0 ;
  assign n29006 = ~n1720 & n12441 ;
  assign n29007 = n29006 ^ n8728 ^ 1'b0 ;
  assign n29008 = n8833 & ~n29007 ;
  assign n29009 = n5051 & ~n5630 ;
  assign n29010 = n29009 ^ n14765 ^ 1'b0 ;
  assign n29011 = n29010 ^ n4536 ^ 1'b0 ;
  assign n29012 = n20685 | n29011 ;
  assign n29013 = n7530 ^ n2928 ^ 1'b0 ;
  assign n29014 = n28960 | n29013 ;
  assign n29015 = n23718 & ~n29014 ;
  assign n29016 = ~n1018 & n3625 ;
  assign n29017 = n13021 ^ n10157 ^ 1'b0 ;
  assign n29018 = n14447 | n29017 ;
  assign n29019 = n29016 | n29018 ;
  assign n29020 = n14418 | n21643 ;
  assign n29021 = n4275 & n24173 ;
  assign n29022 = n6000 & n6925 ;
  assign n29023 = ~n15662 & n29022 ;
  assign n29024 = ~n1812 & n29023 ;
  assign n29025 = n4582 & ~n29024 ;
  assign n29026 = n26948 & n29025 ;
  assign n29027 = ~n6188 & n14258 ;
  assign n29028 = n10400 & n29027 ;
  assign n29029 = n8937 & n29028 ;
  assign n29030 = n29029 ^ n20718 ^ n11751 ;
  assign n29031 = n23247 ^ n19097 ^ n8278 ;
  assign n29032 = n13677 ^ n7115 ^ 1'b0 ;
  assign n29033 = n1611 & n13936 ;
  assign n29034 = n9698 ^ n9276 ^ 1'b0 ;
  assign n29035 = n8262 | n29034 ;
  assign n29036 = n9934 ^ n2765 ^ 1'b0 ;
  assign n29037 = n27880 & ~n29036 ;
  assign n29040 = n8231 ^ n5118 ^ 1'b0 ;
  assign n29041 = ~n4002 & n29040 ;
  assign n29038 = n12737 ^ n11462 ^ n6412 ;
  assign n29039 = ( n46 & n1995 ) | ( n46 & ~n29038 ) | ( n1995 & ~n29038 ) ;
  assign n29042 = n29041 ^ n29039 ^ n26162 ;
  assign n29043 = n6493 ^ n3446 ^ 1'b0 ;
  assign n29044 = ~n25601 & n29043 ;
  assign n29045 = n29044 ^ n15190 ^ 1'b0 ;
  assign n29046 = n14082 & ~n14224 ;
  assign n29047 = n10356 ^ n2678 ^ 1'b0 ;
  assign n29048 = ( n492 & n8310 ) | ( n492 & ~n29047 ) | ( n8310 & ~n29047 ) ;
  assign n29049 = n29048 ^ n16160 ^ n4862 ;
  assign n29050 = n28044 ^ n11036 ^ 1'b0 ;
  assign n29051 = n20781 ^ n7223 ^ 1'b0 ;
  assign n29052 = n340 & ~n29051 ;
  assign n29053 = n3967 & n4869 ;
  assign n29054 = n29053 ^ n1188 ^ 1'b0 ;
  assign n29055 = n2190 & ~n9137 ;
  assign n29056 = n29054 & n29055 ;
  assign n29057 = n1645 & ~n29056 ;
  assign n29058 = n29057 ^ n14095 ^ 1'b0 ;
  assign n29059 = n20217 & ~n23333 ;
  assign n29060 = n29059 ^ n22812 ^ 1'b0 ;
  assign n29061 = n29060 ^ n12494 ^ 1'b0 ;
  assign n29062 = n21312 & n29061 ;
  assign n29063 = n28384 ^ n11130 ^ 1'b0 ;
  assign n29064 = n19065 & n29063 ;
  assign n29065 = ( n1389 & n14246 ) | ( n1389 & n29064 ) | ( n14246 & n29064 ) ;
  assign n29066 = n13439 ^ n4607 ^ 1'b0 ;
  assign n29067 = n22804 | n29066 ;
  assign n29068 = n1263 & n29067 ;
  assign n29069 = ~n5377 & n29068 ;
  assign n29070 = n19646 & ~n29069 ;
  assign n29071 = ~n2995 & n6134 ;
  assign n29072 = ( n6493 & n8349 ) | ( n6493 & ~n19255 ) | ( n8349 & ~n19255 ) ;
  assign n29073 = n29072 ^ n14344 ^ 1'b0 ;
  assign n29074 = n29073 ^ n11962 ^ n1604 ;
  assign n29075 = n2526 | n17661 ;
  assign n29076 = n29074 | n29075 ;
  assign n29079 = n8387 & n24872 ;
  assign n29080 = n29079 ^ n13658 ^ 1'b0 ;
  assign n29077 = n2286 | n11700 ;
  assign n29078 = ( n9958 & n16050 ) | ( n9958 & n29077 ) | ( n16050 & n29077 ) ;
  assign n29081 = n29080 ^ n29078 ^ 1'b0 ;
  assign n29082 = n17963 & ~n28199 ;
  assign n29083 = ~n1875 & n6578 ;
  assign n29084 = n29083 ^ n15692 ^ 1'b0 ;
  assign n29085 = n9479 | n29084 ;
  assign n29086 = ~n8207 & n17578 ;
  assign n29087 = n8207 & n29086 ;
  assign n29088 = n5806 ^ n1727 ^ 1'b0 ;
  assign n29089 = n6962 & n29088 ;
  assign n29090 = n7558 ^ n4688 ^ 1'b0 ;
  assign n29091 = n25910 & ~n29090 ;
  assign n29092 = n29089 & n29091 ;
  assign n29093 = n9211 & n29092 ;
  assign n29094 = n12765 & n14605 ;
  assign n29095 = n29094 ^ n3677 ^ 1'b0 ;
  assign n29096 = n7472 & ~n18954 ;
  assign n29097 = n29096 ^ n8436 ^ 1'b0 ;
  assign n29098 = n15979 & ~n29097 ;
  assign n29099 = n4427 & n29098 ;
  assign n29100 = n15593 ^ n11383 ^ n7626 ;
  assign n29101 = n6547 ^ n1944 ^ 1'b0 ;
  assign n29102 = n352 & ~n29101 ;
  assign n29103 = n4806 & n27997 ;
  assign n29104 = n29103 ^ n16090 ^ 1'b0 ;
  assign n29105 = n1581 & ~n3800 ;
  assign n29106 = ~n12347 & n13117 ;
  assign n29107 = n29106 ^ n23856 ^ 1'b0 ;
  assign n29108 = ~n29105 & n29107 ;
  assign n29109 = n29108 ^ n816 ^ 1'b0 ;
  assign n29110 = n29109 ^ n22161 ^ 1'b0 ;
  assign n29111 = n9003 ^ n4536 ^ 1'b0 ;
  assign n29112 = n16545 | n29111 ;
  assign n29113 = n29112 ^ n14835 ^ 1'b0 ;
  assign n29116 = n2961 ^ n561 ^ 1'b0 ;
  assign n29117 = n6985 | n29116 ;
  assign n29114 = n14144 ^ n1746 ^ 1'b0 ;
  assign n29115 = n12143 & ~n29114 ;
  assign n29118 = n29117 ^ n29115 ^ 1'b0 ;
  assign n29119 = n5033 & ~n11032 ;
  assign n29120 = n3025 & n10747 ;
  assign n29121 = n29120 ^ n16857 ^ 1'b0 ;
  assign n29122 = n29121 ^ n1549 ^ 1'b0 ;
  assign n29123 = n27456 & n29122 ;
  assign n29124 = n2157 | n21315 ;
  assign n29125 = n29124 ^ n21868 ^ 1'b0 ;
  assign n29126 = n19555 ^ n13256 ^ 1'b0 ;
  assign n29127 = n28215 ^ n4123 ^ 1'b0 ;
  assign n29128 = ( n13142 & n16197 ) | ( n13142 & ~n29127 ) | ( n16197 & ~n29127 ) ;
  assign n29129 = n29128 ^ n10681 ^ 1'b0 ;
  assign n29130 = n29126 & ~n29129 ;
  assign n29131 = n17689 ^ n16127 ^ 1'b0 ;
  assign n29132 = ( n313 & n2813 ) | ( n313 & ~n29131 ) | ( n2813 & ~n29131 ) ;
  assign n29134 = ~n7325 & n21387 ;
  assign n29135 = ~n21387 & n29134 ;
  assign n29136 = n16996 & n29135 ;
  assign n29133 = ~n5264 & n20926 ;
  assign n29137 = n29136 ^ n29133 ^ n6412 ;
  assign n29138 = n197 | n5182 ;
  assign n29139 = n18186 | n19429 ;
  assign n29140 = n29139 ^ n7017 ^ 1'b0 ;
  assign n29141 = n7641 & n11180 ;
  assign n29142 = ~n17033 & n29141 ;
  assign n29143 = n12026 & ~n22450 ;
  assign n29144 = n29142 & n29143 ;
  assign n29145 = n12730 & n24743 ;
  assign n29146 = n29145 ^ n25681 ^ 1'b0 ;
  assign n29147 = n18522 & ~n29146 ;
  assign n29148 = ( ~n5702 & n20433 ) | ( ~n5702 & n29147 ) | ( n20433 & n29147 ) ;
  assign n29149 = n28861 ^ n14164 ^ 1'b0 ;
  assign n29150 = ~n16324 & n29149 ;
  assign n29151 = ~n1643 & n22365 ;
  assign n29156 = n23886 ^ n4627 ^ 1'b0 ;
  assign n29152 = n1329 & n17257 ;
  assign n29153 = ~n16080 & n29152 ;
  assign n29154 = n29153 ^ n16278 ^ n4298 ;
  assign n29155 = n3698 | n29154 ;
  assign n29157 = n29156 ^ n29155 ^ 1'b0 ;
  assign n29158 = n2397 & ~n22903 ;
  assign n29159 = n3754 & n4369 ;
  assign n29160 = n29159 ^ n1852 ^ 1'b0 ;
  assign n29161 = n29160 ^ n26451 ^ 1'b0 ;
  assign n29162 = n2463 & n29161 ;
  assign n29163 = n2114 | n15680 ;
  assign n29164 = n29163 ^ n15070 ^ n3985 ;
  assign n29165 = n29164 ^ n16804 ^ 1'b0 ;
  assign n29166 = n13795 & n28494 ;
  assign n29167 = n29166 ^ n14227 ^ 1'b0 ;
  assign n29168 = n1582 & n24406 ;
  assign n29169 = n1762 & ~n18171 ;
  assign n29170 = ~n27120 & n29169 ;
  assign n29171 = n14913 & n23628 ;
  assign n29172 = n29171 ^ n22940 ^ 1'b0 ;
  assign n29173 = n8337 & n12810 ;
  assign n29174 = n29173 ^ n3519 ^ 1'b0 ;
  assign n29175 = ~n3314 & n29174 ;
  assign n29176 = ~n6957 & n29175 ;
  assign n29177 = ~n14481 & n29176 ;
  assign n29178 = n17599 & n21828 ;
  assign n29179 = n29177 & n29178 ;
  assign n29180 = n18765 ^ n7749 ^ 1'b0 ;
  assign n29181 = n17468 & n29180 ;
  assign n29184 = n9293 & n10294 ;
  assign n29185 = n29184 ^ n15349 ^ 1'b0 ;
  assign n29182 = n11805 | n27159 ;
  assign n29183 = n28600 & ~n29182 ;
  assign n29186 = n29185 ^ n29183 ^ 1'b0 ;
  assign n29187 = n4319 ^ n1013 ^ 1'b0 ;
  assign n29188 = n8707 ^ n1456 ^ 1'b0 ;
  assign n29189 = n29187 & n29188 ;
  assign n29190 = ( n2341 & n12393 ) | ( n2341 & n29189 ) | ( n12393 & n29189 ) ;
  assign n29191 = n10527 ^ n2882 ^ 1'b0 ;
  assign n29192 = n24842 ^ n237 ^ 1'b0 ;
  assign n29193 = n29192 ^ n7860 ^ 1'b0 ;
  assign n29194 = n13916 & ~n29193 ;
  assign n29195 = n10915 | n29194 ;
  assign n29196 = ~n2928 & n4308 ;
  assign n29197 = n27429 ^ n4540 ^ 1'b0 ;
  assign n29198 = n176 | n7222 ;
  assign n29199 = n24456 & n29198 ;
  assign n29200 = n1525 & n10118 ;
  assign n29201 = ~n16005 & n29200 ;
  assign n29202 = n1001 & n29201 ;
  assign n29207 = n4260 & ~n15421 ;
  assign n29203 = n654 & ~n10667 ;
  assign n29204 = n29203 ^ n3000 ^ 1'b0 ;
  assign n29205 = n9496 & ~n29204 ;
  assign n29206 = n22127 & n29205 ;
  assign n29208 = n29207 ^ n29206 ^ 1'b0 ;
  assign n29209 = n29208 ^ n3142 ^ 1'b0 ;
  assign n29210 = n6789 ^ n3722 ^ 1'b0 ;
  assign n29211 = n23313 & n29210 ;
  assign n29212 = n9036 & ~n10339 ;
  assign n29213 = ~n4861 & n20871 ;
  assign n29214 = ~n29212 & n29213 ;
  assign n29215 = n29214 ^ n23393 ^ n7354 ;
  assign n29216 = n29215 ^ n19342 ^ n1589 ;
  assign n29217 = n12688 & ~n27295 ;
  assign n29218 = ~n7708 & n29217 ;
  assign n29219 = ~n51 & n29218 ;
  assign n29220 = n29216 | n29219 ;
  assign n29221 = n29220 ^ n9409 ^ 1'b0 ;
  assign n29222 = n26094 ^ n5446 ^ n3710 ;
  assign n29223 = ( n7892 & n20869 ) | ( n7892 & n29222 ) | ( n20869 & n29222 ) ;
  assign n29224 = n6700 ^ n4516 ^ 1'b0 ;
  assign n29225 = ~n24633 & n29224 ;
  assign n29226 = n5224 & n29225 ;
  assign n29227 = n29226 ^ n533 ^ 1'b0 ;
  assign n29228 = n29227 ^ n11867 ^ 1'b0 ;
  assign n29229 = n16124 & ~n29228 ;
  assign n29230 = n861 & ~n29229 ;
  assign n29231 = n29230 ^ n12626 ^ 1'b0 ;
  assign n29232 = n26298 ^ n3240 ^ 1'b0 ;
  assign n29233 = n7280 & ~n29232 ;
  assign n29234 = ( n3221 & n6618 ) | ( n3221 & n9024 ) | ( n6618 & n9024 ) ;
  assign n29235 = ~n7925 & n29234 ;
  assign n29236 = ( n25329 & n28414 ) | ( n25329 & n29235 ) | ( n28414 & n29235 ) ;
  assign n29237 = ~n11420 & n14968 ;
  assign n29238 = n29237 ^ n14587 ^ 1'b0 ;
  assign n29239 = ( n14121 & ~n15338 ) | ( n14121 & n29238 ) | ( ~n15338 & n29238 ) ;
  assign n29240 = n3191 & n12658 ;
  assign n29241 = ( n5694 & n9335 ) | ( n5694 & n15670 ) | ( n9335 & n15670 ) ;
  assign n29242 = ( ~n5054 & n29240 ) | ( ~n5054 & n29241 ) | ( n29240 & n29241 ) ;
  assign n29243 = n3923 & n15389 ;
  assign n29244 = n29243 ^ n2496 ^ 1'b0 ;
  assign n29245 = n29244 ^ n27919 ^ 1'b0 ;
  assign n29246 = n27922 | n28006 ;
  assign n29247 = n23492 | n29246 ;
  assign n29248 = n29247 ^ n18280 ^ 1'b0 ;
  assign n29249 = n21078 ^ n3429 ^ 1'b0 ;
  assign n29250 = n6317 & ~n8176 ;
  assign n29251 = n1745 ^ n1428 ^ 1'b0 ;
  assign n29252 = n1058 & ~n6152 ;
  assign n29253 = n6886 | n29252 ;
  assign n29254 = n29251 & ~n29253 ;
  assign n29255 = n1545 | n4123 ;
  assign n29256 = n1832 | n29255 ;
  assign n29257 = n2616 | n5654 ;
  assign n29258 = n29256 & ~n29257 ;
  assign n29259 = ( n8145 & n26651 ) | ( n8145 & ~n29258 ) | ( n26651 & ~n29258 ) ;
  assign n29260 = ~n7008 & n17455 ;
  assign n29261 = ~n3260 & n29260 ;
  assign n29262 = n29261 ^ n13378 ^ n12314 ;
  assign n29263 = n29262 ^ n23018 ^ 1'b0 ;
  assign n29264 = ( n738 & n12177 ) | ( n738 & ~n16187 ) | ( n12177 & ~n16187 ) ;
  assign n29265 = n2790 | n15299 ;
  assign n29266 = n8212 ^ n7580 ^ 1'b0 ;
  assign n29267 = n18847 & n29266 ;
  assign n29268 = ( ~n301 & n362 ) | ( ~n301 & n29267 ) | ( n362 & n29267 ) ;
  assign n29269 = n2094 & ~n29268 ;
  assign n29270 = ~n29265 & n29269 ;
  assign n29271 = n10987 ^ n9955 ^ 1'b0 ;
  assign n29272 = ~n2960 & n29271 ;
  assign n29273 = n22258 ^ n6242 ^ 1'b0 ;
  assign n29274 = n17576 | n23285 ;
  assign n29275 = n3773 | n29274 ;
  assign n29276 = ( n575 & n3983 ) | ( n575 & n23126 ) | ( n3983 & n23126 ) ;
  assign n29277 = n29276 ^ n14197 ^ 1'b0 ;
  assign n29278 = ~n19492 & n29277 ;
  assign n29279 = ~n3909 & n4629 ;
  assign n29280 = n24337 | n29279 ;
  assign n29281 = n29189 ^ n1064 ^ 1'b0 ;
  assign n29282 = ~n25159 & n29281 ;
  assign n29283 = n7219 & ~n11473 ;
  assign n29284 = ~n1010 & n6247 ;
  assign n29285 = n29284 ^ n9876 ^ 1'b0 ;
  assign n29286 = n29285 ^ n13603 ^ 1'b0 ;
  assign n29287 = n7357 | n15564 ;
  assign n29288 = n8157 ^ n7368 ^ 1'b0 ;
  assign n29289 = n29287 | n29288 ;
  assign n29290 = n21770 ^ n17742 ^ 1'b0 ;
  assign n29291 = ~n29289 & n29290 ;
  assign n29292 = n27469 ^ n2694 ^ n170 ;
  assign n29293 = n2831 & n3985 ;
  assign n29294 = ~n15708 & n29293 ;
  assign n29295 = n16714 & n25661 ;
  assign n29296 = n29294 & n29295 ;
  assign n29297 = ~n126 & n417 ;
  assign n29298 = n29297 ^ n11266 ^ 1'b0 ;
  assign n29299 = n5711 & ~n29298 ;
  assign n29300 = n29299 ^ n3140 ^ 1'b0 ;
  assign n29301 = n3420 ^ n3305 ^ n2883 ;
  assign n29302 = ( n9127 & n13863 ) | ( n9127 & n29301 ) | ( n13863 & n29301 ) ;
  assign n29303 = ( ~n3773 & n8665 ) | ( ~n3773 & n10007 ) | ( n8665 & n10007 ) ;
  assign n29304 = n29302 | n29303 ;
  assign n29305 = n12746 & n22678 ;
  assign n29306 = ~n26190 & n29305 ;
  assign n29307 = ( n4568 & n12425 ) | ( n4568 & ~n22846 ) | ( n12425 & ~n22846 ) ;
  assign n29308 = n29307 ^ n16768 ^ 1'b0 ;
  assign n29309 = n9912 | n22631 ;
  assign n29310 = n10265 & n16326 ;
  assign n29311 = ~n9380 & n29310 ;
  assign n29312 = ~n2333 & n29311 ;
  assign n29313 = n24187 ^ n18152 ^ 1'b0 ;
  assign n29314 = n6581 & n29313 ;
  assign n29315 = n29314 ^ n28070 ^ 1'b0 ;
  assign n29316 = n29312 | n29315 ;
  assign n29318 = n6541 & n20666 ;
  assign n29317 = n14170 ^ n2939 ^ 1'b0 ;
  assign n29319 = n29318 ^ n29317 ^ n7790 ;
  assign n29320 = n4775 ^ n3004 ^ 1'b0 ;
  assign n29321 = n29319 & ~n29320 ;
  assign n29322 = n12400 ^ n10178 ^ 1'b0 ;
  assign n29323 = n5100 & ~n11642 ;
  assign n29324 = n29323 ^ n9040 ^ 1'b0 ;
  assign n29325 = n20910 ^ n12304 ^ 1'b0 ;
  assign n29326 = n13941 ^ n8604 ^ 1'b0 ;
  assign n29328 = n40 & ~n7579 ;
  assign n29329 = n23563 & n29328 ;
  assign n29330 = n20518 & ~n29329 ;
  assign n29331 = n8450 & n29330 ;
  assign n29332 = n16051 & n29331 ;
  assign n29327 = ~n9962 & n13081 ;
  assign n29333 = n29332 ^ n29327 ^ 1'b0 ;
  assign n29334 = n10269 ^ n7872 ^ 1'b0 ;
  assign n29335 = ~n1081 & n11771 ;
  assign n29336 = n2294 ^ n63 ^ 1'b0 ;
  assign n29337 = n29335 & ~n29336 ;
  assign n29338 = ~n11514 & n29337 ;
  assign n29339 = n7925 & n29338 ;
  assign n29340 = n22573 ^ n9857 ^ 1'b0 ;
  assign n29341 = n5344 & ~n29340 ;
  assign n29342 = n12754 ^ n3190 ^ 1'b0 ;
  assign n29343 = n29342 ^ n7213 ^ 1'b0 ;
  assign n29344 = n29341 & n29343 ;
  assign n29345 = n2697 | n19865 ;
  assign n29346 = n29345 ^ n13722 ^ 1'b0 ;
  assign n29347 = ( ~n4699 & n25631 ) | ( ~n4699 & n27851 ) | ( n25631 & n27851 ) ;
  assign n29348 = n19940 & n28292 ;
  assign n29349 = n20748 | n24368 ;
  assign n29350 = n11300 & ~n18142 ;
  assign n29351 = n11131 & n29350 ;
  assign n29352 = n13660 ^ n4257 ^ n3950 ;
  assign n29353 = n17490 | n27044 ;
  assign n29354 = ( n2402 & n14595 ) | ( n2402 & n21571 ) | ( n14595 & n21571 ) ;
  assign n29355 = ~n9614 & n19041 ;
  assign n29356 = n5958 ^ n4127 ^ 1'b0 ;
  assign n29357 = ~n29355 & n29356 ;
  assign n29358 = ~n22829 & n22927 ;
  assign n29359 = n2288 | n29358 ;
  assign n29360 = n29359 ^ n13511 ^ 1'b0 ;
  assign n29361 = n230 & n891 ;
  assign n29362 = n2083 & n29361 ;
  assign n29363 = n9390 ^ n5353 ^ 1'b0 ;
  assign n29364 = n14813 ^ n12070 ^ n499 ;
  assign n29365 = n19348 | n27136 ;
  assign n29366 = n909 | n29365 ;
  assign n29367 = ~n2451 & n10147 ;
  assign n29368 = n29367 ^ n4228 ^ 1'b0 ;
  assign n29369 = n26126 & n29368 ;
  assign n29370 = n14498 & ~n16824 ;
  assign n29371 = ~n11950 & n29370 ;
  assign n29372 = n19270 ^ n1587 ^ 1'b0 ;
  assign n29373 = n14730 & ~n29372 ;
  assign n29374 = n17373 & n20458 ;
  assign n29375 = ~n29373 & n29374 ;
  assign n29376 = n12685 & ~n22508 ;
  assign n29377 = n29375 | n29376 ;
  assign n29378 = n29377 ^ n7808 ^ 1'b0 ;
  assign n29379 = n247 | n24670 ;
  assign n29380 = ( ~n13201 & n18951 ) | ( ~n13201 & n29379 ) | ( n18951 & n29379 ) ;
  assign n29381 = n13616 ^ n5164 ^ 1'b0 ;
  assign n29382 = n3738 & ~n13567 ;
  assign n29383 = n29382 ^ n3035 ^ 1'b0 ;
  assign n29384 = ( n2250 & n22776 ) | ( n2250 & ~n23731 ) | ( n22776 & ~n23731 ) ;
  assign n29385 = ~n647 & n8912 ;
  assign n29386 = ( ~n11875 & n29384 ) | ( ~n11875 & n29385 ) | ( n29384 & n29385 ) ;
  assign n29387 = n7090 ^ n7035 ^ n2209 ;
  assign n29388 = n29387 ^ n15977 ^ 1'b0 ;
  assign n29389 = ( n1311 & n2523 ) | ( n1311 & ~n24633 ) | ( n2523 & ~n24633 ) ;
  assign n29390 = ~n59 & n9337 ;
  assign n29391 = n18932 ^ n11227 ^ n2114 ;
  assign n29392 = n213 | n6183 ;
  assign n29393 = n29392 ^ n11138 ^ 1'b0 ;
  assign n29394 = n17278 | n29393 ;
  assign n29395 = n29394 ^ n20024 ^ n11030 ;
  assign n29396 = n29395 ^ n3229 ^ 1'b0 ;
  assign n29397 = n20946 ^ n3043 ^ 1'b0 ;
  assign n29398 = n15584 & n29397 ;
  assign n29399 = n17278 ^ n7017 ^ n2177 ;
  assign n29400 = n29399 ^ n16462 ^ n4511 ;
  assign n29401 = n21867 ^ n7278 ^ 1'b0 ;
  assign n29402 = ( n9753 & n15097 ) | ( n9753 & n29401 ) | ( n15097 & n29401 ) ;
  assign n29403 = ( n27118 & n28529 ) | ( n27118 & n29402 ) | ( n28529 & n29402 ) ;
  assign n29404 = ( ~n5465 & n13377 ) | ( ~n5465 & n29403 ) | ( n13377 & n29403 ) ;
  assign n29405 = n19410 ^ n6510 ^ 1'b0 ;
  assign n29406 = n9160 & ~n11905 ;
  assign n29407 = ~n4288 & n15384 ;
  assign n29408 = n5415 | n8635 ;
  assign n29409 = n3151 & ~n29408 ;
  assign n29410 = n10457 & n29409 ;
  assign n29411 = n29410 ^ n8506 ^ n4859 ;
  assign n29412 = n1517 | n10159 ;
  assign n29413 = n10393 & ~n29412 ;
  assign n29414 = n29413 ^ n5716 ^ 1'b0 ;
  assign n29415 = n9816 | n29414 ;
  assign n29416 = n13632 ^ n7715 ^ 1'b0 ;
  assign n29417 = ~n6131 & n10426 ;
  assign n29418 = n29417 ^ n582 ^ 1'b0 ;
  assign n29419 = ~n3426 & n6581 ;
  assign n29420 = n29419 ^ n18758 ^ 1'b0 ;
  assign n29421 = n15809 ^ n3196 ^ 1'b0 ;
  assign n29422 = n14471 ^ n4742 ^ 1'b0 ;
  assign n29423 = n7133 & ~n29422 ;
  assign n29424 = n29423 ^ n25818 ^ n17204 ;
  assign n29425 = n2569 & ~n10299 ;
  assign n29426 = n29425 ^ n415 ^ 1'b0 ;
  assign n29427 = n4892 & ~n19363 ;
  assign n29428 = n12091 & n16316 ;
  assign n29429 = n29428 ^ n5004 ^ 1'b0 ;
  assign n29430 = n29429 ^ n25028 ^ n10326 ;
  assign n29431 = n18100 ^ n17153 ^ 1'b0 ;
  assign n29432 = n9545 ^ n6175 ^ 1'b0 ;
  assign n29433 = n14974 | n17389 ;
  assign n29434 = n29432 | n29433 ;
  assign n29435 = ~n9293 & n29434 ;
  assign n29438 = ~n4605 & n7542 ;
  assign n29436 = n4307 | n12127 ;
  assign n29437 = n8606 | n29436 ;
  assign n29439 = n29438 ^ n29437 ^ 1'b0 ;
  assign n29440 = n13040 ^ n2928 ^ 1'b0 ;
  assign n29441 = n13155 & n29440 ;
  assign n29442 = n1487 & n29441 ;
  assign n29443 = n29442 ^ n12675 ^ 1'b0 ;
  assign n29444 = ~n10723 & n18320 ;
  assign n29445 = n1024 & n29444 ;
  assign n29446 = n6511 ^ n3578 ^ 1'b0 ;
  assign n29447 = n1429 & ~n29446 ;
  assign n29448 = n29447 ^ n8821 ^ n769 ;
  assign n29449 = n29448 ^ n17720 ^ 1'b0 ;
  assign n29450 = n6263 & ~n29449 ;
  assign n29451 = n5783 & n29450 ;
  assign n29452 = n24059 ^ n10040 ^ 1'b0 ;
  assign n29453 = ~n29451 & n29452 ;
  assign n29454 = n1382 & n13329 ;
  assign n29455 = ~n7483 & n9583 ;
  assign n29456 = n29454 & n29455 ;
  assign n29457 = n18024 ^ n12243 ^ n7916 ;
  assign n29461 = n8563 ^ n7979 ^ n1051 ;
  assign n29458 = n25453 ^ n16509 ^ 1'b0 ;
  assign n29459 = n29458 ^ n4187 ^ 1'b0 ;
  assign n29460 = n28138 | n29459 ;
  assign n29462 = n29461 ^ n29460 ^ n15647 ;
  assign n29463 = ( n9423 & n29457 ) | ( n9423 & ~n29462 ) | ( n29457 & ~n29462 ) ;
  assign n29464 = n29463 ^ n17162 ^ n3544 ;
  assign n29465 = n22230 ^ n962 ^ 1'b0 ;
  assign n29466 = n7023 ^ n177 ^ 1'b0 ;
  assign n29467 = n17109 | n29466 ;
  assign n29468 = n29467 ^ n26885 ^ 1'b0 ;
  assign n29469 = n28922 ^ n9923 ^ 1'b0 ;
  assign n29470 = n3153 & n17264 ;
  assign n29471 = ~n13234 & n29470 ;
  assign n29472 = n20320 ^ n11433 ^ n8101 ;
  assign n29473 = ( n5242 & ~n8382 ) | ( n5242 & n21833 ) | ( ~n8382 & n21833 ) ;
  assign n29474 = n20724 ^ n5377 ^ 1'b0 ;
  assign n29475 = n29474 ^ n10002 ^ n216 ;
  assign n29476 = n490 ^ n381 ^ 1'b0 ;
  assign n29477 = n29476 ^ n25039 ^ 1'b0 ;
  assign n29478 = n24101 & ~n29477 ;
  assign n29479 = n22481 ^ n6817 ^ 1'b0 ;
  assign n29480 = ~n5112 & n29479 ;
  assign n29481 = ~n29478 & n29480 ;
  assign n29482 = n494 | n3512 ;
  assign n29483 = n7354 | n29482 ;
  assign n29485 = n29241 ^ n16027 ^ 1'b0 ;
  assign n29484 = n14146 & ~n24019 ;
  assign n29486 = n29485 ^ n29484 ^ 1'b0 ;
  assign n29487 = ( n17976 & n29483 ) | ( n17976 & ~n29486 ) | ( n29483 & ~n29486 ) ;
  assign n29488 = ( ~n261 & n3051 ) | ( ~n261 & n11871 ) | ( n3051 & n11871 ) ;
  assign n29489 = n1801 & ~n24260 ;
  assign n29490 = ~n7025 & n29489 ;
  assign n29491 = n18581 ^ n3991 ^ 1'b0 ;
  assign n29492 = ( n8994 & n12537 ) | ( n8994 & n14137 ) | ( n12537 & n14137 ) ;
  assign n29493 = n5661 & ~n29492 ;
  assign n29494 = ~n23456 & n29493 ;
  assign n29495 = n2615 & ~n9261 ;
  assign n29496 = n16641 | n20496 ;
  assign n29497 = n11084 & ~n14246 ;
  assign n29498 = n2005 & n29497 ;
  assign n29499 = n17894 & ~n29498 ;
  assign n29500 = n861 & n25648 ;
  assign n29501 = ~n25648 & n29500 ;
  assign n29502 = n23778 ^ n14725 ^ 1'b0 ;
  assign n29503 = n89 & n29404 ;
  assign n29504 = n113 & n29503 ;
  assign n29505 = n29349 ^ n833 ^ 1'b0 ;
  assign n29506 = n20306 & ~n29505 ;
  assign n29508 = n24872 ^ n1052 ^ 1'b0 ;
  assign n29509 = n668 | n29508 ;
  assign n29510 = n29509 ^ n13188 ^ 1'b0 ;
  assign n29511 = n14790 & n29510 ;
  assign n29507 = ~n5195 & n22876 ;
  assign n29512 = n29511 ^ n29507 ^ 1'b0 ;
  assign n29513 = n29512 ^ n21749 ^ 1'b0 ;
  assign n29516 = n5205 & ~n7113 ;
  assign n29514 = n16027 & n24777 ;
  assign n29515 = n29514 ^ n3120 ^ 1'b0 ;
  assign n29517 = n29516 ^ n29515 ^ n9406 ;
  assign n29518 = ( ~n2435 & n8220 ) | ( ~n2435 & n29517 ) | ( n8220 & n29517 ) ;
  assign n29519 = ( n7201 & n7338 ) | ( n7201 & n19770 ) | ( n7338 & n19770 ) ;
  assign n29520 = n9996 | n12950 ;
  assign n29521 = n974 | n29520 ;
  assign n29522 = ~n12053 & n14898 ;
  assign n29523 = n11152 ^ n7817 ^ 1'b0 ;
  assign n29524 = n29523 ^ n9598 ^ 1'b0 ;
  assign n29525 = ( n6205 & n15889 ) | ( n6205 & n29524 ) | ( n15889 & n29524 ) ;
  assign n29526 = n1791 & n9120 ;
  assign n29527 = n10574 & n29526 ;
  assign n29528 = n29527 ^ n188 ^ 1'b0 ;
  assign n29529 = n8731 & n29528 ;
  assign n29530 = n27035 ^ n26679 ^ 1'b0 ;
  assign n29531 = n9702 & ~n29530 ;
  assign n29532 = n29531 ^ n14381 ^ 1'b0 ;
  assign n29533 = ~n13348 & n29334 ;
  assign n29534 = n29533 ^ n19675 ^ 1'b0 ;
  assign n29535 = ( n263 & n3696 ) | ( n263 & n8842 ) | ( n3696 & n8842 ) ;
  assign n29536 = n21552 ^ n7854 ^ 1'b0 ;
  assign n29537 = n22699 ^ n21213 ^ 1'b0 ;
  assign n29538 = n29537 ^ n12395 ^ 1'b0 ;
  assign n29539 = ~n2994 & n29538 ;
  assign n29540 = n29539 ^ n10798 ^ 1'b0 ;
  assign n29541 = n13034 ^ n6557 ^ 1'b0 ;
  assign n29542 = n26946 ^ n754 ^ 1'b0 ;
  assign n29543 = ~n29541 & n29542 ;
  assign n29544 = n2377 ^ n1431 ^ 1'b0 ;
  assign n29545 = n29543 & n29544 ;
  assign n29546 = ~n9789 & n16912 ;
  assign n29548 = n1889 & ~n20810 ;
  assign n29549 = n12022 & n29548 ;
  assign n29547 = ~n22897 & n27515 ;
  assign n29550 = n29549 ^ n29547 ^ 1'b0 ;
  assign n29551 = n17621 ^ n9806 ^ n4342 ;
  assign n29552 = n6121 | n29551 ;
  assign n29553 = n29552 ^ n19763 ^ 1'b0 ;
  assign n29554 = n14628 ^ n5570 ^ 1'b0 ;
  assign n29555 = n24011 & ~n29554 ;
  assign n29556 = n29553 & n29555 ;
  assign n29557 = ~n20542 & n21206 ;
  assign n29558 = n29557 ^ n17125 ^ 1'b0 ;
  assign n29559 = n6668 | n17220 ;
  assign n29560 = n4471 & n13265 ;
  assign n29561 = ~n29559 & n29560 ;
  assign n29562 = n655 & n4681 ;
  assign n29563 = n29562 ^ n3260 ^ 1'b0 ;
  assign n29564 = n29563 ^ n19387 ^ n14595 ;
  assign n29565 = n4992 ^ n3236 ^ n524 ;
  assign n29566 = n5494 ^ n871 ^ 1'b0 ;
  assign n29567 = ~n6584 & n29566 ;
  assign n29568 = n29565 & n29567 ;
  assign n29569 = n29568 ^ n19710 ^ 1'b0 ;
  assign n29571 = n20036 ^ n12617 ^ n11653 ;
  assign n29570 = n13421 & ~n18681 ;
  assign n29572 = n29571 ^ n29570 ^ 1'b0 ;
  assign n29573 = n1542 | n10729 ;
  assign n29574 = n24209 & ~n29573 ;
  assign n29575 = n29574 ^ n29375 ^ n2528 ;
  assign n29576 = ~n4671 & n29575 ;
  assign n29577 = ~n29572 & n29576 ;
  assign n29578 = ~n9885 & n24841 ;
  assign n29579 = n21982 & n29578 ;
  assign n29580 = n694 & ~n10630 ;
  assign n29581 = n29580 ^ n4985 ^ 1'b0 ;
  assign n29582 = ~n3274 & n24173 ;
  assign n29583 = ( n2599 & ~n3505 ) | ( n2599 & n29582 ) | ( ~n3505 & n29582 ) ;
  assign n29584 = n3435 & ~n17855 ;
  assign n29585 = ~n4196 & n9436 ;
  assign n29586 = n29585 ^ n1279 ^ 1'b0 ;
  assign n29587 = n29586 ^ n13987 ^ 1'b0 ;
  assign n29588 = n29584 | n29587 ;
  assign n29589 = n29588 ^ n26148 ^ 1'b0 ;
  assign n29590 = n8712 | n19230 ;
  assign n29591 = n6667 & ~n10956 ;
  assign n29592 = n2986 & n19277 ;
  assign n29593 = n29592 ^ n9473 ^ 1'b0 ;
  assign n29594 = n29593 ^ n6076 ^ n4941 ;
  assign n29595 = n6611 ^ n3345 ^ 1'b0 ;
  assign n29596 = n13896 | n29595 ;
  assign n29597 = ( n15770 & ~n29594 ) | ( n15770 & n29596 ) | ( ~n29594 & n29596 ) ;
  assign n29600 = n19066 ^ n3501 ^ 1'b0 ;
  assign n29601 = ~n6979 & n29600 ;
  assign n29598 = n4695 & ~n5180 ;
  assign n29599 = ~n5280 & n29598 ;
  assign n29602 = n29601 ^ n29599 ^ 1'b0 ;
  assign n29603 = n11873 & ~n19178 ;
  assign n29604 = n6890 & ~n18242 ;
  assign n29605 = n19347 ^ n10764 ^ n1179 ;
  assign n29606 = ~n26250 & n29605 ;
  assign n29607 = ~n29604 & n29606 ;
  assign n29608 = n16828 ^ n4240 ^ 1'b0 ;
  assign n29613 = n11393 ^ n2949 ^ 1'b0 ;
  assign n29614 = n25655 & n29613 ;
  assign n29609 = ~n9872 & n14102 ;
  assign n29610 = n16934 ^ x3 ^ 1'b0 ;
  assign n29611 = n29609 & n29610 ;
  assign n29612 = n29611 ^ n27267 ^ n27085 ;
  assign n29615 = n29614 ^ n29612 ^ 1'b0 ;
  assign n29616 = n10228 & n17706 ;
  assign n29617 = n15666 & n29616 ;
  assign n29618 = n19665 | n29617 ;
  assign n29619 = n29618 ^ n19429 ^ 1'b0 ;
  assign n29620 = n22134 ^ n15562 ^ 1'b0 ;
  assign n29621 = ( n14164 & ~n14700 ) | ( n14164 & n29620 ) | ( ~n14700 & n29620 ) ;
  assign n29622 = n18019 & n29621 ;
  assign n29623 = n9811 & n29622 ;
  assign n29625 = n24649 ^ n19389 ^ 1'b0 ;
  assign n29626 = ~n6255 & n29625 ;
  assign n29624 = n6670 & ~n13600 ;
  assign n29627 = n29626 ^ n29624 ^ 1'b0 ;
  assign n29629 = n1962 & ~n24736 ;
  assign n29628 = ~n12006 & n13129 ;
  assign n29630 = n29629 ^ n29628 ^ 1'b0 ;
  assign n29631 = n17042 & n29630 ;
  assign n29633 = n4851 ^ n903 ^ 1'b0 ;
  assign n29634 = ( ~n3867 & n4338 ) | ( ~n3867 & n29633 ) | ( n4338 & n29633 ) ;
  assign n29635 = n29634 ^ n16415 ^ 1'b0 ;
  assign n29632 = n11445 & n17590 ;
  assign n29636 = n29635 ^ n29632 ^ 1'b0 ;
  assign n29637 = ~n4502 & n10273 ;
  assign n29638 = n7988 ^ n7682 ^ 1'b0 ;
  assign n29639 = ~n23261 & n29638 ;
  assign n29640 = ~n4032 & n13228 ;
  assign n29641 = n29639 & n29640 ;
  assign n29642 = n29424 ^ n10881 ^ 1'b0 ;
  assign n29643 = n25345 | n29642 ;
  assign n29644 = n28589 | n29643 ;
  assign n29645 = n23248 | n29644 ;
  assign n29646 = ~n6608 & n15349 ;
  assign n29647 = ~n29645 & n29646 ;
  assign n29648 = n15956 ^ n11782 ^ 1'b0 ;
  assign n29649 = ( n2776 & n12328 ) | ( n2776 & ~n20622 ) | ( n12328 & ~n20622 ) ;
  assign n29650 = n2222 ^ n1011 ^ 1'b0 ;
  assign n29651 = n15535 & n29650 ;
  assign n29652 = n570 | n4729 ;
  assign n29653 = n17099 ^ n2416 ^ 1'b0 ;
  assign n29654 = ( n11400 & n15274 ) | ( n11400 & ~n29653 ) | ( n15274 & ~n29653 ) ;
  assign n29655 = n29654 ^ n7653 ^ 1'b0 ;
  assign n29656 = n29652 & n29655 ;
  assign n29657 = n962 & ~n5491 ;
  assign n29658 = n11028 ^ n5717 ^ n231 ;
  assign n29659 = n29658 ^ n17614 ^ 1'b0 ;
  assign n29660 = ~n7393 & n29659 ;
  assign n29661 = n29660 ^ n16218 ^ 1'b0 ;
  assign n29662 = n29657 & n29661 ;
  assign n29663 = ( n7717 & n16585 ) | ( n7717 & n29662 ) | ( n16585 & n29662 ) ;
  assign n29664 = n14965 ^ n8785 ^ 1'b0 ;
  assign n29665 = ( n7467 & n9713 ) | ( n7467 & ~n29664 ) | ( n9713 & ~n29664 ) ;
  assign n29666 = ~n17142 & n26243 ;
  assign n29667 = ~n8758 & n29666 ;
  assign n29668 = n13243 ^ n3409 ^ n1432 ;
  assign n29669 = n2148 & ~n29668 ;
  assign n29670 = n16796 ^ n3801 ^ 1'b0 ;
  assign n29671 = n12593 ^ n5876 ^ 1'b0 ;
  assign n29672 = n15626 ^ n8227 ^ 1'b0 ;
  assign n29673 = n27904 & ~n29672 ;
  assign n29674 = n10507 ^ n9271 ^ 1'b0 ;
  assign n29675 = n1789 & n5809 ;
  assign n29676 = ~n6909 & n29675 ;
  assign n29677 = n29676 ^ n8866 ^ n7658 ;
  assign n29678 = n22085 ^ n15362 ^ 1'b0 ;
  assign n29679 = n6771 | n23622 ;
  assign n29680 = n29679 ^ n13823 ^ 1'b0 ;
  assign n29681 = n29678 & ~n29680 ;
  assign n29682 = n15297 & n24854 ;
  assign n29683 = n10500 ^ n639 ^ 1'b0 ;
  assign n29684 = ~n8164 & n9849 ;
  assign n29685 = n29684 ^ n2545 ^ 1'b0 ;
  assign n29686 = n4840 & n29685 ;
  assign n29687 = n29683 & n29686 ;
  assign n29688 = ~n19886 & n29687 ;
  assign n29689 = ~n205 & n29688 ;
  assign n29690 = n28867 ^ n9009 ^ 1'b0 ;
  assign n29691 = n4267 & n29690 ;
  assign n29692 = n8086 & ~n18256 ;
  assign n29693 = n29692 ^ n3255 ^ 1'b0 ;
  assign n29694 = n29693 ^ n2397 ^ n1810 ;
  assign n29695 = n16234 ^ n1775 ^ 1'b0 ;
  assign n29696 = n29695 ^ n14316 ^ 1'b0 ;
  assign n29697 = n8056 ^ n4541 ^ 1'b0 ;
  assign n29698 = n5799 & n29438 ;
  assign n29699 = n29697 & n29698 ;
  assign n29701 = n4201 ^ n171 ^ 1'b0 ;
  assign n29704 = n22575 ^ n12767 ^ 1'b0 ;
  assign n29702 = n12631 ^ n11040 ^ 1'b0 ;
  assign n29703 = n11349 | n29702 ;
  assign n29705 = n29704 ^ n29703 ^ 1'b0 ;
  assign n29706 = n29705 ^ n20324 ^ 1'b0 ;
  assign n29707 = n29701 | n29706 ;
  assign n29700 = n8184 & ~n9997 ;
  assign n29708 = n29707 ^ n29700 ^ 1'b0 ;
  assign n29709 = ( n7106 & ~n8903 ) | ( n7106 & n29708 ) | ( ~n8903 & n29708 ) ;
  assign n29710 = n8349 ^ n3835 ^ n2198 ;
  assign n29711 = n6316 & ~n29710 ;
  assign n29712 = ~n29709 & n29711 ;
  assign n29713 = n5118 ^ n5004 ^ 1'b0 ;
  assign n29714 = n3420 & n29713 ;
  assign n29715 = n5241 & n29714 ;
  assign n29716 = n21169 | n28929 ;
  assign n29717 = n10565 ^ n5111 ^ 1'b0 ;
  assign n29718 = ~n29716 & n29717 ;
  assign n29719 = n3156 & ~n11818 ;
  assign n29720 = n29719 ^ n10202 ^ 1'b0 ;
  assign n29721 = n9409 | n10279 ;
  assign n29722 = ( n4628 & ~n5921 ) | ( n4628 & n29721 ) | ( ~n5921 & n29721 ) ;
  assign n29723 = n20049 | n25812 ;
  assign n29724 = n29723 ^ n6215 ^ 1'b0 ;
  assign n29725 = ~n59 & n29408 ;
  assign n29726 = n29725 ^ n19560 ^ n5494 ;
  assign n29727 = n29726 ^ n1178 ^ 1'b0 ;
  assign n29728 = n18063 & ~n21123 ;
  assign n29729 = n29728 ^ n14723 ^ 1'b0 ;
  assign n29730 = n25791 ^ n2028 ^ 1'b0 ;
  assign n29731 = ~n19867 & n29730 ;
  assign n29732 = ~n29729 & n29731 ;
  assign n29733 = n29727 & n29732 ;
  assign n29734 = n4980 | n23064 ;
  assign n29735 = n13743 ^ n508 ^ 1'b0 ;
  assign n29736 = n29735 ^ n16084 ^ 1'b0 ;
  assign n29737 = n13270 ^ n3615 ^ 1'b0 ;
  assign n29738 = n8490 & n29737 ;
  assign n29739 = ~n12537 & n16594 ;
  assign n29740 = n7186 | n20748 ;
  assign n29741 = n29740 ^ n247 ^ 1'b0 ;
  assign n29742 = n12539 & n29741 ;
  assign n29743 = n11069 ^ n9932 ^ 1'b0 ;
  assign n29744 = ~n461 & n29743 ;
  assign n29745 = n13078 & ~n29744 ;
  assign n29746 = n15228 ^ n8392 ^ n3321 ;
  assign n29747 = ~n8656 & n15963 ;
  assign n29748 = n29747 ^ n19791 ^ n612 ;
  assign n29749 = n17590 ^ n13677 ^ n11795 ;
  assign n29750 = n5266 & n16112 ;
  assign n29751 = n7649 & ~n10939 ;
  assign n29752 = n8976 & n29751 ;
  assign n29753 = n16770 ^ n2776 ^ 1'b0 ;
  assign n29754 = n256 & n29753 ;
  assign n29755 = n29754 ^ n17973 ^ 1'b0 ;
  assign n29756 = n29752 | n29755 ;
  assign n29757 = n17299 ^ n8884 ^ 1'b0 ;
  assign n29758 = n21553 ^ n691 ^ 1'b0 ;
  assign n29759 = n5853 | n29758 ;
  assign n29760 = n23588 ^ n11201 ^ 1'b0 ;
  assign n29761 = n1156 & n29760 ;
  assign n29762 = n29759 & n29761 ;
  assign n29763 = ~n6076 & n10236 ;
  assign n29764 = n27407 & n29763 ;
  assign n29765 = n5662 & ~n16785 ;
  assign n29766 = n29765 ^ n15759 ^ 1'b0 ;
  assign n29771 = n15310 | n24482 ;
  assign n29772 = n29771 ^ n5607 ^ 1'b0 ;
  assign n29767 = n7347 | n13382 ;
  assign n29768 = n21851 & n29767 ;
  assign n29769 = ~n9033 & n29768 ;
  assign n29770 = n6399 | n29769 ;
  assign n29773 = n29772 ^ n29770 ^ 1'b0 ;
  assign n29774 = ~n1563 & n7146 ;
  assign n29775 = n10396 ^ n1944 ^ 1'b0 ;
  assign n29776 = ~n29774 & n29775 ;
  assign n29777 = n29776 ^ n14533 ^ 1'b0 ;
  assign n29779 = n13708 ^ n8472 ^ 1'b0 ;
  assign n29780 = ~n12991 & n29779 ;
  assign n29778 = n10598 ^ n1876 ^ n885 ;
  assign n29781 = n29780 ^ n29778 ^ 1'b0 ;
  assign n29782 = n7037 & ~n21037 ;
  assign n29783 = n21403 ^ n8304 ^ 1'b0 ;
  assign n29784 = n25890 ^ n7665 ^ 1'b0 ;
  assign n29785 = n29783 & ~n29784 ;
  assign n29786 = n16805 & ~n20691 ;
  assign n29787 = n600 & n14902 ;
  assign n29788 = n3926 ^ n1577 ^ 1'b0 ;
  assign n29789 = n29788 ^ n20217 ^ n17966 ;
  assign n29790 = n29789 ^ n15874 ^ 1'b0 ;
  assign n29792 = n5941 | n7902 ;
  assign n29793 = n29792 ^ n3128 ^ 1'b0 ;
  assign n29794 = ~n9503 & n27322 ;
  assign n29795 = ~n29793 & n29794 ;
  assign n29791 = n4008 & ~n16591 ;
  assign n29796 = n29795 ^ n29791 ^ 1'b0 ;
  assign n29797 = n5906 ^ n1569 ^ 1'b0 ;
  assign n29798 = n3246 | n13771 ;
  assign n29799 = n7395 & ~n29798 ;
  assign n29800 = n29799 ^ n8153 ^ 1'b0 ;
  assign n29802 = n22324 ^ n11682 ^ 1'b0 ;
  assign n29803 = n9116 & n29802 ;
  assign n29801 = n8156 ^ n2273 ^ 1'b0 ;
  assign n29804 = n29803 ^ n29801 ^ n16168 ;
  assign n29805 = n14145 ^ n11598 ^ n4400 ;
  assign n29806 = ~n15912 & n29805 ;
  assign n29807 = n22985 ^ n7500 ^ 1'b0 ;
  assign n29808 = n6217 | n13109 ;
  assign n29809 = n22812 | n29808 ;
  assign n29810 = n9117 & n29809 ;
  assign n29811 = n18522 ^ n2591 ^ 1'b0 ;
  assign n29812 = n10953 ^ n4294 ^ n2667 ;
  assign n29813 = n10958 & n23294 ;
  assign n29814 = n960 & n965 ;
  assign n29815 = n20609 | n26362 ;
  assign n29816 = n29815 ^ n16572 ^ 1'b0 ;
  assign n29817 = n15729 ^ n5793 ^ 1'b0 ;
  assign n29818 = n8440 & n11862 ;
  assign n29819 = n29818 ^ n4034 ^ 1'b0 ;
  assign n29820 = n2196 & ~n4383 ;
  assign n29821 = n29820 ^ n9160 ^ 1'b0 ;
  assign n29822 = n29819 | n29821 ;
  assign n29823 = n10786 ^ n9377 ^ 1'b0 ;
  assign n29824 = n15439 | n29823 ;
  assign n29825 = n29824 ^ n688 ^ 1'b0 ;
  assign n29826 = n7163 | n29825 ;
  assign n29827 = n10589 ^ n3120 ^ n1630 ;
  assign n29828 = n29826 & n29827 ;
  assign n29829 = n54 & ~n9882 ;
  assign n29830 = n29829 ^ n12748 ^ 1'b0 ;
  assign n29831 = ( ~n3131 & n18539 ) | ( ~n3131 & n29830 ) | ( n18539 & n29830 ) ;
  assign n29832 = ~n11581 & n29831 ;
  assign n29833 = n19567 | n20767 ;
  assign n29834 = n1099 | n29833 ;
  assign n29835 = n5108 | n8577 ;
  assign n29836 = n18912 & n29835 ;
  assign n29837 = n2006 & ~n3760 ;
  assign n29838 = n29837 ^ n7875 ^ n7601 ;
  assign n29839 = n24444 ^ n10333 ^ n7579 ;
  assign n29840 = n29838 & n29839 ;
  assign n29842 = ( ~n6227 & n9879 ) | ( ~n6227 & n12850 ) | ( n9879 & n12850 ) ;
  assign n29841 = ( n7925 & ~n8630 ) | ( n7925 & n11683 ) | ( ~n8630 & n11683 ) ;
  assign n29843 = n29842 ^ n29841 ^ 1'b0 ;
  assign n29844 = n10399 & ~n29843 ;
  assign n29845 = ~n2073 & n4972 ;
  assign n29846 = n29845 ^ n4091 ^ 1'b0 ;
  assign n29847 = n1835 | n29846 ;
  assign n29848 = ~n6460 & n21430 ;
  assign n29849 = n29847 & n29848 ;
  assign n29850 = n18651 | n29849 ;
  assign n29851 = n25706 | n29850 ;
  assign n29852 = ~n5788 & n29851 ;
  assign n29853 = n10633 | n19529 ;
  assign n29854 = n26669 ^ n1071 ^ 1'b0 ;
  assign n29855 = ~n17005 & n29854 ;
  assign n29856 = n4048 & ~n12929 ;
  assign n29857 = n29856 ^ n12222 ^ 1'b0 ;
  assign n29858 = ( n28602 & n29855 ) | ( n28602 & ~n29857 ) | ( n29855 & ~n29857 ) ;
  assign n29859 = n25151 ^ n19909 ^ 1'b0 ;
  assign n29860 = ( n1762 & n3081 ) | ( n1762 & n3630 ) | ( n3081 & n3630 ) ;
  assign n29861 = n4747 & ~n29860 ;
  assign n29862 = n23763 & n29861 ;
  assign n29863 = n25097 ^ n9907 ^ 1'b0 ;
  assign n29864 = n29863 ^ n13539 ^ 1'b0 ;
  assign n29865 = ~n16796 & n29864 ;
  assign n29866 = n13738 ^ n8326 ^ n2987 ;
  assign n29867 = ( n2048 & n6309 ) | ( n2048 & n8204 ) | ( n6309 & n8204 ) ;
  assign n29868 = ( n19068 & n29866 ) | ( n19068 & ~n29867 ) | ( n29866 & ~n29867 ) ;
  assign n29869 = n15617 ^ n1652 ^ 1'b0 ;
  assign n29870 = ( n25159 & n28850 ) | ( n25159 & ~n29869 ) | ( n28850 & ~n29869 ) ;
  assign n29871 = n4142 & ~n6073 ;
  assign n29872 = n29871 ^ n5717 ^ 1'b0 ;
  assign n29873 = n24084 & ~n29872 ;
  assign n29874 = n24567 ^ n20210 ^ 1'b0 ;
  assign n29879 = ~n11517 & n16796 ;
  assign n29875 = n11161 ^ n8911 ^ n7991 ;
  assign n29876 = n29875 ^ n5997 ^ 1'b0 ;
  assign n29877 = n2731 & ~n29876 ;
  assign n29878 = n6521 & ~n29877 ;
  assign n29880 = n29879 ^ n29878 ^ n4242 ;
  assign n29881 = n492 | n1571 ;
  assign n29882 = n16497 | n29881 ;
  assign n29883 = ( n6852 & ~n15097 ) | ( n6852 & n15308 ) | ( ~n15097 & n15308 ) ;
  assign n29884 = n11269 ^ n6811 ^ 1'b0 ;
  assign n29885 = n29883 | n29884 ;
  assign n29886 = n20964 & ~n29885 ;
  assign n29887 = ~n29882 & n29886 ;
  assign n29888 = ( n993 & ~n3540 ) | ( n993 & n16164 ) | ( ~n3540 & n16164 ) ;
  assign n29889 = n12810 ^ n8792 ^ n1204 ;
  assign n29890 = n29889 ^ n10665 ^ 1'b0 ;
  assign n29891 = n18334 | n29890 ;
  assign n29892 = n29888 | n29891 ;
  assign n29893 = n542 | n7534 ;
  assign n29894 = n29893 ^ n6825 ^ 1'b0 ;
  assign n29899 = n5685 | n22084 ;
  assign n29900 = n29899 ^ n23986 ^ n5594 ;
  assign n29895 = n16935 ^ n13025 ^ n4498 ;
  assign n29896 = n11105 ^ n1842 ^ 1'b0 ;
  assign n29897 = ~n29895 & n29896 ;
  assign n29898 = n29897 ^ n26219 ^ 1'b0 ;
  assign n29901 = n29900 ^ n29898 ^ n18289 ;
  assign n29902 = ~n29894 & n29901 ;
  assign n29903 = n29902 ^ n3087 ^ 1'b0 ;
  assign n29905 = n4180 ^ n1175 ^ n23 ;
  assign n29904 = n3466 & ~n5285 ;
  assign n29906 = n29905 ^ n29904 ^ 1'b0 ;
  assign n29907 = n15726 ^ n9372 ^ 1'b0 ;
  assign n29908 = ~n73 & n20695 ;
  assign n29909 = ~n3588 & n12086 ;
  assign n29910 = n3127 & n29909 ;
  assign n29911 = n316 & ~n18453 ;
  assign n29912 = n29911 ^ n3420 ^ 1'b0 ;
  assign n29913 = ~n3459 & n5040 ;
  assign n29914 = n29912 & n29913 ;
  assign n29915 = n29910 & ~n29914 ;
  assign n29916 = ~n12736 & n29915 ;
  assign n29917 = n16010 ^ n7199 ^ 1'b0 ;
  assign n29918 = n20513 ^ n12391 ^ 1'b0 ;
  assign n29919 = n2456 & n29918 ;
  assign n29920 = n1230 | n15065 ;
  assign n29921 = ( n3530 & n4908 ) | ( n3530 & n11914 ) | ( n4908 & n11914 ) ;
  assign n29922 = n9360 & ~n17484 ;
  assign n29923 = ~n25347 & n29922 ;
  assign n29924 = ( n23204 & n29270 ) | ( n23204 & ~n29923 ) | ( n29270 & ~n29923 ) ;
  assign n29926 = n10829 & n24438 ;
  assign n29925 = n1295 & ~n25341 ;
  assign n29927 = n29926 ^ n29925 ^ 1'b0 ;
  assign n29928 = n12964 | n24496 ;
  assign n29929 = n16 & n5614 ;
  assign n29930 = n10120 ^ n5610 ^ 1'b0 ;
  assign n29931 = x0 | n29930 ;
  assign n29933 = n12037 ^ n8508 ^ 1'b0 ;
  assign n29934 = n7472 & n29933 ;
  assign n29935 = n29934 ^ n6656 ^ n230 ;
  assign n29932 = ~n8130 & n11897 ;
  assign n29936 = n29935 ^ n29932 ^ 1'b0 ;
  assign n29937 = n9489 & ~n29936 ;
  assign n29938 = ( ~n4126 & n12690 ) | ( ~n4126 & n14363 ) | ( n12690 & n14363 ) ;
  assign n29939 = n8438 & n8529 ;
  assign n29940 = ~n6212 & n29939 ;
  assign n29941 = n3950 & ~n29940 ;
  assign n29942 = ~n29938 & n29941 ;
  assign n29943 = n29942 ^ n4587 ^ 1'b0 ;
  assign n29944 = n9986 | n28670 ;
  assign n29945 = n6345 ^ n3767 ^ 1'b0 ;
  assign n29946 = n3330 & n12852 ;
  assign n29947 = n6221 & ~n10425 ;
  assign n29948 = ~n20027 & n29947 ;
  assign n29949 = ( n18226 & n19894 ) | ( n18226 & ~n29948 ) | ( n19894 & ~n29948 ) ;
  assign n29950 = n13248 & ~n16034 ;
  assign n29951 = ~n7890 & n25206 ;
  assign n29952 = ~n1891 & n29951 ;
  assign n29953 = ~n28432 & n29952 ;
  assign n29954 = n28380 ^ n9858 ^ 1'b0 ;
  assign n29955 = n18634 & n29954 ;
  assign n29956 = n1560 & n7361 ;
  assign n29957 = n29956 ^ n7055 ^ 1'b0 ;
  assign n29958 = n9624 & ~n23388 ;
  assign n29959 = n3005 ^ n2677 ^ 1'b0 ;
  assign n29960 = n12051 | n29959 ;
  assign n29961 = n3568 & n16060 ;
  assign n29962 = ~n29960 & n29961 ;
  assign n29963 = n1292 & n24355 ;
  assign n29964 = n29963 ^ n8177 ^ 1'b0 ;
  assign n29965 = n6051 ^ n5061 ^ 1'b0 ;
  assign n29966 = n5697 | n29965 ;
  assign n29967 = n10559 | n29966 ;
  assign n29968 = n29474 & ~n29967 ;
  assign n29969 = n8490 ^ n183 ^ 1'b0 ;
  assign n29970 = n6240 & ~n20444 ;
  assign n29971 = n1424 | n29970 ;
  assign n29972 = n29971 ^ n23674 ^ 1'b0 ;
  assign n29973 = n19613 ^ n8106 ^ 1'b0 ;
  assign n29974 = n8318 ^ n1143 ^ 1'b0 ;
  assign n29975 = n1160 & ~n29974 ;
  assign n29976 = n29975 ^ n29558 ^ n11190 ;
  assign n29977 = n11997 ^ n4421 ^ 1'b0 ;
  assign n29978 = n5064 | n15850 ;
  assign n29979 = n9755 ^ n3464 ^ 1'b0 ;
  assign n29980 = n12898 & ~n29872 ;
  assign n29983 = n2798 & n7580 ;
  assign n29981 = ~n9201 & n23211 ;
  assign n29982 = n29981 ^ n24852 ^ 1'b0 ;
  assign n29984 = n29983 ^ n29982 ^ 1'b0 ;
  assign n29985 = n12937 & ~n29984 ;
  assign n29986 = n12967 ^ n475 ^ 1'b0 ;
  assign n29987 = n14369 & n29986 ;
  assign n29988 = ~n4637 & n29987 ;
  assign n29989 = ( n13865 & ~n22421 ) | ( n13865 & n29988 ) | ( ~n22421 & n29988 ) ;
  assign n29990 = n29989 ^ n12817 ^ 1'b0 ;
  assign n29991 = n18519 ^ n2050 ^ n1296 ;
  assign n29992 = n1006 & ~n29991 ;
  assign n29993 = n8888 & ~n9020 ;
  assign n29994 = n29993 ^ n24285 ^ n6245 ;
  assign n29995 = ( n11314 & n15009 ) | ( n11314 & n15029 ) | ( n15009 & n15029 ) ;
  assign n29996 = n1154 | n7149 ;
  assign n29997 = n28223 & ~n29996 ;
  assign n29998 = n27180 | n29997 ;
  assign n29999 = n24493 | n29998 ;
  assign n30000 = n465 & ~n3137 ;
  assign n30001 = ~n5127 & n21525 ;
  assign n30002 = n4788 & n30001 ;
  assign n30003 = n30002 ^ n1201 ^ 1'b0 ;
  assign n30004 = n23695 ^ n5963 ^ 1'b0 ;
  assign n30005 = n563 & n18048 ;
  assign n30006 = n2770 ^ n1081 ^ 1'b0 ;
  assign n30007 = n13211 & ~n30006 ;
  assign n30008 = n30007 ^ n24032 ^ n18841 ;
  assign n30009 = ( n10422 & n12658 ) | ( n10422 & ~n22097 ) | ( n12658 & ~n22097 ) ;
  assign n30010 = n16399 & ~n30009 ;
  assign n30011 = n30010 ^ n5546 ^ 1'b0 ;
  assign n30015 = ~n15209 & n17036 ;
  assign n30016 = n18311 & n30015 ;
  assign n30017 = n18701 & n30016 ;
  assign n30012 = n19656 ^ n3941 ^ 1'b0 ;
  assign n30013 = n191 | n30012 ;
  assign n30014 = n2352 & ~n30013 ;
  assign n30018 = n30017 ^ n30014 ^ 1'b0 ;
  assign n30019 = n21936 ^ n19884 ^ n2170 ;
  assign n30020 = n3628 | n6353 ;
  assign n30021 = n4858 ^ n1779 ^ 1'b0 ;
  assign n30022 = n1936 & n26162 ;
  assign n30023 = n14858 ^ n8407 ^ 1'b0 ;
  assign n30024 = n10662 | n13695 ;
  assign n30025 = n30024 ^ n6511 ^ 1'b0 ;
  assign n30026 = n5477 & n30025 ;
  assign n30027 = n4508 & ~n30026 ;
  assign n30028 = n7354 ^ n7225 ^ 1'b0 ;
  assign n30029 = ~n4530 & n6163 ;
  assign n30030 = n30029 ^ n572 ^ 1'b0 ;
  assign n30031 = n2354 & ~n30030 ;
  assign n30032 = n30031 ^ n3932 ^ x6 ;
  assign n30033 = n30028 & ~n30032 ;
  assign n30034 = n12858 & ~n24168 ;
  assign n30037 = n3739 & n6810 ;
  assign n30035 = n9339 & n18981 ;
  assign n30036 = ( n6082 & n14335 ) | ( n6082 & ~n30035 ) | ( n14335 & ~n30035 ) ;
  assign n30038 = n30037 ^ n30036 ^ n7354 ;
  assign n30039 = n19946 ^ n2064 ^ 1'b0 ;
  assign n30040 = n5225 | n12090 ;
  assign n30041 = n14692 ^ n12460 ^ 1'b0 ;
  assign n30042 = n16321 | n30041 ;
  assign n30043 = ~n1100 & n14981 ;
  assign n30044 = n11116 | n30043 ;
  assign n30050 = n6699 ^ n1094 ^ 1'b0 ;
  assign n30045 = n6352 | n15344 ;
  assign n30046 = n30045 ^ n9843 ^ 1'b0 ;
  assign n30047 = n3260 | n30046 ;
  assign n30048 = ~n4203 & n30047 ;
  assign n30049 = n30048 ^ n4313 ^ 1'b0 ;
  assign n30051 = n30050 ^ n30049 ^ 1'b0 ;
  assign n30052 = n2797 & ~n30051 ;
  assign n30053 = n2618 & n30052 ;
  assign n30054 = n30053 ^ n13671 ^ 1'b0 ;
  assign n30057 = n3455 ^ n2837 ^ 1'b0 ;
  assign n30058 = n9376 ^ n5924 ^ n1928 ;
  assign n30059 = n8663 & n30058 ;
  assign n30060 = ~n30057 & n30059 ;
  assign n30055 = n23806 ^ n21474 ^ n18239 ;
  assign n30056 = ~n23027 & n30055 ;
  assign n30061 = n30060 ^ n30056 ^ 1'b0 ;
  assign n30062 = n388 & ~n15340 ;
  assign n30063 = n16001 ^ n49 ^ 1'b0 ;
  assign n30064 = n30062 | n30063 ;
  assign n30065 = n30064 ^ n15930 ^ 1'b0 ;
  assign n30066 = n7631 | n9416 ;
  assign n30067 = n11356 | n30066 ;
  assign n30071 = n4272 & n7098 ;
  assign n30068 = n11025 & ~n25792 ;
  assign n30069 = ~n27353 & n30068 ;
  assign n30070 = n30069 ^ n3747 ^ 1'b0 ;
  assign n30072 = n30071 ^ n30070 ^ n25601 ;
  assign n30073 = n10163 ^ n9787 ^ 1'b0 ;
  assign n30074 = n7150 & n30073 ;
  assign n30075 = ~n3957 & n30074 ;
  assign n30076 = n1183 & ~n14295 ;
  assign n30077 = n281 & n30076 ;
  assign n30078 = n30077 ^ n10576 ^ 1'b0 ;
  assign n30079 = n2740 & n30078 ;
  assign n30080 = n30079 ^ n21640 ^ n11628 ;
  assign n30081 = ~n30075 & n30080 ;
  assign n30082 = n30081 ^ n1214 ^ 1'b0 ;
  assign n30083 = n3968 ^ n670 ^ 1'b0 ;
  assign n30084 = n14786 & ~n27267 ;
  assign n30085 = ~n30083 & n30084 ;
  assign n30086 = n4308 | n15916 ;
  assign n30087 = n30086 ^ n15207 ^ 1'b0 ;
  assign n30088 = n25812 ^ n2070 ^ 1'b0 ;
  assign n30089 = n40 & n5828 ;
  assign n30090 = n30089 ^ n5061 ^ 1'b0 ;
  assign n30091 = ( n15078 & n15420 ) | ( n15078 & n30090 ) | ( n15420 & n30090 ) ;
  assign n30092 = ( n4164 & n30088 ) | ( n4164 & ~n30091 ) | ( n30088 & ~n30091 ) ;
  assign n30093 = ( n850 & n19987 ) | ( n850 & n22950 ) | ( n19987 & n22950 ) ;
  assign n30094 = n5683 & ~n23606 ;
  assign n30095 = n3595 & n3835 ;
  assign n30096 = n30095 ^ n3949 ^ 1'b0 ;
  assign n30097 = ~n30094 & n30096 ;
  assign n30098 = n30097 ^ n30087 ^ 1'b0 ;
  assign n30099 = n14356 | n18500 ;
  assign n30100 = ~n19775 & n30099 ;
  assign n30101 = n3897 & ~n28534 ;
  assign n30102 = ( n15263 & n15573 ) | ( n15263 & n30101 ) | ( n15573 & n30101 ) ;
  assign n30103 = n12992 & n14646 ;
  assign n30104 = n30103 ^ n2617 ^ 1'b0 ;
  assign n30105 = n3043 | n4359 ;
  assign n30106 = n5688 | n10443 ;
  assign n30107 = n7678 & ~n30106 ;
  assign n30108 = n10511 ^ n6289 ^ n3690 ;
  assign n30109 = n15443 & n30108 ;
  assign n30110 = n30107 & n30109 ;
  assign n30111 = n3351 | n30110 ;
  assign n30112 = n30105 & ~n30111 ;
  assign n30115 = n3885 | n10361 ;
  assign n30116 = n1091 | n30115 ;
  assign n30113 = n5557 ^ n2911 ^ 1'b0 ;
  assign n30114 = n27107 | n30113 ;
  assign n30117 = n30116 ^ n30114 ^ 1'b0 ;
  assign n30118 = n8242 & n30117 ;
  assign n30119 = n30118 ^ n11231 ^ 1'b0 ;
  assign n30120 = n2382 | n3884 ;
  assign n30121 = n30120 ^ n1125 ^ 1'b0 ;
  assign n30122 = n14918 & ~n23607 ;
  assign n30123 = ~n10068 & n30122 ;
  assign n30124 = ~n9162 & n18089 ;
  assign n30125 = n15056 & n30124 ;
  assign n30126 = ~n30123 & n30125 ;
  assign n30127 = n352 | n7273 ;
  assign n30128 = n890 & n30127 ;
  assign n30129 = n30128 ^ n22263 ^ n4825 ;
  assign n30130 = ~n3691 & n6815 ;
  assign n30131 = n3899 & n4555 ;
  assign n30132 = n2294 & n30131 ;
  assign n30133 = n30132 ^ n14872 ^ 1'b0 ;
  assign n30134 = n11154 | n16136 ;
  assign n30135 = n20428 ^ n12596 ^ 1'b0 ;
  assign n30136 = n1079 | n30135 ;
  assign n30137 = n29688 ^ n5253 ^ 1'b0 ;
  assign n30138 = n10507 | n20269 ;
  assign n30139 = ( ~n11667 & n16070 ) | ( ~n11667 & n30138 ) | ( n16070 & n30138 ) ;
  assign n30140 = ( n11128 & n14622 ) | ( n11128 & ~n30139 ) | ( n14622 & ~n30139 ) ;
  assign n30141 = ( n179 & n1781 ) | ( n179 & ~n10088 ) | ( n1781 & ~n10088 ) ;
  assign n30142 = ~n18761 & n24918 ;
  assign n30143 = n30142 ^ n16828 ^ 1'b0 ;
  assign n30144 = n9146 & n30143 ;
  assign n30145 = n30144 ^ n26069 ^ 1'b0 ;
  assign n30146 = n13670 | n27600 ;
  assign n30147 = n2469 & ~n6319 ;
  assign n30148 = n15036 & ~n30147 ;
  assign n30149 = n10400 & n17401 ;
  assign n30150 = ~n30047 & n30149 ;
  assign n30151 = n3505 & ~n13335 ;
  assign n30152 = n1201 & n30151 ;
  assign n30153 = n3899 ^ n1779 ^ 1'b0 ;
  assign n30154 = n30153 ^ n17364 ^ n12637 ;
  assign n30155 = ~n1940 & n11009 ;
  assign n30156 = n30155 ^ n1447 ^ 1'b0 ;
  assign n30157 = n30156 ^ n6381 ^ 1'b0 ;
  assign n30158 = n30154 & n30157 ;
  assign n30159 = n30158 ^ n24538 ^ n21266 ;
  assign n30160 = n9311 ^ n1412 ^ 1'b0 ;
  assign n30161 = ~n6032 & n28118 ;
  assign n30162 = ~n11329 & n30161 ;
  assign n30163 = n30162 ^ n3879 ^ 1'b0 ;
  assign n30164 = ~n29448 & n30163 ;
  assign n30165 = ~n30160 & n30164 ;
  assign n30166 = n26672 ^ n5806 ^ 1'b0 ;
  assign n30167 = n14208 ^ n1842 ^ 1'b0 ;
  assign n30168 = n29586 & n30167 ;
  assign n30169 = n8408 & ~n30168 ;
  assign n30170 = n30169 ^ n20662 ^ n5074 ;
  assign n30171 = x1 & ~n14731 ;
  assign n30172 = n30170 & ~n30171 ;
  assign n30173 = n16233 & ~n29302 ;
  assign n30174 = n25633 ^ n5716 ^ n923 ;
  assign n30175 = n1013 | n14606 ;
  assign n30176 = n647 | n30175 ;
  assign n30177 = n30176 ^ n10591 ^ 1'b0 ;
  assign n30178 = n24444 | n30177 ;
  assign n30179 = n27303 ^ n15781 ^ n913 ;
  assign n30180 = n28308 & ~n30179 ;
  assign n30181 = ( n3793 & ~n14972 ) | ( n3793 & n26537 ) | ( ~n14972 & n26537 ) ;
  assign n30182 = n18421 ^ n15958 ^ 1'b0 ;
  assign n30183 = n14445 & ~n30182 ;
  assign n30184 = n17520 | n24117 ;
  assign n30185 = n27560 ^ n15513 ^ n607 ;
  assign n30186 = n9811 & ~n30185 ;
  assign n30187 = ~n21755 & n29131 ;
  assign n30188 = n30187 ^ n1679 ^ 1'b0 ;
  assign n30189 = n29077 ^ n20984 ^ n20931 ;
  assign n30190 = x10 & ~n13654 ;
  assign n30191 = ~n174 & n30190 ;
  assign n30192 = n30191 ^ n18115 ^ 1'b0 ;
  assign n30193 = ( ~n11443 & n13015 ) | ( ~n11443 & n18888 ) | ( n13015 & n18888 ) ;
  assign n30194 = ~n23578 & n26766 ;
  assign n30195 = n13712 ^ n2070 ^ 1'b0 ;
  assign n30196 = n6968 & ~n30195 ;
  assign n30197 = n6805 & ~n12091 ;
  assign n30198 = ~n30196 & n30197 ;
  assign n30199 = n30198 ^ n20279 ^ 1'b0 ;
  assign n30200 = n3464 & n12536 ;
  assign n30201 = n30200 ^ n6804 ^ 1'b0 ;
  assign n30202 = n30201 ^ n19135 ^ n13677 ;
  assign n30203 = n16164 ^ n287 ^ 1'b0 ;
  assign n30204 = ~n30202 & n30203 ;
  assign n30205 = n6802 & n12691 ;
  assign n30206 = ~n30204 & n30205 ;
  assign n30207 = n4180 | n8638 ;
  assign n30208 = n2716 & n12214 ;
  assign n30209 = ( n7055 & n14112 ) | ( n7055 & n17640 ) | ( n14112 & n17640 ) ;
  assign n30210 = n30209 ^ n9552 ^ n2617 ;
  assign n30211 = n2076 & ~n19283 ;
  assign n30213 = n18711 ^ n230 ^ 1'b0 ;
  assign n30214 = n12606 | n30213 ;
  assign n30212 = ~n23980 & n25833 ;
  assign n30215 = n30214 ^ n30212 ^ 1'b0 ;
  assign n30216 = n4086 | n8514 ;
  assign n30217 = n30216 ^ n17023 ^ 1'b0 ;
  assign n30218 = n5925 & ~n6205 ;
  assign n30219 = ~n63 & n30218 ;
  assign n30220 = ~n30217 & n30219 ;
  assign n30221 = n7137 ^ n1825 ^ 1'b0 ;
  assign n30222 = n30220 & ~n30221 ;
  assign n30223 = ~n17169 & n24772 ;
  assign n30224 = n5581 & n30223 ;
  assign n30225 = n11956 | n30224 ;
  assign n30226 = ~n12267 & n29548 ;
  assign n30229 = n1439 & ~n2631 ;
  assign n30230 = ~n3245 & n30229 ;
  assign n30227 = n4377 & ~n9126 ;
  assign n30228 = ~n5803 & n30227 ;
  assign n30231 = n30230 ^ n30228 ^ n13945 ;
  assign n30232 = n30226 & ~n30231 ;
  assign n30233 = n14606 & n30232 ;
  assign n30234 = ~n481 & n5420 ;
  assign n30235 = n30234 ^ n4918 ^ 1'b0 ;
  assign n30236 = n30235 ^ n18237 ^ n10326 ;
  assign n30237 = n11844 | n30236 ;
  assign n30238 = ( n10777 & n12155 ) | ( n10777 & n13538 ) | ( n12155 & n13538 ) ;
  assign n30239 = n25042 ^ n15592 ^ 1'b0 ;
  assign n30240 = ( ~n21667 & n26630 ) | ( ~n21667 & n30239 ) | ( n26630 & n30239 ) ;
  assign n30241 = n9765 ^ n1296 ^ 1'b0 ;
  assign n30242 = ~n13258 & n30241 ;
  assign n30243 = n22739 ^ n1088 ^ 1'b0 ;
  assign n30244 = n30242 & n30243 ;
  assign n30245 = ~n23387 & n29455 ;
  assign n30246 = ~n11360 & n30245 ;
  assign n30247 = n19632 & ~n29203 ;
  assign n30248 = n30247 ^ n13473 ^ 1'b0 ;
  assign n30251 = ( ~n95 & n524 ) | ( ~n95 & n3998 ) | ( n524 & n3998 ) ;
  assign n30249 = n11273 & ~n23239 ;
  assign n30250 = n26162 & n30249 ;
  assign n30252 = n30251 ^ n30250 ^ 1'b0 ;
  assign n30253 = n22776 ^ n478 ^ 1'b0 ;
  assign n30254 = n24162 & n30253 ;
  assign n30255 = n11936 & ~n16605 ;
  assign n30256 = n9832 & n30255 ;
  assign n30257 = n30256 ^ n9875 ^ 1'b0 ;
  assign n30258 = n24412 ^ n1563 ^ 1'b0 ;
  assign n30259 = n22539 ^ n6657 ^ 1'b0 ;
  assign n30260 = n373 & n30259 ;
  assign n30261 = n5997 & ~n28492 ;
  assign n30262 = n30260 & n30261 ;
  assign n30263 = n16618 | n30262 ;
  assign n30264 = n7226 | n9905 ;
  assign n30265 = n30264 ^ n6596 ^ 1'b0 ;
  assign n30266 = n7233 & ~n10539 ;
  assign n30267 = n30266 ^ n29121 ^ 1'b0 ;
  assign n30268 = n24462 | n30267 ;
  assign n30269 = n30268 ^ n3020 ^ 1'b0 ;
  assign n30270 = n18076 & ~n26699 ;
  assign n30271 = ~n3062 & n30270 ;
  assign n30272 = ( n6831 & n18263 ) | ( n6831 & n21057 ) | ( n18263 & n21057 ) ;
  assign n30273 = n24380 ^ n5581 ^ 1'b0 ;
  assign n30274 = ~n176 & n8733 ;
  assign n30275 = n30274 ^ n16378 ^ 1'b0 ;
  assign n30276 = ( n17057 & n30273 ) | ( n17057 & n30275 ) | ( n30273 & n30275 ) ;
  assign n30277 = n30276 ^ n13987 ^ n4275 ;
  assign n30278 = ~n4987 & n26481 ;
  assign n30279 = ~n1578 & n30278 ;
  assign n30280 = n2296 & ~n9826 ;
  assign n30281 = ~n8383 & n30280 ;
  assign n30282 = n30281 ^ n16118 ^ 1'b0 ;
  assign n30283 = ~n1068 & n2734 ;
  assign n30284 = n18982 ^ n2060 ^ 1'b0 ;
  assign n30285 = ~n1853 & n2785 ;
  assign n30286 = n30285 ^ n28301 ^ 1'b0 ;
  assign n30287 = n9100 | n18124 ;
  assign n30288 = n9852 & ~n20896 ;
  assign n30289 = ~n11864 & n30288 ;
  assign n30290 = n30289 ^ n7315 ^ 1'b0 ;
  assign n30291 = n12668 ^ n9325 ^ 1'b0 ;
  assign n30292 = n5012 & n30291 ;
  assign n30293 = ~n29596 & n30292 ;
  assign n30298 = ~n2440 & n13881 ;
  assign n30299 = n321 & n30298 ;
  assign n30294 = n164 & n12304 ;
  assign n30295 = ~n2504 & n30294 ;
  assign n30296 = n30295 ^ n536 ^ 1'b0 ;
  assign n30297 = n263 | n30296 ;
  assign n30300 = n30299 ^ n30297 ^ n24200 ;
  assign n30301 = n30300 ^ n4536 ^ 1'b0 ;
  assign n30302 = n8625 | n30301 ;
  assign n30303 = ~n17449 & n22785 ;
  assign n30304 = ~n20638 & n30303 ;
  assign n30305 = n8629 & n10118 ;
  assign n30306 = n2650 | n27303 ;
  assign n30307 = n5691 | n30306 ;
  assign n30308 = n111 | n8291 ;
  assign n30309 = n30307 | n30308 ;
  assign n30310 = n3469 | n22362 ;
  assign n30311 = n30310 ^ n10120 ^ 1'b0 ;
  assign n30312 = n29513 & ~n30311 ;
  assign n30313 = n15904 ^ n4690 ^ 1'b0 ;
  assign n30314 = n2674 & n20097 ;
  assign n30315 = n30314 ^ n9325 ^ 1'b0 ;
  assign n30316 = n3508 & n11791 ;
  assign n30317 = ~n9576 & n30316 ;
  assign n30318 = n15984 | n30317 ;
  assign n30319 = n9011 & ~n30318 ;
  assign n30320 = n30319 ^ n6435 ^ 1'b0 ;
  assign n30321 = ~n2986 & n30320 ;
  assign n30322 = ( ~n7896 & n24703 ) | ( ~n7896 & n30321 ) | ( n24703 & n30321 ) ;
  assign n30323 = ~n6902 & n26708 ;
  assign n30324 = n30323 ^ n8376 ^ 1'b0 ;
  assign n30325 = n203 & n30324 ;
  assign n30326 = n30325 ^ n5707 ^ 1'b0 ;
  assign n30327 = n30326 ^ n48 ^ 1'b0 ;
  assign n30328 = n30322 & n30327 ;
  assign n30329 = n29704 ^ n18681 ^ 1'b0 ;
  assign n30330 = ( n19553 & n22951 ) | ( n19553 & ~n30329 ) | ( n22951 & ~n30329 ) ;
  assign n30333 = ( n10801 & ~n11475 ) | ( n10801 & n23964 ) | ( ~n11475 & n23964 ) ;
  assign n30331 = n11949 ^ n3704 ^ 1'b0 ;
  assign n30332 = ( ~n7762 & n8644 ) | ( ~n7762 & n30331 ) | ( n8644 & n30331 ) ;
  assign n30334 = n30333 ^ n30332 ^ 1'b0 ;
  assign n30336 = ~n5251 & n5622 ;
  assign n30337 = n7214 | n30336 ;
  assign n30338 = n21723 & ~n30337 ;
  assign n30335 = n22750 & n29107 ;
  assign n30339 = n30338 ^ n30335 ^ 1'b0 ;
  assign n30340 = n30334 & n30339 ;
  assign n30341 = n10350 ^ n3375 ^ 1'b0 ;
  assign n30342 = n30341 ^ n22892 ^ n18981 ;
  assign n30343 = n29324 ^ n19159 ^ 1'b0 ;
  assign n30344 = n28118 & n30343 ;
  assign n30345 = ( n8429 & n17364 ) | ( n8429 & n26789 ) | ( n17364 & n26789 ) ;
  assign n30346 = n30345 ^ n24894 ^ 1'b0 ;
  assign n30347 = n17130 ^ n15955 ^ n4941 ;
  assign n30348 = ( ~n6380 & n27149 ) | ( ~n6380 & n30347 ) | ( n27149 & n30347 ) ;
  assign n30349 = n27390 ^ n10737 ^ 1'b0 ;
  assign n30350 = n19186 ^ n2648 ^ 1'b0 ;
  assign n30351 = n30350 ^ n2335 ^ 1'b0 ;
  assign n30352 = n11756 | n30351 ;
  assign n30353 = n25760 ^ n1964 ^ 1'b0 ;
  assign n30354 = n6221 & ~n30353 ;
  assign n30355 = n10397 | n14598 ;
  assign n30356 = n2067 & ~n30355 ;
  assign n30357 = n13481 | n30356 ;
  assign n30358 = n2583 | n28373 ;
  assign n30359 = n30358 ^ n21425 ^ 1'b0 ;
  assign n30360 = n8878 & n21001 ;
  assign n30361 = n7831 & ~n30360 ;
  assign n30362 = n27035 & n30361 ;
  assign n30363 = n30362 ^ n25279 ^ n7544 ;
  assign n30374 = n10229 ^ n6487 ^ n6052 ;
  assign n30371 = n17614 ^ n2977 ^ 1'b0 ;
  assign n30372 = n30371 ^ n2657 ^ 1'b0 ;
  assign n30373 = ~n18190 & n30372 ;
  assign n30368 = n17488 & n25760 ;
  assign n30369 = n30368 ^ n3554 ^ 1'b0 ;
  assign n30364 = n18002 ^ n11781 ^ n1300 ;
  assign n30365 = ~n18461 & n30364 ;
  assign n30366 = n8063 & n30365 ;
  assign n30367 = n2517 | n30366 ;
  assign n30370 = n30369 ^ n30367 ^ 1'b0 ;
  assign n30375 = n30374 ^ n30373 ^ n30370 ;
  assign n30377 = ( n3214 & n3459 ) | ( n3214 & n24841 ) | ( n3459 & n24841 ) ;
  assign n30376 = n5331 & ~n25397 ;
  assign n30378 = n30377 ^ n30376 ^ 1'b0 ;
  assign n30380 = ~n10452 & n15512 ;
  assign n30381 = n29987 & ~n30380 ;
  assign n30382 = n4815 & n30381 ;
  assign n30379 = n797 | n25159 ;
  assign n30383 = n30382 ^ n30379 ^ 1'b0 ;
  assign n30384 = n5479 ^ n1315 ^ 1'b0 ;
  assign n30385 = n7770 & n30384 ;
  assign n30386 = ~n14509 & n30385 ;
  assign n30387 = n25421 | n30386 ;
  assign n30388 = n28774 & ~n30387 ;
  assign n30389 = n9086 & n13141 ;
  assign n30390 = n6957 & n19199 ;
  assign n30391 = n6398 ^ n4569 ^ 1'b0 ;
  assign n30392 = n30391 ^ n16168 ^ 1'b0 ;
  assign n30393 = n10163 & ~n30392 ;
  assign n30394 = n30393 ^ n12727 ^ 1'b0 ;
  assign n30395 = n26518 ^ n2581 ^ 1'b0 ;
  assign n30396 = n30394 & ~n30395 ;
  assign n30397 = n12921 ^ n1043 ^ 1'b0 ;
  assign n30398 = n8789 ^ n102 ^ n55 ;
  assign n30399 = n14232 ^ n5109 ^ 1'b0 ;
  assign n30400 = n3531 & ~n30399 ;
  assign n30401 = ~n11961 & n30400 ;
  assign n30402 = n30401 ^ n24189 ^ 1'b0 ;
  assign n30403 = n30398 & n30402 ;
  assign n30404 = ~n1154 & n2961 ;
  assign n30405 = x10 & n30404 ;
  assign n30406 = n1160 | n30405 ;
  assign n30407 = ( ~n1078 & n2770 ) | ( ~n1078 & n29034 ) | ( n2770 & n29034 ) ;
  assign n30408 = n30406 & ~n30407 ;
  assign n30409 = n28195 & n30408 ;
  assign n30410 = n19267 ^ n4447 ^ n431 ;
  assign n30411 = n21417 ^ n8721 ^ 1'b0 ;
  assign n30412 = n22661 & ~n30411 ;
  assign n30413 = n24485 & ~n27538 ;
  assign n30414 = n22797 ^ n10939 ^ n4305 ;
  assign n30415 = n6100 ^ n5373 ^ 1'b0 ;
  assign n30416 = n10741 & ~n30415 ;
  assign n30417 = n30416 ^ n27979 ^ 1'b0 ;
  assign n30419 = ( ~n10411 & n14175 ) | ( ~n10411 & n14350 ) | ( n14175 & n14350 ) ;
  assign n30420 = n3878 & ~n30419 ;
  assign n30418 = n17034 & n24327 ;
  assign n30421 = n30420 ^ n30418 ^ n22372 ;
  assign n30422 = n6417 ^ n3069 ^ 1'b0 ;
  assign n30423 = n30422 ^ n6498 ^ 1'b0 ;
  assign n30424 = n9631 & ~n28929 ;
  assign n30425 = n2558 & n30424 ;
  assign n30426 = ~n15867 & n30425 ;
  assign n30427 = n5736 & ~n12010 ;
  assign n30428 = n11974 & ~n15876 ;
  assign n30429 = ~n30427 & n30428 ;
  assign n30430 = n8451 | n13056 ;
  assign n30431 = n4852 & ~n30430 ;
  assign n30432 = n29767 ^ n3345 ^ 1'b0 ;
  assign n30433 = ( n2050 & n3703 ) | ( n2050 & n30432 ) | ( n3703 & n30432 ) ;
  assign n30434 = n4987 ^ n2472 ^ 1'b0 ;
  assign n30435 = ~n5885 & n30434 ;
  assign n30436 = ( n30431 & ~n30433 ) | ( n30431 & n30435 ) | ( ~n30433 & n30435 ) ;
  assign n30438 = n15933 ^ n12233 ^ 1'b0 ;
  assign n30437 = n16616 & ~n18924 ;
  assign n30439 = n30438 ^ n30437 ^ 1'b0 ;
  assign n30440 = n8725 | n30439 ;
  assign n30441 = n27048 ^ n23565 ^ n10465 ;
  assign n30442 = n30441 ^ n2457 ^ 1'b0 ;
  assign n30443 = n26852 & n30442 ;
  assign n30444 = n30443 ^ n29302 ^ 1'b0 ;
  assign n30445 = n4432 & ~n30444 ;
  assign n30446 = n20971 | n30445 ;
  assign n30447 = n2466 & ~n30446 ;
  assign n30448 = n7479 ^ n3667 ^ 1'b0 ;
  assign n30449 = n22094 & n30448 ;
  assign n30450 = n27208 | n30449 ;
  assign n30456 = ( n442 & n5594 ) | ( n442 & n17818 ) | ( n5594 & n17818 ) ;
  assign n30451 = n10551 ^ n1300 ^ 1'b0 ;
  assign n30452 = n16864 & ~n23760 ;
  assign n30453 = ~n30451 & n30452 ;
  assign n30454 = n24715 & ~n30453 ;
  assign n30455 = n30454 ^ n17089 ^ 1'b0 ;
  assign n30457 = n30456 ^ n30455 ^ 1'b0 ;
  assign n30458 = n30450 & ~n30457 ;
  assign n30460 = ~n5274 & n11002 ;
  assign n30461 = ~n16092 & n30460 ;
  assign n30459 = n99 | n216 ;
  assign n30462 = n30461 ^ n30459 ^ 1'b0 ;
  assign n30463 = n11134 & n29458 ;
  assign n30464 = ~n594 & n30463 ;
  assign n30465 = ( n4536 & ~n10670 ) | ( n4536 & n28795 ) | ( ~n10670 & n28795 ) ;
  assign n30466 = n30465 ^ n14593 ^ n1024 ;
  assign n30467 = n15932 ^ n14089 ^ 1'b0 ;
  assign n30468 = n30466 & ~n30467 ;
  assign n30469 = ( ~n2940 & n5037 ) | ( ~n2940 & n25041 ) | ( n5037 & n25041 ) ;
  assign n30470 = n13729 ^ n13377 ^ n285 ;
  assign n30471 = ~n12116 & n20450 ;
  assign n30472 = n12139 ^ n10077 ^ n6498 ;
  assign n30473 = ~n1628 & n13007 ;
  assign n30474 = n13025 ^ n11609 ^ 1'b0 ;
  assign n30475 = n29910 | n30474 ;
  assign n30476 = ~n9377 & n30475 ;
  assign n30477 = n30476 ^ n7580 ^ 1'b0 ;
  assign n30478 = n9823 & ~n18240 ;
  assign n30479 = n30139 ^ n8557 ^ 1'b0 ;
  assign n30480 = n10181 & n23227 ;
  assign n30482 = n4574 & ~n10273 ;
  assign n30483 = n30482 ^ n26624 ^ 1'b0 ;
  assign n30481 = ~n9626 & n25221 ;
  assign n30484 = n30483 ^ n30481 ^ 1'b0 ;
  assign n30485 = ~n20341 & n23806 ;
  assign n30486 = n10108 & n30485 ;
  assign n30487 = n17552 | n22651 ;
  assign n30488 = n18541 ^ n7253 ^ n4219 ;
  assign n30489 = n10122 ^ n6411 ^ 1'b0 ;
  assign n30490 = ( n8359 & n30488 ) | ( n8359 & ~n30489 ) | ( n30488 & ~n30489 ) ;
  assign n30491 = n14324 ^ n5813 ^ 1'b0 ;
  assign n30492 = n15592 | n26125 ;
  assign n30493 = n30492 ^ n11944 ^ 1'b0 ;
  assign n30494 = n25968 ^ n14997 ^ 1'b0 ;
  assign n30495 = ( n1081 & ~n9017 ) | ( n1081 & n29298 ) | ( ~n9017 & n29298 ) ;
  assign n30496 = n6924 & n12369 ;
  assign n30497 = ~n4710 & n30496 ;
  assign n30498 = n7260 & n7807 ;
  assign n30499 = ~n7807 & n30498 ;
  assign n30500 = n2246 | n30499 ;
  assign n30501 = n29462 | n30500 ;
  assign n30502 = n29880 ^ n24311 ^ n9279 ;
  assign n30503 = n6288 & ~n23552 ;
  assign n30504 = ~n20540 & n30503 ;
  assign n30505 = ( n8590 & ~n19347 ) | ( n8590 & n22584 ) | ( ~n19347 & n22584 ) ;
  assign n30506 = n6628 & ~n16234 ;
  assign n30507 = n29638 | n30506 ;
  assign n30508 = n16691 & n25624 ;
  assign n30509 = ~n30507 & n30508 ;
  assign n30510 = n30509 ^ n28839 ^ n5506 ;
  assign n30511 = n14603 ^ n8203 ^ 1'b0 ;
  assign n30515 = n18961 ^ n16217 ^ 1'b0 ;
  assign n30512 = n6531 & ~n10232 ;
  assign n30513 = n5130 & n30512 ;
  assign n30514 = n30513 ^ n25559 ^ n488 ;
  assign n30516 = n30515 ^ n30514 ^ n24841 ;
  assign n30517 = n8420 & ~n15885 ;
  assign n30518 = ~n617 & n29486 ;
  assign n30519 = ~n26994 & n30518 ;
  assign n30520 = n17267 ^ n15535 ^ 1'b0 ;
  assign n30521 = ~n2979 & n30520 ;
  assign n30522 = n24793 ^ n19811 ^ 1'b0 ;
  assign n30523 = n11440 & n26246 ;
  assign n30524 = n2119 | n27937 ;
  assign n30525 = n30524 ^ n1118 ^ 1'b0 ;
  assign n30526 = n25056 & n25538 ;
  assign n30527 = n30526 ^ n25627 ^ 1'b0 ;
  assign n30528 = n22603 & ~n29128 ;
  assign n30529 = n25791 ^ n3279 ^ 1'b0 ;
  assign n30530 = ( n8534 & ~n11777 ) | ( n8534 & n20526 ) | ( ~n11777 & n20526 ) ;
  assign n30531 = ( n3156 & n30529 ) | ( n3156 & ~n30530 ) | ( n30529 & ~n30530 ) ;
  assign n30532 = ( n2946 & ~n16402 ) | ( n2946 & n21573 ) | ( ~n16402 & n21573 ) ;
  assign n30533 = n20349 ^ n2534 ^ 1'b0 ;
  assign n30534 = n2606 & n30533 ;
  assign n30535 = n30534 ^ n3209 ^ 1'b0 ;
  assign n30536 = n14983 ^ n14488 ^ 1'b0 ;
  assign n30537 = ~n628 & n4552 ;
  assign n30538 = ~n8058 & n30537 ;
  assign n30539 = n10938 & ~n30538 ;
  assign n30540 = n29039 ^ n15160 ^ 1'b0 ;
  assign n30541 = n19352 | n30540 ;
  assign n30542 = n609 & n3053 ;
  assign n30543 = n5145 & n10103 ;
  assign n30544 = ~n4631 & n30543 ;
  assign n30545 = n6115 & ~n17621 ;
  assign n30546 = n30545 ^ n15018 ^ 1'b0 ;
  assign n30547 = n28304 & ~n30546 ;
  assign n30548 = n3847 & ~n7173 ;
  assign n30549 = n6360 & ~n22245 ;
  assign n30550 = n22735 ^ n33 ^ 1'b0 ;
  assign n30551 = ~n19060 & n30550 ;
  assign n30552 = ~n3035 & n6511 ;
  assign n30553 = ( n8253 & ~n9538 ) | ( n8253 & n30552 ) | ( ~n9538 & n30552 ) ;
  assign n30554 = ~n15418 & n30553 ;
  assign n30555 = ~n15021 & n30554 ;
  assign n30556 = ( n5732 & n26448 ) | ( n5732 & ~n30555 ) | ( n26448 & ~n30555 ) ;
  assign n30557 = n22879 ^ n5888 ^ 1'b0 ;
  assign n30558 = n3044 & ~n18849 ;
  assign n30559 = n30558 ^ n19969 ^ 1'b0 ;
  assign n30560 = n23548 & ~n30559 ;
  assign n30561 = n10051 ^ n7438 ^ 1'b0 ;
  assign n30562 = n30560 & n30561 ;
  assign n30563 = n6052 & ~n16917 ;
  assign n30564 = n9420 | n30563 ;
  assign n30565 = n21052 ^ x3 ^ 1'b0 ;
  assign n30566 = n9989 ^ n8025 ^ 1'b0 ;
  assign n30567 = n1767 & ~n30566 ;
  assign n30568 = n13093 ^ n1063 ^ 1'b0 ;
  assign n30569 = ~n3738 & n30568 ;
  assign n30570 = ~n27133 & n30569 ;
  assign n30571 = n18565 & n24283 ;
  assign n30572 = ~n13162 & n30571 ;
  assign n30573 = n13811 ^ n7450 ^ 1'b0 ;
  assign n30574 = n14459 & n30573 ;
  assign n30575 = n30574 ^ n436 ^ 1'b0 ;
  assign n30576 = n27613 ^ n8630 ^ 1'b0 ;
  assign n30577 = n4980 | n5892 ;
  assign n30578 = n2995 | n30577 ;
  assign n30579 = n18174 ^ n6539 ^ 1'b0 ;
  assign n30580 = n11453 | n30579 ;
  assign n30581 = n30580 ^ n15761 ^ 1'b0 ;
  assign n30582 = n30581 ^ n16858 ^ 1'b0 ;
  assign n30583 = n15323 & ~n28600 ;
  assign n30585 = n7364 ^ n712 ^ 1'b0 ;
  assign n30586 = n7154 | n30585 ;
  assign n30584 = n1569 & ~n18052 ;
  assign n30587 = n30586 ^ n30584 ^ 1'b0 ;
  assign n30588 = ~n13550 & n20650 ;
  assign n30589 = ~n26518 & n30588 ;
  assign n30590 = n1547 & ~n30589 ;
  assign n30591 = n14864 | n30590 ;
  assign n30592 = n8800 & ~n22158 ;
  assign n30593 = n30592 ^ n22996 ^ 1'b0 ;
  assign n30594 = n30593 ^ n1893 ^ 1'b0 ;
  assign n30595 = n4271 ^ n493 ^ 1'b0 ;
  assign n30596 = n2816 & ~n12722 ;
  assign n30597 = n30596 ^ n29189 ^ 1'b0 ;
  assign n30598 = n1826 & n28737 ;
  assign n30599 = n29339 ^ n7867 ^ 1'b0 ;
  assign n30600 = ~n3430 & n30599 ;
  assign n30601 = n2074 ^ n2032 ^ 1'b0 ;
  assign n30602 = ~n5987 & n30601 ;
  assign n30603 = n1846 & ~n30602 ;
  assign n30604 = n30603 ^ n1666 ^ 1'b0 ;
  assign n30605 = n5402 & n30604 ;
  assign n30606 = n23780 & n24502 ;
  assign n30607 = n10708 | n11760 ;
  assign n30608 = n16070 & ~n30607 ;
  assign n30609 = n9716 & ~n30608 ;
  assign n30610 = ~n4316 & n30609 ;
  assign n30611 = ~n8869 & n30610 ;
  assign n30612 = ( n12159 & n26261 ) | ( n12159 & ~n30611 ) | ( n26261 & ~n30611 ) ;
  assign n30613 = n2485 | n9713 ;
  assign n30614 = n30613 ^ n6234 ^ 1'b0 ;
  assign n30615 = n13199 | n30614 ;
  assign n30616 = n11283 | n30615 ;
  assign n30617 = n10962 & n30616 ;
  assign n30618 = n3246 | n30617 ;
  assign n30619 = n6266 & n28790 ;
  assign n30620 = n30619 ^ n3542 ^ 1'b0 ;
  assign n30621 = n10832 ^ n349 ^ 1'b0 ;
  assign n30622 = n2716 & ~n30621 ;
  assign n30623 = ~n30620 & n30622 ;
  assign n30624 = n21654 ^ n852 ^ 1'b0 ;
  assign n30625 = n13202 & ~n30624 ;
  assign n30626 = n7071 ^ n1287 ^ 1'b0 ;
  assign n30627 = n23497 ^ n17663 ^ 1'b0 ;
  assign n30628 = n30626 | n30627 ;
  assign n30629 = n30628 ^ n16169 ^ n8720 ;
  assign n30631 = ( n3002 & n11893 ) | ( n3002 & ~n20343 ) | ( n11893 & ~n20343 ) ;
  assign n30630 = n3711 | n27403 ;
  assign n30632 = n30631 ^ n30630 ^ 1'b0 ;
  assign n30636 = n108 & n8096 ;
  assign n30633 = n2214 & ~n19509 ;
  assign n30634 = n6808 & n30633 ;
  assign n30635 = n21296 | n30634 ;
  assign n30637 = n30636 ^ n30635 ^ 1'b0 ;
  assign n30654 = ~n811 & n2327 ;
  assign n30655 = n811 & n30654 ;
  assign n30656 = n30655 ^ n2992 ^ 1'b0 ;
  assign n30638 = n10885 ^ n8840 ^ n7097 ;
  assign n30639 = n684 | n23245 ;
  assign n30640 = n23245 & ~n30639 ;
  assign n30641 = n30638 | n30640 ;
  assign n30642 = n30638 & ~n30641 ;
  assign n30643 = n23113 | n30642 ;
  assign n30644 = ~n156 & n1296 ;
  assign n30645 = n156 & n30644 ;
  assign n30646 = ~n923 & n30645 ;
  assign n30647 = n3638 & ~n30646 ;
  assign n30648 = ~n3638 & n30647 ;
  assign n30649 = n3187 & n6286 ;
  assign n30650 = ~n3187 & n30649 ;
  assign n30651 = n30648 | n30650 ;
  assign n30652 = n1977 | n30651 ;
  assign n30653 = n30643 & n30652 ;
  assign n30657 = n30656 ^ n30653 ^ 1'b0 ;
  assign n30658 = n985 ^ n154 ^ 1'b0 ;
  assign n30659 = n30657 & n30658 ;
  assign n30676 = n22185 ^ n3998 ^ 1'b0 ;
  assign n30661 = n3818 & n5562 ;
  assign n30662 = n30661 ^ n9084 ^ 1'b0 ;
  assign n30663 = ~n8289 & n30662 ;
  assign n30664 = n14093 & n30663 ;
  assign n30660 = n7400 | n9778 ;
  assign n30665 = n30664 ^ n30660 ^ 1'b0 ;
  assign n30666 = ~n1287 & n12812 ;
  assign n30667 = n30666 ^ n1010 ^ 1'b0 ;
  assign n30668 = ~n5551 & n30667 ;
  assign n30669 = n30668 ^ n14593 ^ 1'b0 ;
  assign n30670 = n5770 ^ n4543 ^ 1'b0 ;
  assign n30671 = n30669 | n30670 ;
  assign n30672 = n30665 | n30671 ;
  assign n30673 = n11298 & ~n30672 ;
  assign n30674 = n4072 & ~n30673 ;
  assign n30675 = ~n22526 & n30674 ;
  assign n30677 = n30676 ^ n30675 ^ 1'b0 ;
  assign n30678 = n16038 | n27142 ;
  assign n30679 = n26159 | n30678 ;
  assign n30680 = n6712 ^ n3004 ^ 1'b0 ;
  assign n30681 = ( n13230 & n23258 ) | ( n13230 & ~n30680 ) | ( n23258 & ~n30680 ) ;
  assign n30682 = n30681 ^ n12663 ^ 1'b0 ;
  assign n30683 = ( n25064 & ~n30679 ) | ( n25064 & n30682 ) | ( ~n30679 & n30682 ) ;
  assign n30684 = n22605 ^ n1894 ^ 1'b0 ;
  assign n30685 = n1168 & n11137 ;
  assign n30686 = n28543 & ~n30685 ;
  assign n30687 = n5098 | n7408 ;
  assign n30688 = n30687 ^ n22346 ^ 1'b0 ;
  assign n30689 = n1791 & ~n13708 ;
  assign n30690 = n30689 ^ n2194 ^ 1'b0 ;
  assign n30691 = n11307 | n15252 ;
  assign n30692 = n15252 & ~n30691 ;
  assign n30693 = n5589 & ~n30692 ;
  assign n30694 = n5713 & n30693 ;
  assign n30695 = n20526 ^ n3577 ^ 1'b0 ;
  assign n30696 = n4997 ^ n2449 ^ 1'b0 ;
  assign n30697 = ~n9788 & n15589 ;
  assign n30698 = n5822 & n26227 ;
  assign n30699 = n5545 & n30698 ;
  assign n30700 = n21713 ^ n10593 ^ 1'b0 ;
  assign n30701 = ( n3461 & n4723 ) | ( n3461 & ~n30700 ) | ( n4723 & ~n30700 ) ;
  assign n30702 = n22261 ^ n16590 ^ n3957 ;
  assign n30703 = n30702 ^ n35 ^ 1'b0 ;
  assign n30704 = ~n16583 & n22383 ;
  assign n30705 = n2743 & ~n8318 ;
  assign n30706 = n30705 ^ n22564 ^ 1'b0 ;
  assign n30707 = ( n3877 & ~n7021 ) | ( n3877 & n17287 ) | ( ~n7021 & n17287 ) ;
  assign n30708 = n6521 & ~n30707 ;
  assign n30709 = n30706 & n30708 ;
  assign n30710 = ~n4009 & n6375 ;
  assign n30711 = n30710 ^ n11483 ^ 1'b0 ;
  assign n30712 = n3985 ^ n2223 ^ 1'b0 ;
  assign n30713 = n1384 & ~n21176 ;
  assign n30714 = n30712 & n30713 ;
  assign n30715 = n23214 ^ n12002 ^ 1'b0 ;
  assign n30716 = ~n30714 & n30715 ;
  assign n30717 = n8350 ^ n3203 ^ 1'b0 ;
  assign n30718 = ~n4502 & n30717 ;
  assign n30719 = n30718 ^ n8173 ^ 1'b0 ;
  assign n30720 = n21271 & n30719 ;
  assign n30721 = ( n141 & n15016 ) | ( n141 & ~n22918 ) | ( n15016 & ~n22918 ) ;
  assign n30722 = n16700 ^ n8168 ^ 1'b0 ;
  assign n30723 = n11418 ^ n10333 ^ n2636 ;
  assign n30724 = n16670 & ~n30723 ;
  assign n30725 = ~n8427 & n30724 ;
  assign n30726 = ~n4977 & n30725 ;
  assign n30727 = n13509 & n14052 ;
  assign n30728 = n30727 ^ n9161 ^ 1'b0 ;
  assign n30729 = ~n68 & n30728 ;
  assign n30730 = n4142 & ~n30729 ;
  assign n30731 = n30730 ^ n18963 ^ 1'b0 ;
  assign n30732 = ~n4320 & n18841 ;
  assign n30733 = ~n6231 & n30732 ;
  assign n30734 = ~n6987 & n9516 ;
  assign n30735 = n2726 & n30734 ;
  assign n30736 = ~n1630 & n3531 ;
  assign n30737 = ~n3531 & n30736 ;
  assign n30738 = ~n25315 & n30737 ;
  assign n30739 = n7762 & n14706 ;
  assign n30740 = n30738 & n30739 ;
  assign n30741 = ( ~n29153 & n30735 ) | ( ~n29153 & n30740 ) | ( n30735 & n30740 ) ;
  assign n30742 = n6107 | n20112 ;
  assign n30743 = n10105 | n30742 ;
  assign n30744 = n2546 | n30743 ;
  assign n30745 = ( ~n89 & n4804 ) | ( ~n89 & n7719 ) | ( n4804 & n7719 ) ;
  assign n30746 = n30745 ^ n962 ^ 1'b0 ;
  assign n30747 = n30746 ^ n20264 ^ 1'b0 ;
  assign n30749 = n10779 & ~n30727 ;
  assign n30748 = n8731 & ~n9594 ;
  assign n30750 = n30749 ^ n30748 ^ 1'b0 ;
  assign n30751 = n15345 & ~n16301 ;
  assign n30754 = ( n2447 & n13740 ) | ( n2447 & n26489 ) | ( n13740 & n26489 ) ;
  assign n30753 = n6069 | n23308 ;
  assign n30752 = n11893 ^ n8015 ^ 1'b0 ;
  assign n30755 = n30754 ^ n30753 ^ n30752 ;
  assign n30756 = n2619 & ~n25222 ;
  assign n30757 = n30756 ^ n5459 ^ 1'b0 ;
  assign n30758 = ( n11908 & ~n12213 ) | ( n11908 & n23742 ) | ( ~n12213 & n23742 ) ;
  assign n30759 = n26434 | n30758 ;
  assign n30760 = n30759 ^ n13810 ^ 1'b0 ;
  assign n30761 = n30760 ^ n18299 ^ 1'b0 ;
  assign n30762 = n2350 | n30761 ;
  assign n30763 = n13283 | n17932 ;
  assign n30764 = n30763 ^ n6666 ^ 1'b0 ;
  assign n30765 = ~n4686 & n30764 ;
  assign n30766 = n9959 ^ n3603 ^ 1'b0 ;
  assign n30767 = n6042 | n30766 ;
  assign n30768 = ( n1175 & n17233 ) | ( n1175 & ~n30767 ) | ( n17233 & ~n30767 ) ;
  assign n30769 = n17222 | n24118 ;
  assign n30770 = n18107 & ~n30769 ;
  assign n30771 = ~n3833 & n14600 ;
  assign n30772 = n16776 & n30771 ;
  assign n30773 = n30772 ^ n12460 ^ 1'b0 ;
  assign n30774 = ~n15222 & n30773 ;
  assign n30775 = n8754 ^ n976 ^ 1'b0 ;
  assign n30776 = n7654 & n30775 ;
  assign n30777 = n10294 & n30776 ;
  assign n30778 = n1411 & n29652 ;
  assign n30779 = n8811 & n30778 ;
  assign n30780 = n8991 | n12251 ;
  assign n30781 = n30780 ^ n8884 ^ 1'b0 ;
  assign n30782 = n30781 ^ n648 ^ 1'b0 ;
  assign n30783 = n30782 ^ n27490 ^ 1'b0 ;
  assign n30784 = n30036 ^ n6799 ^ n989 ;
  assign n30785 = n22405 & n30784 ;
  assign n30786 = n12301 & n30785 ;
  assign n30787 = n16331 ^ n5898 ^ 1'b0 ;
  assign n30788 = n13812 ^ n12083 ^ 1'b0 ;
  assign n30789 = ~n30787 & n30788 ;
  assign n30790 = ~n14144 & n27860 ;
  assign n30791 = n30790 ^ n21506 ^ 1'b0 ;
  assign n30792 = n6199 & n30791 ;
  assign n30793 = ~n14936 & n16430 ;
  assign n30794 = n30793 ^ n12931 ^ 1'b0 ;
  assign n30795 = ~n18720 & n28209 ;
  assign n30798 = n9543 & ~n14831 ;
  assign n30799 = n10384 ^ n723 ^ 1'b0 ;
  assign n30800 = n8490 | n30799 ;
  assign n30801 = n30798 & ~n30800 ;
  assign n30796 = n13947 | n16549 ;
  assign n30797 = n21206 & n30796 ;
  assign n30802 = n30801 ^ n30797 ^ 1'b0 ;
  assign n30803 = ~n26392 & n30802 ;
  assign n30804 = n4674 & n30803 ;
  assign n30805 = n15712 ^ n13984 ^ 1'b0 ;
  assign n30806 = n30805 ^ n29830 ^ 1'b0 ;
  assign n30807 = n30806 ^ n13695 ^ n5764 ;
  assign n30808 = n21337 & ~n30807 ;
  assign n30809 = n7091 ^ n6380 ^ 1'b0 ;
  assign n30810 = ~n16168 & n18929 ;
  assign n30811 = ( n20411 & ~n30809 ) | ( n20411 & n30810 ) | ( ~n30809 & n30810 ) ;
  assign n30812 = ~n14580 & n24121 ;
  assign n30813 = n30812 ^ n8547 ^ 1'b0 ;
  assign n30814 = ~n15588 & n30813 ;
  assign n30815 = n3918 & ~n29766 ;
  assign n30816 = ~n1151 & n30815 ;
  assign n30818 = n7495 & ~n29774 ;
  assign n30817 = n500 | n11922 ;
  assign n30819 = n30818 ^ n30817 ^ 1'b0 ;
  assign n30820 = n6477 & n17432 ;
  assign n30821 = ~n4201 & n12663 ;
  assign n30822 = n4201 & n30821 ;
  assign n30823 = n2977 & ~n6597 ;
  assign n30824 = ~n2977 & n30823 ;
  assign n30825 = n7707 & n30824 ;
  assign n30826 = n23537 | n30825 ;
  assign n30827 = n30822 | n30826 ;
  assign n30828 = n28773 ^ n3135 ^ 1'b0 ;
  assign n30829 = ~n30827 & n30828 ;
  assign n30830 = ~n10123 & n30829 ;
  assign n30832 = n9021 & ~n25614 ;
  assign n30833 = ~n2082 & n30832 ;
  assign n30834 = n30833 ^ n27385 ^ 1'b0 ;
  assign n30831 = n2702 & ~n8588 ;
  assign n30835 = n30834 ^ n30831 ^ 1'b0 ;
  assign n30836 = ( n4447 & n6383 ) | ( n4447 & n6437 ) | ( n6383 & n6437 ) ;
  assign n30837 = n30836 ^ n8967 ^ 1'b0 ;
  assign n30838 = n26883 | n30837 ;
  assign n30839 = n7233 ^ n1655 ^ 1'b0 ;
  assign n30841 = n26400 ^ n16278 ^ 1'b0 ;
  assign n30842 = n7724 & ~n30841 ;
  assign n30840 = n1118 & n24751 ;
  assign n30843 = n30842 ^ n30840 ^ 1'b0 ;
  assign n30844 = n28872 ^ n23838 ^ 1'b0 ;
  assign n30845 = n8953 & n10113 ;
  assign n30846 = n30845 ^ n6202 ^ 1'b0 ;
  assign n30847 = n10235 & ~n12155 ;
  assign n30848 = n30846 | n30847 ;
  assign n30849 = n26715 ^ n15251 ^ 1'b0 ;
  assign n30850 = ( n6727 & n27417 ) | ( n6727 & ~n30849 ) | ( n27417 & ~n30849 ) ;
  assign n30851 = n17153 ^ n11088 ^ 1'b0 ;
  assign n30852 = n30851 ^ n18556 ^ n10318 ;
  assign n30853 = n28255 & n30852 ;
  assign n30854 = n18649 & n20136 ;
  assign n30855 = n30854 ^ n21495 ^ 1'b0 ;
  assign n30856 = n25283 ^ n2773 ^ n923 ;
  assign n30857 = n8827 & n30856 ;
  assign n30858 = n30857 ^ n838 ^ 1'b0 ;
  assign n30859 = n30858 ^ n23665 ^ n22134 ;
  assign n30860 = ( n126 & n13363 ) | ( n126 & ~n13904 ) | ( n13363 & ~n13904 ) ;
  assign n30861 = n125 | n30860 ;
  assign n30862 = n30861 ^ n1964 ^ 1'b0 ;
  assign n30863 = n30862 ^ n24465 ^ n7915 ;
  assign n30864 = n30863 ^ n7238 ^ 1'b0 ;
  assign n30865 = n17487 & n30864 ;
  assign n30866 = ~n1170 & n14164 ;
  assign n30867 = n8008 | n30866 ;
  assign n30868 = n14227 & n30867 ;
  assign n30869 = n16650 ^ n10555 ^ n1220 ;
  assign n30870 = n9588 & ~n14709 ;
  assign n30871 = n30870 ^ n22706 ^ n21647 ;
  assign n30872 = n260 | n22488 ;
  assign n30873 = n30872 ^ n18600 ^ 1'b0 ;
  assign n30874 = n6383 & n6846 ;
  assign n30875 = n28511 & n30874 ;
  assign n30876 = n19529 ^ n16302 ^ 1'b0 ;
  assign n30877 = ~n11854 & n30876 ;
  assign n30878 = ~n2045 & n30877 ;
  assign n30879 = n8337 & ~n30461 ;
  assign n30880 = n27623 ^ n18601 ^ 1'b0 ;
  assign n30881 = n1612 ^ n1489 ^ 1'b0 ;
  assign n30882 = ( n13018 & ~n13653 ) | ( n13018 & n30881 ) | ( ~n13653 & n30881 ) ;
  assign n30883 = n30882 ^ n14365 ^ 1'b0 ;
  assign n30884 = n24737 & n30883 ;
  assign n30885 = n1579 & ~n4620 ;
  assign n30886 = n17220 & n30885 ;
  assign n30887 = n30886 ^ n13111 ^ 1'b0 ;
  assign n30888 = n30887 ^ n24742 ^ n20685 ;
  assign n30889 = n7516 & ~n30888 ;
  assign n30890 = n30889 ^ n28895 ^ 1'b0 ;
  assign n30891 = n8008 ^ n987 ^ 1'b0 ;
  assign n30892 = n30891 ^ n1909 ^ n1525 ;
  assign n30893 = n11608 ^ n8010 ^ 1'b0 ;
  assign n30894 = n3985 & ~n30893 ;
  assign n30895 = ( n4587 & n8820 ) | ( n4587 & ~n30894 ) | ( n8820 & ~n30894 ) ;
  assign n30896 = n12815 & ~n30895 ;
  assign n30897 = n536 | n21474 ;
  assign n30898 = n30897 ^ n8463 ^ 1'b0 ;
  assign n30899 = n3634 & n12857 ;
  assign n30900 = n30898 & n30899 ;
  assign n30901 = n3648 & n7490 ;
  assign n30902 = n30901 ^ n4252 ^ 1'b0 ;
  assign n30903 = n19373 | n30902 ;
  assign n30904 = n19007 ^ n15767 ^ 1'b0 ;
  assign n30905 = n14709 ^ n10741 ^ n6877 ;
  assign n30906 = n30905 ^ n1043 ^ 1'b0 ;
  assign n30907 = n15776 & ~n30906 ;
  assign n30908 = n28798 | n30907 ;
  assign n30909 = n30908 ^ n11091 ^ 1'b0 ;
  assign n30910 = ~n30904 & n30909 ;
  assign n30911 = n24348 ^ n6497 ^ 1'b0 ;
  assign n30912 = n22206 ^ n2259 ^ 1'b0 ;
  assign n30913 = n30912 ^ n29772 ^ n13823 ;
  assign n30914 = n14981 ^ n2995 ^ 1'b0 ;
  assign n30915 = n728 & ~n30914 ;
  assign n30916 = n18745 ^ n2134 ^ 1'b0 ;
  assign n30917 = n24846 & n30916 ;
  assign n30918 = n16038 & n25363 ;
  assign n30919 = n10391 & ~n30918 ;
  assign n30920 = n30919 ^ n20984 ^ 1'b0 ;
  assign n30921 = ~n5044 & n18148 ;
  assign n30922 = n30921 ^ n30415 ^ 1'b0 ;
  assign n30923 = ~n13752 & n30922 ;
  assign n30924 = n7228 ^ n362 ^ 1'b0 ;
  assign n30925 = n30924 ^ n7839 ^ 1'b0 ;
  assign n30926 = n27049 & n30925 ;
  assign n30927 = n3626 & n12119 ;
  assign n30928 = n12540 & n30927 ;
  assign n30929 = n20277 & n30928 ;
  assign n30930 = n11880 ^ n3483 ^ 1'b0 ;
  assign n30931 = n4331 & ~n30930 ;
  assign n30932 = n7092 & ~n20836 ;
  assign n30933 = n16441 | n20705 ;
  assign n30934 = ~n6601 & n14524 ;
  assign n30935 = n8489 ^ n8130 ^ 1'b0 ;
  assign n30936 = ~n30934 & n30935 ;
  assign n30937 = n30936 ^ n19826 ^ 1'b0 ;
  assign n30938 = n6098 | n11892 ;
  assign n30939 = n25254 ^ n6152 ^ 1'b0 ;
  assign n30940 = n3510 & n30939 ;
  assign n30944 = n6821 | n11171 ;
  assign n30941 = n16641 | n17520 ;
  assign n30942 = n9110 ^ n3877 ^ 1'b0 ;
  assign n30943 = n30941 & n30942 ;
  assign n30945 = n30944 ^ n30943 ^ 1'b0 ;
  assign n30946 = n30940 & ~n30945 ;
  assign n30947 = n22631 & n30569 ;
  assign n30948 = n24456 & n30947 ;
  assign n30949 = n4231 & n16622 ;
  assign n30950 = n1709 & n30949 ;
  assign n30951 = n30948 | n30950 ;
  assign n30952 = n30951 ^ n4243 ^ 1'b0 ;
  assign n30953 = n13274 ^ n4923 ^ 1'b0 ;
  assign n30954 = n30953 ^ n30235 ^ 1'b0 ;
  assign n30955 = n2746 & n10498 ;
  assign n30956 = ~n1751 & n30955 ;
  assign n30957 = n13023 | n26266 ;
  assign n30958 = ~n5709 & n30957 ;
  assign n30960 = n887 & n16858 ;
  assign n30959 = n1549 & n10648 ;
  assign n30961 = n30960 ^ n30959 ^ 1'b0 ;
  assign n30962 = ~n9199 & n25479 ;
  assign n30963 = ~n5130 & n30962 ;
  assign n30964 = ( n6305 & n15060 ) | ( n6305 & ~n25337 ) | ( n15060 & ~n25337 ) ;
  assign n30965 = n9128 ^ n3691 ^ 1'b0 ;
  assign n30966 = n2882 & ~n30965 ;
  assign n30967 = n7279 ^ n483 ^ 1'b0 ;
  assign n30968 = n14148 & n30967 ;
  assign n30969 = n30966 & n30968 ;
  assign n30970 = n21363 ^ n3856 ^ 1'b0 ;
  assign n30971 = ~n7295 & n30970 ;
  assign n30972 = ~n20950 & n30971 ;
  assign n30973 = n4468 | n30972 ;
  assign n30974 = n9889 | n30973 ;
  assign n30975 = n17865 & n30974 ;
  assign n30976 = ~n14279 & n17923 ;
  assign n30977 = ( n1542 & n23183 ) | ( n1542 & ~n27586 ) | ( n23183 & ~n27586 ) ;
  assign n30978 = n23067 ^ n22503 ^ 1'b0 ;
  assign n30979 = n4590 & n7600 ;
  assign n30980 = n8182 & ~n30979 ;
  assign n30981 = n30980 ^ n12499 ^ 1'b0 ;
  assign n30983 = n2482 | n12975 ;
  assign n30982 = n2898 | n8794 ;
  assign n30984 = n30983 ^ n30982 ^ 1'b0 ;
  assign n30985 = n28486 ^ n11969 ^ 1'b0 ;
  assign n30986 = n7945 | n30985 ;
  assign n30987 = n30986 ^ n29467 ^ 1'b0 ;
  assign n30990 = n10830 ^ n8395 ^ 1'b0 ;
  assign n30991 = n20129 & n30990 ;
  assign n30992 = n4427 & ~n30991 ;
  assign n30988 = n12196 ^ n6180 ^ 1'b0 ;
  assign n30989 = n3833 | n30988 ;
  assign n30993 = n30992 ^ n30989 ^ 1'b0 ;
  assign n30994 = n17993 | n30993 ;
  assign n30995 = n10951 ^ n4072 ^ 1'b0 ;
  assign n30996 = ( n3939 & n6010 ) | ( n3939 & n11626 ) | ( n6010 & n11626 ) ;
  assign n30997 = ( ~n2381 & n12053 ) | ( ~n2381 & n30996 ) | ( n12053 & n30996 ) ;
  assign n30998 = n30997 ^ n9823 ^ 1'b0 ;
  assign n30999 = n2622 | n19102 ;
  assign n31000 = n3625 & ~n30999 ;
  assign n31001 = n14915 | n16142 ;
  assign n31002 = ( n2156 & ~n5091 ) | ( n2156 & n31001 ) | ( ~n5091 & n31001 ) ;
  assign n31003 = ( ~n11077 & n11786 ) | ( ~n11077 & n31002 ) | ( n11786 & n31002 ) ;
  assign n31004 = ( ~n2499 & n31000 ) | ( ~n2499 & n31003 ) | ( n31000 & n31003 ) ;
  assign n31005 = n8648 ^ n4804 ^ n2436 ;
  assign n31006 = n23556 ^ n1489 ^ 1'b0 ;
  assign n31007 = n31005 & ~n31006 ;
  assign n31008 = ~n12306 & n31007 ;
  assign n31009 = n16023 | n31008 ;
  assign n31010 = n20910 ^ n3603 ^ 1'b0 ;
  assign n31011 = ( ~n169 & n3968 ) | ( ~n169 & n5675 ) | ( n3968 & n5675 ) ;
  assign n31012 = n31010 | n31011 ;
  assign n31013 = n260 | n19018 ;
  assign n31014 = n31013 ^ n22786 ^ 1'b0 ;
  assign n31015 = n20545 & n25365 ;
  assign n31016 = n15025 | n31015 ;
  assign n31017 = n16256 & ~n31016 ;
  assign n31018 = ( n5781 & n6558 ) | ( n5781 & ~n21013 ) | ( n6558 & ~n21013 ) ;
  assign n31019 = n3341 ^ n3170 ^ 1'b0 ;
  assign n31020 = n6100 & n31019 ;
  assign n31021 = n1532 | n31020 ;
  assign n31022 = ( ~n8265 & n14491 ) | ( ~n8265 & n31021 ) | ( n14491 & n31021 ) ;
  assign n31023 = n1848 & ~n19925 ;
  assign n31024 = n10639 & n31023 ;
  assign n31025 = n31024 ^ n4371 ^ 1'b0 ;
  assign n31026 = n8615 & n31025 ;
  assign n31027 = ~n18899 & n31026 ;
  assign n31028 = ~n31022 & n31027 ;
  assign n31029 = n7488 & n7746 ;
  assign n31030 = ~n8508 & n31029 ;
  assign n31031 = n7641 & ~n31030 ;
  assign n31032 = n29225 ^ n12103 ^ 1'b0 ;
  assign n31033 = n31031 & ~n31032 ;
  assign n31034 = ~n23522 & n24097 ;
  assign n31035 = n12904 ^ n9081 ^ 1'b0 ;
  assign n31036 = n6069 & ~n23168 ;
  assign n31037 = n31036 ^ n19420 ^ 1'b0 ;
  assign n31038 = n31035 & ~n31037 ;
  assign n31039 = n4391 ^ n3626 ^ 1'b0 ;
  assign n31040 = ( n11227 & n19212 ) | ( n11227 & ~n31039 ) | ( n19212 & ~n31039 ) ;
  assign n31041 = n8451 | n17018 ;
  assign n31042 = n12974 & ~n31041 ;
  assign n31043 = n10952 | n12772 ;
  assign n31044 = n20002 | n24093 ;
  assign n31045 = ~n9939 & n31044 ;
  assign n31046 = ( ~n1760 & n2535 ) | ( ~n1760 & n14364 ) | ( n2535 & n14364 ) ;
  assign n31047 = n2281 & n11424 ;
  assign n31048 = n28664 & ~n31047 ;
  assign n31049 = ( n15210 & ~n31046 ) | ( n15210 & n31048 ) | ( ~n31046 & n31048 ) ;
  assign n31050 = n166 & n7860 ;
  assign n31051 = n17324 & n31050 ;
  assign n31052 = ~n774 & n9443 ;
  assign n31053 = n31052 ^ n3655 ^ 1'b0 ;
  assign n31054 = n8303 | n31053 ;
  assign n31055 = n28297 ^ n17520 ^ 1'b0 ;
  assign n31056 = ~n12995 & n31055 ;
  assign n31057 = n5632 & ~n20727 ;
  assign n31058 = n7319 & n31057 ;
  assign n31059 = ( n24044 & ~n26409 ) | ( n24044 & n31058 ) | ( ~n26409 & n31058 ) ;
  assign n31060 = n3699 ^ n1285 ^ 1'b0 ;
  assign n31061 = n7696 & n31060 ;
  assign n31062 = n21019 ^ n3609 ^ 1'b0 ;
  assign n31063 = n31061 & ~n31062 ;
  assign n31064 = n31063 ^ n22747 ^ 1'b0 ;
  assign n31065 = ~n10591 & n28543 ;
  assign n31066 = n19597 & ~n20199 ;
  assign n31067 = ~n17201 & n31066 ;
  assign n31068 = n1660 ^ n1296 ^ 1'b0 ;
  assign n31069 = n3120 & n31068 ;
  assign n31070 = n1367 ^ n245 ^ 1'b0 ;
  assign n31071 = n31070 ^ n11410 ^ 1'b0 ;
  assign n31072 = n31071 ^ n23065 ^ 1'b0 ;
  assign n31073 = n8711 | n31072 ;
  assign n31074 = n685 | n4227 ;
  assign n31075 = n31074 ^ n20805 ^ n9509 ;
  assign n31079 = n7249 ^ n6082 ^ 1'b0 ;
  assign n31080 = n7286 | n31079 ;
  assign n31076 = ~n5617 & n9193 ;
  assign n31077 = n31076 ^ n22588 ^ 1'b0 ;
  assign n31078 = n5632 & n31077 ;
  assign n31081 = n31080 ^ n31078 ^ 1'b0 ;
  assign n31082 = ~n17438 & n20686 ;
  assign n31083 = n31082 ^ n15114 ^ 1'b0 ;
  assign n31089 = n16850 & ~n18221 ;
  assign n31090 = n31089 ^ n7103 ^ 1'b0 ;
  assign n31084 = n2213 & n7612 ;
  assign n31085 = n8054 | n31084 ;
  assign n31086 = n31085 ^ n15030 ^ n3908 ;
  assign n31087 = ~n8517 & n24467 ;
  assign n31088 = n31086 & n31087 ;
  assign n31091 = n31090 ^ n31088 ^ 1'b0 ;
  assign n31092 = n24834 ^ n5535 ^ 1'b0 ;
  assign n31093 = n31092 ^ n2889 ^ 1'b0 ;
  assign n31094 = n22638 & ~n31093 ;
  assign n31095 = ( ~n24621 & n27899 ) | ( ~n24621 & n31094 ) | ( n27899 & n31094 ) ;
  assign n31096 = n5102 ^ n5039 ^ n4156 ;
  assign n31097 = n4502 ^ n3645 ^ 1'b0 ;
  assign n31098 = n6656 & ~n31097 ;
  assign n31099 = n31096 & n31098 ;
  assign n31100 = n31099 ^ n14392 ^ 1'b0 ;
  assign n31101 = n29894 | n31100 ;
  assign n31102 = ~n13684 & n21394 ;
  assign n31103 = ~n2434 & n31102 ;
  assign n31104 = ~n8871 & n31103 ;
  assign n31105 = n15251 ^ n10164 ^ 1'b0 ;
  assign n31106 = ( n2234 & ~n28087 ) | ( n2234 & n31105 ) | ( ~n28087 & n31105 ) ;
  assign n31107 = n6630 & n21323 ;
  assign n31108 = n3512 | n15849 ;
  assign n31109 = n5029 & ~n31108 ;
  assign n31110 = n13987 & ~n31109 ;
  assign n31111 = n2405 & ~n13919 ;
  assign n31112 = ~n8799 & n31111 ;
  assign n31113 = n19165 ^ n9110 ^ n6804 ;
  assign n31114 = n31113 ^ n11727 ^ 1'b0 ;
  assign n31115 = n31114 ^ n16827 ^ 1'b0 ;
  assign n31116 = n28550 & n31115 ;
  assign n31117 = n31116 ^ n14508 ^ 1'b0 ;
  assign n31118 = n8086 & ~n10292 ;
  assign n31119 = n5191 & ~n21564 ;
  assign n31120 = n25239 & n31119 ;
  assign n31121 = ~n11295 & n11988 ;
  assign n31122 = ( n15079 & n21443 ) | ( n15079 & n31121 ) | ( n21443 & n31121 ) ;
  assign n31123 = ( n21982 & n22038 ) | ( n21982 & n25483 ) | ( n22038 & n25483 ) ;
  assign n31125 = n4183 & n13598 ;
  assign n31126 = n3797 & n31125 ;
  assign n31124 = n4454 & ~n30246 ;
  assign n31127 = n31126 ^ n31124 ^ 1'b0 ;
  assign n31128 = ( ~n5033 & n14489 ) | ( ~n5033 & n19367 ) | ( n14489 & n19367 ) ;
  assign n31129 = n2616 | n11309 ;
  assign n31130 = n31129 ^ n11753 ^ 1'b0 ;
  assign n31131 = ( n3002 & n27959 ) | ( n3002 & ~n31130 ) | ( n27959 & ~n31130 ) ;
  assign n31132 = n23168 ^ n12936 ^ n2625 ;
  assign n31133 = n6240 | n31132 ;
  assign n31134 = n5262 | n31133 ;
  assign n31135 = n8985 | n18146 ;
  assign n31136 = ~n21755 & n31135 ;
  assign n31137 = n6710 & n12708 ;
  assign n31138 = n31137 ^ n7586 ^ 1'b0 ;
  assign n31139 = n7642 | n12066 ;
  assign n31140 = n15388 | n31139 ;
  assign n31141 = n31140 ^ n28606 ^ 1'b0 ;
  assign n31142 = n10468 & ~n15571 ;
  assign n31143 = n31142 ^ n19292 ^ 1'b0 ;
  assign n31144 = n31143 ^ n645 ^ 1'b0 ;
  assign n31145 = n3465 ^ n329 ^ 1'b0 ;
  assign n31146 = n3575 & n31145 ;
  assign n31147 = ( n15122 & ~n17951 ) | ( n15122 & n31146 ) | ( ~n17951 & n31146 ) ;
  assign n31148 = n10017 ^ n3170 ^ n2884 ;
  assign n31149 = ~n14555 & n31148 ;
  assign n31150 = n31149 ^ n3368 ^ 1'b0 ;
  assign n31151 = n6037 | n31150 ;
  assign n31152 = n9591 | n14275 ;
  assign n31153 = n17331 & ~n31152 ;
  assign n31154 = n22918 & n31153 ;
  assign n31155 = ~n4725 & n4947 ;
  assign n31156 = n31155 ^ n3195 ^ 1'b0 ;
  assign n31157 = n14229 ^ n6885 ^ n5311 ;
  assign n31158 = n10796 | n16521 ;
  assign n31159 = n1525 | n31158 ;
  assign n31160 = ~n16990 & n30057 ;
  assign n31161 = ~n4937 & n15800 ;
  assign n31162 = ~n25045 & n31161 ;
  assign n31163 = n1694 & n4354 ;
  assign n31164 = ~n12307 & n31163 ;
  assign n31165 = n14980 | n31164 ;
  assign n31166 = n7940 ^ n6076 ^ 1'b0 ;
  assign n31167 = n27601 & ~n31166 ;
  assign n31168 = n1416 | n15167 ;
  assign n31169 = ( n2332 & ~n4114 ) | ( n2332 & n12785 ) | ( ~n4114 & n12785 ) ;
  assign n31170 = n17700 | n23188 ;
  assign n31171 = n31170 ^ n3114 ^ 1'b0 ;
  assign n31172 = n31169 | n31171 ;
  assign n31173 = n18297 ^ n8143 ^ 1'b0 ;
  assign n31174 = n3037 | n12435 ;
  assign n31175 = n15769 & ~n31174 ;
  assign n31176 = n31175 ^ n7462 ^ 1'b0 ;
  assign n31177 = n19013 ^ n18843 ^ 1'b0 ;
  assign n31178 = n10414 | n31177 ;
  assign n31179 = n1841 | n10361 ;
  assign n31180 = n31179 ^ n16652 ^ 1'b0 ;
  assign n31181 = n13938 | n31180 ;
  assign n31182 = n25814 & ~n31181 ;
  assign n31183 = ( n3641 & n3666 ) | ( n3641 & n31182 ) | ( n3666 & n31182 ) ;
  assign n31184 = n31183 ^ n20771 ^ n4416 ;
  assign n31185 = n15228 & ~n21948 ;
  assign n31186 = ~n20593 & n31185 ;
  assign n31187 = n22776 ^ n9764 ^ n3466 ;
  assign n31188 = n31187 ^ n14485 ^ 1'b0 ;
  assign n31189 = n8759 ^ n4283 ^ 1'b0 ;
  assign n31190 = n2190 & n6477 ;
  assign n31191 = n26168 ^ n21529 ^ n13289 ;
  assign n31192 = n3387 ^ n332 ^ 1'b0 ;
  assign n31193 = ~n9341 & n31192 ;
  assign n31194 = ( n4200 & n9465 ) | ( n4200 & n15775 ) | ( n9465 & n15775 ) ;
  assign n31195 = ~n15976 & n31194 ;
  assign n31197 = ( ~n15461 & n17961 ) | ( ~n15461 & n27576 ) | ( n17961 & n27576 ) ;
  assign n31196 = n4659 | n29413 ;
  assign n31198 = n31197 ^ n31196 ^ 1'b0 ;
  assign n31199 = n6551 & ~n9034 ;
  assign n31200 = n19675 | n31199 ;
  assign n31201 = n19317 & n31200 ;
  assign n31202 = n5511 & n31201 ;
  assign n31203 = n12642 & ~n18324 ;
  assign n31204 = n31202 & n31203 ;
  assign n31206 = n1055 & ~n27040 ;
  assign n31205 = ~n5186 & n20711 ;
  assign n31207 = n31206 ^ n31205 ^ 1'b0 ;
  assign n31208 = n13344 ^ n784 ^ 1'b0 ;
  assign n31209 = n11450 & n31208 ;
  assign n31210 = n14071 ^ n2186 ^ n78 ;
  assign n31211 = n18498 ^ n6976 ^ 1'b0 ;
  assign n31212 = ( n13448 & n31210 ) | ( n13448 & ~n31211 ) | ( n31210 & ~n31211 ) ;
  assign n31213 = n20198 ^ n3473 ^ 1'b0 ;
  assign n31214 = n31213 ^ n27631 ^ 1'b0 ;
  assign n31215 = n30078 & n31214 ;
  assign n31216 = n19079 ^ n10418 ^ 1'b0 ;
  assign n31217 = n15706 & ~n31216 ;
  assign n31218 = n9638 ^ n9228 ^ 1'b0 ;
  assign n31219 = ( n1658 & n5564 ) | ( n1658 & n8267 ) | ( n5564 & n8267 ) ;
  assign n31220 = n15199 ^ n5645 ^ 1'b0 ;
  assign n31221 = ( n334 & ~n12742 ) | ( n334 & n31220 ) | ( ~n12742 & n31220 ) ;
  assign n31222 = n10550 ^ n2645 ^ 1'b0 ;
  assign n31223 = ~n17708 & n31222 ;
  assign n31224 = n1198 & ~n9886 ;
  assign n31225 = n24951 ^ n6996 ^ n3818 ;
  assign n31226 = n1104 ^ n922 ^ 1'b0 ;
  assign n31227 = n1368 & n31226 ;
  assign n31228 = n31227 ^ n2090 ^ 1'b0 ;
  assign n31229 = n12837 & ~n31228 ;
  assign n31230 = ~n10376 & n27684 ;
  assign n31231 = n31229 & n31230 ;
  assign n31232 = n21991 & n23143 ;
  assign n31234 = n772 & ~n1642 ;
  assign n31233 = n22334 ^ n20385 ^ 1'b0 ;
  assign n31235 = n31234 ^ n31233 ^ 1'b0 ;
  assign n31236 = ~n5594 & n31235 ;
  assign n31237 = ~n3642 & n29351 ;
  assign n31238 = n14332 ^ n760 ^ n490 ;
  assign n31241 = ~n601 & n26569 ;
  assign n31239 = n10054 ^ n2835 ^ 1'b0 ;
  assign n31240 = n23676 & n31239 ;
  assign n31242 = n31241 ^ n31240 ^ n2810 ;
  assign n31243 = n5781 ^ n4807 ^ n842 ;
  assign n31244 = ( n191 & n6049 ) | ( n191 & ~n29461 ) | ( n6049 & ~n29461 ) ;
  assign n31245 = n31244 ^ n21387 ^ n7621 ;
  assign n31246 = n3532 & ~n31245 ;
  assign n31247 = n31246 ^ n26685 ^ 1'b0 ;
  assign n31248 = n17795 & ~n25436 ;
  assign n31249 = n31248 ^ n22584 ^ 1'b0 ;
  assign n31250 = n31249 ^ n24824 ^ 1'b0 ;
  assign n31251 = ~n20829 & n31250 ;
  assign n31252 = ( ~n1842 & n12335 ) | ( ~n1842 & n13705 ) | ( n12335 & n13705 ) ;
  assign n31253 = n1280 & n26073 ;
  assign n31254 = n18132 ^ n247 ^ 1'b0 ;
  assign n31255 = n30070 & ~n31254 ;
  assign n31256 = n4177 ^ n730 ^ 1'b0 ;
  assign n31257 = n31256 ^ n7324 ^ 1'b0 ;
  assign n31258 = n13400 ^ n8084 ^ n3671 ;
  assign n31259 = ~n24219 & n31258 ;
  assign n31260 = ( n9208 & ~n22662 ) | ( n9208 & n31259 ) | ( ~n22662 & n31259 ) ;
  assign n31261 = n31260 ^ n2397 ^ 1'b0 ;
  assign n31262 = n5638 & ~n7366 ;
  assign n31263 = ~n3704 & n11614 ;
  assign n31264 = n25930 & n31263 ;
  assign n31265 = n31264 ^ n17761 ^ 1'b0 ;
  assign n31266 = ( n39 & n174 ) | ( n39 & n1815 ) | ( n174 & n1815 ) ;
  assign n31267 = n6953 & ~n31266 ;
  assign n31268 = n13860 & n31267 ;
  assign n31269 = n15868 ^ n8519 ^ 1'b0 ;
  assign n31270 = n31268 | n31269 ;
  assign n31271 = n23487 ^ n2885 ^ 1'b0 ;
  assign n31272 = n20299 & ~n31271 ;
  assign n31273 = n31272 ^ n4262 ^ 1'b0 ;
  assign n31274 = ~n10093 & n26026 ;
  assign n31275 = ~n1319 & n10171 ;
  assign n31276 = n31275 ^ n4928 ^ 1'b0 ;
  assign n31277 = ( n27673 & n29471 ) | ( n27673 & ~n31276 ) | ( n29471 & ~n31276 ) ;
  assign n31278 = n6101 | n24482 ;
  assign n31279 = n31278 ^ n1568 ^ 1'b0 ;
  assign n31281 = ( ~n2864 & n13107 ) | ( ~n2864 & n23376 ) | ( n13107 & n23376 ) ;
  assign n31280 = n18174 & ~n25775 ;
  assign n31282 = n31281 ^ n31280 ^ 1'b0 ;
  assign n31283 = n1296 | n1305 ;
  assign n31284 = n4222 | n12241 ;
  assign n31285 = n1177 | n31284 ;
  assign n31286 = n263 & ~n553 ;
  assign n31287 = ~n13778 & n31286 ;
  assign n31288 = ~n31285 & n31287 ;
  assign n31289 = ~n5461 & n15130 ;
  assign n31290 = n7254 | n25318 ;
  assign n31291 = n4086 & ~n31290 ;
  assign n31292 = n31289 | n31291 ;
  assign n31293 = n2702 & ~n14381 ;
  assign n31294 = n24266 ^ n6263 ^ 1'b0 ;
  assign n31295 = ~n21733 & n31294 ;
  assign n31296 = n15466 ^ n7065 ^ 1'b0 ;
  assign n31297 = n26975 | n31296 ;
  assign n31301 = n21057 ^ n12044 ^ 1'b0 ;
  assign n31298 = ~n2207 & n10420 ;
  assign n31299 = n31298 ^ n2569 ^ 1'b0 ;
  assign n31300 = n5339 & n31299 ;
  assign n31302 = n31301 ^ n31300 ^ 1'b0 ;
  assign n31303 = ( n9973 & ~n15228 ) | ( n9973 & n31302 ) | ( ~n15228 & n31302 ) ;
  assign n31304 = n7180 & n13719 ;
  assign n31305 = n31304 ^ n16040 ^ 1'b0 ;
  assign n31306 = ( n13078 & ~n13940 ) | ( n13078 & n31305 ) | ( ~n13940 & n31305 ) ;
  assign n31307 = ( n6111 & n13099 ) | ( n6111 & ~n15388 ) | ( n13099 & ~n15388 ) ;
  assign n31308 = ~n6335 & n31307 ;
  assign n31309 = ~n1142 & n11167 ;
  assign n31310 = n23783 & n31309 ;
  assign n31311 = ( n7106 & n11346 ) | ( n7106 & n30017 ) | ( n11346 & n30017 ) ;
  assign n31312 = n8340 & ~n16644 ;
  assign n31313 = n514 & n31312 ;
  assign n31314 = n31313 ^ n30225 ^ 1'b0 ;
  assign n31315 = n1572 & ~n3534 ;
  assign n31316 = n22940 & ~n31315 ;
  assign n31317 = n31316 ^ n156 ^ 1'b0 ;
  assign n31318 = n31317 ^ n30991 ^ n4160 ;
  assign n31319 = n6027 | n16963 ;
  assign n31320 = n31319 ^ n26149 ^ 1'b0 ;
  assign n31321 = n9483 | n31320 ;
  assign n31322 = n31321 ^ n2570 ^ 1'b0 ;
  assign n31323 = n4457 | n27602 ;
  assign n31324 = n2129 & n10819 ;
  assign n31325 = ~n26489 & n31324 ;
  assign n31326 = ( n6789 & n17881 ) | ( n6789 & ~n31325 ) | ( n17881 & ~n31325 ) ;
  assign n31327 = n5685 ^ n5430 ^ 1'b0 ;
  assign n31328 = ( n11599 & n17771 ) | ( n11599 & ~n31327 ) | ( n17771 & ~n31327 ) ;
  assign n31329 = ~n16295 & n31328 ;
  assign n31330 = n3940 & ~n15130 ;
  assign n31333 = n3176 ^ n269 ^ 1'b0 ;
  assign n31334 = ~n9083 & n31333 ;
  assign n31332 = n4185 & n20740 ;
  assign n31335 = n31334 ^ n31332 ^ 1'b0 ;
  assign n31331 = ~n12623 & n17780 ;
  assign n31336 = n31335 ^ n31331 ^ 1'b0 ;
  assign n31337 = n31336 ^ n21803 ^ 1'b0 ;
  assign n31338 = n31330 | n31337 ;
  assign n31339 = n31338 ^ n14295 ^ n12976 ;
  assign n31340 = n396 | n1076 ;
  assign n31341 = n29344 ^ n21318 ^ n20795 ;
  assign n31342 = n8231 ^ n162 ^ 1'b0 ;
  assign n31343 = n21251 & ~n31342 ;
  assign n31344 = n31343 ^ n14283 ^ 1'b0 ;
  assign n31345 = ~n5975 & n28354 ;
  assign n31346 = n636 & n31345 ;
  assign n31347 = n21863 ^ n19987 ^ 1'b0 ;
  assign n31348 = n29047 | n31347 ;
  assign n31349 = n31348 ^ n43 ^ 1'b0 ;
  assign n31350 = n10348 | n17299 ;
  assign n31352 = n13505 ^ n2714 ^ 1'b0 ;
  assign n31351 = ( n2889 & n11260 ) | ( n2889 & ~n17809 ) | ( n11260 & ~n17809 ) ;
  assign n31353 = n31352 ^ n31351 ^ n8392 ;
  assign n31354 = n7963 & ~n28454 ;
  assign n31355 = n31354 ^ n11809 ^ 1'b0 ;
  assign n31356 = n26665 ^ n4572 ^ n3496 ;
  assign n31357 = ~n11314 & n29303 ;
  assign n31358 = n15612 ^ n12269 ^ 1'b0 ;
  assign n31359 = n5167 & ~n31358 ;
  assign n31360 = n17369 & n31359 ;
  assign n31362 = n6451 ^ n1993 ^ 1'b0 ;
  assign n31361 = n644 & ~n24562 ;
  assign n31363 = n31362 ^ n31361 ^ n17202 ;
  assign n31364 = n27608 & n31363 ;
  assign n31365 = n102 & ~n230 ;
  assign n31366 = n15804 & ~n31365 ;
  assign n31367 = n5099 & ~n31366 ;
  assign n31368 = ~n722 & n8407 ;
  assign n31369 = n31367 & n31368 ;
  assign n31370 = ~n8145 & n31369 ;
  assign n31371 = ~n536 & n31370 ;
  assign n31372 = n31371 ^ n23134 ^ 1'b0 ;
  assign n31373 = n1464 | n6953 ;
  assign n31374 = n7494 ^ n4237 ^ 1'b0 ;
  assign n31375 = ~n7586 & n31374 ;
  assign n31376 = n6167 & n18363 ;
  assign n31377 = n2882 & n3255 ;
  assign n31378 = n27272 ^ n19090 ^ n18022 ;
  assign n31379 = n31377 & n31378 ;
  assign n31380 = ( ~n3687 & n4681 ) | ( ~n3687 & n13240 ) | ( n4681 & n13240 ) ;
  assign n31381 = ~n3039 & n3736 ;
  assign n31382 = n17053 | n17897 ;
  assign n31383 = n31381 & n31382 ;
  assign n31384 = n2544 ^ n814 ^ 1'b0 ;
  assign n31385 = n3038 & n23004 ;
  assign n31386 = n156 & n31385 ;
  assign n31387 = n31386 ^ n23 ^ 1'b0 ;
  assign n31388 = n2586 & ~n11882 ;
  assign n31389 = n31388 ^ n4124 ^ 1'b0 ;
  assign n31390 = ~n7568 & n31389 ;
  assign n31391 = n31387 & n31390 ;
  assign n31392 = n20842 ^ n3174 ^ 1'b0 ;
  assign n31393 = n11558 ^ n2790 ^ 1'b0 ;
  assign n31394 = n31393 ^ n31071 ^ n1364 ;
  assign n31395 = ~n31392 & n31394 ;
  assign n31396 = n1169 & n12470 ;
  assign n31397 = n31396 ^ n23529 ^ 1'b0 ;
  assign n31398 = ( n10812 & ~n27888 ) | ( n10812 & n31397 ) | ( ~n27888 & n31397 ) ;
  assign n31399 = ~n5511 & n26012 ;
  assign n31400 = n213 | n8291 ;
  assign n31401 = ( n8091 & n31399 ) | ( n8091 & ~n31400 ) | ( n31399 & ~n31400 ) ;
  assign n31402 = ( n7505 & n9060 ) | ( n7505 & ~n12593 ) | ( n9060 & ~n12593 ) ;
  assign n31403 = n31402 ^ n12551 ^ n3286 ;
  assign n31404 = n31401 & ~n31403 ;
  assign n31405 = n22688 | n27689 ;
  assign n31406 = n4252 | n31405 ;
  assign n31407 = n19775 ^ n4189 ^ n949 ;
  assign n31408 = n14043 | n31407 ;
  assign n31409 = n24240 ^ n9649 ^ 1'b0 ;
  assign n31413 = n2582 | n4226 ;
  assign n31410 = n7443 & n8256 ;
  assign n31411 = ~n6544 & n20487 ;
  assign n31412 = ( n20661 & n31410 ) | ( n20661 & n31411 ) | ( n31410 & n31411 ) ;
  assign n31414 = n31413 ^ n31412 ^ 1'b0 ;
  assign n31415 = n11365 ^ n2523 ^ 1'b0 ;
  assign n31416 = n28580 | n31415 ;
  assign n31417 = n8889 | n31416 ;
  assign n31418 = n31417 ^ n15520 ^ 1'b0 ;
  assign n31419 = n13738 | n21311 ;
  assign n31420 = n6675 & ~n31419 ;
  assign n31421 = n3922 & ~n14373 ;
  assign n31422 = n31420 & ~n31421 ;
  assign n31423 = n22878 ^ n12527 ^ 1'b0 ;
  assign n31424 = n30953 & ~n31423 ;
  assign n31425 = n20322 ^ n13249 ^ 1'b0 ;
  assign n31426 = n11570 ^ n10125 ^ n5097 ;
  assign n31427 = n17842 | n18458 ;
  assign n31428 = n23229 ^ n17912 ^ n2831 ;
  assign n31429 = n10390 & n24513 ;
  assign n31430 = n906 | n23756 ;
  assign n31431 = n31430 ^ n6953 ^ 1'b0 ;
  assign n31432 = n31431 ^ n11253 ^ 1'b0 ;
  assign n31433 = n4337 | n31432 ;
  assign n31434 = n6671 & n11006 ;
  assign n31435 = n31434 ^ n4703 ^ 1'b0 ;
  assign n31436 = n3577 & ~n30782 ;
  assign n31437 = n25276 ^ n17881 ^ 1'b0 ;
  assign n31438 = n7074 | n15177 ;
  assign n31439 = n43 & ~n31438 ;
  assign n31440 = ( n17710 & n28179 ) | ( n17710 & ~n31439 ) | ( n28179 & ~n31439 ) ;
  assign n31445 = n6623 & ~n7404 ;
  assign n31441 = n12573 | n25543 ;
  assign n31442 = n4093 | n31441 ;
  assign n31443 = n31442 ^ n27063 ^ 1'b0 ;
  assign n31444 = n5870 | n31443 ;
  assign n31446 = n31445 ^ n31444 ^ 1'b0 ;
  assign n31447 = n8140 | n30380 ;
  assign n31448 = n17325 | n31447 ;
  assign n31450 = n4572 & ~n10741 ;
  assign n31451 = n10741 & n31450 ;
  assign n31449 = n8574 ^ n3261 ^ n1487 ;
  assign n31452 = n31451 ^ n31449 ^ n19238 ;
  assign n31453 = n6712 | n30295 ;
  assign n31454 = ~n7006 & n11974 ;
  assign n31455 = n17062 ^ n13682 ^ n5580 ;
  assign n31456 = n5199 & ~n31455 ;
  assign n31457 = n23193 & n24481 ;
  assign n31458 = n31457 ^ n17809 ^ 1'b0 ;
  assign n31468 = n18377 | n20374 ;
  assign n31462 = ~n1515 & n2524 ;
  assign n31463 = n1515 & n31462 ;
  assign n31464 = n31463 ^ n1003 ^ 1'b0 ;
  assign n31465 = n9152 | n31464 ;
  assign n31466 = n31464 & ~n31465 ;
  assign n31459 = n4122 ^ n1193 ^ 1'b0 ;
  assign n31460 = n31459 ^ n23607 ^ 1'b0 ;
  assign n31461 = n31460 ^ n23315 ^ n15100 ;
  assign n31467 = n31466 ^ n31461 ^ n24227 ;
  assign n31469 = n31468 ^ n31467 ^ 1'b0 ;
  assign n31470 = n15130 & n31344 ;
  assign n31471 = n31470 ^ n7358 ^ 1'b0 ;
  assign n31472 = n957 | n8933 ;
  assign n31473 = n31472 ^ n101 ^ 1'b0 ;
  assign n31474 = n31473 ^ n16339 ^ n11919 ;
  assign n31475 = n20137 ^ n10265 ^ 1'b0 ;
  assign n31476 = ~n31474 & n31475 ;
  assign n31477 = n5737 | n30870 ;
  assign n31478 = n6554 | n8205 ;
  assign n31479 = n2180 & ~n2846 ;
  assign n31480 = ~n24905 & n31479 ;
  assign n31481 = ~n31478 & n31480 ;
  assign n31482 = n7900 ^ n6411 ^ 1'b0 ;
  assign n31483 = ~n16334 & n31482 ;
  assign n31484 = ~n28133 & n31483 ;
  assign n31485 = n31484 ^ n26643 ^ 1'b0 ;
  assign n31486 = n30307 ^ n6175 ^ 1'b0 ;
  assign n31487 = n15012 ^ n628 ^ 1'b0 ;
  assign n31488 = n31486 | n31487 ;
  assign n31489 = n664 & n20059 ;
  assign n31490 = ~n10428 & n31489 ;
  assign n31491 = n31490 ^ n3294 ^ 1'b0 ;
  assign n31492 = n3825 & n30128 ;
  assign n31495 = ( n4243 & ~n9150 ) | ( n4243 & n23040 ) | ( ~n9150 & n23040 ) ;
  assign n31493 = n3987 | n9663 ;
  assign n31494 = n4422 & ~n31493 ;
  assign n31496 = n31495 ^ n31494 ^ 1'b0 ;
  assign n31497 = n27013 | n31166 ;
  assign n31498 = n31497 ^ n15375 ^ 1'b0 ;
  assign n31499 = n216 | n15290 ;
  assign n31500 = n29091 | n31499 ;
  assign n31501 = n7921 ^ n3892 ^ 1'b0 ;
  assign n31502 = n31501 ^ n23761 ^ n9197 ;
  assign n31503 = n31500 | n31502 ;
  assign n31504 = n1921 | n6016 ;
  assign n31505 = n22131 & ~n31504 ;
  assign n31506 = n19894 & n22202 ;
  assign n31507 = n31505 & ~n31506 ;
  assign n31508 = n24350 & n26600 ;
  assign n31509 = n420 & ~n27753 ;
  assign n31510 = n23676 ^ n14539 ^ 1'b0 ;
  assign n31511 = n13018 & ~n24655 ;
  assign n31514 = n430 & n7156 ;
  assign n31512 = n2839 & n10125 ;
  assign n31513 = ~n21441 & n31512 ;
  assign n31515 = n31514 ^ n31513 ^ n17114 ;
  assign n31516 = n27739 ^ n272 ^ 1'b0 ;
  assign n31517 = ~n8004 & n14190 ;
  assign n31518 = n22130 ^ n10356 ^ 1'b0 ;
  assign n31519 = n19813 ^ n14777 ^ 1'b0 ;
  assign n31520 = ( n62 & ~n1238 ) | ( n62 & n7779 ) | ( ~n1238 & n7779 ) ;
  assign n31521 = n23904 | n31520 ;
  assign n31522 = n31521 ^ n26113 ^ 1'b0 ;
  assign n31523 = n3630 ^ n2131 ^ 1'b0 ;
  assign n31524 = ~n3394 & n31523 ;
  assign n31525 = ~n1660 & n31524 ;
  assign n31526 = n29448 & n31525 ;
  assign n31527 = ~n2230 & n10755 ;
  assign n31528 = n31527 ^ n1545 ^ 1'b0 ;
  assign n31530 = n7402 ^ n524 ^ 1'b0 ;
  assign n31531 = n31530 ^ n15675 ^ 1'b0 ;
  assign n31529 = n11378 | n14897 ;
  assign n31532 = n31531 ^ n31529 ^ 1'b0 ;
  assign n31535 = n14211 ^ n1768 ^ n1310 ;
  assign n31534 = n9113 & n21394 ;
  assign n31536 = n31535 ^ n31534 ^ 1'b0 ;
  assign n31533 = n12022 ^ n10442 ^ n5638 ;
  assign n31537 = n31536 ^ n31533 ^ 1'b0 ;
  assign n31538 = n1110 | n31537 ;
  assign n31539 = ~n184 & n1715 ;
  assign n31540 = n31539 ^ n8382 ^ 1'b0 ;
  assign n31541 = ( n381 & n8695 ) | ( n381 & ~n10240 ) | ( n8695 & ~n10240 ) ;
  assign n31542 = ~n2827 & n3401 ;
  assign n31543 = n8448 & n31542 ;
  assign n31544 = n10285 | n15499 ;
  assign n31545 = ~n31543 & n31544 ;
  assign n31546 = n31545 ^ n10236 ^ 1'b0 ;
  assign n31549 = n8032 ^ n940 ^ 1'b0 ;
  assign n31547 = n6981 & n10329 ;
  assign n31548 = n12033 & ~n31547 ;
  assign n31550 = n31549 ^ n31548 ^ 1'b0 ;
  assign n31551 = n11709 & n31550 ;
  assign n31552 = n31551 ^ n838 ^ 1'b0 ;
  assign n31553 = n1344 | n14898 ;
  assign n31554 = n26462 ^ n13448 ^ 1'b0 ;
  assign n31555 = n3732 | n14893 ;
  assign n31556 = n4239 & ~n31555 ;
  assign n31557 = n11503 | n31556 ;
  assign n31558 = n31557 ^ n17732 ^ 1'b0 ;
  assign n31559 = n31558 ^ n19232 ^ 1'b0 ;
  assign n31560 = ~n15568 & n31559 ;
  assign n31561 = n22249 ^ n19407 ^ 1'b0 ;
  assign n31562 = n24044 ^ n14177 ^ 1'b0 ;
  assign n31563 = n7087 ^ n5748 ^ n13 ;
  assign n31564 = n3650 & n31563 ;
  assign n31565 = n18531 ^ n17788 ^ 1'b0 ;
  assign n31566 = n17018 | n31565 ;
  assign n31567 = ~n11450 & n18585 ;
  assign n31568 = ( ~n14305 & n15324 ) | ( ~n14305 & n18639 ) | ( n15324 & n18639 ) ;
  assign n31569 = n6523 ^ n1822 ^ 1'b0 ;
  assign n31570 = n7507 & n31569 ;
  assign n31571 = n11277 ^ n10208 ^ 1'b0 ;
  assign n31572 = n1288 & ~n31571 ;
  assign n31573 = n31570 & n31572 ;
  assign n31574 = ~n7750 & n31573 ;
  assign n31575 = n4974 ^ n351 ^ 1'b0 ;
  assign n31576 = n5702 | n31575 ;
  assign n31577 = ~n9909 & n31576 ;
  assign n31578 = n10441 & n31577 ;
  assign n31579 = n19798 & n21466 ;
  assign n31580 = n21813 ^ n572 ^ 1'b0 ;
  assign n31581 = n19829 & n31580 ;
  assign n31584 = n10042 & n21682 ;
  assign n31582 = n12416 | n30681 ;
  assign n31583 = n28845 & n31582 ;
  assign n31585 = n31584 ^ n31583 ^ 1'b0 ;
  assign n31586 = n3203 & n25620 ;
  assign n31587 = n31586 ^ n4435 ^ 1'b0 ;
  assign n31588 = n25061 ^ n12617 ^ 1'b0 ;
  assign n31589 = n26449 | n31588 ;
  assign n31593 = n1811 & n5799 ;
  assign n31594 = ~n1811 & n31593 ;
  assign n31590 = n2621 | n6473 ;
  assign n31591 = n31590 ^ n2307 ^ 1'b0 ;
  assign n31592 = n31591 ^ n9752 ^ 1'b0 ;
  assign n31595 = n31594 ^ n31592 ^ 1'b0 ;
  assign n31596 = n19598 ^ n16768 ^ n12406 ;
  assign n31597 = ( ~n3863 & n14204 ) | ( ~n3863 & n31596 ) | ( n14204 & n31596 ) ;
  assign n31598 = n5182 & ~n9598 ;
  assign n31599 = ~n9147 & n31598 ;
  assign n31600 = n31599 ^ n1876 ^ n994 ;
  assign n31601 = ( n5048 & n25326 ) | ( n5048 & ~n31600 ) | ( n25326 & ~n31600 ) ;
  assign n31602 = n1853 | n5228 ;
  assign n31603 = n31602 ^ n14593 ^ 1'b0 ;
  assign n31604 = ~n3904 & n31603 ;
  assign n31605 = n31604 ^ n10465 ^ 1'b0 ;
  assign n31606 = n3717 & ~n31605 ;
  assign n31607 = n19409 ^ n16750 ^ n4803 ;
  assign n31608 = n10849 & n31607 ;
  assign n31609 = ~n695 & n3112 ;
  assign n31610 = n1969 & ~n17174 ;
  assign n31611 = ~n1066 & n2226 ;
  assign n31612 = n384 ^ n43 ^ 1'b0 ;
  assign n31613 = n2338 & n31612 ;
  assign n31614 = n5229 & n9260 ;
  assign n31615 = ~n5635 & n31614 ;
  assign n31616 = ( n5924 & n16527 ) | ( n5924 & n31615 ) | ( n16527 & n31615 ) ;
  assign n31617 = n7329 | n21694 ;
  assign n31618 = n850 & n31617 ;
  assign n31619 = ~n17162 & n31618 ;
  assign n31620 = n31616 | n31619 ;
  assign n31621 = n1993 & ~n31620 ;
  assign n31622 = ( n863 & ~n4498 ) | ( n863 & n31621 ) | ( ~n4498 & n31621 ) ;
  assign n31623 = ( n15205 & ~n31613 ) | ( n15205 & n31622 ) | ( ~n31613 & n31622 ) ;
  assign n31624 = n31623 ^ n4915 ^ 1'b0 ;
  assign n31625 = n19012 & ~n21968 ;
  assign n31626 = n31625 ^ n3658 ^ 1'b0 ;
  assign n31627 = n14057 | n17906 ;
  assign n31628 = n6454 & n22831 ;
  assign n31629 = n20288 | n31628 ;
  assign n31630 = n31628 & ~n31629 ;
  assign n31631 = n31138 ^ n17813 ^ 1'b0 ;
  assign n31632 = n11178 & ~n12309 ;
  assign n31633 = n9642 & ~n12505 ;
  assign n31634 = n2221 ^ n2092 ^ 1'b0 ;
  assign n31635 = ( n1818 & n5406 ) | ( n1818 & n31634 ) | ( n5406 & n31634 ) ;
  assign n31636 = n647 & n2495 ;
  assign n31637 = n31636 ^ n2186 ^ 1'b0 ;
  assign n31638 = ~n8101 & n22661 ;
  assign n31639 = ~n15751 & n31638 ;
  assign n31640 = ~n8303 & n20689 ;
  assign n31641 = n31640 ^ n1625 ^ 1'b0 ;
  assign n31642 = n15009 & n23143 ;
  assign n31643 = ~n16385 & n31642 ;
  assign n31644 = n8193 ^ n6583 ^ n3531 ;
  assign n31645 = n1120 & n31644 ;
  assign n31647 = n1787 & n13284 ;
  assign n31646 = n10362 & ~n20902 ;
  assign n31648 = n31647 ^ n31646 ^ 1'b0 ;
  assign n31649 = ( n12124 & n13415 ) | ( n12124 & ~n31648 ) | ( n13415 & ~n31648 ) ;
  assign n31650 = n28085 ^ n16050 ^ n7490 ;
  assign n31651 = ~n10079 & n31650 ;
  assign n31652 = n6078 | n6835 ;
  assign n31653 = n2365 & ~n31652 ;
  assign n31654 = ~n8158 & n31653 ;
  assign n31655 = n22582 ^ n3232 ^ 1'b0 ;
  assign n31656 = ( n3642 & n28494 ) | ( n3642 & ~n31655 ) | ( n28494 & ~n31655 ) ;
  assign n31657 = n15172 ^ n7144 ^ 1'b0 ;
  assign n31658 = ~n10669 & n21514 ;
  assign n31659 = ~n31657 & n31658 ;
  assign n31660 = ~n14677 & n16356 ;
  assign n31661 = ~n12053 & n31660 ;
  assign n31662 = n31661 ^ n11824 ^ 1'b0 ;
  assign n31663 = n23795 & ~n28760 ;
  assign n31664 = ( n4493 & ~n24789 ) | ( n4493 & n31663 ) | ( ~n24789 & n31663 ) ;
  assign n31665 = n11753 & n22796 ;
  assign n31666 = ~n3828 & n16625 ;
  assign n31667 = ~n31665 & n31666 ;
  assign n31668 = n8138 | n9357 ;
  assign n31669 = n29017 & ~n31668 ;
  assign n31670 = ~n5891 & n12426 ;
  assign n31671 = n18843 | n31670 ;
  assign n31672 = n31671 ^ n8248 ^ 1'b0 ;
  assign n31674 = n25509 ^ n8000 ^ 1'b0 ;
  assign n31673 = ( n3214 & ~n5824 ) | ( n3214 & n17408 ) | ( ~n5824 & n17408 ) ;
  assign n31675 = n31674 ^ n31673 ^ n24215 ;
  assign n31676 = n15706 ^ n14833 ^ n3634 ;
  assign n31677 = n16826 ^ n12258 ^ n6787 ;
  assign n31678 = n31677 ^ n6109 ^ n575 ;
  assign n31679 = n16738 & n31678 ;
  assign n31680 = n31679 ^ n14641 ^ n5967 ;
  assign n31681 = n8314 | n23998 ;
  assign n31682 = n31681 ^ n14332 ^ 1'b0 ;
  assign n31683 = n11980 ^ n6091 ^ 1'b0 ;
  assign n31684 = ~n31682 & n31683 ;
  assign n31685 = n7766 & n26794 ;
  assign n31687 = ~n6375 & n12060 ;
  assign n31688 = n5009 | n31687 ;
  assign n31686 = n1287 | n16232 ;
  assign n31689 = n31688 ^ n31686 ^ 1'b0 ;
  assign n31690 = n31689 ^ n29827 ^ 1'b0 ;
  assign n31691 = n22494 | n31690 ;
  assign n31692 = n31691 ^ n28253 ^ 1'b0 ;
  assign n31693 = n200 & ~n2940 ;
  assign n31694 = n5557 ^ n5549 ^ 1'b0 ;
  assign n31695 = n31694 ^ n30602 ^ 1'b0 ;
  assign n31696 = n31695 ^ n14300 ^ n10342 ;
  assign n31697 = n31696 ^ n22613 ^ 1'b0 ;
  assign n31698 = n21017 & n22210 ;
  assign n31699 = n31698 ^ n4473 ^ 1'b0 ;
  assign n31700 = n192 & ~n31699 ;
  assign n31701 = n17916 & ~n20460 ;
  assign n31702 = ~n9191 & n31701 ;
  assign n31703 = n3397 & n17165 ;
  assign n31704 = n23480 ^ n7847 ^ 1'b0 ;
  assign n31705 = ~n5412 & n18278 ;
  assign n31706 = ~n18278 & n31705 ;
  assign n31707 = n2741 | n23760 ;
  assign n31708 = n29910 | n31707 ;
  assign n31709 = n36 & n31708 ;
  assign n31710 = ~n31706 & n31709 ;
  assign n31711 = n17366 ^ n1868 ^ 1'b0 ;
  assign n31712 = n26929 & ~n31711 ;
  assign n31713 = n5078 | n5197 ;
  assign n31714 = n31713 ^ n3240 ^ 1'b0 ;
  assign n31715 = ~n14943 & n15865 ;
  assign n31716 = n13942 & ~n31715 ;
  assign n31717 = n31716 ^ n7739 ^ 1'b0 ;
  assign n31718 = n31717 ^ n7121 ^ n4704 ;
  assign n31722 = n22228 ^ n4582 ^ n3526 ;
  assign n31723 = n31722 ^ n23432 ^ 1'b0 ;
  assign n31724 = n14183 ^ n5072 ^ 1'b0 ;
  assign n31725 = ~n31723 & n31724 ;
  assign n31726 = n31725 ^ n16369 ^ 1'b0 ;
  assign n31727 = n31726 ^ n14526 ^ 1'b0 ;
  assign n31719 = n3693 & ~n28153 ;
  assign n31720 = n31719 ^ n3345 ^ 1'b0 ;
  assign n31721 = n12395 & ~n31720 ;
  assign n31728 = n31727 ^ n31721 ^ 1'b0 ;
  assign n31729 = n19795 ^ n19463 ^ 1'b0 ;
  assign n31730 = n15290 & n31729 ;
  assign n31731 = n29683 ^ n24676 ^ 1'b0 ;
  assign n31732 = n11162 & n31731 ;
  assign n31733 = ( ~n15003 & n19544 ) | ( ~n15003 & n31732 ) | ( n19544 & n31732 ) ;
  assign n31734 = n13065 ^ n6670 ^ n5461 ;
  assign n31735 = n6839 & ~n31734 ;
  assign n31736 = n13123 ^ n7039 ^ 1'b0 ;
  assign n31737 = n7801 & n31736 ;
  assign n31738 = n31737 ^ n14204 ^ 1'b0 ;
  assign n31739 = n6345 & n29663 ;
  assign n31740 = n31623 ^ n11782 ^ 1'b0 ;
  assign n31741 = n17357 ^ n42 ^ 1'b0 ;
  assign n31742 = ~n14278 & n31741 ;
  assign n31743 = n21352 ^ n11519 ^ n5322 ;
  assign n31744 = n27064 & n31743 ;
  assign n31745 = n29140 & n31744 ;
  assign n31746 = n13059 & n30461 ;
  assign n31747 = n15975 ^ n5254 ^ 1'b0 ;
  assign n31748 = n18121 ^ n17614 ^ n740 ;
  assign n31749 = n9070 | n31010 ;
  assign n31750 = n31457 ^ n11531 ^ n8833 ;
  assign n31751 = n2029 & ~n10729 ;
  assign n31752 = n31751 ^ n1889 ^ 1'b0 ;
  assign n31753 = n6221 ^ n5735 ^ n1484 ;
  assign n31754 = n31753 ^ n18601 ^ 1'b0 ;
  assign n31755 = n3628 | n12239 ;
  assign n31756 = n21416 ^ n8560 ^ 1'b0 ;
  assign n31757 = ~n20609 & n31756 ;
  assign n31758 = n31757 ^ n1374 ^ 1'b0 ;
  assign n31759 = n31755 | n31758 ;
  assign n31760 = n19013 | n20399 ;
  assign n31761 = ~n2186 & n27525 ;
  assign n31762 = n31761 ^ n22227 ^ 1'b0 ;
  assign n31763 = ~n1080 & n7402 ;
  assign n31764 = n31763 ^ n11055 ^ 1'b0 ;
  assign n31765 = n31764 ^ n9490 ^ n1094 ;
  assign n31766 = n30957 | n31765 ;
  assign n31767 = n18 | n31766 ;
  assign n31768 = n2431 & n22369 ;
  assign n31769 = n2735 | n6947 ;
  assign n31770 = n31769 ^ n10727 ^ n5073 ;
  assign n31771 = n14572 & n31770 ;
  assign n31772 = n3650 & n18099 ;
  assign n31773 = n19964 ^ n10448 ^ 1'b0 ;
  assign n31774 = n31772 & n31773 ;
  assign n31775 = n220 & ~n31774 ;
  assign n31776 = n8114 ^ n4508 ^ 1'b0 ;
  assign n31777 = n18581 ^ n6317 ^ 1'b0 ;
  assign n31778 = n31776 & ~n31777 ;
  assign n31779 = n3067 & n10543 ;
  assign n31780 = n31779 ^ n23445 ^ 1'b0 ;
  assign n31781 = n7634 & n20053 ;
  assign n31782 = n29997 ^ n11102 ^ 1'b0 ;
  assign n31783 = n5533 & n31782 ;
  assign n31784 = n2414 & ~n7605 ;
  assign n31785 = n9012 ^ n578 ^ 1'b0 ;
  assign n31786 = n709 | n31785 ;
  assign n31787 = n12823 & n15017 ;
  assign n31788 = n31786 & n31787 ;
  assign n31789 = n676 | n31788 ;
  assign n31790 = n31789 ^ n29863 ^ 1'b0 ;
  assign n31791 = n13522 ^ n6069 ^ n2373 ;
  assign n31792 = n9584 & n31791 ;
  assign n31793 = ~n8253 & n31792 ;
  assign n31794 = ~n10261 & n10282 ;
  assign n31795 = ( n3114 & n15976 ) | ( n3114 & ~n31794 ) | ( n15976 & ~n31794 ) ;
  assign n31796 = ~n5241 & n31795 ;
  assign n31797 = n31796 ^ n20188 ^ 1'b0 ;
  assign n31798 = n31797 ^ n22378 ^ n21313 ;
  assign n31799 = n14438 & n20715 ;
  assign n31800 = ( ~n752 & n12571 ) | ( ~n752 & n31799 ) | ( n12571 & n31799 ) ;
  assign n31801 = n10520 | n18684 ;
  assign n31802 = n31801 ^ n14363 ^ 1'b0 ;
  assign n31803 = n4911 & n31802 ;
  assign n31804 = n27123 & n31803 ;
  assign n31805 = n24282 & n31256 ;
  assign n31806 = n4892 & n8784 ;
  assign n31807 = n31806 ^ n12271 ^ 1'b0 ;
  assign n31808 = n969 & ~n29358 ;
  assign n31809 = n31808 ^ n6611 ^ 1'b0 ;
  assign n31810 = n31807 | n31809 ;
  assign n31811 = n21241 ^ n15685 ^ n324 ;
  assign n31812 = n5653 ^ n3793 ^ 1'b0 ;
  assign n31813 = n9833 & n31812 ;
  assign n31814 = n22318 & n31813 ;
  assign n31815 = n31814 ^ n24748 ^ n14226 ;
  assign n31816 = ~n1891 & n19695 ;
  assign n31817 = n13761 ^ n318 ^ 1'b0 ;
  assign n31818 = n31816 | n31817 ;
  assign n31819 = ( ~n8204 & n12878 ) | ( ~n8204 & n14104 ) | ( n12878 & n14104 ) ;
  assign n31820 = n24046 | n31819 ;
  assign n31821 = n31820 ^ n5704 ^ 1'b0 ;
  assign n31822 = n5545 | n29668 ;
  assign n31823 = n3781 & ~n31822 ;
  assign n31824 = n4413 | n31823 ;
  assign n31825 = n31824 ^ n15490 ^ 1'b0 ;
  assign n31826 = n3503 | n19695 ;
  assign n31827 = n31826 ^ n28347 ^ 1'b0 ;
  assign n31828 = ~n14059 & n22542 ;
  assign n31829 = n16158 & n24612 ;
  assign n31830 = n31829 ^ n6496 ^ 1'b0 ;
  assign n31831 = n31830 ^ n27744 ^ n5913 ;
  assign n31833 = n14797 ^ n4341 ^ 1'b0 ;
  assign n31832 = n13308 & n19979 ;
  assign n31834 = n31833 ^ n31832 ^ 1'b0 ;
  assign n31835 = n19572 ^ n14878 ^ n8982 ;
  assign n31836 = n31835 ^ n974 ^ 1'b0 ;
  assign n31837 = n31834 & ~n31836 ;
  assign n31838 = n18695 ^ n10261 ^ 1'b0 ;
  assign n31839 = ~n1050 & n31838 ;
  assign n31841 = n11307 | n31129 ;
  assign n31842 = n12931 | n31841 ;
  assign n31843 = n31842 ^ n26711 ^ 1'b0 ;
  assign n31840 = n21396 & n30465 ;
  assign n31844 = n31843 ^ n31840 ^ n3785 ;
  assign n31845 = n15280 ^ n8497 ^ 1'b0 ;
  assign n31846 = n3073 | n31845 ;
  assign n31847 = n558 | n31174 ;
  assign n31848 = n969 & ~n31847 ;
  assign n31849 = n6027 | n31848 ;
  assign n31850 = n13697 ^ n9999 ^ 1'b0 ;
  assign n31852 = n6550 | n20147 ;
  assign n31853 = n20977 & ~n31852 ;
  assign n31854 = ( n10962 & n11037 ) | ( n10962 & ~n31853 ) | ( n11037 & ~n31853 ) ;
  assign n31851 = n21323 & ~n27925 ;
  assign n31855 = n31854 ^ n31851 ^ 1'b0 ;
  assign n31856 = n263 & ~n15112 ;
  assign n31857 = ~n11437 & n31856 ;
  assign n31858 = ( n5339 & n6211 ) | ( n5339 & ~n31857 ) | ( n6211 & ~n31857 ) ;
  assign n31859 = ~n5430 & n31858 ;
  assign n31860 = n31859 ^ n9626 ^ 1'b0 ;
  assign n31861 = n5430 ^ n1172 ^ n1003 ;
  assign n31862 = n6557 & ~n31861 ;
  assign n31863 = n9059 | n29905 ;
  assign n31864 = n31863 ^ n22244 ^ 1'b0 ;
  assign n31865 = n12903 ^ n2139 ^ 1'b0 ;
  assign n31867 = n5585 & n7707 ;
  assign n31868 = n31867 ^ n1156 ^ 1'b0 ;
  assign n31869 = ~n11318 & n31868 ;
  assign n31866 = ~n7411 & n8241 ;
  assign n31870 = n31869 ^ n31866 ^ 1'b0 ;
  assign n31871 = n23113 & ~n31870 ;
  assign n31872 = n31865 & ~n31871 ;
  assign n31873 = n31864 & n31872 ;
  assign n31874 = n5537 | n14614 ;
  assign n31875 = n5592 & n31874 ;
  assign n31876 = n2704 & n31875 ;
  assign n31877 = n18138 ^ n15972 ^ 1'b0 ;
  assign n31880 = x10 | n18277 ;
  assign n31881 = n7392 & ~n31880 ;
  assign n31878 = ~n966 & n7169 ;
  assign n31879 = n185 & n31878 ;
  assign n31882 = n31881 ^ n31879 ^ n17324 ;
  assign n31883 = n15224 | n22607 ;
  assign n31884 = n2256 ^ n687 ^ 1'b0 ;
  assign n31885 = n13850 & ~n26408 ;
  assign n31886 = n31884 & n31885 ;
  assign n31887 = n31886 ^ n12759 ^ 1'b0 ;
  assign n31889 = n11277 & ~n11824 ;
  assign n31890 = n31889 ^ n24735 ^ 1'b0 ;
  assign n31888 = ~n19066 & n31727 ;
  assign n31891 = n31890 ^ n31888 ^ 1'b0 ;
  assign n31895 = ~n1360 & n5280 ;
  assign n31896 = n1360 & n31895 ;
  assign n31892 = n9552 | n10461 ;
  assign n31893 = n9552 & ~n31892 ;
  assign n31894 = n11955 | n31893 ;
  assign n31897 = n31896 ^ n31894 ^ 1'b0 ;
  assign n31898 = n31897 ^ n23285 ^ 1'b0 ;
  assign n31899 = ~n14379 & n31898 ;
  assign n31900 = n7026 ^ n5702 ^ n426 ;
  assign n31901 = n11609 ^ n6098 ^ 1'b0 ;
  assign n31902 = ( n408 & ~n15965 ) | ( n408 & n31901 ) | ( ~n15965 & n31901 ) ;
  assign n31903 = n15641 ^ n9506 ^ 1'b0 ;
  assign n31904 = ~n408 & n31903 ;
  assign n31905 = n31904 ^ n1400 ^ 1'b0 ;
  assign n31906 = n8745 & n31905 ;
  assign n31907 = n21172 | n31906 ;
  assign n31908 = ( n6422 & n12901 ) | ( n6422 & n14246 ) | ( n12901 & n14246 ) ;
  assign n31909 = n30057 ^ n21652 ^ 1'b0 ;
  assign n31910 = n23194 | n31909 ;
  assign n31911 = n31908 | n31910 ;
  assign n31912 = n31911 ^ n28526 ^ 1'b0 ;
  assign n31913 = ~n890 & n1357 ;
  assign n31914 = ~n1357 & n31913 ;
  assign n31915 = n3027 | n31914 ;
  assign n31916 = n13572 | n31915 ;
  assign n31917 = n31915 & ~n31916 ;
  assign n31918 = n27033 & ~n31917 ;
  assign n31919 = n31917 & n31918 ;
  assign n31920 = n23134 ^ n13863 ^ 1'b0 ;
  assign n31921 = n10935 & ~n15079 ;
  assign n31922 = n4967 ^ n3508 ^ 1'b0 ;
  assign n31923 = n22862 & n31922 ;
  assign n31925 = n14593 ^ n3460 ^ 1'b0 ;
  assign n31926 = n13608 | n31925 ;
  assign n31924 = n16 & ~n1818 ;
  assign n31927 = n31926 ^ n31924 ^ 1'b0 ;
  assign n31928 = n22200 ^ n6699 ^ n452 ;
  assign n31930 = n5229 & n6211 ;
  assign n31929 = n15838 ^ n13854 ^ n1409 ;
  assign n31931 = n31930 ^ n31929 ^ 1'b0 ;
  assign n31932 = n31928 | n31931 ;
  assign n31933 = n29517 ^ n2064 ^ 1'b0 ;
  assign n31934 = ( n853 & n31932 ) | ( n853 & n31933 ) | ( n31932 & n31933 ) ;
  assign n31935 = n7413 ^ n41 ^ 1'b0 ;
  assign n31936 = n31935 ^ n31393 ^ 1'b0 ;
  assign n31937 = n15796 ^ n10884 ^ 1'b0 ;
  assign n31938 = ( ~n14807 & n16032 ) | ( ~n14807 & n31937 ) | ( n16032 & n31937 ) ;
  assign n31939 = n23217 & n29704 ;
  assign n31940 = n8764 | n31939 ;
  assign n31941 = n11549 & ~n15233 ;
  assign n31942 = n14914 ^ n645 ^ 1'b0 ;
  assign n31943 = ~n31281 & n31942 ;
  assign n31944 = n9463 | n20811 ;
  assign n31945 = ( n6693 & n31334 ) | ( n6693 & n31944 ) | ( n31334 & n31944 ) ;
  assign n31946 = n31945 ^ n4093 ^ 1'b0 ;
  assign n31947 = n11533 & n31946 ;
  assign n31948 = n18126 ^ n7094 ^ 1'b0 ;
  assign n31949 = n31948 ^ n28327 ^ 1'b0 ;
  assign n31950 = ~n2871 & n24961 ;
  assign n31951 = ~n2259 & n31950 ;
  assign n31952 = n17973 ^ n8832 ^ 1'b0 ;
  assign n31954 = n6733 & ~n21136 ;
  assign n31955 = n31954 ^ n12677 ^ 1'b0 ;
  assign n31953 = n7864 & n28077 ;
  assign n31956 = n31955 ^ n31953 ^ n14026 ;
  assign n31957 = n947 & ~n31956 ;
  assign n31958 = n31957 ^ n31460 ^ n811 ;
  assign n31959 = n31958 ^ n23851 ^ 1'b0 ;
  assign n31960 = n6238 ^ n22 ^ 1'b0 ;
  assign n31961 = n31026 ^ n19213 ^ 1'b0 ;
  assign n31964 = n26276 ^ n9814 ^ 1'b0 ;
  assign n31962 = n8767 ^ n8321 ^ 1'b0 ;
  assign n31963 = n31962 ^ n962 ^ 1'b0 ;
  assign n31965 = n31964 ^ n31963 ^ 1'b0 ;
  assign n31966 = n31961 & ~n31965 ;
  assign n31967 = n9284 & n15244 ;
  assign n31968 = ( n755 & ~n5535 ) | ( n755 & n22210 ) | ( ~n5535 & n22210 ) ;
  assign n31969 = n31968 ^ n23979 ^ n1105 ;
  assign n31970 = n28243 ^ n352 ^ n283 ;
  assign n31971 = ~n5469 & n29027 ;
  assign n31972 = n31971 ^ n350 ^ 1'b0 ;
  assign n31974 = n8097 & n10656 ;
  assign n31975 = n31974 ^ n11635 ^ 1'b0 ;
  assign n31973 = n3932 & ~n28428 ;
  assign n31976 = n31975 ^ n31973 ^ 1'b0 ;
  assign n31977 = n31976 ^ n25998 ^ 1'b0 ;
  assign n31978 = n30991 ^ n2161 ^ 1'b0 ;
  assign n31979 = n19991 | n31978 ;
  assign n31980 = n12482 | n31979 ;
  assign n31981 = n31980 ^ n23047 ^ 1'b0 ;
  assign n31982 = n27477 ^ n17201 ^ 1'b0 ;
  assign n31983 = n15042 ^ n7124 ^ 1'b0 ;
  assign n31984 = ~n12921 & n24378 ;
  assign n31985 = ( n1003 & n31983 ) | ( n1003 & ~n31984 ) | ( n31983 & ~n31984 ) ;
  assign n31986 = n1948 | n31985 ;
  assign n31987 = n17123 & n29946 ;
  assign n31988 = n13218 | n30863 ;
  assign n31992 = n9052 ^ n4643 ^ 1'b0 ;
  assign n31989 = n10224 | n13538 ;
  assign n31990 = n31989 ^ n15543 ^ 1'b0 ;
  assign n31991 = n23480 | n31990 ;
  assign n31993 = n31992 ^ n31991 ^ n725 ;
  assign n31995 = ~n360 & n5004 ;
  assign n31996 = n31995 ^ n2434 ^ 1'b0 ;
  assign n31997 = ~n25522 & n31996 ;
  assign n31998 = n31997 ^ n1472 ^ 1'b0 ;
  assign n31999 = n31998 ^ n738 ^ 1'b0 ;
  assign n31994 = n1247 | n9820 ;
  assign n32000 = n31999 ^ n31994 ^ 1'b0 ;
  assign n32001 = n2589 & n25253 ;
  assign n32002 = n10579 & n32001 ;
  assign n32003 = n4976 & ~n13716 ;
  assign n32004 = n22185 & n32003 ;
  assign n32005 = n1179 & ~n3707 ;
  assign n32006 = n32005 ^ n15855 ^ 1'b0 ;
  assign n32007 = n32006 ^ n9084 ^ n5469 ;
  assign n32008 = ~n31549 & n32007 ;
  assign n32009 = n32008 ^ n18419 ^ 1'b0 ;
  assign n32010 = n32009 ^ n897 ^ 1'b0 ;
  assign n32011 = ~n32004 & n32010 ;
  assign n32012 = n8323 ^ n188 ^ 1'b0 ;
  assign n32013 = n8206 & ~n8597 ;
  assign n32014 = ~n5010 & n32013 ;
  assign n32015 = n23326 ^ n14347 ^ n10780 ;
  assign n32016 = n20496 ^ n2889 ^ 1'b0 ;
  assign n32017 = n27340 & n32016 ;
  assign n32018 = n8567 & n32017 ;
  assign n32019 = n32015 & n32018 ;
  assign n32020 = n24699 ^ n23023 ^ n17586 ;
  assign n32021 = n17648 ^ n1263 ^ n829 ;
  assign n32022 = n7978 | n32021 ;
  assign n32023 = n27699 & ~n32022 ;
  assign n32024 = n12235 | n32023 ;
  assign n32025 = ( n10634 & ~n15173 ) | ( n10634 & n24896 ) | ( ~n15173 & n24896 ) ;
  assign n32026 = n16549 & ~n32025 ;
  assign n32027 = n7547 & n12166 ;
  assign n32028 = n18102 ^ n4892 ^ 1'b0 ;
  assign n32029 = n12632 & n32028 ;
  assign n32030 = n5042 & n32029 ;
  assign n32031 = n32030 ^ n3853 ^ 1'b0 ;
  assign n32032 = n32027 & n32031 ;
  assign n32033 = n14873 | n21528 ;
  assign n32034 = n32033 ^ n13887 ^ 1'b0 ;
  assign n32035 = n6846 | n29712 ;
  assign n32036 = ~n32034 & n32035 ;
  assign n32037 = n4551 | n6551 ;
  assign n32038 = n32037 ^ n3305 ^ 1'b0 ;
  assign n32039 = n6827 | n17082 ;
  assign n32040 = n32039 ^ n10118 ^ 1'b0 ;
  assign n32041 = n32040 ^ n13603 ^ 1'b0 ;
  assign n32042 = n6885 & n17570 ;
  assign n32043 = n32042 ^ n5872 ^ 1'b0 ;
  assign n32044 = ~n131 & n26484 ;
  assign n32045 = ( n991 & n10816 ) | ( n991 & n28735 ) | ( n10816 & n28735 ) ;
  assign n32046 = n25257 ^ n6230 ^ 1'b0 ;
  assign n32047 = ~n32045 & n32046 ;
  assign n32048 = n32047 ^ n28202 ^ 1'b0 ;
  assign n32052 = n20169 & ~n29611 ;
  assign n32049 = n16861 & n30882 ;
  assign n32050 = ~n11446 & n32049 ;
  assign n32051 = n299 & ~n32050 ;
  assign n32053 = n32052 ^ n32051 ^ 1'b0 ;
  assign n32055 = n6147 & ~n24900 ;
  assign n32056 = n32055 ^ n6144 ^ 1'b0 ;
  assign n32054 = ( n3156 & ~n6703 ) | ( n3156 & n11438 ) | ( ~n6703 & n11438 ) ;
  assign n32057 = n32056 ^ n32054 ^ 1'b0 ;
  assign n32058 = n17652 ^ n2815 ^ 1'b0 ;
  assign n32059 = n3548 & n32058 ;
  assign n32060 = n10399 & n29335 ;
  assign n32061 = n32060 ^ n19996 ^ 1'b0 ;
  assign n32062 = n3218 | n13112 ;
  assign n32063 = n32062 ^ n12803 ^ 1'b0 ;
  assign n32064 = n6008 | n16983 ;
  assign n32065 = n32064 ^ n14476 ^ 1'b0 ;
  assign n32066 = ~n12081 & n15516 ;
  assign n32067 = n15993 ^ n12472 ^ 1'b0 ;
  assign n32068 = n30451 ^ n172 ^ 1'b0 ;
  assign n32070 = n9151 & n15537 ;
  assign n32069 = n2544 ^ n2278 ^ 1'b0 ;
  assign n32071 = n32070 ^ n32069 ^ 1'b0 ;
  assign n32072 = ~n2946 & n30608 ;
  assign n32073 = n32072 ^ n11154 ^ 1'b0 ;
  assign n32074 = n26220 ^ n9631 ^ 1'b0 ;
  assign n32075 = n10856 ^ n6847 ^ 1'b0 ;
  assign n32076 = ( n1733 & n26588 ) | ( n1733 & n32075 ) | ( n26588 & n32075 ) ;
  assign n32078 = n19672 ^ n3329 ^ 1'b0 ;
  assign n32077 = n5073 & ~n13137 ;
  assign n32079 = n32078 ^ n32077 ^ n20274 ;
  assign n32080 = n2882 | n26010 ;
  assign n32081 = n2882 & ~n32080 ;
  assign n32082 = n2752 | n7869 ;
  assign n32083 = n32081 & ~n32082 ;
  assign n32084 = n209 & n570 ;
  assign n32085 = ~n570 & n32084 ;
  assign n32086 = n6146 & n11480 ;
  assign n32087 = n32085 & n32086 ;
  assign n32088 = n2731 & ~n3500 ;
  assign n32089 = n32087 & n32088 ;
  assign n32090 = n32089 ^ n9241 ^ 1'b0 ;
  assign n32091 = n16616 & n32090 ;
  assign n32092 = n32083 & n32091 ;
  assign n32093 = n13785 & ~n22695 ;
  assign n32094 = n10991 ^ n6298 ^ 1'b0 ;
  assign n32095 = n23342 ^ n4667 ^ 1'b0 ;
  assign n32096 = n8234 ^ n1201 ^ n131 ;
  assign n32097 = n32096 ^ n27995 ^ 1'b0 ;
  assign n32098 = n7242 & n32097 ;
  assign n32099 = n22507 ^ n800 ^ 1'b0 ;
  assign n32100 = n3166 & ~n32099 ;
  assign n32101 = n28032 ^ n19742 ^ n14876 ;
  assign n32102 = n9796 ^ n2337 ^ 1'b0 ;
  assign n32103 = n25139 & n27237 ;
  assign n32104 = n23802 ^ n2561 ^ 1'b0 ;
  assign n32105 = n12854 | n32104 ;
  assign n32106 = n3826 & ~n15568 ;
  assign n32107 = n23014 ^ n9417 ^ 1'b0 ;
  assign n32108 = n32106 & n32107 ;
  assign n32109 = n26246 ^ n17109 ^ 1'b0 ;
  assign n32110 = ~n8604 & n32109 ;
  assign n32111 = n7004 & n32110 ;
  assign n32112 = n4410 | n10157 ;
  assign n32113 = n32112 ^ n17616 ^ 1'b0 ;
  assign n32114 = n22997 & ~n32113 ;
  assign n32115 = ~n3778 & n32114 ;
  assign n32116 = ( n458 & n919 ) | ( n458 & ~n1485 ) | ( n919 & ~n1485 ) ;
  assign n32117 = n7141 & n32116 ;
  assign n32118 = n32117 ^ n11653 ^ n7510 ;
  assign n32119 = ( n2845 & n6498 ) | ( n2845 & n19698 ) | ( n6498 & n19698 ) ;
  assign n32120 = n3823 & ~n20360 ;
  assign n32121 = ~n1216 & n32120 ;
  assign n32122 = n3084 ^ n220 ^ 1'b0 ;
  assign n32123 = n16969 & ~n22185 ;
  assign n32124 = n29927 ^ n12018 ^ 1'b0 ;
  assign n32125 = n604 & ~n10391 ;
  assign n32126 = n10962 & ~n21000 ;
  assign n32127 = ~n570 & n3060 ;
  assign n32128 = n5102 | n32127 ;
  assign n32129 = n18107 ^ n6915 ^ 1'b0 ;
  assign n32130 = ( ~n15839 & n32128 ) | ( ~n15839 & n32129 ) | ( n32128 & n32129 ) ;
  assign n32131 = ( ~n408 & n1800 ) | ( ~n408 & n14962 ) | ( n1800 & n14962 ) ;
  assign n32132 = ( n418 & n3290 ) | ( n418 & n5254 ) | ( n3290 & n5254 ) ;
  assign n32133 = ( n8806 & n32131 ) | ( n8806 & ~n32132 ) | ( n32131 & ~n32132 ) ;
  assign n32134 = n32133 ^ n17822 ^ 1'b0 ;
  assign n32135 = n108 | n32134 ;
  assign n32136 = n32135 ^ n8552 ^ 1'b0 ;
  assign n32137 = n29548 & ~n32136 ;
  assign n32138 = n32137 ^ n11269 ^ 1'b0 ;
  assign n32139 = n12810 & n21443 ;
  assign n32140 = n32139 ^ n26631 ^ 1'b0 ;
  assign n32141 = n6531 ^ n1395 ^ 1'b0 ;
  assign n32142 = n9635 | n32141 ;
  assign n32143 = n2135 & n23441 ;
  assign n32144 = ~n1151 & n26298 ;
  assign n32145 = n23766 & n32144 ;
  assign n32146 = n4200 | n18619 ;
  assign n32147 = ~n20199 & n32146 ;
  assign n32148 = n6119 ^ n3415 ^ 1'b0 ;
  assign n32149 = n11925 | n20444 ;
  assign n32150 = n32148 & ~n32149 ;
  assign n32151 = n24246 & n32150 ;
  assign n32152 = n8334 ^ n5124 ^ 1'b0 ;
  assign n32153 = n881 & n3750 ;
  assign n32154 = ~n289 & n32153 ;
  assign n32155 = ( n3754 & ~n10523 ) | ( n3754 & n15456 ) | ( ~n10523 & n15456 ) ;
  assign n32156 = n32155 ^ n3578 ^ 1'b0 ;
  assign n32157 = n11322 | n32156 ;
  assign n32158 = n6249 ^ n5965 ^ n3923 ;
  assign n32159 = ( n780 & ~n4226 ) | ( n780 & n32158 ) | ( ~n4226 & n32158 ) ;
  assign n32160 = n4725 | n21484 ;
  assign n32161 = n21148 ^ n4558 ^ n543 ;
  assign n32162 = n32160 & n32161 ;
  assign n32163 = n12692 ^ n7771 ^ n4463 ;
  assign n32164 = n30373 ^ n24212 ^ 1'b0 ;
  assign n32165 = ~n21990 & n32164 ;
  assign n32166 = n17614 ^ n9324 ^ 1'b0 ;
  assign n32167 = n32166 ^ n25151 ^ 1'b0 ;
  assign n32168 = n5098 & n32167 ;
  assign n32170 = n20563 ^ n20281 ^ n6423 ;
  assign n32169 = n22692 & n28761 ;
  assign n32171 = n32170 ^ n32169 ^ 1'b0 ;
  assign n32172 = n15777 ^ n12839 ^ 1'b0 ;
  assign n32173 = n32171 | n32172 ;
  assign n32174 = n28191 ^ n1820 ^ 1'b0 ;
  assign n32175 = n32174 ^ n12490 ^ 1'b0 ;
  assign n32176 = n32173 & ~n32175 ;
  assign n32177 = n25208 ^ n9973 ^ 1'b0 ;
  assign n32178 = n11114 & n32177 ;
  assign n32179 = n16440 ^ n15244 ^ 1'b0 ;
  assign n32180 = n22639 & n32179 ;
  assign n32181 = n32180 ^ n27998 ^ n16441 ;
  assign n32182 = n17952 ^ n6478 ^ 1'b0 ;
  assign n32183 = ~n3059 & n32182 ;
  assign n32184 = n32183 ^ n21393 ^ n5683 ;
  assign n32185 = n3312 | n23810 ;
  assign n32186 = ~n668 & n1704 ;
  assign n32187 = n12171 & n32186 ;
  assign n32188 = n3088 & n7037 ;
  assign n32189 = n11131 | n32188 ;
  assign n32190 = n32189 ^ n1754 ^ 1'b0 ;
  assign n32191 = n10960 & ~n32190 ;
  assign n32192 = ~n3636 & n17999 ;
  assign n32193 = n5493 & ~n32192 ;
  assign n32194 = ( n21895 & n32191 ) | ( n21895 & n32193 ) | ( n32191 & n32193 ) ;
  assign n32195 = ~n2560 & n4114 ;
  assign n32196 = n32195 ^ n22694 ^ 1'b0 ;
  assign n32197 = n10088 | n25297 ;
  assign n32198 = n17075 & ~n23217 ;
  assign n32199 = ( n3740 & n9167 ) | ( n3740 & n11656 ) | ( n9167 & n11656 ) ;
  assign n32200 = n30031 & n30406 ;
  assign n32201 = n11954 & ~n32200 ;
  assign n32202 = ( n10366 & n12585 ) | ( n10366 & n32201 ) | ( n12585 & n32201 ) ;
  assign n32203 = n32202 ^ n2967 ^ 1'b0 ;
  assign n32204 = ~n32199 & n32203 ;
  assign n32205 = ~n17534 & n31483 ;
  assign n32206 = n19393 | n32205 ;
  assign n32207 = n32206 ^ n3632 ^ 1'b0 ;
  assign n32208 = n5679 & ~n32207 ;
  assign n32209 = n32208 ^ n2619 ^ 1'b0 ;
  assign n32210 = n1517 & n6462 ;
  assign n32211 = ~n16635 & n20859 ;
  assign n32212 = n32211 ^ n2039 ^ 1'b0 ;
  assign n32213 = n32210 | n32212 ;
  assign n32214 = n15702 & ~n24405 ;
  assign n32215 = n18880 & n25078 ;
  assign n32216 = n32215 ^ n4132 ^ 1'b0 ;
  assign n32217 = n706 | n22726 ;
  assign n32218 = n25247 & ~n32217 ;
  assign n32219 = ~n15074 & n29423 ;
  assign n32220 = n32219 ^ n5115 ^ 1'b0 ;
  assign n32221 = n3053 | n17507 ;
  assign n32222 = n12668 & ~n20648 ;
  assign n32223 = n1276 & n32222 ;
  assign n32224 = n19102 | n20047 ;
  assign n32225 = n32224 ^ n22836 ^ n12263 ;
  assign n32230 = n5495 ^ n3161 ^ n1992 ;
  assign n32226 = n4911 & ~n9130 ;
  assign n32227 = n32226 ^ n2670 ^ 1'b0 ;
  assign n32228 = n32227 ^ n6408 ^ 1'b0 ;
  assign n32229 = n11197 | n32228 ;
  assign n32231 = n32230 ^ n32229 ^ n20668 ;
  assign n32232 = n16154 & ~n21217 ;
  assign n32233 = n32232 ^ n3744 ^ 1'b0 ;
  assign n32234 = n7262 ^ n3941 ^ 1'b0 ;
  assign n32235 = n6601 & n32234 ;
  assign n32236 = n21597 ^ n11518 ^ n3007 ;
  assign n32237 = n4439 & ~n13440 ;
  assign n32238 = n32237 ^ n2584 ^ 1'b0 ;
  assign n32239 = n27897 ^ n7976 ^ 1'b0 ;
  assign n32240 = n32239 ^ n11575 ^ 1'b0 ;
  assign n32241 = n1506 & n29859 ;
  assign n32242 = n32240 & n32241 ;
  assign n32243 = n5533 ^ n4082 ^ 1'b0 ;
  assign n32244 = n15585 & ~n32243 ;
  assign n32245 = n32244 ^ n4849 ^ n3175 ;
  assign n32246 = ~n603 & n1877 ;
  assign n32247 = n32246 ^ n11114 ^ 1'b0 ;
  assign n32248 = n11722 | n22976 ;
  assign n32249 = n1836 & ~n32248 ;
  assign n32250 = n30099 ^ n1175 ^ 1'b0 ;
  assign n32251 = n18342 & n32250 ;
  assign n32252 = ( n432 & n3532 ) | ( n432 & ~n21770 ) | ( n3532 & ~n21770 ) ;
  assign n32253 = n3351 | n14381 ;
  assign n32254 = n9005 & n32253 ;
  assign n32255 = n2076 & ~n23364 ;
  assign n32256 = n23960 ^ n10435 ^ n6539 ;
  assign n32257 = n24970 ^ n14557 ^ 1'b0 ;
  assign n32262 = n23908 & n24462 ;
  assign n32263 = n21596 | n32262 ;
  assign n32264 = n32263 ^ n7640 ^ 1'b0 ;
  assign n32259 = n16491 ^ n14425 ^ n2142 ;
  assign n32260 = n32259 ^ n16440 ^ 1'b0 ;
  assign n32261 = n6811 & n32260 ;
  assign n32265 = n32264 ^ n32261 ^ n1031 ;
  assign n32258 = ~n6225 & n24363 ;
  assign n32266 = n32265 ^ n32258 ^ 1'b0 ;
  assign n32267 = n32266 ^ n2352 ^ 1'b0 ;
  assign n32268 = n32257 & n32267 ;
  assign n32269 = n32256 & ~n32268 ;
  assign n32270 = n9780 | n10949 ;
  assign n32271 = ~n23966 & n32270 ;
  assign n32272 = n9162 & n28158 ;
  assign n32273 = n32272 ^ n19308 ^ 1'b0 ;
  assign n32274 = n2432 & ~n32273 ;
  assign n32275 = ( n13605 & n15194 ) | ( n13605 & n16925 ) | ( n15194 & n16925 ) ;
  assign n32276 = ( n408 & n5543 ) | ( n408 & n8218 ) | ( n5543 & n8218 ) ;
  assign n32277 = n17471 | n30350 ;
  assign n32278 = n17471 & ~n32277 ;
  assign n32279 = n32276 | n32278 ;
  assign n32280 = n32276 & ~n32279 ;
  assign n32281 = n30011 ^ n13062 ^ 1'b0 ;
  assign n32282 = n29774 | n32281 ;
  assign n32283 = n25747 ^ n10657 ^ n9578 ;
  assign n32284 = ~n25829 & n32283 ;
  assign n32285 = n32284 ^ n14757 ^ 1'b0 ;
  assign n32286 = n17844 & ~n32285 ;
  assign n32287 = n30888 ^ n16913 ^ n15246 ;
  assign n32290 = n29498 ^ n16837 ^ n10285 ;
  assign n32288 = n18680 ^ n9779 ^ 1'b0 ;
  assign n32289 = n32288 ^ n14981 ^ n4376 ;
  assign n32291 = n32290 ^ n32289 ^ 1'b0 ;
  assign n32292 = n27877 ^ n8584 ^ 1'b0 ;
  assign n32293 = ~n2937 & n9075 ;
  assign n32294 = n32293 ^ n14100 ^ 1'b0 ;
  assign n32295 = n9072 | n32294 ;
  assign n32296 = n15552 & n32295 ;
  assign n32297 = n32292 & n32296 ;
  assign n32298 = n21848 ^ n9402 ^ 1'b0 ;
  assign n32299 = n5418 ^ n261 ^ 1'b0 ;
  assign n32300 = n15316 ^ n712 ^ 1'b0 ;
  assign n32301 = n10117 & n12317 ;
  assign n32302 = n32301 ^ n1526 ^ 1'b0 ;
  assign n32303 = n2558 & n6596 ;
  assign n32304 = ( ~n11581 & n18428 ) | ( ~n11581 & n32303 ) | ( n18428 & n32303 ) ;
  assign n32305 = n29047 & n30521 ;
  assign n32306 = n30219 ^ n8847 ^ 1'b0 ;
  assign n32307 = n13400 ^ n4903 ^ 1'b0 ;
  assign n32308 = n5634 | n32307 ;
  assign n32309 = n32308 ^ n12787 ^ 1'b0 ;
  assign n32310 = n2609 | n32309 ;
  assign n32311 = n32310 ^ n6181 ^ 1'b0 ;
  assign n32312 = n3630 | n32311 ;
  assign n32313 = n32306 & ~n32312 ;
  assign n32314 = n9184 | n27854 ;
  assign n32315 = n7473 & ~n32314 ;
  assign n32316 = n2836 & n3133 ;
  assign n32318 = ~n6620 & n8939 ;
  assign n32319 = ~n8606 & n32318 ;
  assign n32317 = n2297 | n9528 ;
  assign n32320 = n32319 ^ n32317 ^ 1'b0 ;
  assign n32321 = n22372 ^ n15993 ^ 1'b0 ;
  assign n32322 = n4710 ^ n575 ^ 1'b0 ;
  assign n32323 = n9933 & n32322 ;
  assign n32324 = ( n15811 & ~n23801 ) | ( n15811 & n32323 ) | ( ~n23801 & n32323 ) ;
  assign n32325 = n2225 | n32324 ;
  assign n32326 = n2676 & ~n32325 ;
  assign n32327 = ~n2427 & n24482 ;
  assign n32328 = n12723 | n32327 ;
  assign n32329 = n32328 ^ n19965 ^ n853 ;
  assign n32331 = n18389 ^ n10441 ^ 1'b0 ;
  assign n32332 = n12159 ^ n9184 ^ 1'b0 ;
  assign n32333 = n13073 | n32332 ;
  assign n32334 = ( n22061 & ~n32331 ) | ( n22061 & n32333 ) | ( ~n32331 & n32333 ) ;
  assign n32335 = n32334 ^ n24485 ^ 1'b0 ;
  assign n32336 = ~n10118 & n32335 ;
  assign n32330 = ( n4990 & n8552 ) | ( n4990 & n14023 ) | ( n8552 & n14023 ) ;
  assign n32337 = n32336 ^ n32330 ^ n29537 ;
  assign n32340 = ~x3 & n9041 ;
  assign n32341 = n99 & n32340 ;
  assign n32338 = n8721 & n19182 ;
  assign n32339 = n32338 ^ n19269 ^ 1'b0 ;
  assign n32342 = n32341 ^ n32339 ^ 1'b0 ;
  assign n32343 = n28714 ^ n21571 ^ 1'b0 ;
  assign n32344 = ~n147 & n32343 ;
  assign n32345 = n32344 ^ n28470 ^ 1'b0 ;
  assign n32346 = n5099 & n14872 ;
  assign n32347 = n32346 ^ n9195 ^ 1'b0 ;
  assign n32348 = n31500 ^ n12128 ^ 1'b0 ;
  assign n32349 = ~n25540 & n32348 ;
  assign n32350 = ~n5554 & n32349 ;
  assign n32352 = ~n7149 & n32112 ;
  assign n32353 = ( n6356 & n31415 ) | ( n6356 & ~n32352 ) | ( n31415 & ~n32352 ) ;
  assign n32351 = n20226 | n28026 ;
  assign n32354 = n32353 ^ n32351 ^ 1'b0 ;
  assign n32355 = n12206 ^ n10998 ^ 1'b0 ;
  assign n32356 = n8856 ^ n5707 ^ 1'b0 ;
  assign n32357 = n32355 | n32356 ;
  assign n32358 = n10379 | n32357 ;
  assign n32359 = n32358 ^ n26156 ^ n18176 ;
  assign n32360 = n18223 | n32359 ;
  assign n32361 = n32360 ^ n6115 ^ 1'b0 ;
  assign n32362 = n875 & n18729 ;
  assign n32363 = ~n2484 & n8824 ;
  assign n32364 = n32363 ^ n726 ^ 1'b0 ;
  assign n32365 = ~n5672 & n32364 ;
  assign n32366 = n19364 ^ n2203 ^ 1'b0 ;
  assign n32367 = n23200 ^ n8493 ^ 1'b0 ;
  assign n32369 = n3326 ^ n1232 ^ 1'b0 ;
  assign n32368 = ~n884 & n14991 ;
  assign n32370 = n32369 ^ n32368 ^ 1'b0 ;
  assign n32371 = n32370 ^ n3153 ^ 1'b0 ;
  assign n32372 = ~n32367 & n32371 ;
  assign n32373 = n15353 & n24684 ;
  assign n32374 = n19322 ^ n6851 ^ 1'b0 ;
  assign n32375 = n7641 ^ n6667 ^ 1'b0 ;
  assign n32376 = n23975 | n32375 ;
  assign n32377 = n15380 ^ n11429 ^ 1'b0 ;
  assign n32378 = n32376 & n32377 ;
  assign n32381 = n23025 ^ n3271 ^ 1'b0 ;
  assign n32382 = ~n15249 & n32381 ;
  assign n32379 = ~n9533 & n17809 ;
  assign n32380 = ~n17809 & n32379 ;
  assign n32383 = n32382 ^ n32380 ^ 1'b0 ;
  assign n32384 = n32383 ^ n7622 ^ 1'b0 ;
  assign n32385 = n640 | n21307 ;
  assign n32386 = n450 & ~n2074 ;
  assign n32387 = n2916 & n8294 ;
  assign n32388 = ~n25795 & n32387 ;
  assign n32389 = n32388 ^ n15350 ^ 1'b0 ;
  assign n32390 = n23606 ^ n15271 ^ n5676 ;
  assign n32391 = n32390 ^ n13045 ^ 1'b0 ;
  assign n32392 = n26421 | n32391 ;
  assign n32393 = n5144 & n7276 ;
  assign n32394 = ~n4044 & n32393 ;
  assign n32395 = ~n18251 & n32394 ;
  assign n32396 = n7134 ^ n3256 ^ 1'b0 ;
  assign n32397 = n32396 ^ n24187 ^ 1'b0 ;
  assign n32398 = n6229 & n32397 ;
  assign n32399 = n32398 ^ n29385 ^ 1'b0 ;
  assign n32400 = ~n7074 & n31129 ;
  assign n32401 = n15759 & ~n32400 ;
  assign n32402 = ~n10779 & n32401 ;
  assign n32403 = n4010 & ~n7060 ;
  assign n32404 = n32403 ^ n30885 ^ 1'b0 ;
  assign n32405 = ( ~n7494 & n12923 ) | ( ~n7494 & n21997 ) | ( n12923 & n21997 ) ;
  assign n32410 = n17818 ^ n10697 ^ 1'b0 ;
  assign n32408 = ( n3122 & n3817 ) | ( n3122 & ~n4120 ) | ( n3817 & ~n4120 ) ;
  assign n32409 = ( n6149 & n9849 ) | ( n6149 & n32408 ) | ( n9849 & n32408 ) ;
  assign n32406 = n9258 ^ n5357 ^ 1'b0 ;
  assign n32407 = n7832 & n32406 ;
  assign n32411 = n32410 ^ n32409 ^ n32407 ;
  assign n32412 = ~n44 & n7605 ;
  assign n32413 = ~n12500 & n32412 ;
  assign n32414 = n32413 ^ n3238 ^ 1'b0 ;
  assign n32415 = n11418 & n32414 ;
  assign n32416 = ( n16652 & ~n21254 ) | ( n16652 & n32415 ) | ( ~n21254 & n32415 ) ;
  assign n32417 = ~n5806 & n26096 ;
  assign n32418 = ~n2306 & n12413 ;
  assign n32419 = n32418 ^ n12357 ^ 1'b0 ;
  assign n32420 = n32419 ^ n8074 ^ 1'b0 ;
  assign n32421 = ~n32417 & n32420 ;
  assign n32422 = n19613 ^ n1716 ^ 1'b0 ;
  assign n32423 = n2322 & n31116 ;
  assign n32424 = n10381 & ~n27410 ;
  assign n32425 = n32424 ^ n1190 ^ 1'b0 ;
  assign n32426 = n17813 ^ n5433 ^ n5270 ;
  assign n32427 = n32426 ^ n15040 ^ n9975 ;
  assign n32428 = n24754 ^ n11628 ^ 1'b0 ;
  assign n32429 = ~n4211 & n5503 ;
  assign n32430 = n17805 & ~n32429 ;
  assign n32431 = n32430 ^ n2819 ^ 1'b0 ;
  assign n32432 = n20897 & n25560 ;
  assign n32433 = n32432 ^ n12875 ^ 1'b0 ;
  assign n32434 = ~n32431 & n32433 ;
  assign n32435 = n24355 & n32434 ;
  assign n32436 = n32428 & n32435 ;
  assign n32437 = n29801 ^ n1162 ^ 1'b0 ;
  assign n32438 = n17520 ^ n17020 ^ n8143 ;
  assign n32439 = ~n28070 & n32438 ;
  assign n32440 = ~n5996 & n24844 ;
  assign n32441 = n32440 ^ n27594 ^ 1'b0 ;
  assign n32442 = n185 | n7481 ;
  assign n32443 = n1131 & ~n28138 ;
  assign n32444 = ~n5861 & n32443 ;
  assign n32445 = n8260 & ~n32444 ;
  assign n32446 = n32442 & n32445 ;
  assign n32447 = n2678 | n6686 ;
  assign n32448 = ( ~n18080 & n30431 ) | ( ~n18080 & n32447 ) | ( n30431 & n32447 ) ;
  assign n32449 = ( ~n3115 & n19207 ) | ( ~n3115 & n21940 ) | ( n19207 & n21940 ) ;
  assign n32450 = n3395 & n23762 ;
  assign n32451 = n32450 ^ n221 ^ 1'b0 ;
  assign n32452 = n25281 ^ n22464 ^ 1'b0 ;
  assign n32453 = ~n1848 & n17085 ;
  assign n32454 = n30033 ^ n3070 ^ 1'b0 ;
  assign n32456 = n8115 ^ n6330 ^ 1'b0 ;
  assign n32455 = n3769 | n22806 ;
  assign n32457 = n32456 ^ n32455 ^ 1'b0 ;
  assign n32458 = n32457 ^ n21808 ^ 1'b0 ;
  assign n32459 = n10328 & ~n11573 ;
  assign n32460 = n21569 ^ n20153 ^ 1'b0 ;
  assign n32461 = n20896 | n32460 ;
  assign n32463 = n9929 ^ n8029 ^ 1'b0 ;
  assign n32464 = ~n13943 & n32463 ;
  assign n32465 = n32464 ^ n9887 ^ 1'b0 ;
  assign n32462 = n6107 & ~n17478 ;
  assign n32466 = n32465 ^ n32462 ^ 1'b0 ;
  assign n32473 = ( n1234 & ~n5652 ) | ( n1234 & n19456 ) | ( ~n5652 & n19456 ) ;
  assign n32467 = ~n3962 & n22605 ;
  assign n32468 = n32467 ^ n10187 ^ 1'b0 ;
  assign n32469 = n15895 & ~n32468 ;
  assign n32470 = n5880 & n32469 ;
  assign n32471 = n37 & ~n32470 ;
  assign n32472 = n2808 & n32471 ;
  assign n32474 = n32473 ^ n32472 ^ n30260 ;
  assign n32475 = n22669 ^ n13995 ^ n1746 ;
  assign n32476 = n13963 & n32475 ;
  assign n32477 = n9658 & n24068 ;
  assign n32478 = n6451 & n32477 ;
  assign n32479 = n1586 & n10016 ;
  assign n32480 = n22559 & ~n30806 ;
  assign n32481 = n32480 ^ n31239 ^ 1'b0 ;
  assign n32482 = n22918 ^ n21107 ^ 1'b0 ;
  assign n32484 = n734 & n17752 ;
  assign n32485 = n8445 & n32484 ;
  assign n32483 = n7059 | n7216 ;
  assign n32486 = n32485 ^ n32483 ^ 1'b0 ;
  assign n32487 = n32482 & ~n32486 ;
  assign n32488 = ~n32482 & n32487 ;
  assign n32489 = n28140 ^ n3111 ^ 1'b0 ;
  assign n32490 = ~n6226 & n17753 ;
  assign n32491 = n20317 ^ n9805 ^ 1'b0 ;
  assign n32492 = n14236 & ~n32491 ;
  assign n32493 = ~n32490 & n32492 ;
  assign n32494 = n9476 & n32493 ;
  assign n32495 = n5704 ^ n4851 ^ n4146 ;
  assign n32496 = n32495 ^ n14875 ^ 1'b0 ;
  assign n32497 = ~n11546 & n17324 ;
  assign n32498 = n32497 ^ n15349 ^ 1'b0 ;
  assign n32499 = n11542 | n32498 ;
  assign n32500 = n32499 ^ n11751 ^ 1'b0 ;
  assign n32501 = n15552 ^ n10393 ^ 1'b0 ;
  assign n32502 = n32501 ^ n9309 ^ n471 ;
  assign n32503 = n10352 & ~n26611 ;
  assign n32504 = n18023 ^ n8608 ^ 1'b0 ;
  assign n32505 = n32503 | n32504 ;
  assign n32506 = ~n4280 & n19341 ;
  assign n32507 = n20351 ^ n7920 ^ 1'b0 ;
  assign n32508 = n9281 | n32507 ;
  assign n32509 = n32508 ^ n20924 ^ n9446 ;
  assign n32510 = n10719 & ~n32509 ;
  assign n32511 = n1326 | n13554 ;
  assign n32512 = n12335 ^ n5225 ^ 1'b0 ;
  assign n32513 = ~n17747 & n32512 ;
  assign n32514 = ~n4275 & n9168 ;
  assign n32515 = n4257 & n16590 ;
  assign n32516 = n28457 ^ n7153 ^ 1'b0 ;
  assign n32517 = ~n51 & n1890 ;
  assign n32518 = n32179 | n32517 ;
  assign n32519 = n29660 | n32518 ;
  assign n32520 = n32519 ^ n4232 ^ 1'b0 ;
  assign n32526 = n19976 ^ n17954 ^ 1'b0 ;
  assign n32527 = ~n3908 & n32526 ;
  assign n32521 = n1004 & n12506 ;
  assign n32522 = ~n14670 & n32521 ;
  assign n32523 = ~n32521 & n32522 ;
  assign n32524 = n32523 ^ n22243 ^ 1'b0 ;
  assign n32525 = ~n15576 & n32524 ;
  assign n32528 = n32527 ^ n32525 ^ 1'b0 ;
  assign n32529 = n6322 | n21361 ;
  assign n32530 = n16138 & ~n32529 ;
  assign n32531 = n11114 & ~n32530 ;
  assign n32532 = n10919 & n32531 ;
  assign n32533 = n32532 ^ n10348 ^ 1'b0 ;
  assign n32534 = ~n19924 & n32533 ;
  assign n32535 = n32534 ^ n11065 ^ 1'b0 ;
  assign n32536 = ( n953 & n1201 ) | ( n953 & n3242 ) | ( n1201 & n3242 ) ;
  assign n32537 = n10264 ^ n7058 ^ n6682 ;
  assign n32538 = n32014 | n32537 ;
  assign n32539 = ~n19342 & n19541 ;
  assign n32540 = n30866 ^ n11921 ^ n2060 ;
  assign n32541 = n10952 | n31520 ;
  assign n32542 = n19917 | n32541 ;
  assign n32543 = ~n10951 & n17276 ;
  assign n32544 = n15401 & n32543 ;
  assign n32545 = ( ~n628 & n13112 ) | ( ~n628 & n32544 ) | ( n13112 & n32544 ) ;
  assign n32546 = n32542 | n32545 ;
  assign n32547 = n23937 & n26778 ;
  assign n32548 = n7361 | n24240 ;
  assign n32549 = n32548 ^ n4404 ^ 1'b0 ;
  assign n32550 = n6014 | n10888 ;
  assign n32551 = n4977 | n32550 ;
  assign n32552 = ~n6451 & n18820 ;
  assign n32553 = ~n18587 & n32552 ;
  assign n32554 = n7227 | n13276 ;
  assign n32555 = ~n20896 & n32554 ;
  assign n32556 = ( n25163 & n32553 ) | ( n25163 & n32555 ) | ( n32553 & n32555 ) ;
  assign n32557 = n18758 | n27321 ;
  assign n32558 = n6890 & ~n10792 ;
  assign n32559 = n23729 ^ n1706 ^ 1'b0 ;
  assign n32560 = n24756 ^ n22393 ^ n11904 ;
  assign n32561 = n18586 | n19574 ;
  assign n32562 = ~n3744 & n25016 ;
  assign n32563 = n6902 | n26674 ;
  assign n32564 = n19650 & ~n32563 ;
  assign n32565 = n3712 & n21818 ;
  assign n32566 = n32565 ^ n13162 ^ 1'b0 ;
  assign n32567 = n4019 & ~n32566 ;
  assign n32568 = n32567 ^ n6365 ^ n2566 ;
  assign n32569 = ~n8526 & n18465 ;
  assign n32570 = n32569 ^ n184 ^ 1'b0 ;
  assign n32571 = n1762 & ~n32570 ;
  assign n32572 = n722 | n11676 ;
  assign n32573 = n6579 | n32572 ;
  assign n32574 = ( n3816 & n5845 ) | ( n3816 & ~n10583 ) | ( n5845 & ~n10583 ) ;
  assign n32575 = n16347 ^ n9122 ^ 1'b0 ;
  assign n32576 = n32574 & ~n32575 ;
  assign n32577 = ~n15180 & n32576 ;
  assign n32578 = ~n32573 & n32577 ;
  assign n32583 = n188 & n4663 ;
  assign n32584 = ~n32183 & n32583 ;
  assign n32585 = n32584 ^ n846 ^ 1'b0 ;
  assign n32586 = n13331 ^ n1628 ^ 1'b0 ;
  assign n32587 = n32585 & ~n32586 ;
  assign n32580 = ~n5975 & n7114 ;
  assign n32579 = n24157 ^ n8793 ^ n3671 ;
  assign n32581 = n32580 ^ n32579 ^ n12449 ;
  assign n32582 = n31170 & ~n32581 ;
  assign n32588 = n32587 ^ n32582 ^ 1'b0 ;
  assign n32589 = ~n5366 & n10638 ;
  assign n32590 = n24961 ^ n3505 ^ 1'b0 ;
  assign n32591 = n3607 & ~n28953 ;
  assign n32592 = n32591 ^ n12731 ^ 1'b0 ;
  assign n32593 = n26453 ^ n5797 ^ 1'b0 ;
  assign n32594 = n14112 & ~n31543 ;
  assign n32595 = n696 & ~n4966 ;
  assign n32596 = n32595 ^ n15955 ^ 1'b0 ;
  assign n32597 = n7140 & ~n13965 ;
  assign n32598 = n14737 | n29591 ;
  assign n32599 = n32597 | n32598 ;
  assign n32600 = ~n18688 & n27952 ;
  assign n32601 = n32600 ^ n30083 ^ 1'b0 ;
  assign n32602 = n6198 & n8830 ;
  assign n32603 = n513 | n32602 ;
  assign n32604 = n2022 | n32603 ;
  assign n32605 = n7977 | n31536 ;
  assign n32606 = n4629 | n32605 ;
  assign n32607 = n32606 ^ n3662 ^ 1'b0 ;
  assign n32608 = n11197 & ~n24110 ;
  assign n32609 = n32608 ^ n25421 ^ n12283 ;
  assign n32610 = n11813 & n19662 ;
  assign n32611 = n32610 ^ n18849 ^ n12755 ;
  assign n32612 = n6877 & n22776 ;
  assign n32615 = n22253 ^ n18383 ^ 1'b0 ;
  assign n32616 = n28618 | n32615 ;
  assign n32613 = n16864 & ~n21202 ;
  assign n32614 = n6739 | n32613 ;
  assign n32617 = n32616 ^ n32614 ^ 1'b0 ;
  assign n32618 = n2321 | n6294 ;
  assign n32619 = n32618 ^ n7419 ^ 1'b0 ;
  assign n32620 = n32619 ^ n12574 ^ 1'b0 ;
  assign n32621 = n1192 & n3968 ;
  assign n32622 = n32621 ^ n32180 ^ 1'b0 ;
  assign n32623 = ~n8690 & n9539 ;
  assign n32624 = n236 & n9895 ;
  assign n32625 = n32624 ^ n13934 ^ 1'b0 ;
  assign n32626 = n32623 | n32625 ;
  assign n32627 = n14786 | n32626 ;
  assign n32628 = ~n1709 & n13823 ;
  assign n32629 = n15700 ^ n9313 ^ 1'b0 ;
  assign n32630 = ~n16103 & n32629 ;
  assign n32632 = n2070 & ~n18784 ;
  assign n32633 = n32632 ^ n14350 ^ 1'b0 ;
  assign n32631 = n11505 | n32023 ;
  assign n32634 = n32633 ^ n32631 ^ 1'b0 ;
  assign n32635 = n6518 ^ n4204 ^ 1'b0 ;
  assign n32636 = ( n6114 & ~n18619 ) | ( n6114 & n32635 ) | ( ~n18619 & n32635 ) ;
  assign n32637 = n12010 ^ n4668 ^ n1287 ;
  assign n32638 = n25736 ^ n14771 ^ 1'b0 ;
  assign n32639 = n25921 & ~n32638 ;
  assign n32640 = n15788 ^ n10676 ^ 1'b0 ;
  assign n32641 = n32639 & n32640 ;
  assign n32642 = n7943 & n14583 ;
  assign n32643 = ~n615 & n32642 ;
  assign n32644 = n32643 ^ n21803 ^ n7055 ;
  assign n32645 = n26465 ^ n17659 ^ 1'b0 ;
  assign n32646 = n32645 ^ n19149 ^ n12611 ;
  assign n32647 = ~n3573 & n10360 ;
  assign n32648 = n13019 & n31213 ;
  assign n32649 = n32648 ^ n20835 ^ 1'b0 ;
  assign n32650 = ( n845 & ~n3491 ) | ( n845 & n21624 ) | ( ~n3491 & n21624 ) ;
  assign n32651 = ~n4153 & n11698 ;
  assign n32652 = n32651 ^ n16168 ^ 1'b0 ;
  assign n32653 = n32650 & ~n32652 ;
  assign n32654 = n2818 ^ n2428 ^ 1'b0 ;
  assign n32655 = n29789 & ~n32654 ;
  assign n32656 = n6377 | n23872 ;
  assign n32657 = n15083 & n32656 ;
  assign n32658 = n32657 ^ n22735 ^ 1'b0 ;
  assign n32659 = n29256 & ~n29948 ;
  assign n32660 = n32659 ^ n24260 ^ 1'b0 ;
  assign n32661 = n4767 | n7757 ;
  assign n32662 = n15406 | n32661 ;
  assign n32663 = n32660 | n32662 ;
  assign n32664 = n21724 ^ n14768 ^ 1'b0 ;
  assign n32666 = n688 | n31220 ;
  assign n32667 = n32666 ^ n7407 ^ n3457 ;
  assign n32665 = n12679 | n16935 ;
  assign n32668 = n32667 ^ n32665 ^ 1'b0 ;
  assign n32669 = n28984 | n32668 ;
  assign n32670 = n11717 & ~n32669 ;
  assign n32671 = ~n2047 & n3949 ;
  assign n32672 = ( n13479 & ~n20614 ) | ( n13479 & n32671 ) | ( ~n20614 & n32671 ) ;
  assign n32673 = n4773 | n24389 ;
  assign n32674 = n32673 ^ n9160 ^ 1'b0 ;
  assign n32675 = n16251 ^ n3626 ^ n1772 ;
  assign n32676 = n32675 ^ n11805 ^ 1'b0 ;
  assign n32677 = n29450 & ~n32676 ;
  assign n32678 = n15269 & n17653 ;
  assign n32679 = n32678 ^ n20576 ^ n9877 ;
  assign n32683 = n301 & n12302 ;
  assign n32684 = n32683 ^ n9773 ^ 1'b0 ;
  assign n32685 = n32684 ^ n8516 ^ 1'b0 ;
  assign n32686 = n13112 | n32685 ;
  assign n32687 = n32686 ^ n17985 ^ 1'b0 ;
  assign n32688 = ~n5936 & n32687 ;
  assign n32680 = n1073 & ~n9497 ;
  assign n32681 = n823 & n32680 ;
  assign n32682 = ~n14450 & n32681 ;
  assign n32689 = n32688 ^ n32682 ^ 1'b0 ;
  assign n32690 = ( n672 & n885 ) | ( n672 & n32689 ) | ( n885 & n32689 ) ;
  assign n32691 = n7112 | n10720 ;
  assign n32694 = n23401 & ~n30918 ;
  assign n32695 = n8774 & n32694 ;
  assign n32696 = n32695 ^ n19996 ^ n3195 ;
  assign n32692 = n3564 | n17100 ;
  assign n32693 = n25155 & n32692 ;
  assign n32697 = n32696 ^ n32693 ^ n2569 ;
  assign n32698 = n4750 | n9110 ;
  assign n32699 = n7646 ^ n6386 ^ 1'b0 ;
  assign n32700 = ~n32698 & n32699 ;
  assign n32701 = n32700 ^ n3532 ^ 1'b0 ;
  assign n32702 = n24658 & ~n32701 ;
  assign n32703 = n32702 ^ n2157 ^ 1'b0 ;
  assign n32704 = ~n19513 & n32703 ;
  assign n32705 = ~n29897 & n32704 ;
  assign n32706 = n18894 ^ n10252 ^ 1'b0 ;
  assign n32707 = n17039 | n32706 ;
  assign n32708 = ( ~n145 & n22506 ) | ( ~n145 & n32707 ) | ( n22506 & n32707 ) ;
  assign n32709 = n752 & n5189 ;
  assign n32710 = ( n8703 & n10382 ) | ( n8703 & n17525 ) | ( n10382 & n17525 ) ;
  assign n32711 = n18770 & ~n32710 ;
  assign n32712 = n32711 ^ n15421 ^ 1'b0 ;
  assign n32713 = n18264 | n32712 ;
  assign n32714 = n21345 ^ n2327 ^ 1'b0 ;
  assign n32715 = n19714 & n20458 ;
  assign n32716 = n570 & n23168 ;
  assign n32717 = n32716 ^ n23870 ^ 1'b0 ;
  assign n32718 = n7644 & ~n32717 ;
  assign n32719 = n32715 & n32718 ;
  assign n32720 = n283 & ~n25482 ;
  assign n32721 = n7927 | n18451 ;
  assign n32722 = n32720 & ~n32721 ;
  assign n32723 = ~n2422 & n18853 ;
  assign n32724 = n32723 ^ n9481 ^ 1'b0 ;
  assign n32725 = ( n1444 & n17080 ) | ( n1444 & ~n17966 ) | ( n17080 & ~n17966 ) ;
  assign n32726 = n22576 & n30667 ;
  assign n32728 = ~n3479 & n11852 ;
  assign n32727 = n1729 & ~n31689 ;
  assign n32729 = n32728 ^ n32727 ^ 1'b0 ;
  assign n32731 = ~n7243 & n30729 ;
  assign n32732 = n17420 & n25682 ;
  assign n32733 = ~n32731 & n32732 ;
  assign n32730 = ~n2389 & n13210 ;
  assign n32734 = n32733 ^ n32730 ^ 1'b0 ;
  assign n32735 = n24193 | n25479 ;
  assign n32736 = n27761 ^ n7551 ^ 1'b0 ;
  assign n32737 = ~n22420 & n32736 ;
  assign n32738 = n17948 & ~n28301 ;
  assign n32739 = n12925 | n23765 ;
  assign n32740 = n32739 ^ n31809 ^ 1'b0 ;
  assign n32741 = n9787 | n11917 ;
  assign n32742 = n32741 ^ n1348 ^ 1'b0 ;
  assign n32743 = ~n4852 & n32742 ;
  assign n32744 = n580 & n2986 ;
  assign n32745 = n32743 & n32744 ;
  assign n32746 = n24022 ^ n22536 ^ n16025 ;
  assign n32747 = n31912 & n32746 ;
  assign n32748 = n20334 & n32747 ;
  assign n32749 = n22419 ^ n1632 ^ 1'b0 ;
  assign n32750 = n30851 ^ n8500 ^ 1'b0 ;
  assign n32751 = n15375 | n32750 ;
  assign n32752 = n15876 & ~n32751 ;
  assign n32753 = ( n2284 & n3014 ) | ( n2284 & n5261 ) | ( n3014 & n5261 ) ;
  assign n32754 = n779 & ~n2131 ;
  assign n32755 = n19976 & n32754 ;
  assign n32756 = n25890 & n32755 ;
  assign n32757 = n13848 ^ n11544 ^ 1'b0 ;
  assign n32758 = n25807 & ~n32757 ;
  assign n32761 = n8537 ^ n5654 ^ 1'b0 ;
  assign n32759 = n32438 ^ n11952 ^ n9721 ;
  assign n32760 = n14218 | n32759 ;
  assign n32762 = n32761 ^ n32760 ^ 1'b0 ;
  assign n32763 = n32762 ^ n28589 ^ n3084 ;
  assign n32764 = ( n18509 & n23469 ) | ( n18509 & ~n27995 ) | ( n23469 & ~n27995 ) ;
  assign n32765 = n30517 ^ n5627 ^ 1'b0 ;
  assign n32766 = n28529 & n32765 ;
  assign n32767 = n18707 ^ n7062 ^ 1'b0 ;
  assign n32768 = n32056 ^ n7958 ^ 1'b0 ;
  assign n32769 = n7998 | n9011 ;
  assign n32770 = n5834 & ~n32769 ;
  assign n32771 = ~n6227 & n22442 ;
  assign n32772 = n32771 ^ n7020 ^ 1'b0 ;
  assign n32773 = ~n33 & n23922 ;
  assign n32774 = n8780 & n32773 ;
  assign n32775 = n32774 ^ n25187 ^ 1'b0 ;
  assign n32776 = n55 | n9213 ;
  assign n32777 = n32776 ^ n1974 ^ 1'b0 ;
  assign n32778 = n55 | n1311 ;
  assign n32779 = ~n24308 & n32778 ;
  assign n32780 = n9956 ^ n3181 ^ 1'b0 ;
  assign n32781 = n10339 | n32780 ;
  assign n32782 = ~n734 & n32781 ;
  assign n32783 = ( n32777 & ~n32779 ) | ( n32777 & n32782 ) | ( ~n32779 & n32782 ) ;
  assign n32784 = ~n6993 & n23120 ;
  assign n32785 = n5747 ^ n3755 ^ 1'b0 ;
  assign n32786 = n14255 ^ n2350 ^ 1'b0 ;
  assign n32787 = n14756 | n32786 ;
  assign n32788 = n10292 | n19533 ;
  assign n32789 = ( ~n3959 & n17484 ) | ( ~n3959 & n32788 ) | ( n17484 & n32788 ) ;
  assign n32796 = n15709 ^ n1312 ^ 1'b0 ;
  assign n32793 = ~n5822 & n11006 ;
  assign n32794 = n1841 & n32793 ;
  assign n32795 = ( ~n10056 & n15504 ) | ( ~n10056 & n32794 ) | ( n15504 & n32794 ) ;
  assign n32790 = n13586 ^ n8860 ^ 1'b0 ;
  assign n32791 = n16473 ^ n7977 ^ 1'b0 ;
  assign n32792 = n32790 | n32791 ;
  assign n32797 = n32796 ^ n32795 ^ n32792 ;
  assign n32798 = n9226 & ~n27277 ;
  assign n32799 = n20778 ^ n18240 ^ n12758 ;
  assign n32800 = n14207 ^ n5908 ^ 1'b0 ;
  assign n32801 = n16664 & n32800 ;
  assign n32802 = n29492 ^ n2507 ^ 1'b0 ;
  assign n32803 = n32801 & ~n32802 ;
  assign n32804 = n11497 & n32803 ;
  assign n32805 = n32804 ^ n18408 ^ 1'b0 ;
  assign n32806 = ~n4730 & n5399 ;
  assign n32807 = ~n18404 & n26369 ;
  assign n32808 = n32807 ^ n32795 ^ n15728 ;
  assign n32809 = n20007 & ~n32808 ;
  assign n32810 = x0 & ~n23824 ;
  assign n32811 = ~n3430 & n21570 ;
  assign n32813 = n3685 & ~n10630 ;
  assign n32814 = n32813 ^ n3146 ^ 1'b0 ;
  assign n32815 = ~n8691 & n32814 ;
  assign n32812 = n10664 & n15259 ;
  assign n32816 = n32815 ^ n32812 ^ 1'b0 ;
  assign n32817 = ~n1437 & n29716 ;
  assign n32818 = n17311 ^ n14771 ^ n9208 ;
  assign n32819 = n32817 & ~n32818 ;
  assign n32820 = ~n7596 & n18723 ;
  assign n32821 = n26910 | n32820 ;
  assign n32826 = n11060 & n23531 ;
  assign n32827 = n12363 | n32826 ;
  assign n32822 = n376 | n15041 ;
  assign n32823 = n32822 ^ n3461 ^ 1'b0 ;
  assign n32824 = n11993 & ~n32823 ;
  assign n32825 = n10133 & n32824 ;
  assign n32828 = n32827 ^ n32825 ^ 1'b0 ;
  assign n32829 = ~n32821 & n32828 ;
  assign n32830 = ~n1100 & n32829 ;
  assign n32831 = n32830 ^ n19244 ^ 1'b0 ;
  assign n32832 = n22363 ^ n11564 ^ 1'b0 ;
  assign n32833 = n32831 & n32832 ;
  assign n32834 = n27967 & n32833 ;
  assign n32835 = ( n4338 & n10956 ) | ( n4338 & n17050 ) | ( n10956 & n17050 ) ;
  assign n32836 = n709 | n2695 ;
  assign n32837 = n2695 & ~n32836 ;
  assign n32838 = ~n4785 & n32837 ;
  assign n32839 = ( n30029 & ~n31102 ) | ( n30029 & n32838 ) | ( ~n31102 & n32838 ) ;
  assign n32840 = n11238 ^ n647 ^ 1'b0 ;
  assign n32841 = n29154 & n32840 ;
  assign n32842 = n9659 & n17490 ;
  assign n32843 = ~n8150 & n16794 ;
  assign n32844 = n32843 ^ n10233 ^ 1'b0 ;
  assign n32845 = n16189 ^ n15761 ^ n12734 ;
  assign n32846 = n32845 ^ n17548 ^ 1'b0 ;
  assign n32847 = n19034 ^ n18150 ^ n7636 ;
  assign n32848 = ( n5910 & n11510 ) | ( n5910 & ~n32847 ) | ( n11510 & ~n32847 ) ;
  assign n32849 = ~n24383 & n32848 ;
  assign n32850 = n6299 & ~n10066 ;
  assign n32851 = ~n3263 & n32850 ;
  assign n32852 = n32851 ^ n5529 ^ 1'b0 ;
  assign n32853 = n32852 ^ n29040 ^ 1'b0 ;
  assign n32854 = ~n9337 & n16859 ;
  assign n32855 = n32854 ^ n17226 ^ 1'b0 ;
  assign n32856 = ~n7000 & n7405 ;
  assign n32857 = ~n32855 & n32856 ;
  assign n32858 = n32857 ^ n29783 ^ n2382 ;
  assign n32859 = ( n795 & n24672 ) | ( n795 & ~n32858 ) | ( n24672 & ~n32858 ) ;
  assign n32860 = ~n897 & n8353 ;
  assign n32861 = n32860 ^ n1105 ^ 1'b0 ;
  assign n32862 = ~n10756 & n32861 ;
  assign n32863 = n11465 & n32862 ;
  assign n32864 = n32863 ^ n18177 ^ n17123 ;
  assign n32865 = ~n2425 & n29192 ;
  assign n32866 = n11162 & ~n17592 ;
  assign n32867 = n4477 & n32866 ;
  assign n32868 = n32867 ^ n10469 ^ 1'b0 ;
  assign n32869 = n3560 & ~n4884 ;
  assign n32870 = n694 & n32869 ;
  assign n32871 = ~n3313 & n9605 ;
  assign n32873 = n13860 ^ n4543 ^ 1'b0 ;
  assign n32872 = ~n3141 & n7839 ;
  assign n32874 = n32873 ^ n32872 ^ 1'b0 ;
  assign n32875 = n32871 & n32874 ;
  assign n32876 = ~n9019 & n32875 ;
  assign n32877 = n25908 & ~n31042 ;
  assign n32878 = n32877 ^ n29678 ^ 1'b0 ;
  assign n32879 = n6008 | n32878 ;
  assign n32880 = n6181 & n14532 ;
  assign n32881 = n32880 ^ n8902 ^ 1'b0 ;
  assign n32882 = n26030 & n32881 ;
  assign n32883 = ~n18824 & n23550 ;
  assign n32884 = ~n32882 & n32883 ;
  assign n32887 = n7180 & ~n12755 ;
  assign n32888 = n32887 ^ n4368 ^ 1'b0 ;
  assign n32885 = n16374 | n18438 ;
  assign n32886 = n32885 ^ n32444 ^ 1'b0 ;
  assign n32889 = n32888 ^ n32886 ^ n21562 ;
  assign n32891 = ~n765 & n6199 ;
  assign n32890 = x10 & ~n18169 ;
  assign n32892 = n32891 ^ n32890 ^ 1'b0 ;
  assign n32893 = ( n966 & n18583 ) | ( n966 & n32892 ) | ( n18583 & n32892 ) ;
  assign n32894 = n13605 | n25680 ;
  assign n32895 = n8638 & ~n32894 ;
  assign n32896 = ( n8311 & ~n12574 ) | ( n8311 & n32895 ) | ( ~n12574 & n32895 ) ;
  assign n32897 = n32896 ^ n5822 ^ 1'b0 ;
  assign n32898 = n15674 ^ n15533 ^ 1'b0 ;
  assign n32899 = n32897 & ~n32898 ;
  assign n32905 = n15582 ^ n15488 ^ n6470 ;
  assign n32900 = ~n628 & n12802 ;
  assign n32901 = ~n3250 & n32900 ;
  assign n32902 = n14193 ^ n13455 ^ 1'b0 ;
  assign n32903 = ~n32901 & n32902 ;
  assign n32904 = ~n17868 & n32903 ;
  assign n32906 = n32905 ^ n32904 ^ 1'b0 ;
  assign n32907 = n962 & ~n6639 ;
  assign n32908 = ~n10798 & n12395 ;
  assign n32909 = n3056 & ~n32908 ;
  assign n32910 = n8231 & ~n24649 ;
  assign n32911 = n2955 & n32910 ;
  assign n32912 = n802 | n3144 ;
  assign n32913 = n16127 ^ n829 ^ 1'b0 ;
  assign n32914 = n4322 & ~n32913 ;
  assign n32917 = n3312 | n3392 ;
  assign n32918 = n554 | n32917 ;
  assign n32915 = n5338 ^ n2226 ^ n829 ;
  assign n32916 = n554 & ~n32915 ;
  assign n32919 = n32918 ^ n32916 ^ 1'b0 ;
  assign n32920 = ( n26013 & ~n32914 ) | ( n26013 & n32919 ) | ( ~n32914 & n32919 ) ;
  assign n32921 = n4221 & ~n10786 ;
  assign n32922 = n3912 ^ n1597 ^ 1'b0 ;
  assign n32923 = ~n711 & n32922 ;
  assign n32924 = n32921 & n32923 ;
  assign n32925 = n32924 ^ n1864 ^ 1'b0 ;
  assign n32926 = ~n8466 & n32925 ;
  assign n32928 = ~n7527 & n11533 ;
  assign n32927 = n6259 & n26565 ;
  assign n32929 = n32928 ^ n32927 ^ 1'b0 ;
  assign n32930 = n12545 & ~n14665 ;
  assign n32931 = n13063 & n32930 ;
  assign n32932 = n10326 & ~n30614 ;
  assign n32933 = ~n8724 & n32932 ;
  assign n32934 = n32931 & n32933 ;
  assign n32935 = ( n98 & n9039 ) | ( n98 & n10734 ) | ( n9039 & n10734 ) ;
  assign n32936 = n16259 ^ n13265 ^ 1'b0 ;
  assign n32937 = n9716 & n32936 ;
  assign n32938 = n22187 ^ n5791 ^ 1'b0 ;
  assign n32939 = n32937 & ~n32938 ;
  assign n32940 = n32939 ^ n10414 ^ n5114 ;
  assign n32941 = ~n8743 & n11065 ;
  assign n32942 = n10960 | n19964 ;
  assign n32943 = n3313 & ~n9441 ;
  assign n32944 = ~n17683 & n32943 ;
  assign n32945 = n838 & n32944 ;
  assign n32946 = n315 ^ n141 ^ 1'b0 ;
  assign n32947 = n4769 | n12051 ;
  assign n32948 = n32946 & ~n32947 ;
  assign n32949 = n22495 ^ n10851 ^ 1'b0 ;
  assign n32950 = n9606 ^ n3855 ^ 1'b0 ;
  assign n32951 = ~n4104 & n32950 ;
  assign n32952 = n3269 | n20763 ;
  assign n32953 = n11950 | n32952 ;
  assign n32954 = ~n20897 & n32953 ;
  assign n32955 = n2408 & n7641 ;
  assign n32956 = n32955 ^ n24077 ^ 1'b0 ;
  assign n32957 = n23 & n777 ;
  assign n32958 = n32957 ^ n18513 ^ 1'b0 ;
  assign n32959 = n19969 ^ n13832 ^ 1'b0 ;
  assign n32960 = n13457 & ~n32959 ;
  assign n32961 = n25032 & n30870 ;
  assign n32962 = n6131 ^ n398 ^ 1'b0 ;
  assign n32963 = ( ~n403 & n3868 ) | ( ~n403 & n32962 ) | ( n3868 & n32962 ) ;
  assign n32964 = n22456 & n24836 ;
  assign n32965 = ~n32963 & n32964 ;
  assign n32966 = n25592 ^ n20385 ^ n390 ;
  assign n32967 = ~n32143 & n32966 ;
  assign n32968 = n22205 & n32967 ;
  assign n32969 = n6029 | n10942 ;
  assign n32970 = n20019 ^ n13722 ^ n3445 ;
  assign n32971 = n5353 & ~n5834 ;
  assign n32972 = n13172 & n32971 ;
  assign n32973 = n32972 ^ n15420 ^ n2813 ;
  assign n32974 = n25459 ^ n4888 ^ n57 ;
  assign n32975 = ( ~n14426 & n20397 ) | ( ~n14426 & n20467 ) | ( n20397 & n20467 ) ;
  assign n32976 = n27897 & n32975 ;
  assign n32977 = n32976 ^ n4161 ^ 1'b0 ;
  assign n32978 = n2124 & n13522 ;
  assign n32979 = n868 & n32978 ;
  assign n32980 = n572 & n3209 ;
  assign n32981 = n13689 & n32980 ;
  assign n32982 = n15472 | n32981 ;
  assign n32983 = n32982 ^ n23227 ^ 1'b0 ;
  assign n32984 = n32979 | n32983 ;
  assign n32985 = n32984 ^ n25625 ^ 1'b0 ;
  assign n32986 = n612 & ~n32985 ;
  assign n32987 = n17659 ^ n16590 ^ 1'b0 ;
  assign n32988 = n184 | n2825 ;
  assign n32989 = n14358 | n32988 ;
  assign n32990 = n32989 ^ n8979 ^ 1'b0 ;
  assign n32991 = ~n772 & n7543 ;
  assign n32992 = n29752 ^ n22981 ^ n6951 ;
  assign n32993 = n32992 ^ n26722 ^ 1'b0 ;
  assign n32994 = n2051 & ~n32993 ;
  assign n32995 = n8184 ^ n5113 ^ 1'b0 ;
  assign n32996 = n32995 ^ n6348 ^ 1'b0 ;
  assign n32997 = n7320 & n32996 ;
  assign n33001 = n9474 ^ n9070 ^ n4975 ;
  assign n32998 = n3575 | n6178 ;
  assign n32999 = n32998 ^ n23500 ^ n2019 ;
  assign n33000 = ( n5357 & n5797 ) | ( n5357 & n32999 ) | ( n5797 & n32999 ) ;
  assign n33002 = n33001 ^ n33000 ^ n21370 ;
  assign n33003 = n11025 & ~n12407 ;
  assign n33004 = ~n24450 & n33003 ;
  assign n33005 = n11300 ^ n6618 ^ 1'b0 ;
  assign n33006 = n2022 & n10846 ;
  assign n33007 = n15266 | n33006 ;
  assign n33008 = n33007 ^ n22353 ^ 1'b0 ;
  assign n33009 = n3149 & n29746 ;
  assign n33010 = n31410 ^ n8948 ^ 1'b0 ;
  assign n33011 = n30723 ^ n11488 ^ 1'b0 ;
  assign n33012 = ~n20024 & n33011 ;
  assign n33017 = n10764 ^ n1327 ^ 1'b0 ;
  assign n33018 = ~n5756 & n33017 ;
  assign n33013 = n1017 & ~n5062 ;
  assign n33014 = ~n1017 & n33013 ;
  assign n33015 = n33014 ^ n8211 ^ 1'b0 ;
  assign n33016 = n395 & ~n33015 ;
  assign n33019 = n33018 ^ n33016 ^ 1'b0 ;
  assign n33020 = n572 | n16839 ;
  assign n33021 = n2818 & n19372 ;
  assign n33022 = n8626 ^ n7822 ^ 1'b0 ;
  assign n33023 = n17945 ^ n709 ^ 1'b0 ;
  assign n33024 = n12040 & ~n33023 ;
  assign n33025 = n33024 ^ n21251 ^ n2622 ;
  assign n33026 = ( n33021 & n33022 ) | ( n33021 & ~n33025 ) | ( n33022 & ~n33025 ) ;
  assign n33027 = n12451 & n25489 ;
  assign n33028 = n33027 ^ n27619 ^ 1'b0 ;
  assign n33029 = n2696 | n15401 ;
  assign n33030 = n33029 ^ n19799 ^ 1'b0 ;
  assign n33031 = n7159 ^ n612 ^ 1'b0 ;
  assign n33032 = n9218 & n33031 ;
  assign n33033 = n33032 ^ n23050 ^ 1'b0 ;
  assign n33034 = n4316 & n33033 ;
  assign n33035 = n16622 & n19468 ;
  assign n33036 = ~n6025 & n8901 ;
  assign n33037 = ~n15177 & n20608 ;
  assign n33038 = n33037 ^ n11769 ^ 1'b0 ;
  assign n33039 = n19209 | n33038 ;
  assign n33040 = n26683 & ~n33039 ;
  assign n33041 = n30957 ^ n15392 ^ 1'b0 ;
  assign n33042 = n5045 & n29297 ;
  assign n33043 = ( n6167 & ~n7675 ) | ( n6167 & n12134 ) | ( ~n7675 & n12134 ) ;
  assign n33044 = n33043 ^ n12868 ^ 1'b0 ;
  assign n33045 = n6564 ^ n1405 ^ 1'b0 ;
  assign n33046 = n6551 & n33045 ;
  assign n33047 = ~n24534 & n33046 ;
  assign n33048 = n8962 & ~n33047 ;
  assign n33049 = n47 & n33048 ;
  assign n33050 = n2395 & n6340 ;
  assign n33051 = n21624 & n33050 ;
  assign n33057 = n11558 ^ n177 ^ 1'b0 ;
  assign n33056 = ~n1241 & n4196 ;
  assign n33058 = n33057 ^ n33056 ^ 1'b0 ;
  assign n33059 = ( n15063 & n24640 ) | ( n15063 & ~n33058 ) | ( n24640 & ~n33058 ) ;
  assign n33052 = n4430 & n10405 ;
  assign n33053 = n33052 ^ n23399 ^ 1'b0 ;
  assign n33054 = n18465 ^ n16006 ^ 1'b0 ;
  assign n33055 = n33053 & ~n33054 ;
  assign n33060 = n33059 ^ n33055 ^ n2622 ;
  assign n33061 = n3610 & n20301 ;
  assign n33062 = n33061 ^ n7441 ^ 1'b0 ;
  assign n33064 = n5395 | n16581 ;
  assign n33065 = n8904 | n33064 ;
  assign n33066 = n33065 ^ n27818 ^ 1'b0 ;
  assign n33067 = n30251 & n33066 ;
  assign n33063 = n299 & ~n9961 ;
  assign n33068 = n33067 ^ n33063 ^ 1'b0 ;
  assign n33069 = n30671 ^ n780 ^ 1'b0 ;
  assign n33070 = ~n17238 & n33069 ;
  assign n33071 = n33070 ^ n30425 ^ 1'b0 ;
  assign n33072 = n8265 & ~n33071 ;
  assign n33073 = n33072 ^ n16378 ^ 1'b0 ;
  assign n33074 = n13950 & ~n33073 ;
  assign n33075 = n28835 ^ n7540 ^ 1'b0 ;
  assign n33076 = n17380 ^ n7239 ^ 1'b0 ;
  assign n33077 = n6381 | n33076 ;
  assign n33078 = n30324 ^ n183 ^ 1'b0 ;
  assign n33079 = n17149 ^ n8445 ^ 1'b0 ;
  assign n33080 = n33079 ^ n28176 ^ 1'b0 ;
  assign n33081 = ( ~n33077 & n33078 ) | ( ~n33077 & n33080 ) | ( n33078 & n33080 ) ;
  assign n33082 = n17373 ^ n15101 ^ 1'b0 ;
  assign n33083 = n8049 ^ n7193 ^ 1'b0 ;
  assign n33084 = ( ~n9109 & n23170 ) | ( ~n9109 & n33083 ) | ( n23170 & n33083 ) ;
  assign n33085 = x9 & n889 ;
  assign n33086 = n9231 & n9730 ;
  assign n33087 = n19697 | n33086 ;
  assign n33088 = x0 | n21647 ;
  assign n33091 = n16721 ^ n3500 ^ 1'b0 ;
  assign n33089 = ( ~n1277 & n9612 ) | ( ~n1277 & n26599 ) | ( n9612 & n26599 ) ;
  assign n33090 = n11329 & ~n33089 ;
  assign n33092 = n33091 ^ n33090 ^ 1'b0 ;
  assign n33093 = n10719 ^ n9989 ^ 1'b0 ;
  assign n33094 = n22530 & n33093 ;
  assign n33095 = ~n2545 & n33094 ;
  assign n33096 = ~n7477 & n18046 ;
  assign n33097 = n4992 & n33096 ;
  assign n33098 = n33097 ^ n12895 ^ 1'b0 ;
  assign n33104 = n2094 & ~n13402 ;
  assign n33105 = n33104 ^ n2044 ^ 1'b0 ;
  assign n33099 = n13703 ^ n6985 ^ n4281 ;
  assign n33100 = n4515 | n21041 ;
  assign n33101 = n33100 ^ n13238 ^ 1'b0 ;
  assign n33102 = n33101 ^ n25601 ^ 1'b0 ;
  assign n33103 = n33099 | n33102 ;
  assign n33106 = n33105 ^ n33103 ^ 1'b0 ;
  assign n33107 = n5704 | n15959 ;
  assign n33108 = n30407 & ~n33107 ;
  assign n33109 = n23258 & ~n33108 ;
  assign n33110 = ~n31026 & n33109 ;
  assign n33111 = n27656 & ~n33110 ;
  assign n33112 = n20831 ^ n1628 ^ 1'b0 ;
  assign n33113 = ~n16568 & n33112 ;
  assign n33114 = n33113 ^ n17380 ^ 1'b0 ;
  assign n33115 = n10634 ^ n5531 ^ n3174 ;
  assign n33116 = n33115 ^ n30198 ^ 1'b0 ;
  assign n33117 = n2627 | n7318 ;
  assign n33118 = n33117 ^ n30760 ^ 1'b0 ;
  assign n33119 = ~n2994 & n33118 ;
  assign n33120 = n19577 ^ n7460 ^ 1'b0 ;
  assign n33121 = ~n17037 & n33120 ;
  assign n33122 = n19310 & ~n29439 ;
  assign n33123 = n33122 ^ n6060 ^ 1'b0 ;
  assign n33124 = ( ~n9770 & n20588 ) | ( ~n9770 & n27135 ) | ( n20588 & n27135 ) ;
  assign n33125 = n33124 ^ n16385 ^ 1'b0 ;
  assign n33126 = ~n3330 & n33125 ;
  assign n33127 = n17207 ^ n7957 ^ 1'b0 ;
  assign n33128 = n3007 ^ n870 ^ 1'b0 ;
  assign n33129 = n10239 & ~n33128 ;
  assign n33130 = n33129 ^ n3489 ^ 1'b0 ;
  assign n33131 = ~n32823 & n33130 ;
  assign n33132 = n32823 & n33131 ;
  assign n33133 = ~n2695 & n33132 ;
  assign n33134 = ~n33132 & n33133 ;
  assign n33135 = n18036 ^ n1906 ^ 1'b0 ;
  assign n33136 = n5180 ^ n2006 ^ 1'b0 ;
  assign n33137 = n29455 & n33136 ;
  assign n33138 = ( ~n11956 & n33135 ) | ( ~n11956 & n33137 ) | ( n33135 & n33137 ) ;
  assign n33139 = n33138 ^ n25260 ^ n3802 ;
  assign n33140 = n21315 & n28898 ;
  assign n33141 = ~n139 & n11902 ;
  assign n33142 = ~n27055 & n33141 ;
  assign n33143 = n33142 ^ n12166 ^ 1'b0 ;
  assign n33144 = n1682 | n20897 ;
  assign n33145 = n44 & ~n15272 ;
  assign n33146 = n5533 & n15963 ;
  assign n33147 = n23286 & n33146 ;
  assign n33148 = n33145 & n33147 ;
  assign n33149 = n8936 & ~n19870 ;
  assign n33150 = n21734 | n25208 ;
  assign n33151 = n6954 | n15953 ;
  assign n33152 = n33151 ^ n25076 ^ 1'b0 ;
  assign n33153 = n20205 ^ n6922 ^ n6360 ;
  assign n33154 = n6620 | n12075 ;
  assign n33155 = n19351 & n33154 ;
  assign n33156 = ~n33153 & n33155 ;
  assign n33158 = n5987 | n28070 ;
  assign n33159 = n5987 & ~n33158 ;
  assign n33160 = n8222 | n10938 ;
  assign n33161 = n33160 ^ n2887 ^ 1'b0 ;
  assign n33162 = n33161 ^ n17439 ^ 1'b0 ;
  assign n33163 = n33159 | n33162 ;
  assign n33157 = ~n22717 & n24330 ;
  assign n33164 = n33163 ^ n33157 ^ 1'b0 ;
  assign n33165 = n33164 ^ n5722 ^ 1'b0 ;
  assign n33166 = n9449 & n33165 ;
  assign n33170 = n5106 & n5386 ;
  assign n33167 = n1124 & n13676 ;
  assign n33168 = n33167 ^ n14903 ^ 1'b0 ;
  assign n33169 = n33168 ^ n12227 ^ n162 ;
  assign n33171 = n33170 ^ n33169 ^ n20503 ;
  assign n33172 = ( n1373 & ~n1400 ) | ( n1373 & n9420 ) | ( ~n1400 & n9420 ) ;
  assign n33173 = ~n22996 & n33172 ;
  assign n33174 = ~n14188 & n15350 ;
  assign n33175 = n33174 ^ n23173 ^ 1'b0 ;
  assign n33176 = n11119 ^ n8172 ^ 1'b0 ;
  assign n33177 = n7452 | n33176 ;
  assign n33178 = n23042 ^ n16325 ^ 1'b0 ;
  assign n33179 = n41 & n15191 ;
  assign n33180 = n18479 | n33179 ;
  assign n33181 = ( ~n23483 & n32264 ) | ( ~n23483 & n33180 ) | ( n32264 & n33180 ) ;
  assign n33182 = n132 | n15791 ;
  assign n33183 = n33182 ^ n29983 ^ 1'b0 ;
  assign n33184 = n2917 & n32521 ;
  assign n33185 = n33184 ^ n1084 ^ 1'b0 ;
  assign n33186 = n31184 ^ n25333 ^ 1'b0 ;
  assign n33187 = n3310 | n33186 ;
  assign n33188 = n26287 ^ n8427 ^ n191 ;
  assign n33189 = n33188 ^ n13250 ^ 1'b0 ;
  assign n33190 = n7768 | n33189 ;
  assign n33196 = n18850 & n20281 ;
  assign n33195 = n15751 & ~n16158 ;
  assign n33191 = n16154 & ~n29060 ;
  assign n33192 = ~n1278 & n33191 ;
  assign n33193 = n33192 ^ n16695 ^ 1'b0 ;
  assign n33194 = n14520 | n33193 ;
  assign n33197 = n33196 ^ n33195 ^ n33194 ;
  assign n33198 = ~n5162 & n30068 ;
  assign n33199 = n24021 & n33198 ;
  assign n33200 = ( n4159 & n12707 ) | ( n4159 & ~n33199 ) | ( n12707 & ~n33199 ) ;
  assign n33201 = x10 & n8993 ;
  assign n33202 = n135 & n15007 ;
  assign n33203 = n7794 ^ n763 ^ 1'b0 ;
  assign n33204 = n30211 ^ n1249 ^ 1'b0 ;
  assign n33205 = n33203 & n33204 ;
  assign n33206 = ~n7913 & n22353 ;
  assign n33207 = n20112 ^ n3471 ^ 1'b0 ;
  assign n33208 = n344 & n7927 ;
  assign n33209 = n33208 ^ n9962 ^ 1'b0 ;
  assign n33210 = n14116 & ~n33209 ;
  assign n33211 = ( ~n8714 & n33207 ) | ( ~n8714 & n33210 ) | ( n33207 & n33210 ) ;
  assign n33212 = n17155 ^ n1367 ^ 1'b0 ;
  assign n33213 = n33212 ^ n8897 ^ n6384 ;
  assign n33214 = n1295 & ~n11447 ;
  assign n33215 = n33214 ^ n26573 ^ 1'b0 ;
  assign n33216 = n28346 ^ n10802 ^ 1'b0 ;
  assign n33217 = n3644 & ~n33216 ;
  assign n33218 = ~n3738 & n6229 ;
  assign n33219 = n22052 & n33218 ;
  assign n33220 = n3581 & n22724 ;
  assign n33221 = ~n3229 & n33220 ;
  assign n33222 = n33221 ^ n14115 ^ n4922 ;
  assign n33223 = n20176 ^ n9246 ^ 1'b0 ;
  assign n33224 = ( n5974 & n24644 ) | ( n5974 & n33223 ) | ( n24644 & n33223 ) ;
  assign n33225 = n9224 | n12204 ;
  assign n33226 = n33225 ^ n27735 ^ 1'b0 ;
  assign n33227 = n7925 & n10705 ;
  assign n33228 = ~n1138 & n33227 ;
  assign n33229 = n12177 | n33228 ;
  assign n33230 = n806 | n33229 ;
  assign n33231 = n10219 | n17168 ;
  assign n33232 = n2831 & n33231 ;
  assign n33233 = ~n21056 & n33232 ;
  assign n33234 = ~n1533 & n2022 ;
  assign n33235 = n33234 ^ n6071 ^ 1'b0 ;
  assign n33236 = n7104 ^ n3173 ^ 1'b0 ;
  assign n33237 = n33236 ^ n9968 ^ 1'b0 ;
  assign n33238 = n13091 | n33237 ;
  assign n33239 = n8890 ^ n1900 ^ 1'b0 ;
  assign n33240 = n27886 | n33239 ;
  assign n33241 = n5606 ^ n5374 ^ 1'b0 ;
  assign n33242 = n7641 & n33241 ;
  assign n33243 = n17550 & n33242 ;
  assign n33244 = ~n10812 & n28442 ;
  assign n33245 = n33244 ^ n22854 ^ 1'b0 ;
  assign n33246 = n23674 & n33245 ;
  assign n33247 = n33246 ^ n18884 ^ 1'b0 ;
  assign n33248 = ( ~n25612 & n28495 ) | ( ~n25612 & n33247 ) | ( n28495 & n33247 ) ;
  assign n33249 = n25234 ^ n2139 ^ 1'b0 ;
  assign n33250 = n33248 & ~n33249 ;
  assign n33251 = n33250 ^ n27507 ^ 1'b0 ;
  assign n33254 = n1550 & ~n24996 ;
  assign n33255 = n33254 ^ n9341 ^ 1'b0 ;
  assign n33252 = n16492 ^ n3313 ^ 1'b0 ;
  assign n33253 = n20698 & ~n33252 ;
  assign n33256 = n33255 ^ n33253 ^ n32134 ;
  assign n33257 = n10369 ^ n5527 ^ 1'b0 ;
  assign n33258 = n756 | n7859 ;
  assign n33259 = n10583 & ~n33258 ;
  assign n33260 = n4012 | n10963 ;
  assign n33261 = n33260 ^ n12525 ^ 1'b0 ;
  assign n33263 = ~n5004 & n9285 ;
  assign n33262 = n3409 | n17283 ;
  assign n33264 = n33263 ^ n33262 ^ 1'b0 ;
  assign n33265 = n24202 ^ n11652 ^ 1'b0 ;
  assign n33266 = ( n7652 & ~n20761 ) | ( n7652 & n27877 ) | ( ~n20761 & n27877 ) ;
  assign n33270 = n4549 ^ n4196 ^ 1'b0 ;
  assign n33267 = n1940 | n13218 ;
  assign n33268 = ( ~n13361 & n24665 ) | ( ~n13361 & n33267 ) | ( n24665 & n33267 ) ;
  assign n33269 = n3533 & n33268 ;
  assign n33271 = n33270 ^ n33269 ^ 1'b0 ;
  assign n33272 = n11118 & n12822 ;
  assign n33273 = n9422 ^ n3608 ^ 1'b0 ;
  assign n33274 = n9393 & n33273 ;
  assign n33275 = n28026 ^ n2633 ^ 1'b0 ;
  assign n33276 = n7120 ^ n6614 ^ 1'b0 ;
  assign n33277 = ~n33275 & n33276 ;
  assign n33278 = n33277 ^ n982 ^ 1'b0 ;
  assign n33279 = n15972 & n33278 ;
  assign n33280 = n33274 & n33279 ;
  assign n33281 = n9864 & n33280 ;
  assign n33282 = n3140 | n10296 ;
  assign n33283 = n9117 & ~n14351 ;
  assign n33284 = ~n6337 & n33283 ;
  assign n33285 = n30502 ^ n13747 ^ 1'b0 ;
  assign n33286 = n23 & ~n9655 ;
  assign n33287 = ~n24736 & n33286 ;
  assign n33290 = n2599 ^ n324 ^ 1'b0 ;
  assign n33288 = ~n12883 & n27829 ;
  assign n33289 = n2182 & n33288 ;
  assign n33291 = n33290 ^ n33289 ^ 1'b0 ;
  assign n33292 = n15199 & n33291 ;
  assign n33293 = n14381 | n15607 ;
  assign n33294 = ~n1395 & n33293 ;
  assign n33295 = ~n2230 & n6564 ;
  assign n33296 = n17765 | n33295 ;
  assign n33297 = n13072 ^ n5348 ^ 1'b0 ;
  assign n33298 = n2044 | n10170 ;
  assign n33299 = n33298 ^ n5442 ^ 1'b0 ;
  assign n33300 = n7110 | n33299 ;
  assign n33301 = n29611 & ~n33300 ;
  assign n33302 = n978 & ~n33301 ;
  assign n33303 = n22103 | n25674 ;
  assign n33304 = n33303 ^ n22161 ^ 1'b0 ;
  assign n33305 = n32077 & ~n33304 ;
  assign n33306 = n33305 ^ n1344 ^ 1'b0 ;
  assign n33307 = ( n3602 & n8001 ) | ( n3602 & n8784 ) | ( n8001 & n8784 ) ;
  assign n33308 = ( n21578 & n26453 ) | ( n21578 & ~n33307 ) | ( n26453 & ~n33307 ) ;
  assign n33309 = n5370 | n10418 ;
  assign n33310 = n33308 | n33309 ;
  assign n33311 = n25477 ^ n1837 ^ 1'b0 ;
  assign n33312 = ~n3998 & n13714 ;
  assign n33313 = n33312 ^ n14752 ^ 1'b0 ;
  assign n33314 = n20589 ^ n206 ^ 1'b0 ;
  assign n33315 = ~n6471 & n9902 ;
  assign n33316 = n682 & ~n17583 ;
  assign n33317 = n33316 ^ n6614 ^ 1'b0 ;
  assign n33318 = n20250 ^ n7087 ^ n2148 ;
  assign n33319 = n33318 ^ n32707 ^ 1'b0 ;
  assign n33320 = n1173 | n22373 ;
  assign n33321 = n10738 & ~n33320 ;
  assign n33322 = n33321 ^ n21990 ^ 1'b0 ;
  assign n33323 = n27276 & n33322 ;
  assign n33324 = n6451 | n31814 ;
  assign n33325 = n2324 & n2736 ;
  assign n33326 = ~n13570 & n33325 ;
  assign n33327 = ( n228 & ~n8271 ) | ( n228 & n33326 ) | ( ~n8271 & n33326 ) ;
  assign n33328 = n18337 ^ n4105 ^ n158 ;
  assign n33329 = n33328 ^ n1332 ^ 1'b0 ;
  assign n33330 = n33329 ^ n7544 ^ 1'b0 ;
  assign n33331 = n7911 | n33330 ;
  assign n33332 = n4598 & ~n5794 ;
  assign n33333 = n12486 & ~n20134 ;
  assign n33334 = n33332 & n33333 ;
  assign n33335 = n33334 ^ n980 ^ 1'b0 ;
  assign n33336 = ~n17622 & n33335 ;
  assign n33337 = n10241 & n13396 ;
  assign n33338 = n17781 & n33337 ;
  assign n33339 = n3330 & ~n14211 ;
  assign n33340 = n9503 & n33339 ;
  assign n33341 = n12456 & ~n33340 ;
  assign n33342 = n17677 & n21020 ;
  assign n33343 = n19503 ^ n4769 ^ 1'b0 ;
  assign n33344 = n28257 | n33343 ;
  assign n33345 = n33344 ^ n20593 ^ 1'b0 ;
  assign n33346 = n15167 & n15737 ;
  assign n33347 = n33346 ^ n7900 ^ 1'b0 ;
  assign n33349 = n8524 & n23787 ;
  assign n33348 = n4307 | n13748 ;
  assign n33350 = n33349 ^ n33348 ^ 1'b0 ;
  assign n33351 = n33350 ^ n9851 ^ 1'b0 ;
  assign n33352 = n33347 & n33351 ;
  assign n33353 = ~n12810 & n19165 ;
  assign n33354 = ~n3243 & n33353 ;
  assign n33355 = n18945 ^ n7789 ^ 1'b0 ;
  assign n33356 = n13137 ^ n4653 ^ 1'b0 ;
  assign n33357 = n6616 & ~n33356 ;
  assign n33358 = n12806 | n33357 ;
  assign n33359 = n28086 ^ n5389 ^ 1'b0 ;
  assign n33360 = n33359 ^ n30164 ^ 1'b0 ;
  assign n33361 = n25321 | n27697 ;
  assign n33362 = n33361 ^ n2190 ^ 1'b0 ;
  assign n33363 = n514 & ~n771 ;
  assign n33364 = n18761 & n33363 ;
  assign n33365 = n953 & n18063 ;
  assign n33366 = ~n10386 & n33365 ;
  assign n33369 = n14974 | n20518 ;
  assign n33367 = ( n1652 & n1996 ) | ( n1652 & n2732 ) | ( n1996 & n2732 ) ;
  assign n33368 = n33367 ^ n26923 ^ 1'b0 ;
  assign n33370 = n33369 ^ n33368 ^ 1'b0 ;
  assign n33371 = ~n33366 & n33370 ;
  assign n33372 = n20 & ~n26392 ;
  assign n33373 = n33372 ^ n26457 ^ n7821 ;
  assign n33374 = n6678 & n33231 ;
  assign n33375 = n33374 ^ n9020 ^ 1'b0 ;
  assign n33376 = n28149 | n33375 ;
  assign n33377 = n873 & ~n15189 ;
  assign n33378 = n1614 & ~n33377 ;
  assign n33379 = n33378 ^ n29089 ^ 1'b0 ;
  assign n33380 = n11919 & ~n23944 ;
  assign n33381 = n12493 & n12707 ;
  assign n33382 = n1506 & ~n33381 ;
  assign n33383 = n33382 ^ n23089 ^ 1'b0 ;
  assign n33384 = n11658 ^ n6595 ^ 1'b0 ;
  assign n33385 = n1262 & n33384 ;
  assign n33386 = n3519 & n11429 ;
  assign n33387 = n11958 & ~n13164 ;
  assign n33388 = n21862 ^ n18302 ^ 1'b0 ;
  assign n33389 = n13889 | n33388 ;
  assign n33390 = n32955 ^ n18736 ^ 1'b0 ;
  assign n33391 = ~n6892 & n33390 ;
  assign n33392 = n33391 ^ n26769 ^ 1'b0 ;
  assign n33393 = n7544 & ~n12169 ;
  assign n33394 = n10209 ^ n8137 ^ n759 ;
  assign n33395 = n33394 ^ n14774 ^ 1'b0 ;
  assign n33396 = ~n33393 & n33395 ;
  assign n33397 = n4352 | n15504 ;
  assign n33398 = n4607 & ~n33397 ;
  assign n33399 = n10178 ^ n3662 ^ 1'b0 ;
  assign n33400 = n16828 & n33399 ;
  assign n33401 = n33400 ^ n6716 ^ 1'b0 ;
  assign n33402 = n33398 | n33401 ;
  assign n33403 = n5128 & n33402 ;
  assign n33404 = n3713 & n33403 ;
  assign n33405 = n9290 | n12928 ;
  assign n33406 = ~n1980 & n3590 ;
  assign n33407 = ~n33405 & n33406 ;
  assign n33408 = ~n75 & n4345 ;
  assign n33409 = ( n464 & n20343 ) | ( n464 & ~n21052 ) | ( n20343 & ~n21052 ) ;
  assign n33410 = ~n10311 & n26437 ;
  assign n33411 = n33410 ^ n20679 ^ 1'b0 ;
  assign n33412 = n33411 ^ n16898 ^ 1'b0 ;
  assign n33413 = n29946 ^ n14769 ^ 1'b0 ;
  assign n33414 = n32166 & n33413 ;
  assign n33415 = n2271 ^ n2230 ^ 1'b0 ;
  assign n33416 = ( n576 & n27356 ) | ( n576 & n33415 ) | ( n27356 & n33415 ) ;
  assign n33417 = n2790 & ~n6138 ;
  assign n33418 = n7354 & ~n29581 ;
  assign n33419 = n7572 & n33418 ;
  assign n33420 = n10479 | n14749 ;
  assign n33421 = n13785 ^ n5080 ^ 1'b0 ;
  assign n33422 = n15975 | n33421 ;
  assign n33423 = n12129 | n18095 ;
  assign n33424 = n33423 ^ n3393 ^ 1'b0 ;
  assign n33425 = ~n33422 & n33424 ;
  assign n33426 = n33420 & ~n33425 ;
  assign n33427 = n2449 | n8220 ;
  assign n33428 = n14775 ^ n11905 ^ 1'b0 ;
  assign n33429 = n8140 | n33428 ;
  assign n33430 = n33429 ^ n30300 ^ x3 ;
  assign n33431 = n33430 ^ n28436 ^ 1'b0 ;
  assign n33432 = n30809 | n33431 ;
  assign n33433 = n33427 & n33432 ;
  assign n33434 = n4772 | n8565 ;
  assign n33435 = ~n73 & n6097 ;
  assign n33436 = n33435 ^ n9135 ^ 1'b0 ;
  assign n33437 = n13613 & ~n31074 ;
  assign n33438 = ( n4896 & ~n33436 ) | ( n4896 & n33437 ) | ( ~n33436 & n33437 ) ;
  assign n33439 = ~n14381 & n33438 ;
  assign n33440 = ~n17346 & n33439 ;
  assign n33441 = ( n4882 & n22677 ) | ( n4882 & ~n26268 ) | ( n22677 & ~n26268 ) ;
  assign n33442 = n16615 | n33441 ;
  assign n33443 = n619 | n33442 ;
  assign n33444 = n4572 & ~n17614 ;
  assign n33445 = n33444 ^ n1690 ^ 1'b0 ;
  assign n33446 = ( n16940 & n33443 ) | ( n16940 & ~n33445 ) | ( n33443 & ~n33445 ) ;
  assign n33447 = ( n2370 & n5055 ) | ( n2370 & ~n23428 ) | ( n5055 & ~n23428 ) ;
  assign n33448 = n21046 & ~n32423 ;
  assign n33449 = ~n33447 & n33448 ;
  assign n33450 = n23950 | n33449 ;
  assign n33451 = n4729 & ~n26247 ;
  assign n33452 = n33451 ^ n1818 ^ 1'b0 ;
  assign n33453 = n25387 ^ n10543 ^ 1'b0 ;
  assign n33454 = n33452 & ~n33453 ;
  assign n33455 = n2008 | n29663 ;
  assign n33456 = n8698 | n33455 ;
  assign n33457 = n15895 ^ n15197 ^ 1'b0 ;
  assign n33458 = ~n11182 & n33457 ;
  assign n33459 = ~n8195 & n33458 ;
  assign n33460 = n16787 & ~n30863 ;
  assign n33461 = n3428 & ~n4667 ;
  assign n33462 = ~n6274 & n21991 ;
  assign n33463 = ~n28068 & n33462 ;
  assign n33464 = ( ~n110 & n889 ) | ( ~n110 & n4422 ) | ( n889 & n4422 ) ;
  assign n33465 = n8163 & n33464 ;
  assign n33466 = n2008 & n33465 ;
  assign n33467 = n11697 | n33466 ;
  assign n33468 = n1182 & n9947 ;
  assign n33469 = n33468 ^ n10758 ^ 1'b0 ;
  assign n33470 = ~n2205 & n2686 ;
  assign n33471 = ~n33469 & n33470 ;
  assign n33472 = n6166 & n12084 ;
  assign n33473 = n33472 ^ n7254 ^ 1'b0 ;
  assign n33474 = n13838 ^ n9959 ^ 1'b0 ;
  assign n33475 = ~n25406 & n25953 ;
  assign n33476 = n33475 ^ n8631 ^ 1'b0 ;
  assign n33477 = n16715 ^ n1362 ^ 1'b0 ;
  assign n33478 = n16064 & ~n17753 ;
  assign n33479 = ~n6552 & n19917 ;
  assign n33480 = n18505 ^ n4138 ^ 1'b0 ;
  assign n33481 = n33480 ^ n22417 ^ 1'b0 ;
  assign n33483 = n1940 & n5513 ;
  assign n33482 = n16079 ^ n13196 ^ 1'b0 ;
  assign n33484 = n33483 ^ n33482 ^ 1'b0 ;
  assign n33485 = n33481 | n33484 ;
  assign n33486 = n18462 ^ n18030 ^ n2785 ;
  assign n33487 = n29210 | n30816 ;
  assign n33488 = n33487 ^ n11734 ^ 1'b0 ;
  assign n33489 = n5665 | n12933 ;
  assign n33490 = n10161 | n17112 ;
  assign n33491 = n33489 & ~n33490 ;
  assign n33492 = n15864 ^ n12397 ^ 1'b0 ;
  assign n33493 = n27823 ^ n6430 ^ 1'b0 ;
  assign n33495 = ~n1633 & n8279 ;
  assign n33496 = n33495 ^ n7078 ^ 1'b0 ;
  assign n33497 = n11500 | n33496 ;
  assign n33494 = n10684 & n10793 ;
  assign n33498 = n33497 ^ n33494 ^ 1'b0 ;
  assign n33499 = n33498 ^ n17558 ^ n99 ;
  assign n33500 = n4925 & n15271 ;
  assign n33501 = n5193 & n33500 ;
  assign n33502 = n31432 | n33501 ;
  assign n33503 = n1310 & ~n33502 ;
  assign n33504 = n9465 ^ n7069 ^ 1'b0 ;
  assign n33505 = n33504 ^ n10667 ^ n10576 ;
  assign n33508 = n24540 ^ n10068 ^ 1'b0 ;
  assign n33506 = n10898 & ~n15705 ;
  assign n33507 = n33506 ^ n3398 ^ 1'b0 ;
  assign n33509 = n33508 ^ n33507 ^ n3371 ;
  assign n33511 = ~n2986 & n11095 ;
  assign n33510 = n2125 & n6050 ;
  assign n33512 = n33511 ^ n33510 ^ n32684 ;
  assign n33513 = n9583 & n10051 ;
  assign n33514 = n7286 & n33513 ;
  assign n33515 = n17484 | n23084 ;
  assign n33516 = n33515 ^ n19397 ^ 1'b0 ;
  assign n33517 = ~n33514 & n33516 ;
  assign n33518 = n31617 ^ n21226 ^ 1'b0 ;
  assign n33519 = n1822 & ~n6565 ;
  assign n33520 = ~n8215 & n33519 ;
  assign n33521 = ( n9635 & n20250 ) | ( n9635 & ~n33520 ) | ( n20250 & ~n33520 ) ;
  assign n33522 = n694 & ~n15993 ;
  assign n33523 = n33522 ^ n4447 ^ 1'b0 ;
  assign n33524 = n33523 ^ n150 ^ 1'b0 ;
  assign n33525 = n26098 ^ n5272 ^ 1'b0 ;
  assign n33526 = ~n30509 & n33525 ;
  assign n33527 = n33526 ^ n3636 ^ 1'b0 ;
  assign n33528 = n4892 | n9097 ;
  assign n33529 = n15334 & n16852 ;
  assign n33530 = n31795 & n33529 ;
  assign n33531 = n33530 ^ n18730 ^ n12033 ;
  assign n33532 = n15636 ^ n8530 ^ 1'b0 ;
  assign n33533 = n23190 & ~n32684 ;
  assign n33534 = n33533 ^ n28068 ^ 1'b0 ;
  assign n33535 = ~n3968 & n8965 ;
  assign n33536 = n33534 & n33535 ;
  assign n33537 = ~n10229 & n16876 ;
  assign n33538 = n33537 ^ n10546 ^ 1'b0 ;
  assign n33539 = n33538 ^ n23795 ^ 1'b0 ;
  assign n33540 = n20186 ^ n6191 ^ n3399 ;
  assign n33541 = n22496 ^ n2294 ^ 1'b0 ;
  assign n33542 = ~n7108 & n33541 ;
  assign n33543 = n8133 ^ n8129 ^ n5845 ;
  assign n33544 = n326 & ~n3174 ;
  assign n33545 = n11190 & n33544 ;
  assign n33546 = n20600 ^ n1664 ^ 1'b0 ;
  assign n33547 = n8597 & n11836 ;
  assign n33548 = ~n1459 & n23946 ;
  assign n33550 = n6307 | n16519 ;
  assign n33551 = n33550 ^ n6682 ^ 1'b0 ;
  assign n33549 = ( n20954 & ~n21578 ) | ( n20954 & n29156 ) | ( ~n21578 & n29156 ) ;
  assign n33552 = n33551 ^ n33549 ^ n3840 ;
  assign n33553 = n15692 & n29574 ;
  assign n33554 = n10129 & n31582 ;
  assign n33555 = ~n33553 & n33554 ;
  assign n33556 = n25347 ^ n18453 ^ n7101 ;
  assign n33557 = n15654 ^ n8830 ^ 1'b0 ;
  assign n33558 = n33536 ^ n1134 ^ 1'b0 ;
  assign n33559 = n33557 | n33558 ;
  assign n33560 = ~n13782 & n14827 ;
  assign n33561 = n21323 & n30746 ;
  assign n33562 = n4624 & n33561 ;
  assign n33563 = n2195 | n6308 ;
  assign n33564 = n17729 & ~n33563 ;
  assign n33565 = n13034 ^ n3993 ^ 1'b0 ;
  assign n33566 = n11296 | n33565 ;
  assign n33567 = n475 & ~n4990 ;
  assign n33568 = n33567 ^ n863 ^ 1'b0 ;
  assign n33571 = n4947 & n6808 ;
  assign n33572 = n6437 & ~n33571 ;
  assign n33573 = ~n14858 & n33572 ;
  assign n33569 = n4658 | n5823 ;
  assign n33570 = n23983 | n33569 ;
  assign n33574 = n33573 ^ n33570 ^ 1'b0 ;
  assign n33575 = x7 & n11749 ;
  assign n33576 = n33574 & n33575 ;
  assign n33577 = ~n14768 & n22906 ;
  assign n33584 = ~n13059 & n22453 ;
  assign n33583 = n7984 & n10950 ;
  assign n33585 = n33584 ^ n33583 ^ 1'b0 ;
  assign n33578 = n231 ^ n135 ^ 1'b0 ;
  assign n33579 = n10065 | n10430 ;
  assign n33580 = n33579 ^ n7763 ^ 1'b0 ;
  assign n33581 = n16405 & n33580 ;
  assign n33582 = n33578 & n33581 ;
  assign n33586 = n33585 ^ n33582 ^ 1'b0 ;
  assign n33587 = n9181 & ~n33586 ;
  assign n33588 = n10101 ^ n3732 ^ 1'b0 ;
  assign n33589 = n24759 ^ n16917 ^ 1'b0 ;
  assign n33590 = ~n6173 & n33589 ;
  assign n33591 = n33590 ^ n15061 ^ 1'b0 ;
  assign n33592 = n21418 ^ n8120 ^ 1'b0 ;
  assign n33593 = n9075 & ~n33592 ;
  assign n33594 = n29004 ^ n26922 ^ 1'b0 ;
  assign n33598 = ~n113 & n24694 ;
  assign n33599 = n33598 ^ n13404 ^ 1'b0 ;
  assign n33595 = n762 & n2686 ;
  assign n33596 = ~n2872 & n33595 ;
  assign n33597 = n33596 ^ n2568 ^ 1'b0 ;
  assign n33600 = n33599 ^ n33597 ^ 1'b0 ;
  assign n33601 = n3033 & ~n9885 ;
  assign n33602 = n33601 ^ n6316 ^ 1'b0 ;
  assign n33603 = n12145 & n20517 ;
  assign n33604 = n33603 ^ n4719 ^ 1'b0 ;
  assign n33605 = n12348 & ~n13509 ;
  assign n33606 = n33605 ^ n27172 ^ 1'b0 ;
  assign n33607 = ( n4847 & n23592 ) | ( n4847 & n24093 ) | ( n23592 & n24093 ) ;
  assign n33608 = n29218 ^ n7603 ^ 1'b0 ;
  assign n33609 = n8063 & ~n10049 ;
  assign n33610 = ~n17768 & n33609 ;
  assign n33611 = n17107 ^ n3234 ^ 1'b0 ;
  assign n33612 = n22345 & ~n23674 ;
  assign n33613 = n11988 ^ n8019 ^ 1'b0 ;
  assign n33614 = ~n7757 & n33613 ;
  assign n33615 = n33614 ^ n5279 ^ 1'b0 ;
  assign n33616 = n1361 & n32918 ;
  assign n33617 = n4644 ^ n3214 ^ 1'b0 ;
  assign n33618 = n33617 ^ n31250 ^ 1'b0 ;
  assign n33619 = n3101 & n7082 ;
  assign n33620 = n27505 ^ n1529 ^ 1'b0 ;
  assign n33621 = ~n2207 & n33620 ;
  assign n33622 = n7468 & n8843 ;
  assign n33623 = n33622 ^ n10674 ^ 1'b0 ;
  assign n33624 = ( n3176 & n6660 ) | ( n3176 & n33623 ) | ( n6660 & n33623 ) ;
  assign n33625 = n1171 | n33624 ;
  assign n33626 = n33625 ^ n21543 ^ 1'b0 ;
  assign n33627 = n5295 & ~n10391 ;
  assign n33628 = n25349 ^ n4604 ^ n1000 ;
  assign n33629 = n33003 ^ n13703 ^ 1'b0 ;
  assign n33630 = n10315 ^ n8385 ^ 1'b0 ;
  assign n33631 = n12055 | n33630 ;
  assign n33632 = n33631 ^ n12133 ^ n4149 ;
  assign n33633 = n19844 ^ n112 ^ 1'b0 ;
  assign n33634 = n33633 ^ n28235 ^ n2106 ;
  assign n33635 = ~n8244 & n18295 ;
  assign n33636 = ~n9987 & n33635 ;
  assign n33637 = n12644 & ~n14675 ;
  assign n33638 = ~n20598 & n33637 ;
  assign n33639 = n317 & n4253 ;
  assign n33640 = n5252 ^ n750 ^ 1'b0 ;
  assign n33641 = ( n5725 & n14222 ) | ( n5725 & n33640 ) | ( n14222 & n33640 ) ;
  assign n33642 = n33641 ^ n801 ^ 1'b0 ;
  assign n33643 = ~n17956 & n33642 ;
  assign n33644 = n7317 ^ n179 ^ 1'b0 ;
  assign n33645 = n33644 ^ n16887 ^ 1'b0 ;
  assign n33646 = ~n17940 & n33645 ;
  assign n33647 = n7818 & ~n33646 ;
  assign n33648 = n33643 | n33647 ;
  assign n33649 = ~n33443 & n33648 ;
  assign n33650 = n6774 | n6819 ;
  assign n33651 = n11430 & n16761 ;
  assign n33652 = n33651 ^ n4490 ^ 1'b0 ;
  assign n33653 = ( n27342 & ~n33650 ) | ( n27342 & n33652 ) | ( ~n33650 & n33652 ) ;
  assign n33654 = n33653 ^ n18638 ^ n10229 ;
  assign n33655 = n18562 & n25687 ;
  assign n33656 = n21723 & n33655 ;
  assign n33657 = n23208 ^ n8416 ^ 1'b0 ;
  assign n33658 = n7976 & ~n33657 ;
  assign n33659 = n14401 | n25494 ;
  assign n33660 = n12543 | n26392 ;
  assign n33661 = n33660 ^ n21975 ^ 1'b0 ;
  assign n33662 = n22100 | n26463 ;
  assign n33663 = n33662 ^ n19265 ^ 1'b0 ;
  assign n33664 = n7026 ^ n3211 ^ 1'b0 ;
  assign n33665 = n5556 | n33664 ;
  assign n33666 = n33665 ^ n9716 ^ 1'b0 ;
  assign n33667 = ( n2913 & ~n8591 ) | ( n2913 & n16787 ) | ( ~n8591 & n16787 ) ;
  assign n33668 = n6374 & ~n33667 ;
  assign n33669 = n33668 ^ n3319 ^ 1'b0 ;
  assign n33670 = n27419 ^ n7240 ^ 1'b0 ;
  assign n33671 = n137 & ~n6979 ;
  assign n33672 = ~n20658 & n33671 ;
  assign n33673 = ( n10854 & n11567 ) | ( n10854 & ~n33672 ) | ( n11567 & ~n33672 ) ;
  assign n33674 = n24580 ^ n23258 ^ 1'b0 ;
  assign n33675 = n22051 | n33674 ;
  assign n33676 = n19097 ^ n15266 ^ 1'b0 ;
  assign n33678 = ~n8764 & n21495 ;
  assign n33677 = n20290 | n31968 ;
  assign n33679 = n33678 ^ n33677 ^ n3479 ;
  assign n33680 = n9893 & n33679 ;
  assign n33681 = n28475 & ~n29448 ;
  assign n33682 = n33681 ^ n934 ^ 1'b0 ;
  assign n33683 = n18742 ^ n7023 ^ 1'b0 ;
  assign n33684 = n19961 | n33683 ;
  assign n33685 = n23158 ^ n11994 ^ 1'b0 ;
  assign n33686 = n2697 | n19684 ;
  assign n33687 = n33686 ^ n2339 ^ 1'b0 ;
  assign n33689 = n12611 & ~n12682 ;
  assign n33690 = n33689 ^ n7762 ^ 1'b0 ;
  assign n33688 = n10345 & ~n26590 ;
  assign n33691 = n33690 ^ n33688 ^ 1'b0 ;
  assign n33692 = n27846 ^ n20654 ^ 1'b0 ;
  assign n33693 = n8218 ^ n8020 ^ 1'b0 ;
  assign n33694 = n6815 & n6833 ;
  assign n33695 = n1124 & ~n5656 ;
  assign n33696 = n33695 ^ n18242 ^ 1'b0 ;
  assign n33697 = n10366 & ~n33696 ;
  assign n33698 = n33697 ^ n23123 ^ 1'b0 ;
  assign n33699 = n11060 ^ n7001 ^ 1'b0 ;
  assign n33700 = ~n33698 & n33699 ;
  assign n33701 = n21441 ^ n4150 ^ 1'b0 ;
  assign n33702 = n17308 & n33701 ;
  assign n33703 = n15094 & ~n33702 ;
  assign n33704 = n7017 & n11363 ;
  assign n33705 = ~n3512 & n21480 ;
  assign n33706 = n5793 ^ n132 ^ 1'b0 ;
  assign n33707 = n33706 ^ n25590 ^ 1'b0 ;
  assign n33708 = n91 & ~n14775 ;
  assign n33709 = n22213 & n33708 ;
  assign n33710 = n22223 ^ n18109 ^ 1'b0 ;
  assign n33711 = n17249 & n18103 ;
  assign n33712 = n33710 | n33711 ;
  assign n33713 = n33712 ^ n22131 ^ 1'b0 ;
  assign n33714 = n33713 ^ n27348 ^ 1'b0 ;
  assign n33715 = n21568 ^ n19461 ^ 1'b0 ;
  assign n33716 = n4483 | n21529 ;
  assign n33717 = n33715 & ~n33716 ;
  assign n33718 = n5498 & n8780 ;
  assign n33719 = n3165 & ~n8816 ;
  assign n33720 = n21680 & n33719 ;
  assign n33721 = n3998 | n22260 ;
  assign n33722 = n33720 & ~n33721 ;
  assign n33723 = n33722 ^ n12589 ^ 1'b0 ;
  assign n33724 = n3622 | n15597 ;
  assign n33725 = n33724 ^ n20835 ^ n20340 ;
  assign n33726 = ~n23757 & n33725 ;
  assign n33727 = n28576 ^ n3330 ^ 1'b0 ;
  assign n33728 = n12451 & ~n33727 ;
  assign n33729 = ~n30502 & n33728 ;
  assign n33730 = ~n33726 & n33729 ;
  assign n33731 = n5172 & n5570 ;
  assign n33732 = n33731 ^ n17663 ^ 1'b0 ;
  assign n33733 = n21512 & n33732 ;
  assign n33734 = n33733 ^ n29437 ^ 1'b0 ;
  assign n33735 = ~n20529 & n33734 ;
  assign n33736 = n1024 & n20951 ;
  assign n33737 = ~n7882 & n12813 ;
  assign n33738 = ( n5809 & n33736 ) | ( n5809 & n33737 ) | ( n33736 & n33737 ) ;
  assign n33740 = ~n3308 & n12663 ;
  assign n33741 = n33740 ^ n6062 ^ 1'b0 ;
  assign n33742 = ~n4516 & n8215 ;
  assign n33743 = n33742 ^ n3508 ^ 1'b0 ;
  assign n33744 = n33741 & ~n33743 ;
  assign n33745 = n26571 & n33744 ;
  assign n33739 = n21148 ^ n3797 ^ 1'b0 ;
  assign n33746 = n33745 ^ n33739 ^ n17860 ;
  assign n33747 = n22 | n3915 ;
  assign n33748 = n26371 ^ n3097 ^ 1'b0 ;
  assign n33749 = n33747 & ~n33748 ;
  assign n33750 = n1787 & n9676 ;
  assign n33751 = n33749 & n33750 ;
  assign n33752 = n17016 ^ n4743 ^ 1'b0 ;
  assign n33753 = n33751 & n33752 ;
  assign n33755 = n8310 ^ n5975 ^ 1'b0 ;
  assign n33754 = n27916 | n28195 ;
  assign n33756 = n33755 ^ n33754 ^ 1'b0 ;
  assign n33757 = n1586 & ~n11074 ;
  assign n33758 = n33757 ^ n1871 ^ 1'b0 ;
  assign n33759 = ~n6099 & n33758 ;
  assign n33760 = n33759 ^ n6315 ^ 1'b0 ;
  assign n33761 = ~n33756 & n33760 ;
  assign n33762 = n33756 & n33761 ;
  assign n33763 = n998 | n22943 ;
  assign n33764 = n257 | n7129 ;
  assign n33765 = n33764 ^ n21555 ^ 1'b0 ;
  assign n33766 = n6477 & ~n33765 ;
  assign n33767 = ~n5675 & n33766 ;
  assign n33768 = n20389 ^ n11447 ^ 1'b0 ;
  assign n33769 = n18474 & n33768 ;
  assign n33770 = n30898 ^ n4002 ^ 1'b0 ;
  assign n33771 = n25157 | n33770 ;
  assign n33772 = n33769 & ~n33771 ;
  assign n33773 = n33772 ^ n4573 ^ 1'b0 ;
  assign n33774 = ~n957 & n8821 ;
  assign n33775 = n33774 ^ n28252 ^ 1'b0 ;
  assign n33776 = n22532 ^ n4536 ^ n4405 ;
  assign n33777 = n33776 ^ n14023 ^ 1'b0 ;
  assign n33778 = n22313 | n33777 ;
  assign n33779 = ( ~n3127 & n33775 ) | ( ~n3127 & n33778 ) | ( n33775 & n33778 ) ;
  assign n33780 = ( n1603 & n24912 ) | ( n1603 & ~n33779 ) | ( n24912 & ~n33779 ) ;
  assign n33781 = n24814 | n33780 ;
  assign n33782 = n33781 ^ n26243 ^ 1'b0 ;
  assign n33783 = n14644 ^ n11856 ^ x3 ;
  assign n33784 = n33783 ^ n1055 ^ 1'b0 ;
  assign n33785 = n12644 & ~n33784 ;
  assign n33786 = n33785 ^ n28933 ^ 1'b0 ;
  assign n33787 = n2354 ^ n1050 ^ 1'b0 ;
  assign n33788 = n469 | n33787 ;
  assign n33789 = ( n24452 & n33786 ) | ( n24452 & n33788 ) | ( n33786 & n33788 ) ;
  assign n33790 = n6532 & n11072 ;
  assign n33791 = n33790 ^ n5769 ^ 1'b0 ;
  assign n33792 = n33791 ^ n23946 ^ n17578 ;
  assign n33793 = n33003 ^ n29681 ^ n29056 ;
  assign n33794 = n4872 & n24408 ;
  assign n33795 = n33794 ^ n21471 ^ 1'b0 ;
  assign n33796 = ~n13060 & n33795 ;
  assign n33797 = n14811 ^ n7349 ^ 1'b0 ;
  assign n33798 = n296 | n33797 ;
  assign n33799 = ~n16201 & n32195 ;
  assign n33800 = n33799 ^ n32196 ^ 1'b0 ;
  assign n33801 = n22479 ^ n5113 ^ 1'b0 ;
  assign n33802 = n1641 & ~n6211 ;
  assign n33803 = n33802 ^ n10816 ^ 1'b0 ;
  assign n33804 = n33803 ^ n22332 ^ n2823 ;
  assign n33805 = n11769 ^ n10731 ^ 1'b0 ;
  assign n33806 = ( n12554 & n20036 ) | ( n12554 & n25024 ) | ( n20036 & n25024 ) ;
  assign n33807 = n22913 ^ n15403 ^ 1'b0 ;
  assign n33808 = n17024 & n33807 ;
  assign n33809 = n10063 & ~n17743 ;
  assign n33810 = ~n25521 & n33809 ;
  assign n33811 = n33810 ^ n6126 ^ n5387 ;
  assign n33812 = n33811 ^ n18493 ^ n3706 ;
  assign n33813 = n28600 ^ n20646 ^ n725 ;
  assign n33814 = n33813 ^ n15626 ^ 1'b0 ;
  assign n33815 = n21912 ^ n18151 ^ 1'b0 ;
  assign n33816 = n32650 ^ n6099 ^ 1'b0 ;
  assign n33817 = n2528 | n11202 ;
  assign n33818 = n23278 & n28358 ;
  assign n33819 = n29144 & n33818 ;
  assign n33820 = n19919 | n26586 ;
  assign n33821 = n7499 ^ n3130 ^ n928 ;
  assign n33822 = n2747 | n33821 ;
  assign n33823 = n33822 ^ n102 ^ 1'b0 ;
  assign n33824 = n33823 ^ n9075 ^ 1'b0 ;
  assign n33825 = n23446 ^ n17285 ^ 1'b0 ;
  assign n33826 = n17693 & ~n33825 ;
  assign n33827 = n4052 ^ x10 ^ 1'b0 ;
  assign n33828 = ~n7285 & n29091 ;
  assign n33829 = n12728 & ~n30786 ;
  assign n33830 = n33829 ^ n1546 ^ 1'b0 ;
  assign n33831 = n14146 ^ n10436 ^ 1'b0 ;
  assign n33832 = n22677 | n33831 ;
  assign n33833 = n33832 ^ n2841 ^ 1'b0 ;
  assign n33834 = n2330 & ~n12479 ;
  assign n33835 = n33359 ^ n3064 ^ 1'b0 ;
  assign n33836 = n10088 & n33835 ;
  assign n33837 = n33834 & n33836 ;
  assign n33838 = n33441 ^ n24240 ^ n10665 ;
  assign n33839 = n15632 | n17520 ;
  assign n33840 = n17520 & ~n33839 ;
  assign n33841 = n4548 & ~n26289 ;
  assign n33842 = n33841 ^ n2077 ^ 1'b0 ;
  assign n33843 = n33842 ^ n23285 ^ 1'b0 ;
  assign n33844 = ( n4968 & n17085 ) | ( n4968 & n33843 ) | ( n17085 & n33843 ) ;
  assign n33845 = ( ~n20727 & n33840 ) | ( ~n20727 & n33844 ) | ( n33840 & n33844 ) ;
  assign n33846 = n2653 | n9408 ;
  assign n33847 = n33846 ^ n2710 ^ 1'b0 ;
  assign n33848 = n3517 & ~n10181 ;
  assign n33849 = ~n7681 & n33848 ;
  assign n33850 = n33847 & n33849 ;
  assign n33851 = ~n18950 & n33850 ;
  assign n33852 = n20970 ^ n17637 ^ 1'b0 ;
  assign n33853 = ~n15879 & n33852 ;
  assign n33854 = ~n23548 & n33853 ;
  assign n33856 = ~n19190 & n21675 ;
  assign n33855 = ~n12718 & n16339 ;
  assign n33857 = n33856 ^ n33855 ^ 1'b0 ;
  assign n33858 = n7190 | n14226 ;
  assign n33859 = n1307 & n6985 ;
  assign n33860 = n4957 | n12731 ;
  assign n33861 = n33859 & ~n33860 ;
  assign n33862 = n16403 & ~n33861 ;
  assign n33863 = n33858 & n33862 ;
  assign n33864 = n33863 ^ n2432 ^ n431 ;
  assign n33865 = n11854 ^ n3943 ^ 1'b0 ;
  assign n33866 = n33865 ^ n383 ^ 1'b0 ;
  assign n33867 = n4009 | n33866 ;
  assign n33868 = n17384 & ~n33867 ;
  assign n33869 = ~n6790 & n9568 ;
  assign n33870 = n12171 & n33869 ;
  assign n33871 = n33870 ^ n21620 ^ 1'b0 ;
  assign n33872 = n10488 & ~n11919 ;
  assign n33873 = n33872 ^ n5639 ^ 1'b0 ;
  assign n33874 = ~n18600 & n33873 ;
  assign n33875 = n19364 ^ n6951 ^ 1'b0 ;
  assign n33876 = n33875 ^ n13863 ^ n8614 ;
  assign n33877 = n9755 & ~n15993 ;
  assign n33878 = n26983 & n33877 ;
  assign n33879 = ( n5481 & n8356 ) | ( n5481 & ~n22239 ) | ( n8356 & ~n22239 ) ;
  assign n33880 = n17690 | n17983 ;
  assign n33881 = n5599 & ~n33880 ;
  assign n33882 = ( n12794 & n25716 ) | ( n12794 & ~n33881 ) | ( n25716 & ~n33881 ) ;
  assign n33883 = n33882 ^ n5200 ^ 1'b0 ;
  assign n33884 = n33879 & n33883 ;
  assign n33885 = n16818 ^ n9459 ^ n1457 ;
  assign n33886 = n33885 ^ n29898 ^ n10235 ;
  assign n33887 = n15511 ^ n14757 ^ n6644 ;
  assign n33888 = n205 | n26637 ;
  assign n33889 = n33888 ^ n464 ^ 1'b0 ;
  assign n33890 = n16475 ^ n12384 ^ 1'b0 ;
  assign n33891 = ~n2350 & n20713 ;
  assign n33892 = ~n33890 & n33891 ;
  assign n33893 = n2797 | n13143 ;
  assign n33894 = ~n11521 & n33893 ;
  assign n33895 = n33894 ^ n30060 ^ 1'b0 ;
  assign n33896 = ~n2165 & n3950 ;
  assign n33897 = n27001 & ~n33896 ;
  assign n33898 = n33897 ^ n29678 ^ 1'b0 ;
  assign n33899 = n21999 ^ n10260 ^ n1600 ;
  assign n33900 = n33899 ^ n4965 ^ 1'b0 ;
  assign n33901 = ~n33898 & n33900 ;
  assign n33902 = ( n21299 & n29880 ) | ( n21299 & n33901 ) | ( n29880 & n33901 ) ;
  assign n33903 = n11607 ^ n5730 ^ 1'b0 ;
  assign n33904 = n14175 & n19165 ;
  assign n33905 = ~n11128 & n33904 ;
  assign n33906 = n6186 & ~n33905 ;
  assign n33907 = n13663 & n33906 ;
  assign n33908 = n448 & ~n6682 ;
  assign n33909 = n9386 ^ n8327 ^ 1'b0 ;
  assign n33910 = n15946 & ~n33909 ;
  assign n33911 = n33910 ^ n17364 ^ 1'b0 ;
  assign n33912 = n30297 ^ n15737 ^ 1'b0 ;
  assign n33913 = n5583 | n33912 ;
  assign n33914 = n33913 ^ n18315 ^ 1'b0 ;
  assign n33915 = n6102 | n32924 ;
  assign n33918 = n21724 ^ n9195 ^ 1'b0 ;
  assign n33916 = n11984 & ~n22081 ;
  assign n33917 = n22335 | n33916 ;
  assign n33919 = n33918 ^ n33917 ^ 1'b0 ;
  assign n33920 = n8222 ^ n3953 ^ 1'b0 ;
  assign n33921 = ~n33919 & n33920 ;
  assign n33922 = n13206 ^ n1188 ^ 1'b0 ;
  assign n33923 = n15487 | n33922 ;
  assign n33924 = n15173 ^ n7428 ^ 1'b0 ;
  assign n33925 = ~n33923 & n33924 ;
  assign n33926 = n33084 ^ n30427 ^ n4785 ;
  assign n33928 = n445 & ~n448 ;
  assign n33929 = n2896 & n33928 ;
  assign n33930 = n6412 | n7687 ;
  assign n33931 = n33929 & ~n33930 ;
  assign n33932 = n13011 | n33931 ;
  assign n33933 = n33932 ^ n838 ^ 1'b0 ;
  assign n33927 = n28255 & ~n33584 ;
  assign n33934 = n33933 ^ n33927 ^ 1'b0 ;
  assign n33935 = n4915 & n33934 ;
  assign n33936 = n15523 & n26049 ;
  assign n33937 = ~n7753 & n33936 ;
  assign n33938 = n29426 ^ n13937 ^ 1'b0 ;
  assign n33939 = n8274 & ~n33938 ;
  assign n33940 = n33939 ^ n1744 ^ 1'b0 ;
  assign n33941 = n13131 | n13818 ;
  assign n33942 = n33941 ^ n1700 ^ 1'b0 ;
  assign n33943 = ( n2186 & n33443 ) | ( n2186 & n33942 ) | ( n33443 & n33942 ) ;
  assign n33944 = n25777 ^ n4804 ^ 1'b0 ;
  assign n33945 = n10843 ^ n1009 ^ 1'b0 ;
  assign n33946 = n19204 ^ n5394 ^ 1'b0 ;
  assign n33947 = n17134 ^ n4896 ^ n1571 ;
  assign n33948 = n33947 ^ n2738 ^ 1'b0 ;
  assign n33949 = n14949 | n33948 ;
  assign n33950 = n33949 ^ n15136 ^ 1'b0 ;
  assign n33951 = n28763 ^ n18902 ^ 1'b0 ;
  assign n33952 = n33950 | n33951 ;
  assign n33953 = n14917 ^ n14312 ^ 1'b0 ;
  assign n33954 = n33953 ^ n9917 ^ 1'b0 ;
  assign n33955 = n4838 ^ n1121 ^ 1'b0 ;
  assign n33956 = n5913 | n33955 ;
  assign n33957 = n25402 ^ n5509 ^ 1'b0 ;
  assign n33958 = n33957 ^ n22772 ^ 1'b0 ;
  assign n33959 = n33956 & ~n33958 ;
  assign n33960 = n15999 & ~n24539 ;
  assign n33961 = n14832 & n33960 ;
  assign n33962 = n12959 | n33961 ;
  assign n33963 = n6008 & ~n33962 ;
  assign n33964 = ( n4402 & n17895 ) | ( n4402 & n33963 ) | ( n17895 & n33963 ) ;
  assign n33965 = ( n2677 & n5924 ) | ( n2677 & ~n6064 ) | ( n5924 & ~n6064 ) ;
  assign n33966 = n33965 ^ n10772 ^ 1'b0 ;
  assign n33967 = ~n3773 & n31727 ;
  assign n33968 = ~n14483 & n16455 ;
  assign n33969 = n33968 ^ n22700 ^ 1'b0 ;
  assign n33970 = n31881 ^ n15512 ^ n3174 ;
  assign n33971 = ~n20298 & n33970 ;
  assign n33972 = ( n224 & n5966 ) | ( n224 & ~n31992 ) | ( n5966 & ~n31992 ) ;
  assign n33973 = n2571 ^ n37 ^ 1'b0 ;
  assign n33974 = ~n2808 & n33973 ;
  assign n33975 = n18145 ^ n16481 ^ n2114 ;
  assign n33976 = n17366 ^ n3833 ^ 1'b0 ;
  assign n33977 = ~n4964 & n31224 ;
  assign n33978 = ~n3713 & n33977 ;
  assign n33979 = n13277 ^ n6524 ^ 1'b0 ;
  assign n33980 = n33979 ^ n2571 ^ 1'b0 ;
  assign n33981 = ~n21160 & n33980 ;
  assign n33982 = ( n2713 & ~n19642 ) | ( n2713 & n29298 ) | ( ~n19642 & n29298 ) ;
  assign n33983 = n31459 ^ n17675 ^ 1'b0 ;
  assign n33984 = n25983 ^ n17096 ^ 1'b0 ;
  assign n33985 = n16473 & ~n33984 ;
  assign n33986 = n15078 | n31180 ;
  assign n33987 = n10125 | n33986 ;
  assign n33988 = n6490 & ~n23743 ;
  assign n33989 = n33988 ^ n23974 ^ 1'b0 ;
  assign n33990 = n5327 | n23886 ;
  assign n33991 = n27916 ^ n5048 ^ 1'b0 ;
  assign n33992 = n19352 | n33991 ;
  assign n33993 = n3891 | n16832 ;
  assign n33994 = n33993 ^ n3791 ^ 1'b0 ;
  assign n33995 = ( n711 & ~n11288 ) | ( n711 & n33994 ) | ( ~n11288 & n33994 ) ;
  assign n33996 = n13699 ^ n4642 ^ 1'b0 ;
  assign n33997 = n7516 & n33996 ;
  assign n33998 = n4112 ^ n3563 ^ 1'b0 ;
  assign n33999 = n31548 & ~n33998 ;
  assign n34000 = n21052 ^ n1400 ^ 1'b0 ;
  assign n34001 = n9357 & ~n13876 ;
  assign n34002 = ~n22806 & n34001 ;
  assign n34003 = n34000 & n34002 ;
  assign n34004 = n1505 | n20529 ;
  assign n34005 = n34004 ^ n14854 ^ 1'b0 ;
  assign n34006 = n34005 ^ n26593 ^ n11113 ;
  assign n34007 = ~n5808 & n7707 ;
  assign n34008 = n217 & n34007 ;
  assign n34009 = n34008 ^ n18632 ^ n5627 ;
  assign n34010 = n21980 ^ n7392 ^ 1'b0 ;
  assign n34011 = n2811 | n34010 ;
  assign n34012 = n29231 & ~n34011 ;
  assign n34013 = n15277 ^ n10962 ^ 1'b0 ;
  assign n34014 = n1853 & n34013 ;
  assign n34015 = n4095 | n7494 ;
  assign n34016 = n34015 ^ n12682 ^ 1'b0 ;
  assign n34017 = n13945 & ~n34016 ;
  assign n34018 = n6947 & ~n13233 ;
  assign n34019 = ( n2982 & ~n3092 ) | ( n2982 & n5168 ) | ( ~n3092 & n5168 ) ;
  assign n34020 = ( n1522 & ~n34018 ) | ( n1522 & n34019 ) | ( ~n34018 & n34019 ) ;
  assign n34021 = n8683 & ~n19733 ;
  assign n34022 = n34021 ^ n32932 ^ 1'b0 ;
  assign n34023 = ~n17122 & n34022 ;
  assign n34024 = n30110 ^ n11876 ^ n10438 ;
  assign n34025 = n34024 ^ n29154 ^ n13642 ;
  assign n34026 = n13743 & ~n27159 ;
  assign n34027 = ~n8469 & n15072 ;
  assign n34028 = ~n28592 & n34027 ;
  assign n34029 = n34028 ^ n30158 ^ 1'b0 ;
  assign n34030 = n11668 & ~n34029 ;
  assign n34031 = ~n5740 & n16440 ;
  assign n34032 = n12874 & n18420 ;
  assign n34033 = n34032 ^ n493 ^ 1'b0 ;
  assign n34034 = n25157 ^ n21190 ^ 1'b0 ;
  assign n34035 = n22586 ^ n9072 ^ 1'b0 ;
  assign n34036 = n30529 ^ n4079 ^ 1'b0 ;
  assign n34037 = n34035 & n34036 ;
  assign n34038 = n34037 ^ n1569 ^ 1'b0 ;
  assign n34039 = n8203 & n23985 ;
  assign n34040 = n6527 | n8449 ;
  assign n34041 = n1693 & n26105 ;
  assign n34042 = n22854 | n34041 ;
  assign n34043 = ~n3554 & n34042 ;
  assign n34044 = ~n34040 & n34043 ;
  assign n34045 = n13007 ^ n691 ^ 1'b0 ;
  assign n34046 = n12469 & ~n34045 ;
  assign n34047 = ~n19605 & n34046 ;
  assign n34048 = n32661 ^ n18945 ^ n11749 ;
  assign n34049 = n17991 ^ n14419 ^ 1'b0 ;
  assign n34050 = ( ~n1075 & n29072 ) | ( ~n1075 & n30127 ) | ( n29072 & n30127 ) ;
  assign n34051 = ~n7666 & n34050 ;
  assign n34052 = n8655 | n34051 ;
  assign n34053 = n31591 ^ n11593 ^ 1'b0 ;
  assign n34054 = n6029 | n12183 ;
  assign n34055 = n7728 | n34054 ;
  assign n34056 = n8587 | n9790 ;
  assign n34057 = n34056 ^ n18733 ^ 1'b0 ;
  assign n34058 = n1454 & ~n3174 ;
  assign n34059 = n2170 & n34058 ;
  assign n34060 = n12734 | n34059 ;
  assign n34061 = ~n13990 & n32268 ;
  assign n34062 = n34061 ^ n28236 ^ 1'b0 ;
  assign n34063 = ( ~n15918 & n26780 ) | ( ~n15918 & n28398 ) | ( n26780 & n28398 ) ;
  assign n34064 = ( ~n2271 & n28901 ) | ( ~n2271 & n32266 ) | ( n28901 & n32266 ) ;
  assign n34065 = n20336 ^ n10284 ^ n4629 ;
  assign n34066 = n1912 & n10269 ;
  assign n34067 = n2623 ^ n1569 ^ 1'b0 ;
  assign n34068 = n34066 | n34067 ;
  assign n34069 = n34068 ^ n825 ^ 1'b0 ;
  assign n34070 = n19811 & n34069 ;
  assign n34071 = n34070 ^ n31174 ^ 1'b0 ;
  assign n34072 = ~n25413 & n27551 ;
  assign n34073 = n34072 ^ n11321 ^ 1'b0 ;
  assign n34074 = n3430 | n34073 ;
  assign n34075 = n8597 | n15914 ;
  assign n34078 = n252 ^ n213 ^ 1'b0 ;
  assign n34079 = ( n15830 & ~n20221 ) | ( n15830 & n34078 ) | ( ~n20221 & n34078 ) ;
  assign n34076 = n6872 & ~n8166 ;
  assign n34077 = n22610 | n34076 ;
  assign n34080 = n34079 ^ n34077 ^ 1'b0 ;
  assign n34081 = n22321 | n34080 ;
  assign n34082 = n21244 & n32820 ;
  assign n34083 = n34082 ^ n15483 ^ 1'b0 ;
  assign n34084 = n23363 ^ n1688 ^ 1'b0 ;
  assign n34085 = n8341 & n34084 ;
  assign n34086 = n34085 ^ n517 ^ 1'b0 ;
  assign n34087 = n4264 ^ n3284 ^ n1775 ;
  assign n34088 = n30901 ^ n6841 ^ 1'b0 ;
  assign n34089 = ~n4884 & n34088 ;
  assign n34090 = ( n23603 & n34087 ) | ( n23603 & n34089 ) | ( n34087 & n34089 ) ;
  assign n34091 = n2464 | n31853 ;
  assign n34092 = n1234 & ~n14650 ;
  assign n34093 = n28728 ^ n8806 ^ 1'b0 ;
  assign n34094 = n17207 & ~n34093 ;
  assign n34095 = n2357 ^ n1828 ^ 1'b0 ;
  assign n34096 = n34095 ^ n18248 ^ n4428 ;
  assign n34097 = n8458 & n34096 ;
  assign n34098 = n14661 & n32606 ;
  assign n34099 = n34097 & n34098 ;
  assign n34100 = n15733 & n22915 ;
  assign n34101 = ~n17308 & n34100 ;
  assign n34102 = ~n7003 & n34101 ;
  assign n34103 = n680 & ~n11321 ;
  assign n34104 = n14952 ^ n11372 ^ n334 ;
  assign n34105 = n23801 & ~n26791 ;
  assign n34106 = n11789 ^ n4647 ^ 1'b0 ;
  assign n34107 = ( n12715 & n15470 ) | ( n12715 & n22566 ) | ( n15470 & n22566 ) ;
  assign n34108 = n5617 & n13470 ;
  assign n34109 = n32984 & n34108 ;
  assign n34110 = n3146 & ~n4602 ;
  assign n34111 = ~n8746 & n34110 ;
  assign n34112 = ( n4761 & ~n10491 ) | ( n4761 & n14073 ) | ( ~n10491 & n14073 ) ;
  assign n34113 = n34111 & n34112 ;
  assign n34114 = n8271 ^ n6264 ^ 1'b0 ;
  assign n34115 = n23452 | n34114 ;
  assign n34116 = n22950 & ~n34115 ;
  assign n34117 = n8557 ^ n4638 ^ 1'b0 ;
  assign n34118 = n23407 ^ n3671 ^ 1'b0 ;
  assign n34119 = ~n3105 & n8833 ;
  assign n34120 = n25315 & n34119 ;
  assign n34121 = ~n1628 & n7694 ;
  assign n34122 = ~n725 & n34121 ;
  assign n34123 = n20716 | n34122 ;
  assign n34124 = n34120 & ~n34123 ;
  assign n34126 = n16131 ^ n10131 ^ 1'b0 ;
  assign n34127 = n5392 & n34126 ;
  assign n34128 = n2128 & n34127 ;
  assign n34129 = n34128 ^ n7460 ^ 1'b0 ;
  assign n34130 = ~n1689 & n17042 ;
  assign n34131 = ~n34129 & n34130 ;
  assign n34132 = n12752 | n34131 ;
  assign n34125 = ~n9835 & n11292 ;
  assign n34133 = n34132 ^ n34125 ^ 1'b0 ;
  assign n34134 = n32045 ^ n7643 ^ 1'b0 ;
  assign n34135 = n21550 ^ n12901 ^ 1'b0 ;
  assign n34136 = ~n592 & n11402 ;
  assign n34137 = ~n34135 & n34136 ;
  assign n34138 = n34137 ^ n32393 ^ n29069 ;
  assign n34139 = n29316 ^ n11490 ^ 1'b0 ;
  assign n34140 = n33265 ^ n7686 ^ 1'b0 ;
  assign n34141 = n16286 & n34140 ;
  assign n34142 = n26426 ^ n9986 ^ 1'b0 ;
  assign n34143 = n11036 ^ n8616 ^ 1'b0 ;
  assign n34144 = n34143 ^ n26741 ^ n3105 ;
  assign n34145 = n15589 & n23014 ;
  assign n34146 = n24875 & ~n34145 ;
  assign n34147 = ~n34144 & n34146 ;
  assign n34148 = n29658 ^ n25089 ^ 1'b0 ;
  assign n34149 = n25425 & n34148 ;
  assign n34150 = ( n1563 & ~n2986 ) | ( n1563 & n8787 ) | ( ~n2986 & n8787 ) ;
  assign n34151 = n29900 & n34150 ;
  assign n34152 = ~n12438 & n27829 ;
  assign n34153 = ~n9636 & n34152 ;
  assign n34154 = n7019 & n33108 ;
  assign n34155 = n30938 ^ n30092 ^ 1'b0 ;
  assign n34156 = ~n16149 & n21127 ;
  assign n34157 = n1654 & n34156 ;
  assign n34158 = n7347 | n34157 ;
  assign n34159 = n34158 ^ n10284 ^ 1'b0 ;
  assign n34160 = n22085 ^ n7376 ^ 1'b0 ;
  assign n34161 = n30516 & ~n34160 ;
  assign n34162 = ~n13117 & n16716 ;
  assign n34163 = n34162 ^ n31445 ^ 1'b0 ;
  assign n34164 = n5210 & ~n34163 ;
  assign n34165 = ( n21454 & n32521 ) | ( n21454 & ~n34164 ) | ( n32521 & ~n34164 ) ;
  assign n34166 = n850 & n17828 ;
  assign n34167 = n34166 ^ n5626 ^ 1'b0 ;
  assign n34168 = n14385 ^ n70 ^ 1'b0 ;
  assign n34169 = n12310 & ~n34168 ;
  assign n34170 = n10999 ^ n9165 ^ 1'b0 ;
  assign n34171 = n17109 | n34170 ;
  assign n34172 = n4016 & n22760 ;
  assign n34173 = n28532 ^ n11081 ^ 1'b0 ;
  assign n34174 = n10273 ^ n10247 ^ 1'b0 ;
  assign n34175 = n34173 & n34174 ;
  assign n34176 = n16440 & ~n34175 ;
  assign n34177 = n14680 & ~n21990 ;
  assign n34178 = ~n10892 & n20226 ;
  assign n34179 = ( n5628 & n10240 ) | ( n5628 & n34178 ) | ( n10240 & n34178 ) ;
  assign n34180 = n6091 ^ n2243 ^ 1'b0 ;
  assign n34181 = ~n1240 & n34180 ;
  assign n34182 = n34181 ^ n209 ^ 1'b0 ;
  assign n34183 = n34182 ^ n24079 ^ n2994 ;
  assign n34184 = n16691 | n18855 ;
  assign n34185 = n3407 | n34184 ;
  assign n34186 = n578 & ~n24652 ;
  assign n34187 = ~n12317 & n34186 ;
  assign n34188 = n3266 & ~n32661 ;
  assign n34189 = n835 & n34188 ;
  assign n34190 = n3116 & n22788 ;
  assign n34191 = n11774 | n29081 ;
  assign n34192 = n11187 & n24263 ;
  assign n34193 = n34192 ^ n7374 ^ 1'b0 ;
  assign n34194 = n30515 ^ n676 ^ 1'b0 ;
  assign n34195 = n27975 & n34194 ;
  assign n34196 = n18911 | n34157 ;
  assign n34197 = n6992 | n24996 ;
  assign n34198 = n34197 ^ n12644 ^ 1'b0 ;
  assign n34201 = n10974 ^ n1418 ^ n1314 ;
  assign n34199 = ~n16168 & n23364 ;
  assign n34200 = n5042 & n34199 ;
  assign n34202 = n34201 ^ n34200 ^ n17001 ;
  assign n34203 = n16871 & ~n26172 ;
  assign n34204 = n34203 ^ n7441 ^ 1'b0 ;
  assign n34205 = n4742 ^ n26 ^ 1'b0 ;
  assign n34206 = n31097 | n34205 ;
  assign n34207 = n34206 ^ n9492 ^ n7391 ;
  assign n34208 = n15423 & ~n34207 ;
  assign n34209 = n34208 ^ n19072 ^ 1'b0 ;
  assign n34210 = n353 & n29575 ;
  assign n34211 = n34210 ^ n2620 ^ 1'b0 ;
  assign n34212 = n6120 & ~n18631 ;
  assign n34213 = n22088 ^ n11772 ^ 1'b0 ;
  assign n34214 = n34212 & n34213 ;
  assign n34215 = n2245 & ~n10707 ;
  assign n34216 = n34215 ^ n17493 ^ n1521 ;
  assign n34219 = n15176 | n28206 ;
  assign n34217 = n25357 ^ n20453 ^ 1'b0 ;
  assign n34218 = n3461 | n34217 ;
  assign n34220 = n34219 ^ n34218 ^ n965 ;
  assign n34221 = n12530 ^ n823 ^ 1'b0 ;
  assign n34222 = ~n29287 & n34221 ;
  assign n34223 = ~n4367 & n11029 ;
  assign n34224 = n15643 & n34223 ;
  assign n34225 = n15819 ^ n11973 ^ 1'b0 ;
  assign n34226 = n9199 ^ n7406 ^ 1'b0 ;
  assign n34227 = ( n8055 & ~n31570 ) | ( n8055 & n34226 ) | ( ~n31570 & n34226 ) ;
  assign n34228 = n24474 ^ n1511 ^ 1'b0 ;
  assign n34230 = n7763 & ~n8489 ;
  assign n34231 = n34230 ^ n704 ^ 1'b0 ;
  assign n34229 = n22332 ^ n6931 ^ 1'b0 ;
  assign n34232 = n34231 ^ n34229 ^ n8039 ;
  assign n34233 = n7874 & n26124 ;
  assign n34234 = n34232 & n34233 ;
  assign n34235 = n1581 | n26224 ;
  assign n34236 = n9817 & ~n34235 ;
  assign n34237 = n34236 ^ n879 ^ 1'b0 ;
  assign n34238 = n5016 & ~n18401 ;
  assign n34239 = n34238 ^ n3401 ^ 1'b0 ;
  assign n34240 = n5791 ^ n3351 ^ n2609 ;
  assign n34241 = ( n686 & n5878 ) | ( n686 & ~n34240 ) | ( n5878 & ~n34240 ) ;
  assign n34242 = n3079 & ~n4034 ;
  assign n34243 = ~n27738 & n28705 ;
  assign n34244 = ~n26762 & n34243 ;
  assign n34245 = n28191 ^ n25812 ^ 1'b0 ;
  assign n34246 = n12932 & n34245 ;
  assign n34247 = n34246 ^ n16826 ^ n9446 ;
  assign n34248 = n10681 ^ n4205 ^ 1'b0 ;
  assign n34249 = ~n12360 & n34248 ;
  assign n34250 = n9304 & n34249 ;
  assign n34251 = ~n9781 & n34250 ;
  assign n34252 = n13632 | n14459 ;
  assign n34253 = ( n1436 & n34251 ) | ( n1436 & ~n34252 ) | ( n34251 & ~n34252 ) ;
  assign n34254 = n10541 | n30199 ;
  assign n34255 = n4523 & ~n34254 ;
  assign n34256 = n15819 | n19795 ;
  assign n34257 = n16666 & n17923 ;
  assign n34258 = ~n4695 & n34257 ;
  assign n34259 = n22473 ^ n3069 ^ n733 ;
  assign n34263 = ~n285 & n14297 ;
  assign n34264 = n5740 & n34263 ;
  assign n34265 = n20602 | n34264 ;
  assign n34260 = ~n3138 & n20535 ;
  assign n34261 = n34260 ^ n8647 ^ 1'b0 ;
  assign n34262 = n12958 | n34261 ;
  assign n34266 = n34265 ^ n34262 ^ n4932 ;
  assign n34267 = n34266 ^ n7159 ^ 1'b0 ;
  assign n34268 = ~n34259 & n34267 ;
  assign n34269 = ~n2954 & n34268 ;
  assign n34270 = n6771 ^ n6541 ^ 1'b0 ;
  assign n34271 = n28065 ^ n6430 ^ 1'b0 ;
  assign n34272 = ( n10526 & n28118 ) | ( n10526 & n29860 ) | ( n28118 & n29860 ) ;
  assign n34273 = n34272 ^ n23302 ^ 1'b0 ;
  assign n34274 = ~n9580 & n34273 ;
  assign n34275 = n34274 ^ n31439 ^ 1'b0 ;
  assign n34276 = n34271 & ~n34275 ;
  assign n34277 = ~n1312 & n16559 ;
  assign n34278 = ( ~n10383 & n14238 ) | ( ~n10383 & n34277 ) | ( n14238 & n34277 ) ;
  assign n34279 = n12423 & n34278 ;
  assign n34280 = n4982 & n34279 ;
  assign n34281 = n17694 ^ n8232 ^ 1'b0 ;
  assign n34282 = n514 & ~n34281 ;
  assign n34283 = ~n15748 & n34282 ;
  assign n34284 = n9332 & ~n33212 ;
  assign n34285 = ~n34283 & n34284 ;
  assign n34286 = n9346 | n13567 ;
  assign n34287 = n34286 ^ n26833 ^ n18055 ;
  assign n34288 = n13732 ^ n9591 ^ n1602 ;
  assign n34289 = ( ~n7585 & n15579 ) | ( ~n7585 & n34288 ) | ( n15579 & n34288 ) ;
  assign n34290 = n1150 | n10815 ;
  assign n34291 = ( n1969 & ~n5643 ) | ( n1969 & n12672 ) | ( ~n5643 & n12672 ) ;
  assign n34292 = ~n10652 & n25103 ;
  assign n34293 = n34291 & n34292 ;
  assign n34294 = n34290 & n34293 ;
  assign n34295 = n30107 ^ n13102 ^ n3466 ;
  assign n34296 = n34295 ^ n17993 ^ 1'b0 ;
  assign n34297 = n7539 & ~n7965 ;
  assign n34298 = n34297 ^ n13084 ^ 1'b0 ;
  assign n34299 = n10263 & ~n34298 ;
  assign n34300 = n34299 ^ n33083 ^ 1'b0 ;
  assign n34301 = n12180 | n30388 ;
  assign n34303 = n2139 & ~n15136 ;
  assign n34304 = n15136 & n34303 ;
  assign n34302 = ~n14193 & n31426 ;
  assign n34305 = n34304 ^ n34302 ^ 1'b0 ;
  assign n34306 = n16236 | n34305 ;
  assign n34307 = n16282 ^ n15678 ^ n1540 ;
  assign n34308 = n34306 | n34307 ;
  assign n34309 = n34308 ^ n7388 ^ 1'b0 ;
  assign n34310 = n27954 ^ n203 ^ 1'b0 ;
  assign n34311 = n2146 & n12854 ;
  assign n34312 = n3124 & ~n34311 ;
  assign n34313 = ( n21624 & ~n28884 ) | ( n21624 & n34312 ) | ( ~n28884 & n34312 ) ;
  assign n34314 = n14404 & n28270 ;
  assign n34315 = n34314 ^ n29334 ^ 1'b0 ;
  assign n34316 = n28224 | n34315 ;
  assign n34317 = n4810 & n20801 ;
  assign n34318 = n8651 | n8906 ;
  assign n34319 = n34318 ^ n4212 ^ 1'b0 ;
  assign n34320 = n34319 ^ n4339 ^ 1'b0 ;
  assign n34321 = ~n2359 & n34320 ;
  assign n34322 = ~n34317 & n34321 ;
  assign n34323 = n16460 & ~n32437 ;
  assign n34324 = n7404 & n34323 ;
  assign n34327 = n9497 | n13270 ;
  assign n34325 = n12465 & n21730 ;
  assign n34326 = n34325 ^ n6816 ^ 1'b0 ;
  assign n34328 = n34327 ^ n34326 ^ 1'b0 ;
  assign n34329 = ~n5394 & n27092 ;
  assign n34330 = n34329 ^ n31505 ^ n10143 ;
  assign n34331 = n4275 ^ n667 ^ 1'b0 ;
  assign n34332 = ~n25396 & n34331 ;
  assign n34333 = n4459 & n34332 ;
  assign n34335 = ~n5231 & n7404 ;
  assign n34334 = n2262 & ~n3109 ;
  assign n34336 = n34335 ^ n34334 ^ 1'b0 ;
  assign n34337 = n25965 ^ n6076 ^ 1'b0 ;
  assign n34338 = n34337 ^ n3341 ^ 1'b0 ;
  assign n34339 = n3574 | n34338 ;
  assign n34340 = n34339 ^ n21318 ^ 1'b0 ;
  assign n34341 = ~n14100 & n32275 ;
  assign n34342 = ~n6591 & n34341 ;
  assign n34343 = n33696 ^ n8547 ^ 1'b0 ;
  assign n34344 = ~n2306 & n2447 ;
  assign n34345 = n34344 ^ n7801 ^ 1'b0 ;
  assign n34346 = n12608 & n34345 ;
  assign n34347 = ( n8376 & n17680 ) | ( n8376 & ~n21838 ) | ( n17680 & ~n21838 ) ;
  assign n34348 = ( n23281 & ~n34346 ) | ( n23281 & n34347 ) | ( ~n34346 & n34347 ) ;
  assign n34349 = n21633 & ~n34348 ;
  assign n34350 = ~n34343 & n34349 ;
  assign n34351 = ~n3392 & n4016 ;
  assign n34352 = n34351 ^ n12688 ^ 1'b0 ;
  assign n34353 = n28675 | n34352 ;
  assign n34354 = ~n5137 & n34353 ;
  assign n34355 = ~n15632 & n19360 ;
  assign n34356 = n17964 & n34355 ;
  assign n34357 = ~n7822 & n34356 ;
  assign n34358 = n34357 ^ n6703 ^ n2691 ;
  assign n34359 = n3153 & n34358 ;
  assign n34360 = ( n1167 & n7049 ) | ( n1167 & ~n20411 ) | ( n7049 & ~n20411 ) ;
  assign n34361 = n17183 ^ n8218 ^ 1'b0 ;
  assign n34362 = ~n6215 & n34361 ;
  assign n34363 = ( n9578 & ~n12698 ) | ( n9578 & n20643 ) | ( ~n12698 & n20643 ) ;
  assign n34364 = n5675 & n20421 ;
  assign n34365 = n34363 & n34364 ;
  assign n34366 = n7078 | n31688 ;
  assign n34367 = n34366 ^ n13857 ^ 1'b0 ;
  assign n34368 = n3199 & ~n34367 ;
  assign n34369 = n11531 ^ n2918 ^ 1'b0 ;
  assign n34370 = n29563 & n34369 ;
  assign n34371 = n34314 ^ n19497 ^ n2864 ;
  assign n34372 = n5603 | n9155 ;
  assign n34373 = n8912 & ~n31129 ;
  assign n34374 = ( n17223 & n34372 ) | ( n17223 & n34373 ) | ( n34372 & n34373 ) ;
  assign n34375 = ~n14448 & n34374 ;
  assign n34376 = n1904 & n13682 ;
  assign n34377 = ~n10705 & n34376 ;
  assign n34378 = ~n34335 & n34377 ;
  assign n34379 = n10727 ^ n587 ^ 1'b0 ;
  assign n34380 = n34378 & n34379 ;
  assign n34381 = n12817 & n15938 ;
  assign n34382 = n2251 & n11841 ;
  assign n34383 = ~n15220 & n17528 ;
  assign n34384 = n10593 & n34383 ;
  assign n34385 = n25119 ^ n998 ^ 1'b0 ;
  assign n34386 = n18882 ^ n8733 ^ n1617 ;
  assign n34387 = n17465 ^ n7228 ^ 1'b0 ;
  assign n34388 = ( n8929 & n22237 ) | ( n8929 & n34387 ) | ( n22237 & n34387 ) ;
  assign n34389 = ~n18986 & n33427 ;
  assign n34390 = ~n10470 & n34389 ;
  assign n34391 = n34390 ^ n14406 ^ 1'b0 ;
  assign n34392 = n34391 ^ n9086 ^ 1'b0 ;
  assign n34393 = n1459 & ~n11359 ;
  assign n34394 = n34393 ^ n29744 ^ 1'b0 ;
  assign n34395 = n3195 & ~n31143 ;
  assign n34396 = n8105 & n34395 ;
  assign n34397 = n1871 ^ n736 ^ 1'b0 ;
  assign n34398 = n9852 & n34397 ;
  assign n34399 = ~n9533 & n14438 ;
  assign n34400 = n34398 & n34399 ;
  assign n34401 = n17638 & ~n24485 ;
  assign n34402 = n33077 ^ n20717 ^ 1'b0 ;
  assign n34403 = n33899 ^ n578 ^ 1'b0 ;
  assign n34404 = n34403 ^ n30912 ^ n26966 ;
  assign n34408 = n12288 ^ n585 ^ 1'b0 ;
  assign n34405 = ( n411 & n1874 ) | ( n411 & n3192 ) | ( n1874 & n3192 ) ;
  assign n34406 = n13945 & ~n34405 ;
  assign n34407 = n34406 ^ n13470 ^ 1'b0 ;
  assign n34409 = n34408 ^ n34407 ^ n17118 ;
  assign n34414 = ~n3217 & n3779 ;
  assign n34411 = ( n2918 & ~n11466 ) | ( n2918 & n13315 ) | ( ~n11466 & n13315 ) ;
  assign n34410 = n607 & n18741 ;
  assign n34412 = n34411 ^ n34410 ^ 1'b0 ;
  assign n34413 = n6102 & ~n34412 ;
  assign n34415 = n34414 ^ n34413 ^ 1'b0 ;
  assign n34417 = n28828 ^ n21228 ^ n82 ;
  assign n34418 = ( n1802 & n29337 ) | ( n1802 & ~n34417 ) | ( n29337 & ~n34417 ) ;
  assign n34419 = n23695 & n34418 ;
  assign n34416 = n25604 ^ n17183 ^ n10494 ;
  assign n34420 = n34419 ^ n34416 ^ 1'b0 ;
  assign n34421 = n23970 ^ n20660 ^ 1'b0 ;
  assign n34422 = n14415 & ~n23650 ;
  assign n34423 = n6142 ^ n1193 ^ 1'b0 ;
  assign n34424 = n7156 | n34423 ;
  assign n34425 = n13084 & ~n34424 ;
  assign n34426 = n30912 & n34425 ;
  assign n34427 = n4660 & n34426 ;
  assign n34428 = n21784 & n34427 ;
  assign n34429 = ~n7195 & n32244 ;
  assign n34430 = n34429 ^ n13067 ^ 1'b0 ;
  assign n34431 = n1315 & ~n24546 ;
  assign n34432 = ~n31131 & n34431 ;
  assign n34433 = ~n42 & n34432 ;
  assign n34434 = n34016 ^ n5064 ^ 1'b0 ;
  assign n34435 = n5877 & ~n27660 ;
  assign n34436 = n5583 & n34435 ;
  assign n34437 = n3732 ^ n1704 ^ 1'b0 ;
  assign n34438 = n8958 & n19072 ;
  assign n34439 = n6564 & n34438 ;
  assign n34440 = ~n2602 & n4219 ;
  assign n34441 = n34440 ^ n8074 ^ 1'b0 ;
  assign n34442 = n13927 ^ n10352 ^ 1'b0 ;
  assign n34443 = n11962 & n34442 ;
  assign n34444 = n3043 ^ n1677 ^ 1'b0 ;
  assign n34445 = ~n34443 & n34444 ;
  assign n34446 = n34445 ^ n8523 ^ 1'b0 ;
  assign n34447 = n1364 & n8327 ;
  assign n34448 = n8724 & n34447 ;
  assign n34449 = n20038 & ~n24801 ;
  assign n34450 = n34448 & n34449 ;
  assign n34451 = n12588 | n34450 ;
  assign n34452 = n24086 ^ n18410 ^ 1'b0 ;
  assign n34453 = n4782 & n25210 ;
  assign n34454 = n34453 ^ n27638 ^ 1'b0 ;
  assign n34455 = n19165 ^ n14083 ^ 1'b0 ;
  assign n34456 = ~n1332 & n34455 ;
  assign n34457 = ( ~n22670 & n34454 ) | ( ~n22670 & n34456 ) | ( n34454 & n34456 ) ;
  assign n34458 = n15641 | n18353 ;
  assign n34459 = ~n2813 & n33599 ;
  assign n34460 = ~n6712 & n12018 ;
  assign n34461 = n34460 ^ n14665 ^ 1'b0 ;
  assign n34462 = n7805 & n34461 ;
  assign n34463 = n1166 & n34462 ;
  assign n34464 = n34463 ^ n15614 ^ n5149 ;
  assign n34465 = ( n14815 & n21945 ) | ( n14815 & n34464 ) | ( n21945 & n34464 ) ;
  assign n34466 = n10210 & n30119 ;
  assign n34467 = n34466 ^ n17539 ^ 1'b0 ;
  assign n34472 = n4769 | n32684 ;
  assign n34473 = n34472 ^ n22530 ^ 1'b0 ;
  assign n34471 = n10303 ^ n9942 ^ 1'b0 ;
  assign n34468 = n15472 ^ n9208 ^ n4531 ;
  assign n34469 = n34468 ^ n6238 ^ 1'b0 ;
  assign n34470 = n34469 ^ n31259 ^ n24599 ;
  assign n34474 = n34473 ^ n34471 ^ n34470 ;
  assign n34475 = ( ~n1996 & n16160 ) | ( ~n1996 & n34474 ) | ( n16160 & n34474 ) ;
  assign n34476 = ~n16998 & n19869 ;
  assign n34477 = n4112 & n13231 ;
  assign n34478 = n246 & n4490 ;
  assign n34479 = n4016 & ~n11353 ;
  assign n34480 = n1744 & n34479 ;
  assign n34481 = n2980 & ~n23928 ;
  assign n34482 = n34481 ^ n31044 ^ 1'b0 ;
  assign n34483 = ~n24949 & n34482 ;
  assign n34484 = n34483 ^ n21210 ^ 1'b0 ;
  assign n34485 = n11103 & ~n25839 ;
  assign n34486 = n14735 ^ n1853 ^ 1'b0 ;
  assign n34487 = n34486 ^ n1069 ^ 1'b0 ;
  assign n34488 = n4605 | n34487 ;
  assign n34489 = n4928 | n5131 ;
  assign n34490 = n34488 | n34489 ;
  assign n34491 = n34490 ^ n19456 ^ n6704 ;
  assign n34492 = n236 & n12239 ;
  assign n34493 = n7227 ^ n5384 ^ 1'b0 ;
  assign n34494 = n31335 | n34493 ;
  assign n34495 = n34494 ^ n10438 ^ 1'b0 ;
  assign n34496 = n33298 ^ n14508 ^ 1'b0 ;
  assign n34497 = n34496 ^ n19429 ^ 1'b0 ;
  assign n34498 = n19721 ^ n2025 ^ n145 ;
  assign n34499 = ~n4674 & n26340 ;
  assign n34500 = n16865 & n34499 ;
  assign n34501 = ~n27810 & n34500 ;
  assign n34502 = ~n2871 & n11304 ;
  assign n34503 = n4760 & n9781 ;
  assign n34504 = ~n18290 & n34503 ;
  assign n34505 = n34504 ^ n6736 ^ 1'b0 ;
  assign n34513 = n4038 & ~n8911 ;
  assign n34507 = n8279 ^ n349 ^ 1'b0 ;
  assign n34508 = n2414 & ~n34507 ;
  assign n34506 = n5344 ^ n2401 ^ 1'b0 ;
  assign n34509 = n34508 ^ n34506 ^ n16187 ;
  assign n34510 = n390 & ~n34509 ;
  assign n34511 = n34510 ^ n19942 ^ 1'b0 ;
  assign n34512 = n16539 & n34511 ;
  assign n34514 = n34513 ^ n34512 ^ 1'b0 ;
  assign n34516 = n12127 | n24994 ;
  assign n34515 = n8028 & ~n29914 ;
  assign n34517 = n34516 ^ n34515 ^ 1'b0 ;
  assign n34518 = n358 & n9578 ;
  assign n34519 = ~n6466 & n34518 ;
  assign n34520 = n34519 ^ n14454 ^ 1'b0 ;
  assign n34523 = ~n17122 & n17186 ;
  assign n34524 = n27731 & ~n34523 ;
  assign n34525 = ~n20548 & n34524 ;
  assign n34521 = n19239 ^ n9898 ^ 1'b0 ;
  assign n34522 = ~n8722 & n34521 ;
  assign n34526 = n34525 ^ n34522 ^ 1'b0 ;
  assign n34529 = n1089 & ~n26010 ;
  assign n34530 = n34529 ^ n23652 ^ 1'b0 ;
  assign n34527 = n4104 | n11182 ;
  assign n34528 = ~n5129 & n34527 ;
  assign n34531 = n34530 ^ n34528 ^ 1'b0 ;
  assign n34532 = n8414 & n10478 ;
  assign n34533 = n30989 ^ n7536 ^ 1'b0 ;
  assign n34534 = n6535 ^ n3844 ^ 1'b0 ;
  assign n34535 = n4274 | n6034 ;
  assign n34536 = n34535 ^ n16173 ^ n4002 ;
  assign n34537 = ~n6444 & n34536 ;
  assign n34538 = n34537 ^ n18105 ^ 1'b0 ;
  assign n34539 = n1024 & n15274 ;
  assign n34542 = ( ~n20946 & n21654 ) | ( ~n20946 & n25958 ) | ( n21654 & n25958 ) ;
  assign n34540 = n29174 ^ n9683 ^ 1'b0 ;
  assign n34541 = ( n20695 & n21862 ) | ( n20695 & n34540 ) | ( n21862 & n34540 ) ;
  assign n34543 = n34542 ^ n34541 ^ n27078 ;
  assign n34546 = n2953 & n3156 ;
  assign n34547 = ~n10279 & n34546 ;
  assign n34545 = n2665 & ~n17001 ;
  assign n34548 = n34547 ^ n34545 ^ 1'b0 ;
  assign n34544 = n17192 | n25897 ;
  assign n34549 = n34548 ^ n34544 ^ n29879 ;
  assign n34551 = n4028 | n12753 ;
  assign n34552 = n34551 ^ n3174 ^ 1'b0 ;
  assign n34550 = n20691 & ~n32388 ;
  assign n34553 = n34552 ^ n34550 ^ 1'b0 ;
  assign n34554 = n28162 ^ n21720 ^ n7556 ;
  assign n34555 = ~n7468 & n8701 ;
  assign n34556 = ~n14961 & n34555 ;
  assign n34557 = n34554 & ~n34556 ;
  assign n34558 = ( n11495 & ~n20473 ) | ( n11495 & n21794 ) | ( ~n20473 & n21794 ) ;
  assign n34559 = n34558 ^ n3962 ^ 1'b0 ;
  assign n34562 = n9385 ^ n200 ^ 1'b0 ;
  assign n34563 = n9101 & ~n34562 ;
  assign n34560 = ( ~n7705 & n17094 ) | ( ~n7705 & n19809 ) | ( n17094 & n19809 ) ;
  assign n34561 = n16877 & ~n34560 ;
  assign n34564 = n34563 ^ n34561 ^ 1'b0 ;
  assign n34565 = n34564 ^ n13020 ^ n569 ;
  assign n34566 = n23183 ^ n1910 ^ 1'b0 ;
  assign n34567 = n10395 & n34566 ;
  assign n34568 = n2898 & n34567 ;
  assign n34569 = ~n9635 & n24339 ;
  assign n34570 = n34569 ^ n9211 ^ 1'b0 ;
  assign n34571 = n29585 ^ n4904 ^ 1'b0 ;
  assign n34572 = n19385 & ~n34571 ;
  assign n34573 = n34572 ^ n8693 ^ 1'b0 ;
  assign n34574 = n23368 & ~n24340 ;
  assign n34575 = n29080 | n34574 ;
  assign n34576 = n9788 ^ n8674 ^ 1'b0 ;
  assign n34577 = n34576 ^ n14565 ^ n217 ;
  assign n34578 = n13522 ^ n2044 ^ 1'b0 ;
  assign n34579 = ~n34577 & n34578 ;
  assign n34580 = n31772 ^ n13256 ^ n1022 ;
  assign n34582 = n18829 ^ n10407 ^ 1'b0 ;
  assign n34581 = n3581 & ~n27788 ;
  assign n34583 = n34582 ^ n34581 ^ 1'b0 ;
  assign n34584 = n26023 ^ n18169 ^ 1'b0 ;
  assign n34585 = n24165 ^ n1932 ^ n710 ;
  assign n34586 = n9250 ^ n3647 ^ n3176 ;
  assign n34587 = ~n26336 & n34586 ;
  assign n34588 = n6591 | n10548 ;
  assign n34589 = ( n9548 & n11741 ) | ( n9548 & n15279 ) | ( n11741 & n15279 ) ;
  assign n34590 = n34589 ^ n19925 ^ 1'b0 ;
  assign n34591 = n34588 & n34590 ;
  assign n34592 = n7600 & ~n34591 ;
  assign n34593 = n21073 ^ n7040 ^ 1'b0 ;
  assign n34594 = n10258 | n34593 ;
  assign n34595 = n16373 | n26087 ;
  assign n34596 = n34595 ^ n7847 ^ 1'b0 ;
  assign n34597 = n28125 & ~n34596 ;
  assign n34598 = n13907 ^ n1382 ^ 1'b0 ;
  assign n34599 = ~n5978 & n34598 ;
  assign n34600 = n9564 ^ n5292 ^ 1'b0 ;
  assign n34601 = n7255 & ~n34600 ;
  assign n34602 = ( n15832 & n22142 ) | ( n15832 & n34601 ) | ( n22142 & n34601 ) ;
  assign n34603 = ( ~n471 & n7559 ) | ( ~n471 & n14354 ) | ( n7559 & n14354 ) ;
  assign n34604 = n23780 | n34603 ;
  assign n34605 = n6682 & n23825 ;
  assign n34606 = n34605 ^ n4263 ^ 1'b0 ;
  assign n34607 = ~n15267 & n34606 ;
  assign n34608 = ~n26977 & n34607 ;
  assign n34609 = n21001 & ~n28719 ;
  assign n34610 = ~n25716 & n34609 ;
  assign n34611 = n8874 & ~n10090 ;
  assign n34612 = n20191 & n34611 ;
  assign n34613 = n34612 ^ n10417 ^ 1'b0 ;
  assign n34614 = n6404 | n34613 ;
  assign n34615 = n34614 ^ n25058 ^ 1'b0 ;
  assign n34616 = n33081 & ~n34615 ;
  assign n34617 = n20105 ^ n13643 ^ n7658 ;
  assign n34618 = ~n32845 & n34617 ;
  assign n34621 = n6802 ^ n5627 ^ 1'b0 ;
  assign n34619 = n3558 & ~n23363 ;
  assign n34620 = n34619 ^ n11723 ^ 1'b0 ;
  assign n34622 = n34621 ^ n34620 ^ 1'b0 ;
  assign n34623 = n19205 & n34622 ;
  assign n34624 = ( n1234 & n4381 ) | ( n1234 & n7523 ) | ( n4381 & n7523 ) ;
  assign n34625 = n6010 & ~n33711 ;
  assign n34626 = ~n34624 & n34625 ;
  assign n34627 = ( ~n11485 & n13240 ) | ( ~n11485 & n25283 ) | ( n13240 & n25283 ) ;
  assign n34628 = n5541 & ~n34627 ;
  assign n34629 = ~n2393 & n10267 ;
  assign n34630 = ~n1131 & n34629 ;
  assign n34631 = n7146 | n34630 ;
  assign n34632 = n34631 ^ n8277 ^ 1'b0 ;
  assign n34633 = n766 | n9242 ;
  assign n34634 = n34633 ^ n4115 ^ n191 ;
  assign n34635 = n18467 ^ n9603 ^ 1'b0 ;
  assign n34636 = ~n34634 & n34635 ;
  assign n34637 = n6004 & ~n22899 ;
  assign n34638 = n10928 | n21644 ;
  assign n34639 = n34638 ^ n12954 ^ 1'b0 ;
  assign n34640 = n9039 ^ n5748 ^ n1483 ;
  assign n34641 = ( n6570 & n18601 ) | ( n6570 & ~n34640 ) | ( n18601 & ~n34640 ) ;
  assign n34642 = n44 & n24986 ;
  assign n34643 = ~n13121 & n34642 ;
  assign n34644 = n10597 & ~n34643 ;
  assign n34646 = n29633 ^ n20695 ^ 1'b0 ;
  assign n34647 = n8720 | n34646 ;
  assign n34645 = n2273 | n17638 ;
  assign n34648 = n34647 ^ n34645 ^ n24770 ;
  assign n34649 = n5935 | n22398 ;
  assign n34650 = n11919 & n34649 ;
  assign n34651 = n16324 | n27605 ;
  assign n34652 = n20704 ^ n1694 ^ 1'b0 ;
  assign n34653 = n33003 & n34652 ;
  assign n34654 = n23900 ^ n11025 ^ n6623 ;
  assign n34655 = ~n3575 & n13680 ;
  assign n34656 = ~n12127 & n21078 ;
  assign n34657 = ~n34655 & n34656 ;
  assign n34658 = n34657 ^ n20041 ^ 1'b0 ;
  assign n34659 = ~n21365 & n34658 ;
  assign n34660 = n24258 & n30208 ;
  assign n34661 = ~n34659 & n34660 ;
  assign n34662 = ~n2642 & n16134 ;
  assign n34663 = n799 | n13161 ;
  assign n34664 = n22527 ^ n15767 ^ 1'b0 ;
  assign n34665 = n34664 ^ n14760 ^ 1'b0 ;
  assign n34666 = ( n1104 & n34663 ) | ( n1104 & ~n34665 ) | ( n34663 & ~n34665 ) ;
  assign n34667 = n34666 ^ n30450 ^ 1'b0 ;
  assign n34668 = n34662 | n34667 ;
  assign n34669 = n22177 ^ n771 ^ 1'b0 ;
  assign n34670 = ~n3633 & n34669 ;
  assign n34671 = ( n5324 & n26344 ) | ( n5324 & n30475 ) | ( n26344 & n30475 ) ;
  assign n34672 = n11560 ^ n4086 ^ 1'b0 ;
  assign n34673 = n5195 & n34672 ;
  assign n34674 = n4260 & n27405 ;
  assign n34675 = ( n5123 & ~n34673 ) | ( n5123 & n34674 ) | ( ~n34673 & n34674 ) ;
  assign n34676 = n4403 | n9565 ;
  assign n34677 = n34676 ^ n6282 ^ 1'b0 ;
  assign n34678 = n5058 ^ n1983 ^ 1'b0 ;
  assign n34679 = n34677 & ~n34678 ;
  assign n34680 = n3943 & ~n8445 ;
  assign n34681 = n34680 ^ n4186 ^ 1'b0 ;
  assign n34682 = n34679 & ~n34681 ;
  assign n34683 = n7574 | n11952 ;
  assign n34684 = n16735 | n28279 ;
  assign n34685 = n34684 ^ n4250 ^ 1'b0 ;
  assign n34686 = n26179 | n34685 ;
  assign n34687 = ~n18277 & n34686 ;
  assign n34688 = n6446 & ~n34687 ;
  assign n34689 = n34688 ^ n29783 ^ 1'b0 ;
  assign n34690 = n34689 ^ n7124 ^ n5424 ;
  assign n34691 = n34690 ^ n26767 ^ 1'b0 ;
  assign n34692 = n2756 & ~n14578 ;
  assign n34693 = n34692 ^ n7774 ^ 1'b0 ;
  assign n34694 = n22100 | n34693 ;
  assign n34695 = n4084 ^ n3658 ^ 1'b0 ;
  assign n34696 = n34695 ^ n25581 ^ n3184 ;
  assign n34697 = n10928 & ~n24732 ;
  assign n34698 = n34697 ^ n29950 ^ 1'b0 ;
  assign n34699 = ~n34696 & n34698 ;
  assign n34700 = n32671 ^ n17259 ^ 1'b0 ;
  assign n34701 = n34700 ^ n31609 ^ 1'b0 ;
  assign n34702 = n14614 ^ n2781 ^ 1'b0 ;
  assign n34703 = n15443 & ~n34702 ;
  assign n34704 = n5139 & ~n12883 ;
  assign n34705 = n9634 & n34704 ;
  assign n34706 = n19845 | n34705 ;
  assign n34707 = ~n10379 & n34706 ;
  assign n34708 = n34707 ^ n24916 ^ 1'b0 ;
  assign n34709 = n31102 ^ n17257 ^ n3240 ;
  assign n34710 = n21447 | n34709 ;
  assign n34711 = n34708 | n34710 ;
  assign n34713 = n2176 ^ n473 ^ 1'b0 ;
  assign n34712 = n9855 & n15442 ;
  assign n34714 = n34713 ^ n34712 ^ n9601 ;
  assign n34715 = ( ~n7452 & n17667 ) | ( ~n7452 & n34714 ) | ( n17667 & n34714 ) ;
  assign n34716 = ( n5447 & n22127 ) | ( n5447 & n34493 ) | ( n22127 & n34493 ) ;
  assign n34717 = n9504 ^ n2854 ^ 1'b0 ;
  assign n34718 = ~n19947 & n34717 ;
  assign n34719 = n34718 ^ n32272 ^ n645 ;
  assign n34720 = n16080 & ~n27341 ;
  assign n34721 = n13963 & ~n32495 ;
  assign n34722 = ~n34720 & n34721 ;
  assign n34723 = n13887 ^ n9714 ^ 1'b0 ;
  assign n34724 = n13332 & n34723 ;
  assign n34725 = ~n19004 & n34724 ;
  assign n34726 = n34725 ^ n10393 ^ 1'b0 ;
  assign n34730 = n7585 | n32681 ;
  assign n34727 = n17535 ^ n1856 ^ 1'b0 ;
  assign n34728 = n9261 & ~n34727 ;
  assign n34729 = n24875 & n34728 ;
  assign n34731 = n34730 ^ n34729 ^ 1'b0 ;
  assign n34733 = n9401 & n15564 ;
  assign n34732 = ~n4886 & n9736 ;
  assign n34734 = n34733 ^ n34732 ^ 1'b0 ;
  assign n34735 = n4200 | n34734 ;
  assign n34736 = n34735 ^ n19476 ^ 1'b0 ;
  assign n34737 = n23443 ^ n20725 ^ n18818 ;
  assign n34738 = n3471 | n10596 ;
  assign n34739 = n34738 ^ n24089 ^ 1'b0 ;
  assign n34740 = n14609 ^ n6178 ^ 1'b0 ;
  assign n34741 = n9241 & n22127 ;
  assign n34742 = ~n14706 & n34741 ;
  assign n34743 = n28857 ^ n15630 ^ 1'b0 ;
  assign n34744 = ~n5713 & n34743 ;
  assign n34745 = n991 & ~n18638 ;
  assign n34746 = n9926 & n34745 ;
  assign n34747 = n34746 ^ n3581 ^ 1'b0 ;
  assign n34748 = ~n17331 & n24553 ;
  assign n34749 = n34748 ^ n16491 ^ n43 ;
  assign n34750 = n34358 ^ n8769 ^ n6102 ;
  assign n34751 = n20978 ^ n17894 ^ 1'b0 ;
  assign n34752 = n21318 | n34751 ;
  assign n34753 = n25505 ^ n3689 ^ 1'b0 ;
  assign n34754 = ~n17712 & n34753 ;
  assign n34755 = n14247 ^ n378 ^ 1'b0 ;
  assign n34756 = n34755 ^ n25594 ^ n24067 ;
  assign n34757 = ( n914 & ~n4582 ) | ( n914 & n10462 ) | ( ~n4582 & n10462 ) ;
  assign n34758 = n30866 | n34757 ;
  assign n34759 = n34756 | n34758 ;
  assign n34760 = n7019 & n7239 ;
  assign n34761 = n34760 ^ n5740 ^ 1'b0 ;
  assign n34762 = ( n11121 & ~n15199 ) | ( n11121 & n34761 ) | ( ~n15199 & n34761 ) ;
  assign n34763 = n30905 ^ n9068 ^ 1'b0 ;
  assign n34764 = ~n566 & n6328 ;
  assign n34765 = n279 & ~n34764 ;
  assign n34766 = ~n18242 & n21212 ;
  assign n34767 = ~n21193 & n34766 ;
  assign n34768 = n34767 ^ n14083 ^ n1337 ;
  assign n34769 = n15241 & ~n34768 ;
  assign n34770 = ( ~n10062 & n19176 ) | ( ~n10062 & n20743 ) | ( n19176 & n20743 ) ;
  assign n34771 = n25635 & ~n34770 ;
  assign n34772 = ~n7761 & n34771 ;
  assign n34773 = ( n15618 & n18193 ) | ( n15618 & n34772 ) | ( n18193 & n34772 ) ;
  assign n34774 = n9798 & n10811 ;
  assign n34775 = n12003 ^ n5284 ^ n3107 ;
  assign n34776 = n2951 | n34775 ;
  assign n34777 = n34776 ^ n3097 ^ 1'b0 ;
  assign n34778 = n34777 ^ n8821 ^ 1'b0 ;
  assign n34779 = ( ~n4515 & n25877 ) | ( ~n4515 & n31514 ) | ( n25877 & n31514 ) ;
  assign n34780 = n4454 | n34779 ;
  assign n34781 = n2021 & n4994 ;
  assign n34782 = n34781 ^ n11262 ^ 1'b0 ;
  assign n34783 = n34782 ^ n32861 ^ 1'b0 ;
  assign n34784 = n842 & ~n34783 ;
  assign n34785 = ~n1115 & n27319 ;
  assign n34786 = n34785 ^ n9591 ^ 1'b0 ;
  assign n34787 = n2115 | n10181 ;
  assign n34794 = n4143 & n10975 ;
  assign n34795 = n34794 ^ n283 ^ 1'b0 ;
  assign n34793 = n870 & n2053 ;
  assign n34796 = n34795 ^ n34793 ^ n21949 ;
  assign n34790 = ~n876 & n11283 ;
  assign n34788 = ( n1000 & ~n7935 ) | ( n1000 & n8748 ) | ( ~n7935 & n8748 ) ;
  assign n34789 = n4368 | n34788 ;
  assign n34791 = n34790 ^ n34789 ^ 1'b0 ;
  assign n34792 = n16050 | n34791 ;
  assign n34797 = n34796 ^ n34792 ^ 1'b0 ;
  assign n34798 = n12036 ^ n4896 ^ n2334 ;
  assign n34799 = ~n29304 & n34798 ;
  assign n34800 = ( n1410 & ~n3393 ) | ( n1410 & n6509 ) | ( ~n3393 & n6509 ) ;
  assign n34801 = n14507 ^ n11867 ^ 1'b0 ;
  assign n34802 = n17574 & ~n34801 ;
  assign n34804 = n160 & ~n11546 ;
  assign n34805 = n34804 ^ n9982 ^ 1'b0 ;
  assign n34803 = n2436 | n21349 ;
  assign n34806 = n34805 ^ n34803 ^ 1'b0 ;
  assign n34807 = ~n10139 & n34806 ;
  assign n34808 = ~n34802 & n34807 ;
  assign n34809 = n24108 ^ n13725 ^ 1'b0 ;
  assign n34810 = n29244 | n34809 ;
  assign n34811 = n13621 ^ n9739 ^ 1'b0 ;
  assign n34812 = ~n9535 & n34811 ;
  assign n34813 = n5234 & n34812 ;
  assign n34814 = n26941 & ~n34813 ;
  assign n34815 = n34814 ^ n1035 ^ 1'b0 ;
  assign n34816 = n10956 ^ n7780 ^ n5908 ;
  assign n34817 = n19385 & ~n31232 ;
  assign n34818 = n15272 ^ n14988 ^ n4428 ;
  assign n34819 = n1950 & n20593 ;
  assign n34820 = ~n16406 & n31469 ;
  assign n34821 = n34819 & n34820 ;
  assign n34822 = n21741 & n21862 ;
  assign n34823 = n4105 | n9404 ;
  assign n34824 = n1959 | n34823 ;
  assign n34825 = n34824 ^ n3193 ^ 1'b0 ;
  assign n34826 = ~n1040 & n34825 ;
  assign n34827 = n22507 ^ n7634 ^ 1'b0 ;
  assign n34828 = n16261 & ~n34827 ;
  assign n34829 = ~n13062 & n34828 ;
  assign n34830 = n8544 | n9530 ;
  assign n34831 = n34830 ^ n33788 ^ n31904 ;
  assign n34832 = n33139 ^ n20571 ^ 1'b0 ;
  assign n34833 = n5300 & ~n30673 ;
  assign n34834 = ~n4102 & n18935 ;
  assign n34837 = n15441 ^ n12758 ^ 1'b0 ;
  assign n34835 = ~n4338 & n10381 ;
  assign n34836 = n34835 ^ n7556 ^ 1'b0 ;
  assign n34838 = n34837 ^ n34836 ^ n16390 ;
  assign n34839 = n32966 ^ n28282 ^ n554 ;
  assign n34840 = n20218 | n34839 ;
  assign n34841 = n25953 ^ n1118 ^ 1'b0 ;
  assign n34842 = ~n1893 & n14561 ;
  assign n34843 = n34842 ^ n9246 ^ 1'b0 ;
  assign n34844 = n34843 ^ n23910 ^ 1'b0 ;
  assign n34845 = ( n9956 & n20603 ) | ( n9956 & ~n34844 ) | ( n20603 & ~n34844 ) ;
  assign n34846 = ( n2325 & ~n10946 ) | ( n2325 & n31005 ) | ( ~n10946 & n31005 ) ;
  assign n34847 = n32201 & n34846 ;
  assign n34848 = ( n17590 & n27914 ) | ( n17590 & ~n34847 ) | ( n27914 & ~n34847 ) ;
  assign n34850 = n26985 ^ n11567 ^ n10548 ;
  assign n34849 = n27619 & n28320 ;
  assign n34851 = n34850 ^ n34849 ^ 1'b0 ;
  assign n34852 = n31684 ^ n29127 ^ n2051 ;
  assign n34853 = ( n5122 & n11472 ) | ( n5122 & n26708 ) | ( n11472 & n26708 ) ;
  assign n34854 = ~n22157 & n26651 ;
  assign n34855 = n34854 ^ n26071 ^ 1'b0 ;
  assign n34856 = n34853 & n34855 ;
  assign n34857 = n22506 & n34856 ;
  assign n34858 = n34857 ^ n3018 ^ 1'b0 ;
  assign n34861 = ~n8480 & n10716 ;
  assign n34862 = n34679 & n34861 ;
  assign n34863 = n24779 & n34862 ;
  assign n34859 = n14862 ^ n2819 ^ 1'b0 ;
  assign n34860 = ~n11750 & n34859 ;
  assign n34864 = n34863 ^ n34860 ^ 1'b0 ;
  assign n34865 = n12112 & ~n27101 ;
  assign n34866 = n34865 ^ n8608 ^ 1'b0 ;
  assign n34867 = n13846 | n27003 ;
  assign n34868 = n11269 ^ n3096 ^ 1'b0 ;
  assign n34869 = n34867 | n34868 ;
  assign n34870 = n4004 ^ n1350 ^ 1'b0 ;
  assign n34871 = n34870 ^ n33065 ^ 1'b0 ;
  assign n34872 = n12830 ^ n4445 ^ 1'b0 ;
  assign n34873 = n14833 & n34872 ;
  assign n34874 = n34873 ^ n4378 ^ 1'b0 ;
  assign n34875 = n34874 ^ n11111 ^ 1'b0 ;
  assign n34876 = n13151 & ~n14158 ;
  assign n34877 = n3842 & ~n30798 ;
  assign n34878 = n34877 ^ n6743 ^ 1'b0 ;
  assign n34879 = ~n12988 & n14047 ;
  assign n34880 = n7287 ^ n1248 ^ 1'b0 ;
  assign n34881 = n9191 & n34880 ;
  assign n34882 = n34881 ^ n9866 ^ 1'b0 ;
  assign n34883 = n31256 ^ n11571 ^ 1'b0 ;
  assign n34884 = n6431 & n9853 ;
  assign n34885 = ( n6093 & n9921 ) | ( n6093 & ~n34884 ) | ( n9921 & ~n34884 ) ;
  assign n34886 = n34885 ^ n4001 ^ 1'b0 ;
  assign n34887 = ( n2213 & n7565 ) | ( n2213 & n17567 ) | ( n7565 & n17567 ) ;
  assign n34888 = n34887 ^ n30506 ^ 1'b0 ;
  assign n34889 = n8058 & n26443 ;
  assign n34890 = n26428 & n34889 ;
  assign n34891 = n34486 ^ n1143 ^ 1'b0 ;
  assign n34892 = n16025 & n34891 ;
  assign n34893 = n34892 ^ n5399 ^ 1'b0 ;
  assign n34895 = ~n1228 & n6528 ;
  assign n34896 = n68 & n34895 ;
  assign n34897 = n12507 & n34896 ;
  assign n34894 = n4000 & ~n23388 ;
  assign n34898 = n34897 ^ n34894 ^ 1'b0 ;
  assign n34899 = n8684 ^ n4044 ^ n2493 ;
  assign n34900 = n11464 & ~n30377 ;
  assign n34901 = n21017 ^ n6383 ^ 1'b0 ;
  assign n34902 = n12192 & ~n13768 ;
  assign n34903 = n11142 & n34902 ;
  assign n34904 = n34901 | n34903 ;
  assign n34905 = n21932 & n25880 ;
  assign n34906 = n24040 ^ n22562 ^ 1'b0 ;
  assign n34907 = ~n34905 & n34906 ;
  assign n34908 = n5979 & ~n14194 ;
  assign n34909 = n34908 ^ n5302 ^ 1'b0 ;
  assign n34910 = ~n30839 & n31549 ;
  assign n34911 = n12041 ^ n2067 ^ 1'b0 ;
  assign n34912 = ~n6369 & n34911 ;
  assign n34913 = n34912 ^ n21358 ^ 1'b0 ;
  assign n34914 = n34910 & n34913 ;
  assign n34915 = n31336 ^ n3266 ^ 1'b0 ;
  assign n34916 = n34915 ^ n13865 ^ 1'b0 ;
  assign n34917 = n31026 & ~n34916 ;
  assign n34918 = n34917 ^ n25461 ^ n4092 ;
  assign n34919 = ~n12482 & n32671 ;
  assign n34920 = n12536 & n34919 ;
  assign n34921 = n16374 | n34920 ;
  assign n34922 = n16468 & ~n16771 ;
  assign n34923 = n19014 ^ n13528 ^ 1'b0 ;
  assign n34924 = n34922 & n34923 ;
  assign n34925 = n18096 ^ n6155 ^ 1'b0 ;
  assign n34926 = n21952 & ~n34925 ;
  assign n34927 = n18501 ^ n16056 ^ n1812 ;
  assign n34928 = n34926 & n34927 ;
  assign n34929 = ~n13059 & n19292 ;
  assign n34930 = ~n11365 & n11846 ;
  assign n34931 = n34930 ^ n11577 ^ 1'b0 ;
  assign n34932 = ( n34137 & n34929 ) | ( n34137 & ~n34931 ) | ( n34929 & ~n34931 ) ;
  assign n34933 = n21808 ^ n21709 ^ n332 ;
  assign n34934 = n11693 & ~n27020 ;
  assign n34935 = n15870 & n34934 ;
  assign n34936 = n23240 & ~n34935 ;
  assign n34937 = n34936 ^ n6097 ^ 1'b0 ;
  assign n34938 = ~n10076 & n34937 ;
  assign n34939 = n34938 ^ n31045 ^ n16684 ;
  assign n34943 = ~n3266 & n7426 ;
  assign n34940 = n14449 ^ n3031 ^ 1'b0 ;
  assign n34941 = n3478 | n34940 ;
  assign n34942 = n29783 & n34941 ;
  assign n34944 = n34943 ^ n34942 ^ n10839 ;
  assign n34945 = ~n28277 & n28529 ;
  assign n34946 = n608 & n22034 ;
  assign n34947 = n6144 & n14730 ;
  assign n34948 = n5168 & n34947 ;
  assign n34949 = n34948 ^ n27345 ^ 1'b0 ;
  assign n34950 = n22334 & ~n34949 ;
  assign n34951 = n15923 | n18911 ;
  assign n34952 = n34951 ^ n6374 ^ 1'b0 ;
  assign n34955 = n13834 | n22593 ;
  assign n34956 = n6934 & ~n34955 ;
  assign n34953 = ~n13068 & n15059 ;
  assign n34954 = n34953 ^ n31187 ^ 1'b0 ;
  assign n34957 = n34956 ^ n34954 ^ n25702 ;
  assign n34958 = n33755 ^ n24485 ^ 1'b0 ;
  assign n34959 = ~n7052 & n34958 ;
  assign n34960 = n22216 & n34959 ;
  assign n34961 = n6339 & n34960 ;
  assign n34962 = ~n22992 & n24481 ;
  assign n34963 = n6301 & n34962 ;
  assign n34964 = n25793 & ~n34963 ;
  assign n34966 = n1614 | n22410 ;
  assign n34965 = n6044 ^ n5373 ^ 1'b0 ;
  assign n34967 = n34966 ^ n34965 ^ 1'b0 ;
  assign n34968 = n283 & n6609 ;
  assign n34969 = n34968 ^ n4862 ^ 1'b0 ;
  assign n34970 = ~n14721 & n34969 ;
  assign n34971 = n654 & n34970 ;
  assign n34972 = n33 & ~n8277 ;
  assign n34973 = n1170 & n34972 ;
  assign n34974 = n34973 ^ n20599 ^ n13507 ;
  assign n34975 = n20983 & ~n34974 ;
  assign n34976 = n34975 ^ n24631 ^ 1'b0 ;
  assign n34977 = n10260 & n30441 ;
  assign n34978 = n6615 & ~n22556 ;
  assign n34979 = ~n34977 & n34978 ;
  assign n34980 = n2418 | n30557 ;
  assign n34982 = n20892 ^ n18729 ^ 1'b0 ;
  assign n34981 = n27853 ^ n341 ^ 1'b0 ;
  assign n34983 = n34982 ^ n34981 ^ 1'b0 ;
  assign n34984 = n8709 & n15609 ;
  assign n34985 = n29814 ^ n5869 ^ n3060 ;
  assign n34986 = n1886 & n34985 ;
  assign n34987 = n30419 & ~n34588 ;
  assign n34988 = n34987 ^ n25479 ^ n11978 ;
  assign n34989 = n3876 ^ n776 ^ 1'b0 ;
  assign n34990 = n18242 & ~n25929 ;
  assign n34991 = ( n11667 & n34989 ) | ( n11667 & n34990 ) | ( n34989 & n34990 ) ;
  assign n34992 = n25123 | n34991 ;
  assign n34993 = n1742 | n26015 ;
  assign n34996 = n18932 ^ n14760 ^ n1353 ;
  assign n34997 = n29185 & ~n34996 ;
  assign n34994 = n4005 & n29256 ;
  assign n34995 = ~n14100 & n34994 ;
  assign n34998 = n34997 ^ n34995 ^ 1'b0 ;
  assign n34999 = n34993 & ~n34998 ;
  assign n35001 = n27454 & ~n31753 ;
  assign n35000 = ~n776 & n3720 ;
  assign n35002 = n35001 ^ n35000 ^ 1'b0 ;
  assign n35003 = ~n11935 & n33597 ;
  assign n35004 = n8156 ^ n864 ^ 1'b0 ;
  assign n35006 = n5850 ^ n1568 ^ 1'b0 ;
  assign n35005 = n11247 | n34540 ;
  assign n35007 = n35006 ^ n35005 ^ 1'b0 ;
  assign n35008 = n6045 ^ n5466 ^ 1'b0 ;
  assign n35009 = n35007 | n35008 ;
  assign n35010 = n35009 ^ n1591 ^ 1'b0 ;
  assign n35011 = n35004 & n35010 ;
  assign n35012 = n35011 ^ n34895 ^ 1'b0 ;
  assign n35013 = n26711 ^ n17098 ^ n10878 ;
  assign n35014 = ~n2967 & n35013 ;
  assign n35015 = n22180 ^ n10679 ^ n6470 ;
  assign n35016 = n35015 ^ n32196 ^ 1'b0 ;
  assign n35017 = ~n18319 & n35016 ;
  assign n35018 = n19429 ^ n15130 ^ 1'b0 ;
  assign n35019 = n16493 ^ n708 ^ 1'b0 ;
  assign n35020 = ( ~n15119 & n35018 ) | ( ~n15119 & n35019 ) | ( n35018 & n35019 ) ;
  assign n35021 = ~n8140 & n26853 ;
  assign n35022 = n5727 | n15059 ;
  assign n35023 = n35021 & ~n35022 ;
  assign n35024 = n35023 ^ n16735 ^ n14315 ;
  assign n35025 = ( ~n11320 & n13550 ) | ( ~n11320 & n28733 ) | ( n13550 & n28733 ) ;
  assign n35026 = n18534 ^ n8310 ^ 1'b0 ;
  assign n35027 = n11652 & ~n35026 ;
  assign n35028 = n1021 | n8421 ;
  assign n35029 = n35028 ^ n1749 ^ 1'b0 ;
  assign n35030 = n29072 | n35029 ;
  assign n35031 = n10639 & ~n35030 ;
  assign n35032 = n12291 ^ n6868 ^ n255 ;
  assign n35033 = n28003 ^ n3904 ^ 1'b0 ;
  assign n35034 = n1668 | n16643 ;
  assign n35035 = n35034 ^ n505 ^ 1'b0 ;
  assign n35036 = ( n1250 & ~n20046 ) | ( n1250 & n35035 ) | ( ~n20046 & n35035 ) ;
  assign n35037 = ( n1712 & n20903 ) | ( n1712 & n35036 ) | ( n20903 & n35036 ) ;
  assign n35038 = n16238 | n27003 ;
  assign n35040 = n6951 | n9469 ;
  assign n35041 = n13018 | n35040 ;
  assign n35042 = ( n8207 & n29842 ) | ( n8207 & n35041 ) | ( n29842 & n35041 ) ;
  assign n35039 = n6451 | n15884 ;
  assign n35043 = n35042 ^ n35039 ^ 1'b0 ;
  assign n35044 = n4383 & ~n29579 ;
  assign n35046 = ( ~n9140 & n19149 ) | ( ~n9140 & n27912 ) | ( n19149 & n27912 ) ;
  assign n35045 = n3563 & ~n25904 ;
  assign n35047 = n35046 ^ n35045 ^ 1'b0 ;
  assign n35048 = ( n3756 & ~n8351 ) | ( n3756 & n14883 ) | ( ~n8351 & n14883 ) ;
  assign n35049 = ( n12668 & n14379 ) | ( n12668 & n35048 ) | ( n14379 & n35048 ) ;
  assign n35050 = n35049 ^ n8021 ^ n890 ;
  assign n35051 = n10341 & ~n24030 ;
  assign n35052 = n14979 & ~n19342 ;
  assign n35053 = n35052 ^ n12400 ^ 1'b0 ;
  assign n35054 = ~n517 & n20541 ;
  assign n35055 = n16572 & n35054 ;
  assign n35056 = n3593 & ~n33557 ;
  assign n35057 = n1322 | n4417 ;
  assign n35058 = n28620 | n35057 ;
  assign n35059 = n12666 ^ n7875 ^ 1'b0 ;
  assign n35060 = n13882 | n35059 ;
  assign n35061 = n35060 ^ n26829 ^ 1'b0 ;
  assign n35062 = n3803 & ~n16169 ;
  assign n35063 = ~n11117 & n35062 ;
  assign n35064 = n23757 ^ n7335 ^ 1'b0 ;
  assign n35065 = ~n35063 & n35064 ;
  assign n35066 = n34929 ^ n6102 ^ 1'b0 ;
  assign n35067 = n31739 | n35066 ;
  assign n35068 = n11482 & ~n35067 ;
  assign n35069 = n11683 | n17080 ;
  assign n35070 = n35069 ^ n17104 ^ n542 ;
  assign n35071 = n9546 ^ n2123 ^ 1'b0 ;
  assign n35072 = n11349 | n13939 ;
  assign n35073 = n31623 & ~n35072 ;
  assign n35074 = n11626 & n35073 ;
  assign n35075 = n2686 & ~n35074 ;
  assign n35076 = n35075 ^ n34936 ^ 1'b0 ;
  assign n35077 = n6139 & n32707 ;
  assign n35078 = ~n8711 & n34755 ;
  assign n35079 = n17332 & n32127 ;
  assign n35080 = n16889 & n26227 ;
  assign n35081 = ~n35079 & n35080 ;
  assign n35082 = n26922 ^ n13075 ^ 1'b0 ;
  assign n35083 = n7925 & ~n35082 ;
  assign n35084 = n4862 & n5706 ;
  assign n35085 = n35084 ^ n26620 ^ 1'b0 ;
  assign n35086 = n29078 | n35085 ;
  assign n35087 = n1459 & ~n22996 ;
  assign n35088 = ~n3455 & n35087 ;
  assign n35089 = n35088 ^ n24324 ^ 1'b0 ;
  assign n35090 = n2274 | n35089 ;
  assign n35091 = n12549 ^ n6865 ^ 1'b0 ;
  assign n35092 = ( n29531 & n34569 ) | ( n29531 & n35091 ) | ( n34569 & n35091 ) ;
  assign n35093 = n13555 ^ n7252 ^ 1'b0 ;
  assign n35094 = n4690 | n16225 ;
  assign n35095 = n35093 | n35094 ;
  assign n35096 = ~n6584 & n11104 ;
  assign n35097 = n35096 ^ n9034 ^ 1'b0 ;
  assign n35098 = ~n29847 & n35097 ;
  assign n35099 = ~n24044 & n35098 ;
  assign n35100 = n18193 ^ n17226 ^ 1'b0 ;
  assign n35101 = n30060 ^ n19525 ^ 1'b0 ;
  assign n35102 = n35101 ^ n23189 ^ n10411 ;
  assign n35103 = n35102 ^ n13026 ^ 1'b0 ;
  assign n35104 = ~n5477 & n22545 ;
  assign n35106 = ( n1909 & n5519 ) | ( n1909 & n14183 ) | ( n5519 & n14183 ) ;
  assign n35105 = ( n9612 & n12522 ) | ( n9612 & ~n13327 ) | ( n12522 & ~n13327 ) ;
  assign n35107 = n35106 ^ n35105 ^ n3477 ;
  assign n35108 = ~n26550 & n35107 ;
  assign n35112 = n24828 & n32688 ;
  assign n35109 = n7449 | n8108 ;
  assign n35110 = n16247 ^ n2102 ^ 1'b0 ;
  assign n35111 = n35109 & ~n35110 ;
  assign n35113 = n35112 ^ n35111 ^ n4048 ;
  assign n35114 = n1247 | n35113 ;
  assign n35115 = ( ~n15867 & n33957 ) | ( ~n15867 & n35114 ) | ( n33957 & n35114 ) ;
  assign n35116 = n6239 & n25958 ;
  assign n35117 = n3244 & ~n35116 ;
  assign n35118 = n35117 ^ n15392 ^ 1'b0 ;
  assign n35119 = n8362 | n35118 ;
  assign n35120 = ~n6689 & n17652 ;
  assign n35121 = ~n25103 & n35120 ;
  assign n35122 = n484 | n35121 ;
  assign n35123 = n4189 & ~n35122 ;
  assign n35124 = n23005 ^ n8556 ^ 1'b0 ;
  assign n35125 = ( n22651 & ~n31164 ) | ( n22651 & n35124 ) | ( ~n31164 & n35124 ) ;
  assign n35126 = n13448 | n35125 ;
  assign n35127 = ~n11406 & n35126 ;
  assign n35128 = n15645 | n26767 ;
  assign n35130 = n526 & n3898 ;
  assign n35129 = n12754 | n29517 ;
  assign n35131 = n35130 ^ n35129 ^ n15531 ;
  assign n35132 = ~n15679 & n34843 ;
  assign n35133 = ( n8447 & n35131 ) | ( n8447 & n35132 ) | ( n35131 & n35132 ) ;
  assign n35134 = n35133 ^ n22223 ^ 1'b0 ;
  assign n35135 = n35128 & ~n35134 ;
  assign n35138 = ~n2599 & n30443 ;
  assign n35139 = ~n10532 & n35138 ;
  assign n35136 = n17579 & n26233 ;
  assign n35137 = n8268 & n35136 ;
  assign n35140 = n35139 ^ n35137 ^ n310 ;
  assign n35141 = n21454 ^ n15217 ^ n12614 ;
  assign n35142 = n10903 ^ n4701 ^ 1'b0 ;
  assign n35143 = n15367 & n35142 ;
  assign n35144 = n8957 & n16622 ;
  assign n35145 = n35144 ^ n20665 ^ 1'b0 ;
  assign n35146 = n30139 & n35145 ;
  assign n35147 = ~n35143 & n35146 ;
  assign n35148 = n6578 & ~n35147 ;
  assign n35149 = n1957 | n24573 ;
  assign n35150 = n11544 & ~n35149 ;
  assign n35151 = ~n1930 & n6229 ;
  assign n35152 = n35151 ^ n3359 ^ 1'b0 ;
  assign n35153 = n2292 | n13943 ;
  assign n35154 = n35153 ^ n29885 ^ 1'b0 ;
  assign n35155 = n29164 & n32519 ;
  assign n35156 = n27426 ^ n24222 ^ n1393 ;
  assign n35157 = n1742 & n3731 ;
  assign n35158 = n15854 & n19800 ;
  assign n35159 = n11172 ^ n2277 ^ 1'b0 ;
  assign n35160 = n9459 & n35159 ;
  assign n35161 = n1062 & n6340 ;
  assign n35162 = n35161 ^ n18077 ^ 1'b0 ;
  assign n35163 = n1745 & n27516 ;
  assign n35164 = ~n35162 & n35163 ;
  assign n35165 = ~n21461 & n35164 ;
  assign n35166 = n34981 ^ n32227 ^ 1'b0 ;
  assign n35167 = n8373 ^ n1200 ^ 1'b0 ;
  assign n35169 = n11533 ^ n728 ^ 1'b0 ;
  assign n35168 = n2728 & n5750 ;
  assign n35170 = n35169 ^ n35168 ^ 1'b0 ;
  assign n35171 = n8094 ^ n3708 ^ 1'b0 ;
  assign n35172 = ~n6036 & n20092 ;
  assign n35173 = n2264 & n35172 ;
  assign n35174 = n9357 ^ n5768 ^ 1'b0 ;
  assign n35175 = n19473 & ~n35174 ;
  assign n35176 = n5070 & ~n5284 ;
  assign n35177 = n35176 ^ n16877 ^ 1'b0 ;
  assign n35178 = n35175 & ~n35177 ;
  assign n35179 = n35173 & n35178 ;
  assign n35180 = n2028 | n3229 ;
  assign n35181 = n38 & ~n35180 ;
  assign n35182 = n11063 ^ n10626 ^ n1741 ;
  assign n35185 = ( n2541 & n10108 ) | ( n2541 & ~n10839 ) | ( n10108 & ~n10839 ) ;
  assign n35183 = n30344 & ~n30972 ;
  assign n35184 = n35183 ^ n9116 ^ 1'b0 ;
  assign n35186 = n35185 ^ n35184 ^ n21701 ;
  assign n35196 = ~n3430 & n5750 ;
  assign n35197 = n35196 ^ n11667 ^ 1'b0 ;
  assign n35198 = ~n6462 & n6664 ;
  assign n35199 = ( n2723 & ~n35197 ) | ( n2723 & n35198 ) | ( ~n35197 & n35198 ) ;
  assign n35200 = ( ~n11676 & n25041 ) | ( ~n11676 & n35199 ) | ( n25041 & n35199 ) ;
  assign n35188 = n6678 & ~n7577 ;
  assign n35187 = n10210 & ~n20496 ;
  assign n35189 = n35188 ^ n35187 ^ 1'b0 ;
  assign n35190 = n18695 & ~n35189 ;
  assign n35191 = ~n2322 & n35190 ;
  assign n35192 = n21552 ^ n6296 ^ 1'b0 ;
  assign n35193 = n35192 ^ n18735 ^ 1'b0 ;
  assign n35194 = n23311 & n35193 ;
  assign n35195 = n35191 & n35194 ;
  assign n35201 = n35200 ^ n35195 ^ n14255 ;
  assign n35202 = n1969 & n24755 ;
  assign n35203 = n923 ^ n867 ^ 1'b0 ;
  assign n35204 = ~n4610 & n35203 ;
  assign n35205 = ~n30472 & n35204 ;
  assign n35206 = ~n35202 & n35205 ;
  assign n35207 = n34467 ^ n18406 ^ 1'b0 ;
  assign n35208 = ~n9045 & n35207 ;
  assign n35209 = n16175 ^ n1639 ^ 1'b0 ;
  assign n35210 = ( n1881 & n19529 ) | ( n1881 & ~n19681 ) | ( n19529 & ~n19681 ) ;
  assign n35211 = n35210 ^ n16495 ^ 1'b0 ;
  assign n35212 = n26979 | n35211 ;
  assign n35213 = n19742 ^ n6221 ^ 1'b0 ;
  assign n35214 = ~n749 & n4574 ;
  assign n35215 = n35214 ^ n10265 ^ 1'b0 ;
  assign n35216 = n10347 & n35215 ;
  assign n35217 = n35213 & n35216 ;
  assign n35218 = n21586 | n24326 ;
  assign n35219 = n35218 ^ n4459 ^ 1'b0 ;
  assign n35220 = n694 & ~n3756 ;
  assign n35221 = ~n25103 & n35220 ;
  assign n35222 = n35221 ^ n4773 ^ 1'b0 ;
  assign n35223 = n14249 | n18392 ;
  assign n35224 = n35223 ^ n10106 ^ 1'b0 ;
  assign n35225 = n1882 ^ n1095 ^ 1'b0 ;
  assign n35226 = n3689 | n7713 ;
  assign n35227 = n32643 ^ n17501 ^ 1'b0 ;
  assign n35228 = n356 & ~n13650 ;
  assign n35229 = n35228 ^ n10579 ^ 1'b0 ;
  assign n35230 = ~n809 & n12086 ;
  assign n35231 = ~n35229 & n35230 ;
  assign n35232 = n29289 ^ n15589 ^ 1'b0 ;
  assign n35233 = n35231 | n35232 ;
  assign n35234 = n1881 & ~n34583 ;
  assign n35235 = n21186 & n35234 ;
  assign n35238 = ~n13010 & n26744 ;
  assign n35239 = n35238 ^ n428 ^ 1'b0 ;
  assign n35236 = n17556 ^ n14152 ^ 1'b0 ;
  assign n35237 = n26773 & n35236 ;
  assign n35240 = n35239 ^ n35237 ^ 1'b0 ;
  assign n35241 = n10464 & ~n15884 ;
  assign n35242 = n8294 ^ n2954 ^ 1'b0 ;
  assign n35243 = n25809 & n35242 ;
  assign n35244 = n2062 & ~n35243 ;
  assign n35245 = n226 | n5559 ;
  assign n35246 = ~n19218 & n26465 ;
  assign n35247 = n35246 ^ n19304 ^ 1'b0 ;
  assign n35248 = n35245 & ~n35247 ;
  assign n35249 = n9204 ^ n457 ^ 1'b0 ;
  assign n35250 = ~n9011 & n35249 ;
  assign n35251 = n16731 & n27536 ;
  assign n35252 = n35251 ^ n250 ^ 1'b0 ;
  assign n35253 = n11977 | n35252 ;
  assign n35256 = n11671 ^ n1553 ^ 1'b0 ;
  assign n35257 = ~n1285 & n35256 ;
  assign n35258 = n35257 ^ n23123 ^ n11366 ;
  assign n35254 = n14110 & ~n22851 ;
  assign n35255 = n28683 & ~n35254 ;
  assign n35259 = n35258 ^ n35255 ^ 1'b0 ;
  assign n35260 = n881 & ~n7916 ;
  assign n35261 = n35260 ^ n1464 ^ 1'b0 ;
  assign n35262 = n4870 | n18593 ;
  assign n35263 = n35261 | n35262 ;
  assign n35265 = n8693 & n23985 ;
  assign n35266 = n162 & n35265 ;
  assign n35264 = n7166 | n18145 ;
  assign n35267 = n35266 ^ n35264 ^ n16932 ;
  assign n35268 = n35267 ^ n7443 ^ n578 ;
  assign n35269 = ( n4981 & ~n9919 ) | ( n4981 & n18985 ) | ( ~n9919 & n18985 ) ;
  assign n35270 = ~n20355 & n35084 ;
  assign n35271 = ~n35269 & n35270 ;
  assign n35272 = n1638 & n12666 ;
  assign n35273 = n25078 ^ n16628 ^ 1'b0 ;
  assign n35274 = n34797 ^ n8330 ^ 1'b0 ;
  assign n35275 = n11516 & ~n27123 ;
  assign n35276 = n35275 ^ n19973 ^ 1'b0 ;
  assign n35277 = ~n2986 & n11254 ;
  assign n35279 = n532 & n15725 ;
  assign n35280 = n35279 ^ n9143 ^ 1'b0 ;
  assign n35278 = ~n10304 & n11285 ;
  assign n35281 = n35280 ^ n35278 ^ 1'b0 ;
  assign n35282 = n20598 ^ n15406 ^ 1'b0 ;
  assign n35283 = n10054 & ~n35282 ;
  assign n35284 = ~n4846 & n18469 ;
  assign n35285 = n35284 ^ n5554 ^ 1'b0 ;
  assign n35286 = n4342 ^ n2743 ^ 1'b0 ;
  assign n35287 = n35285 & n35286 ;
  assign n35288 = n23245 ^ n9586 ^ 1'b0 ;
  assign n35289 = n16977 & ~n35288 ;
  assign n35290 = n8521 ^ n3432 ^ 1'b0 ;
  assign n35291 = n3038 & ~n11331 ;
  assign n35292 = ~n30818 & n35291 ;
  assign n35293 = n14915 ^ n10976 ^ 1'b0 ;
  assign n35294 = n35293 ^ n2696 ^ 1'b0 ;
  assign n35295 = ( ~n13344 & n34953 ) | ( ~n13344 & n35294 ) | ( n34953 & n35294 ) ;
  assign n35296 = ( ~n19929 & n35292 ) | ( ~n19929 & n35295 ) | ( n35292 & n35295 ) ;
  assign n35297 = ~n3310 & n27622 ;
  assign n35298 = n30575 ^ n26029 ^ 1'b0 ;
  assign n35299 = n35297 | n35298 ;
  assign n35300 = n1293 & ~n10815 ;
  assign n35301 = n24794 & n35300 ;
  assign n35302 = n1616 & ~n35301 ;
  assign n35303 = n35302 ^ n31044 ^ 1'b0 ;
  assign n35304 = n9386 & ~n13231 ;
  assign n35305 = n9869 ^ n4490 ^ 1'b0 ;
  assign n35306 = n30538 | n35305 ;
  assign n35307 = n35306 ^ n24388 ^ 1'b0 ;
  assign n35308 = ( x0 & n9625 ) | ( x0 & n22369 ) | ( n9625 & n22369 ) ;
  assign n35309 = n27064 & n35308 ;
  assign n35310 = n35307 & ~n35309 ;
  assign n35311 = n6754 | n15277 ;
  assign n35312 = ~n184 & n9122 ;
  assign n35313 = n3742 & n6707 ;
  assign n35314 = ~n35312 & n35313 ;
  assign n35315 = ~n1459 & n35314 ;
  assign n35316 = n12597 | n35315 ;
  assign n35317 = n32676 & ~n35316 ;
  assign n35318 = ~n1175 & n34932 ;
  assign n35319 = n35318 ^ n2502 ^ 1'b0 ;
  assign n35321 = n220 & ~n7009 ;
  assign n35322 = ~n2958 & n35321 ;
  assign n35320 = ~n8672 & n12583 ;
  assign n35323 = n35322 ^ n35320 ^ 1'b0 ;
  assign n35324 = ~n55 & n10647 ;
  assign n35325 = ~n35323 & n35324 ;
  assign n35326 = n35325 ^ n31146 ^ n9716 ;
  assign n35327 = n35326 ^ n35081 ^ 1'b0 ;
  assign n35330 = n26956 | n29565 ;
  assign n35328 = n3464 ^ n3337 ^ n2370 ;
  assign n35329 = n3568 & ~n35328 ;
  assign n35331 = n35330 ^ n35329 ^ n15260 ;
  assign n35332 = ~n3268 & n16132 ;
  assign n35333 = n28534 ^ n6362 ^ n5195 ;
  assign n35334 = n25155 ^ n9150 ^ 1'b0 ;
  assign n35335 = ~n22123 & n35334 ;
  assign n35336 = n13923 | n35335 ;
  assign n35337 = n35336 ^ n7087 ^ 1'b0 ;
  assign n35338 = n24661 ^ n3301 ^ 1'b0 ;
  assign n35339 = n11837 & ~n15595 ;
  assign n35340 = n17194 & n35339 ;
  assign n35341 = n35340 ^ n17475 ^ 1'b0 ;
  assign n35342 = n23239 & ~n35341 ;
  assign n35343 = n12251 ^ n6251 ^ 1'b0 ;
  assign n35344 = n2350 | n35343 ;
  assign n35345 = n14093 | n35344 ;
  assign n35346 = n10042 ^ n7300 ^ n6762 ;
  assign n35347 = ~n33725 & n35346 ;
  assign n35349 = n7404 & n27959 ;
  assign n35348 = n32468 ^ n23355 ^ 1'b0 ;
  assign n35350 = n35349 ^ n35348 ^ n203 ;
  assign n35351 = n5761 ^ n2122 ^ 1'b0 ;
  assign n35352 = ( n2887 & ~n11111 ) | ( n2887 & n20375 ) | ( ~n11111 & n20375 ) ;
  assign n35353 = ( n4845 & n14835 ) | ( n4845 & n22900 ) | ( n14835 & n22900 ) ;
  assign n35354 = n9151 ^ n5781 ^ 1'b0 ;
  assign n35355 = n10288 ^ n397 ^ 1'b0 ;
  assign n35356 = n22785 ^ n18530 ^ 1'b0 ;
  assign n35357 = ( n9141 & n25366 ) | ( n9141 & n35356 ) | ( n25366 & n35356 ) ;
  assign n35358 = n18210 & ~n28835 ;
  assign n35359 = n22025 ^ n2495 ^ 1'b0 ;
  assign n35360 = n35358 & n35359 ;
  assign n35361 = ~n1523 & n35360 ;
  assign n35362 = n4326 | n30339 ;
  assign n35363 = n28136 & ~n35294 ;
  assign n35364 = ( n1552 & n12106 ) | ( n1552 & n12500 ) | ( n12106 & n12500 ) ;
  assign n35365 = n32398 ^ n20189 ^ 1'b0 ;
  assign n35366 = ( n26783 & n35364 ) | ( n26783 & n35365 ) | ( n35364 & n35365 ) ;
  assign n35367 = n21611 & n24340 ;
  assign n35368 = n19898 & n35367 ;
  assign n35369 = ( n11680 & n15263 ) | ( n11680 & n26409 ) | ( n15263 & n26409 ) ;
  assign n35370 = n29200 ^ n11241 ^ 1'b0 ;
  assign n35371 = n2854 | n35370 ;
  assign n35372 = n35371 ^ n24308 ^ 1'b0 ;
  assign n35373 = n23387 ^ n3441 ^ 1'b0 ;
  assign n35374 = n29654 ^ n4631 ^ 1'b0 ;
  assign n35375 = n9347 & ~n35374 ;
  assign n35376 = n35375 ^ n1931 ^ 1'b0 ;
  assign n35377 = n29966 ^ n3410 ^ 1'b0 ;
  assign n35378 = n35376 & ~n35377 ;
  assign n35379 = n35378 ^ n31578 ^ 1'b0 ;
  assign n35380 = n25682 & ~n35379 ;
  assign n35381 = n35380 ^ n4326 ^ 1'b0 ;
  assign n35382 = n30753 ^ n11456 ^ 1'b0 ;
  assign n35383 = n3770 ^ n1068 ^ 1'b0 ;
  assign n35384 = ~n3575 & n35383 ;
  assign n35385 = ~n17226 & n35384 ;
  assign n35386 = n35385 ^ n19041 ^ 1'b0 ;
  assign n35387 = n27876 ^ n5836 ^ 1'b0 ;
  assign n35388 = ~n14960 & n35387 ;
  assign n35389 = n13165 ^ n9218 ^ n947 ;
  assign n35390 = n12849 ^ n5988 ^ n5554 ;
  assign n35391 = n35390 ^ n31384 ^ n13316 ;
  assign n35392 = n25216 ^ n20124 ^ n15980 ;
  assign n35393 = n35392 ^ n11910 ^ n7639 ;
  assign n35394 = n12175 ^ n10588 ^ n7223 ;
  assign n35395 = n6595 & ~n7900 ;
  assign n35396 = ~n35394 & n35395 ;
  assign n35397 = ~n8907 & n35396 ;
  assign n35398 = n4342 & ~n35397 ;
  assign n35399 = n17030 | n18334 ;
  assign n35400 = n18334 & ~n35399 ;
  assign n35401 = ~n25672 & n31485 ;
  assign n35402 = n35401 ^ n21172 ^ 1'b0 ;
  assign n35405 = n5845 & ~n13094 ;
  assign n35403 = n1852 & ~n5309 ;
  assign n35404 = ~n2060 & n35403 ;
  assign n35406 = n35405 ^ n35404 ^ 1'b0 ;
  assign n35407 = n24457 & ~n35406 ;
  assign n35408 = n35407 ^ n21703 ^ 1'b0 ;
  assign n35409 = n18534 ^ n3634 ^ 1'b0 ;
  assign n35410 = n3560 & ~n35409 ;
  assign n35411 = ( n2918 & n33372 ) | ( n2918 & n35410 ) | ( n33372 & n35410 ) ;
  assign n35412 = n26279 ^ n23040 ^ n17925 ;
  assign n35413 = ( n7363 & n10643 ) | ( n7363 & ~n24973 ) | ( n10643 & ~n24973 ) ;
  assign n35414 = n980 & ~n17466 ;
  assign n35415 = ~n10062 & n35414 ;
  assign n35416 = ( n24270 & n35413 ) | ( n24270 & ~n35415 ) | ( n35413 & ~n35415 ) ;
  assign n35417 = ~n1574 & n16755 ;
  assign n35418 = n13062 & ~n31988 ;
  assign n35419 = n35417 & n35418 ;
  assign n35420 = n4298 & ~n22313 ;
  assign n35422 = ~n12658 & n20422 ;
  assign n35423 = n33955 & n35422 ;
  assign n35424 = n35423 ^ n14826 ^ n11968 ;
  assign n35421 = n14294 | n20298 ;
  assign n35425 = n35424 ^ n35421 ^ 1'b0 ;
  assign n35428 = n7535 ^ n7186 ^ 1'b0 ;
  assign n35429 = n688 & n35428 ;
  assign n35430 = n23030 & n35429 ;
  assign n35431 = n20470 & n35430 ;
  assign n35432 = n35431 ^ n12404 ^ 1'b0 ;
  assign n35433 = n8482 & ~n35432 ;
  assign n35426 = n14363 | n20725 ;
  assign n35427 = ~n28303 & n35426 ;
  assign n35434 = n35433 ^ n35427 ^ 1'b0 ;
  assign n35435 = n1666 & ~n16038 ;
  assign n35436 = n35435 ^ n5129 ^ 1'b0 ;
  assign n35437 = n19917 | n35436 ;
  assign n35438 = n35437 ^ n17139 ^ n480 ;
  assign n35439 = n19570 & n35438 ;
  assign n35440 = n35439 ^ n2280 ^ 1'b0 ;
  assign n35445 = ( n4782 & n8785 ) | ( n4782 & n26754 ) | ( n8785 & n26754 ) ;
  assign n35446 = ~n11286 & n35445 ;
  assign n35447 = n1744 & n35446 ;
  assign n35443 = n9895 & n34989 ;
  assign n35441 = ( n5113 & n9110 ) | ( n5113 & n10699 ) | ( n9110 & n10699 ) ;
  assign n35442 = ~n5494 & n35441 ;
  assign n35444 = n35443 ^ n35442 ^ 1'b0 ;
  assign n35448 = n35447 ^ n35444 ^ n2118 ;
  assign n35449 = n16605 | n19758 ;
  assign n35450 = n35449 ^ n7513 ^ 1'b0 ;
  assign n35451 = n7657 & n35450 ;
  assign n35452 = n35451 ^ n16060 ^ 1'b0 ;
  assign n35453 = n12711 | n22956 ;
  assign n35454 = n469 | n35453 ;
  assign n35455 = n35454 ^ n6703 ^ 1'b0 ;
  assign n35456 = n16796 | n17023 ;
  assign n35457 = n3002 ^ n1153 ^ 1'b0 ;
  assign n35458 = ~n5132 & n10617 ;
  assign n35459 = n35458 ^ n3684 ^ 1'b0 ;
  assign n35460 = n33148 | n35459 ;
  assign n35461 = n35457 & n35460 ;
  assign n35462 = ( ~n1023 & n12097 ) | ( ~n1023 & n13524 ) | ( n12097 & n13524 ) ;
  assign n35463 = ~n1024 & n23917 ;
  assign n35464 = ~n9687 & n35463 ;
  assign n35465 = n13067 | n32467 ;
  assign n35466 = n35465 ^ n7503 ^ 1'b0 ;
  assign n35467 = n8203 & ~n18334 ;
  assign n35468 = ~n2460 & n35467 ;
  assign n35469 = n4807 & ~n7008 ;
  assign n35470 = n21646 ^ n6264 ^ 1'b0 ;
  assign n35471 = n9628 ^ n4977 ^ n4497 ;
  assign n35472 = n2177 ^ n381 ^ 1'b0 ;
  assign n35473 = n35472 ^ n6901 ^ 1'b0 ;
  assign n35474 = n30791 ^ n23456 ^ 1'b0 ;
  assign n35475 = n17771 & n18324 ;
  assign n35476 = n35475 ^ n22874 ^ 1'b0 ;
  assign n35477 = n35476 ^ n31260 ^ n14095 ;
  assign n35483 = n263 & n1789 ;
  assign n35484 = n7017 & ~n35483 ;
  assign n35485 = n35484 ^ n6155 ^ 1'b0 ;
  assign n35486 = n6370 | n35485 ;
  assign n35478 = n765 | n1585 ;
  assign n35479 = n765 & ~n35478 ;
  assign n35480 = n17595 | n35479 ;
  assign n35481 = n35479 & ~n35480 ;
  assign n35482 = n4610 | n35481 ;
  assign n35487 = n35486 ^ n35482 ^ 1'b0 ;
  assign n35488 = n6790 | n35487 ;
  assign n35489 = n35488 ^ n22003 ^ 1'b0 ;
  assign n35490 = n14829 ^ n4969 ^ 1'b0 ;
  assign n35491 = ~n5384 & n35490 ;
  assign n35492 = n29423 ^ n1307 ^ 1'b0 ;
  assign n35493 = n35491 & n35492 ;
  assign n35494 = n26559 ^ n20866 ^ 1'b0 ;
  assign n35495 = n8683 & ~n13876 ;
  assign n35496 = n35495 ^ n28068 ^ 1'b0 ;
  assign n35497 = n1213 & ~n35496 ;
  assign n35498 = n35497 ^ n8296 ^ 1'b0 ;
  assign n35499 = n20830 ^ n2014 ^ 1'b0 ;
  assign n35500 = n7248 | n29729 ;
  assign n35501 = n35500 ^ n12759 ^ 1'b0 ;
  assign n35502 = ( ~n20255 & n35499 ) | ( ~n20255 & n35501 ) | ( n35499 & n35501 ) ;
  assign n35503 = n15586 | n28191 ;
  assign n35504 = n35503 ^ n8181 ^ 1'b0 ;
  assign n35505 = n21132 ^ n18240 ^ n16589 ;
  assign n35506 = n2199 & n12852 ;
  assign n35507 = n35506 ^ n28805 ^ 1'b0 ;
  assign n35508 = n19079 & n35507 ;
  assign n35509 = n10775 & ~n18039 ;
  assign n35510 = ~n6846 & n35509 ;
  assign n35511 = n580 & ~n19335 ;
  assign n35512 = ~n6545 & n35511 ;
  assign n35514 = n3773 | n10491 ;
  assign n35515 = n35514 ^ n13725 ^ 1'b0 ;
  assign n35513 = ~n18929 & n29631 ;
  assign n35516 = n35515 ^ n35513 ^ 1'b0 ;
  assign n35517 = ( n14533 & n25293 ) | ( n14533 & n35516 ) | ( n25293 & n35516 ) ;
  assign n35518 = ~n5101 & n17563 ;
  assign n35519 = n12174 | n15029 ;
  assign n35520 = n26560 & n31010 ;
  assign n35521 = n19608 ^ n12754 ^ 1'b0 ;
  assign n35522 = n12438 & n35521 ;
  assign n35523 = ( n609 & ~n24772 ) | ( n609 & n35522 ) | ( ~n24772 & n35522 ) ;
  assign n35524 = n14112 ^ n13011 ^ 1'b0 ;
  assign n35525 = n13071 ^ n11386 ^ 1'b0 ;
  assign n35526 = n10353 & ~n35525 ;
  assign n35527 = ( n10529 & n28213 ) | ( n10529 & n35257 ) | ( n28213 & n35257 ) ;
  assign n35528 = n35527 ^ n18794 ^ 1'b0 ;
  assign n35529 = ~n6390 & n31078 ;
  assign n35530 = n2787 | n22577 ;
  assign n35531 = ( n2180 & n27534 ) | ( n2180 & n29460 ) | ( n27534 & n29460 ) ;
  assign n35532 = n35531 ^ n24762 ^ 1'b0 ;
  assign n35533 = n24183 & ~n35532 ;
  assign n35534 = n8896 ^ n3341 ^ 1'b0 ;
  assign n35535 = n18192 | n20248 ;
  assign n35536 = n1959 | n35535 ;
  assign n35537 = ~n8695 & n35536 ;
  assign n35538 = n35537 ^ n28378 ^ 1'b0 ;
  assign n35539 = n35534 & n35538 ;
  assign n35540 = n20251 & n25462 ;
  assign n35541 = n3365 | n35540 ;
  assign n35542 = ( n2114 & ~n11697 ) | ( n2114 & n15850 ) | ( ~n11697 & n15850 ) ;
  assign n35543 = ~n23152 & n35542 ;
  assign n35544 = n27101 & n35543 ;
  assign n35545 = n30188 | n35544 ;
  assign n35546 = n15801 | n19244 ;
  assign n35547 = n35546 ^ n26307 ^ 1'b0 ;
  assign n35548 = ( n2271 & n12291 ) | ( n2271 & n33648 ) | ( n12291 & n33648 ) ;
  assign n35549 = n9596 ^ n7792 ^ 1'b0 ;
  assign n35550 = n35548 & ~n35549 ;
  assign n35551 = ~n13572 & n26389 ;
  assign n35552 = n35551 ^ n23302 ^ 1'b0 ;
  assign n35553 = n21183 & n35552 ;
  assign n35554 = n18145 & n35553 ;
  assign n35560 = n1642 & ~n29227 ;
  assign n35557 = n464 | n12833 ;
  assign n35555 = n10686 | n18745 ;
  assign n35556 = n1558 | n35555 ;
  assign n35558 = n35557 ^ n35556 ^ n8203 ;
  assign n35559 = n20513 & ~n35558 ;
  assign n35561 = n35560 ^ n35559 ^ 1'b0 ;
  assign n35563 = n23910 ^ n10973 ^ n6166 ;
  assign n35562 = ~n4835 & n11345 ;
  assign n35564 = n35563 ^ n35562 ^ n18831 ;
  assign n35565 = ~n9292 & n35564 ;
  assign n35566 = n35565 ^ n35178 ^ 1'b0 ;
  assign n35567 = ~n9380 & n30814 ;
  assign n35568 = n28199 & n35567 ;
  assign n35569 = n14361 | n27788 ;
  assign n35570 = ( n1561 & ~n23441 ) | ( n1561 & n35569 ) | ( ~n23441 & n35569 ) ;
  assign n35571 = n177 & n2484 ;
  assign n35572 = ~n1153 & n35571 ;
  assign n35573 = n14537 & ~n35572 ;
  assign n35574 = ~n1311 & n35573 ;
  assign n35575 = n35574 ^ n34881 ^ n9928 ;
  assign n35576 = n6981 & ~n7171 ;
  assign n35577 = n35576 ^ n1231 ^ 1'b0 ;
  assign n35580 = n16704 | n31514 ;
  assign n35581 = n31233 | n35580 ;
  assign n35578 = n25011 ^ n6716 ^ 1'b0 ;
  assign n35579 = n10875 & ~n35578 ;
  assign n35582 = n35581 ^ n35579 ^ 1'b0 ;
  assign n35585 = n12845 ^ n961 ^ 1'b0 ;
  assign n35583 = ~n28487 & n29341 ;
  assign n35584 = n35583 ^ n126 ^ 1'b0 ;
  assign n35586 = n35585 ^ n35584 ^ n8638 ;
  assign n35587 = n20401 ^ n861 ^ 1'b0 ;
  assign n35588 = n1888 & n27049 ;
  assign n35589 = n35588 ^ n24074 ^ 1'b0 ;
  assign n35590 = n7763 | n11615 ;
  assign n35591 = n316 & n3909 ;
  assign n35592 = n35591 ^ n14866 ^ 1'b0 ;
  assign n35593 = ~n24482 & n35592 ;
  assign n35594 = n5178 | n15779 ;
  assign n35595 = n35593 | n35594 ;
  assign n35596 = n35595 ^ n4044 ^ 1'b0 ;
  assign n35597 = n12801 & n26344 ;
  assign n35598 = n19541 & n31684 ;
  assign n35599 = ~n21378 & n35598 ;
  assign n35601 = n34407 ^ n2076 ^ 1'b0 ;
  assign n35600 = n24220 ^ n9050 ^ 1'b0 ;
  assign n35602 = n35601 ^ n35600 ^ n22679 ;
  assign n35603 = n4925 & n35602 ;
  assign n35604 = n10830 & n35603 ;
  assign n35605 = n6816 ^ n2434 ^ 1'b0 ;
  assign n35606 = n35605 ^ n31588 ^ n2098 ;
  assign n35607 = n14920 | n34111 ;
  assign n35608 = ~n3191 & n17869 ;
  assign n35611 = n10722 ^ n4584 ^ 1'b0 ;
  assign n35609 = n22682 | n26603 ;
  assign n35610 = n3088 & n35609 ;
  assign n35612 = n35611 ^ n35610 ^ 1'b0 ;
  assign n35613 = n12340 ^ n10541 ^ n3581 ;
  assign n35614 = n3726 & n5295 ;
  assign n35615 = n23302 & n35614 ;
  assign n35616 = n35615 ^ n12088 ^ 1'b0 ;
  assign n35617 = ~n12641 & n35616 ;
  assign n35618 = n13771 ^ n9408 ^ n707 ;
  assign n35619 = n21370 & n35618 ;
  assign n35622 = n31653 ^ n14347 ^ n12611 ;
  assign n35621 = n9528 & n19041 ;
  assign n35623 = n35622 ^ n35621 ^ 1'b0 ;
  assign n35624 = n1522 | n16911 ;
  assign n35625 = n35623 & ~n35624 ;
  assign n35626 = n35625 ^ n27309 ^ 1'b0 ;
  assign n35620 = n10341 | n33585 ;
  assign n35627 = n35626 ^ n35620 ^ 1'b0 ;
  assign n35628 = ~n3329 & n23081 ;
  assign n35629 = n26273 ^ n1976 ^ 1'b0 ;
  assign n35630 = ~n736 & n12375 ;
  assign n35631 = n21753 & n35630 ;
  assign n35632 = n17658 ^ n17365 ^ 1'b0 ;
  assign n35633 = n35631 | n35632 ;
  assign n35634 = n12346 & n35633 ;
  assign n35635 = n16476 | n24305 ;
  assign n35636 = n4936 & n15026 ;
  assign n35637 = n5219 & n35636 ;
  assign n35638 = ~n35635 & n35637 ;
  assign n35639 = n289 & n6784 ;
  assign n35640 = n18438 & n35639 ;
  assign n35641 = n35640 ^ n1490 ^ 1'b0 ;
  assign n35642 = n4588 | n35641 ;
  assign n35643 = n23537 ^ n2148 ^ 1'b0 ;
  assign n35644 = n4055 & n7868 ;
  assign n35646 = n20791 | n31063 ;
  assign n35647 = n35646 ^ n25219 ^ n10139 ;
  assign n35645 = n20399 ^ n17351 ^ n10140 ;
  assign n35648 = n35647 ^ n35645 ^ n31675 ;
  assign n35649 = ~n1766 & n2125 ;
  assign n35650 = n2708 & n35649 ;
  assign n35651 = ( n6129 & n7704 ) | ( n6129 & ~n35650 ) | ( n7704 & ~n35650 ) ;
  assign n35652 = n35651 ^ n2670 ^ 1'b0 ;
  assign n35653 = n35652 ^ n15671 ^ n11266 ;
  assign n35654 = n23726 & ~n35653 ;
  assign n35655 = n35654 ^ n10309 ^ 1'b0 ;
  assign n35656 = n12296 ^ n9631 ^ 1'b0 ;
  assign n35657 = ~n9388 & n35656 ;
  assign n35658 = n5714 | n10598 ;
  assign n35659 = n12060 ^ n6916 ^ 1'b0 ;
  assign n35660 = ( ~n7407 & n11149 ) | ( ~n7407 & n35659 ) | ( n11149 & n35659 ) ;
  assign n35661 = n6328 | n35660 ;
  assign n35662 = n35661 ^ n23745 ^ 1'b0 ;
  assign n35665 = n13352 ^ n12659 ^ n9139 ;
  assign n35666 = n35665 ^ n15257 ^ 1'b0 ;
  assign n35663 = n11170 ^ n1006 ^ 1'b0 ;
  assign n35664 = n6319 | n35663 ;
  assign n35667 = n35666 ^ n35664 ^ 1'b0 ;
  assign n35668 = n21110 & ~n22360 ;
  assign n35669 = n2797 ^ n68 ^ 1'b0 ;
  assign n35670 = n18493 | n35669 ;
  assign n35671 = n3364 | n23457 ;
  assign n35672 = n10329 & ~n35671 ;
  assign n35673 = n15712 | n35672 ;
  assign n35676 = n3967 ^ n1509 ^ 1'b0 ;
  assign n35677 = n7222 | n35676 ;
  assign n35678 = n35677 ^ n8119 ^ 1'b0 ;
  assign n35679 = ~n5973 & n35678 ;
  assign n35674 = n11513 & ~n29991 ;
  assign n35675 = n35674 ^ n5339 ^ 1'b0 ;
  assign n35680 = n35679 ^ n35675 ^ 1'b0 ;
  assign n35684 = n16693 ^ n4558 ^ 1'b0 ;
  assign n35681 = ~n5754 & n14169 ;
  assign n35682 = n35681 ^ n15097 ^ 1'b0 ;
  assign n35683 = ( n1805 & n17388 ) | ( n1805 & ~n35682 ) | ( n17388 & ~n35682 ) ;
  assign n35685 = n35684 ^ n35683 ^ 1'b0 ;
  assign n35686 = n35685 ^ n11764 ^ 1'b0 ;
  assign n35687 = n3447 & n19657 ;
  assign n35688 = n35687 ^ n23550 ^ 1'b0 ;
  assign n35689 = n849 | n1548 ;
  assign n35690 = n849 & ~n35689 ;
  assign n35691 = x9 & ~n49 ;
  assign n35692 = n49 & n35691 ;
  assign n35693 = x3 & ~n35692 ;
  assign n35694 = ~x3 & n35693 ;
  assign n35695 = x9 & n18 ;
  assign n35696 = ~x3 & n35695 ;
  assign n35697 = n23 | n49 ;
  assign n35698 = n35696 & ~n35697 ;
  assign n35699 = n35694 | n35698 ;
  assign n35700 = n35694 & ~n35699 ;
  assign n35701 = n893 | n35700 ;
  assign n35702 = n35700 & ~n35701 ;
  assign n35703 = n46 & n99 ;
  assign n35704 = ~n99 & n35703 ;
  assign n35705 = n26 & ~n35704 ;
  assign n35706 = n35704 & n35705 ;
  assign n35707 = n205 | n35706 ;
  assign n35708 = n205 & ~n35707 ;
  assign n35709 = n35702 | n35708 ;
  assign n35710 = n35702 & ~n35709 ;
  assign n35711 = n473 & ~n686 ;
  assign n35712 = ~n473 & n35711 ;
  assign n35713 = n934 | n35712 ;
  assign n35714 = n35710 & ~n35713 ;
  assign n35715 = n35690 | n35714 ;
  assign n35716 = n35715 ^ n3334 ^ 1'b0 ;
  assign n35717 = n35342 ^ n466 ^ 1'b0 ;
  assign n35718 = n35716 & ~n35717 ;
  assign n35719 = n1837 & ~n5393 ;
  assign n35720 = n35719 ^ n33736 ^ 1'b0 ;
  assign n35721 = n6924 | n13543 ;
  assign n35722 = ~n8387 & n35721 ;
  assign n35723 = n35722 ^ n20129 ^ n14244 ;
  assign n35724 = n10775 ^ n221 ^ 1'b0 ;
  assign n35725 = n14497 ^ n11225 ^ 1'b0 ;
  assign n35726 = n31948 ^ n31199 ^ n11051 ;
  assign n35727 = n20366 ^ n12302 ^ 1'b0 ;
  assign n35728 = n33003 & ~n35727 ;
  assign n35729 = n26082 ^ n5715 ^ 1'b0 ;
  assign n35730 = n2143 | n2610 ;
  assign n35731 = n32691 & ~n35730 ;
  assign n35732 = n4799 & ~n28991 ;
  assign n35733 = n34994 & ~n35732 ;
  assign n35734 = n30338 ^ n4490 ^ 1'b0 ;
  assign n35735 = ( n4587 & ~n20950 ) | ( n4587 & n35734 ) | ( ~n20950 & n35734 ) ;
  assign n35736 = n10430 ^ n162 ^ 1'b0 ;
  assign n35737 = ( ~n15177 & n26316 ) | ( ~n15177 & n30543 ) | ( n26316 & n30543 ) ;
  assign n35738 = n15209 & ~n35737 ;
  assign n35740 = n32393 ^ n10111 ^ n816 ;
  assign n35741 = n35740 ^ n11393 ^ n11082 ;
  assign n35739 = ~n45 & n35358 ;
  assign n35742 = n35741 ^ n35739 ^ 1'b0 ;
  assign n35743 = n1660 | n35742 ;
  assign n35744 = n35743 ^ n4650 ^ 1'b0 ;
  assign n35745 = n4999 & n6640 ;
  assign n35746 = n35745 ^ n15360 ^ 1'b0 ;
  assign n35747 = ( n825 & ~n1506 ) | ( n825 & n35746 ) | ( ~n1506 & n35746 ) ;
  assign n35748 = n16203 & ~n35747 ;
  assign n35749 = n35748 ^ n30636 ^ n21000 ;
  assign n35750 = n26289 ^ n9216 ^ 1'b0 ;
  assign n35753 = n3477 ^ n2249 ^ 1'b0 ;
  assign n35754 = n1072 & ~n35753 ;
  assign n35751 = n28876 ^ n5886 ^ 1'b0 ;
  assign n35752 = n4810 & n35751 ;
  assign n35755 = n35754 ^ n35752 ^ 1'b0 ;
  assign n35756 = n124 | n9917 ;
  assign n35757 = n34448 ^ n26496 ^ n17729 ;
  assign n35758 = n27167 | n35757 ;
  assign n35760 = n7357 | n11321 ;
  assign n35759 = n28333 ^ n22662 ^ n4322 ;
  assign n35761 = n35760 ^ n35759 ^ n32616 ;
  assign n35762 = n25885 ^ n12273 ^ 1'b0 ;
  assign n35763 = n35762 ^ n3819 ^ 1'b0 ;
  assign n35764 = n3075 & ~n9911 ;
  assign n35765 = n8063 & n35764 ;
  assign n35766 = n7119 & ~n24844 ;
  assign n35767 = n5565 & n16077 ;
  assign n35768 = n19807 ^ n11233 ^ 1'b0 ;
  assign n35769 = n23214 & ~n29973 ;
  assign n35770 = n15799 & ~n29471 ;
  assign n35771 = ~n8493 & n30058 ;
  assign n35772 = n35771 ^ n33834 ^ 1'b0 ;
  assign n35773 = n12698 & n29492 ;
  assign n35774 = n27534 ^ n17743 ^ 1'b0 ;
  assign n35775 = n8872 & ~n15739 ;
  assign n35776 = n35775 ^ n33936 ^ 1'b0 ;
  assign n35777 = n3811 & ~n29368 ;
  assign n35778 = n5719 ^ n5233 ^ 1'b0 ;
  assign n35779 = ( ~n177 & n12155 ) | ( ~n177 & n35778 ) | ( n12155 & n35778 ) ;
  assign n35780 = n24260 ^ n23190 ^ 1'b0 ;
  assign n35781 = n17280 & ~n35780 ;
  assign n35782 = n130 | n34008 ;
  assign n35783 = n21529 | n26799 ;
  assign n35784 = n8355 & ~n35783 ;
  assign n35802 = ~n4045 & n4752 ;
  assign n35803 = ~n4752 & n35802 ;
  assign n35804 = ~n6468 & n35803 ;
  assign n35785 = n130 & ~n2806 ;
  assign n35786 = n2806 & n35785 ;
  assign n35787 = ~n4549 & n35786 ;
  assign n35788 = n2651 & ~n35787 ;
  assign n35790 = ~n361 & n3551 ;
  assign n35791 = n361 & n35790 ;
  assign n35792 = n30043 | n35791 ;
  assign n35793 = n30043 & ~n35792 ;
  assign n35794 = n2627 ^ n2441 ^ n1742 ;
  assign n35795 = n2090 & ~n12266 ;
  assign n35796 = n35795 ^ n10250 ^ 1'b0 ;
  assign n35797 = ~n35794 & n35796 ;
  assign n35798 = n35793 & n35797 ;
  assign n35799 = ~n13689 & n35798 ;
  assign n35789 = n33093 ^ n10467 ^ n9823 ;
  assign n35800 = n35799 ^ n35789 ^ n32062 ;
  assign n35801 = n35788 | n35800 ;
  assign n35805 = n35804 ^ n35801 ^ 1'b0 ;
  assign n35806 = n16347 ^ n5864 ^ 1'b0 ;
  assign n35807 = ( n3838 & ~n15086 ) | ( n3838 & n35806 ) | ( ~n15086 & n35806 ) ;
  assign n35808 = n12093 | n35807 ;
  assign n35809 = n25562 ^ n4523 ^ 1'b0 ;
  assign n35810 = ~n17793 & n35809 ;
  assign n35811 = n2876 & n3929 ;
  assign n35812 = n5557 & n14654 ;
  assign n35813 = n31770 & ~n35812 ;
  assign n35814 = ~n2890 & n35813 ;
  assign n35815 = n22546 | n23052 ;
  assign n35816 = n35815 ^ n29217 ^ 1'b0 ;
  assign n35817 = ( ~n4099 & n21713 ) | ( ~n4099 & n23563 ) | ( n21713 & n23563 ) ;
  assign n35818 = n35817 ^ n4656 ^ 1'b0 ;
  assign n35819 = n35818 ^ n435 ^ 1'b0 ;
  assign n35820 = n3864 ^ n1079 ^ 1'b0 ;
  assign n35821 = ( n21813 & ~n22740 ) | ( n21813 & n35820 ) | ( ~n22740 & n35820 ) ;
  assign n35822 = n1402 & n24647 ;
  assign n35823 = ~n27072 & n35822 ;
  assign n35824 = ~n2148 & n14037 ;
  assign n35825 = n35824 ^ n4544 ^ 1'b0 ;
  assign n35826 = n25927 & ~n35825 ;
  assign n35827 = n17099 ^ n12554 ^ 1'b0 ;
  assign n35828 = n13317 & n17738 ;
  assign n35829 = n35828 ^ n14013 ^ 1'b0 ;
  assign n35830 = n35829 ^ n16440 ^ n582 ;
  assign n35831 = n2245 | n10574 ;
  assign n35832 = n34249 | n35831 ;
  assign n35833 = n33273 | n35832 ;
  assign n35834 = n19465 & ~n35833 ;
  assign n35835 = n1274 | n35834 ;
  assign n35836 = n12143 ^ n7717 ^ n982 ;
  assign n35837 = n35836 ^ n22114 ^ 1'b0 ;
  assign n35838 = n25307 ^ n18969 ^ 1'b0 ;
  assign n35839 = n5100 & ~n35838 ;
  assign n35840 = n17077 | n19415 ;
  assign n35841 = n887 | n35840 ;
  assign n35842 = n21844 & n35841 ;
  assign n35843 = ~n35841 & n35842 ;
  assign n35844 = n14214 | n35660 ;
  assign n35845 = n5843 & ~n35844 ;
  assign n35846 = n10631 ^ n6205 ^ n2222 ;
  assign n35847 = n21494 ^ n6125 ^ 1'b0 ;
  assign n35848 = n3006 & n35847 ;
  assign n35849 = n35846 & n35848 ;
  assign n35850 = n7580 & n22013 ;
  assign n35851 = ~n27479 & n35850 ;
  assign n35852 = n1577 & ~n18591 ;
  assign n35853 = n35852 ^ n10240 ^ 1'b0 ;
  assign n35854 = n11273 ^ n1938 ^ 1'b0 ;
  assign n35855 = n11104 & n35854 ;
  assign n35856 = n3066 & n35855 ;
  assign n35857 = n18290 ^ n10356 ^ n3962 ;
  assign n35858 = n9183 ^ n8549 ^ 1'b0 ;
  assign n35859 = n33674 | n35858 ;
  assign n35860 = n34127 ^ n12129 ^ 1'b0 ;
  assign n35861 = n35860 ^ n27256 ^ 1'b0 ;
  assign n35862 = ~n29287 & n35861 ;
  assign n35863 = n14190 & ~n14799 ;
  assign n35864 = n5997 & ~n14286 ;
  assign n35865 = n27699 ^ n22240 ^ n5028 ;
  assign n35866 = n35865 ^ n11134 ^ 1'b0 ;
  assign n35867 = n31420 | n35866 ;
  assign n35868 = n31458 ^ n24699 ^ 1'b0 ;
  assign n35869 = n17468 ^ n6850 ^ 1'b0 ;
  assign n35870 = n27417 & ~n35869 ;
  assign n35871 = n8398 ^ n1172 ^ 1'b0 ;
  assign n35872 = n34943 ^ n4875 ^ 1'b0 ;
  assign n35873 = ~n12463 & n35872 ;
  assign n35874 = n29799 & n35873 ;
  assign n35875 = n18428 & ~n28774 ;
  assign n35876 = n361 & ~n27393 ;
  assign n35878 = n8327 ^ n6016 ^ 1'b0 ;
  assign n35877 = ~n5836 & n14093 ;
  assign n35879 = n35878 ^ n35877 ^ n5337 ;
  assign n35883 = n12439 ^ n6377 ^ n2523 ;
  assign n35880 = ~n1984 & n15315 ;
  assign n35881 = n19632 & ~n23592 ;
  assign n35882 = ~n35880 & n35881 ;
  assign n35884 = n35883 ^ n35882 ^ n25674 ;
  assign n35885 = n13001 & ~n34111 ;
  assign n35886 = n12935 ^ n1131 ^ 1'b0 ;
  assign n35887 = n14580 & ~n35886 ;
  assign n35888 = n23609 & n35887 ;
  assign n35889 = n35888 ^ n34983 ^ 1'b0 ;
  assign n35890 = n32792 ^ n19642 ^ 1'b0 ;
  assign n35891 = n27641 ^ n4799 ^ 1'b0 ;
  assign n35892 = ( n7140 & n25809 ) | ( n7140 & ~n32429 ) | ( n25809 & ~n32429 ) ;
  assign n35893 = n25596 & ~n29789 ;
  assign n35894 = n29801 & n35893 ;
  assign n35895 = n35894 ^ n2311 ^ 1'b0 ;
  assign n35896 = ~n35892 & n35895 ;
  assign n35897 = n21425 ^ n9823 ^ 1'b0 ;
  assign n35898 = n35897 ^ n32119 ^ 1'b0 ;
  assign n35899 = n6699 | n35898 ;
  assign n35900 = n628 | n17223 ;
  assign n35901 = n28641 ^ n12754 ^ 1'b0 ;
  assign n35902 = n10571 & n19444 ;
  assign n35903 = n17336 ^ n7702 ^ 1'b0 ;
  assign n35904 = n19347 ^ n13242 ^ 1'b0 ;
  assign n35905 = n35903 & n35904 ;
  assign n35906 = n8043 & n27607 ;
  assign n35907 = ~n6513 & n35906 ;
  assign n35908 = n35907 ^ n8025 ^ n5794 ;
  assign n35909 = n18519 ^ n13031 ^ n3573 ;
  assign n35910 = n35909 ^ n14112 ^ n5715 ;
  assign n35911 = n35910 ^ n12821 ^ 1'b0 ;
  assign n35912 = n35911 ^ n27135 ^ n15753 ;
  assign n35913 = n2070 | n3807 ;
  assign n35914 = n35913 ^ n23123 ^ 1'b0 ;
  assign n35915 = n31440 ^ n11281 ^ 1'b0 ;
  assign n35916 = n27205 & ~n35915 ;
  assign n35917 = n35579 ^ n11624 ^ 1'b0 ;
  assign n35918 = n7925 | n35917 ;
  assign n35919 = n23458 ^ n635 ^ 1'b0 ;
  assign n35920 = n33018 & n35919 ;
  assign n35921 = n35920 ^ n27936 ^ 1'b0 ;
  assign n35922 = n7037 | n30031 ;
  assign n35923 = ( n9560 & n14112 ) | ( n9560 & n15277 ) | ( n14112 & n15277 ) ;
  assign n35924 = n15776 ^ n9552 ^ 1'b0 ;
  assign n35925 = n18123 & ~n35924 ;
  assign n35926 = n30235 ^ n13951 ^ 1'b0 ;
  assign n35927 = n35926 ^ n26088 ^ 1'b0 ;
  assign n35928 = n16585 ^ n15683 ^ n7169 ;
  assign n35929 = n35928 ^ n15306 ^ 1'b0 ;
  assign n35930 = n28306 ^ n13023 ^ 1'b0 ;
  assign n35931 = n7754 & ~n35930 ;
  assign n35932 = n7040 & n12821 ;
  assign n35936 = n7300 ^ n5818 ^ 1'b0 ;
  assign n35937 = ~n3546 & n35936 ;
  assign n35938 = n35937 ^ n14042 ^ 1'b0 ;
  assign n35933 = ( n2375 & n2655 ) | ( n2375 & n7293 ) | ( n2655 & n7293 ) ;
  assign n35934 = n20375 ^ n7612 ^ n7416 ;
  assign n35935 = ~n35933 & n35934 ;
  assign n35939 = n35938 ^ n35935 ^ n4116 ;
  assign n35941 = n3855 | n4967 ;
  assign n35942 = n620 & n35941 ;
  assign n35940 = n19048 & ~n23837 ;
  assign n35943 = n35942 ^ n35940 ^ 1'b0 ;
  assign n35944 = n13243 ^ n875 ^ 1'b0 ;
  assign n35945 = n10720 & n35944 ;
  assign n35946 = n35945 ^ n33726 ^ 1'b0 ;
  assign n35947 = n34408 ^ n3148 ^ 1'b0 ;
  assign n35948 = n35946 & n35947 ;
  assign n35949 = ~n4287 & n8247 ;
  assign n35950 = n2266 & n13167 ;
  assign n35951 = n35950 ^ n23004 ^ 1'b0 ;
  assign n35952 = n35951 ^ n14878 ^ 1'b0 ;
  assign n35953 = n12164 & ~n31348 ;
  assign n35954 = ~n35952 & n35953 ;
  assign n35955 = n21114 ^ n4548 ^ 1'b0 ;
  assign n35956 = ~n8319 & n35955 ;
  assign n35957 = n34411 ^ n29318 ^ 1'b0 ;
  assign n35960 = n8211 ^ n6477 ^ 1'b0 ;
  assign n35961 = n18951 | n35960 ;
  assign n35958 = n11879 & ~n25151 ;
  assign n35959 = n4008 | n35958 ;
  assign n35962 = n35961 ^ n35959 ^ 1'b0 ;
  assign n35963 = n2791 & n5309 ;
  assign n35964 = n25349 | n35963 ;
  assign n35965 = n35964 ^ n3053 ^ 1'b0 ;
  assign n35966 = n16166 ^ n8891 ^ 1'b0 ;
  assign n35967 = n23565 & ~n25550 ;
  assign n35968 = ~n22374 & n35967 ;
  assign n35969 = n19084 ^ n12707 ^ n2106 ;
  assign n35970 = ~n22213 & n35969 ;
  assign n35971 = n35968 & n35970 ;
  assign n35972 = n13461 | n21724 ;
  assign n35973 = n15407 | n35972 ;
  assign n35974 = n913 & ~n6398 ;
  assign n35975 = n35974 ^ n11386 ^ 1'b0 ;
  assign n35976 = n9066 | n13953 ;
  assign n35977 = n35976 ^ n6212 ^ 1'b0 ;
  assign n35978 = n3404 & ~n9242 ;
  assign n35979 = n35978 ^ n27808 ^ 1'b0 ;
  assign n35980 = n18048 | n32060 ;
  assign n35981 = ~n8729 & n10481 ;
  assign n35982 = n6916 & n27449 ;
  assign n35983 = n35982 ^ n6447 ^ n1518 ;
  assign n35984 = n27855 & ~n35983 ;
  assign n35985 = n25421 & n35984 ;
  assign n35986 = n8248 & ~n35985 ;
  assign n35987 = ~n8697 & n11029 ;
  assign n35988 = ~n11955 & n35987 ;
  assign n35989 = n8449 | n13346 ;
  assign n35990 = n17496 ^ n4334 ^ 1'b0 ;
  assign n35991 = ~n35989 & n35990 ;
  assign n35992 = n29456 | n31786 ;
  assign n35993 = n35992 ^ n14380 ^ 1'b0 ;
  assign n35994 = n34189 ^ n28691 ^ n27690 ;
  assign n35995 = n5859 & ~n24697 ;
  assign n35996 = n35995 ^ n30091 ^ 1'b0 ;
  assign n35997 = n5394 ^ n1689 ^ 1'b0 ;
  assign n35998 = n14131 | n35997 ;
  assign n35999 = n8334 | n35998 ;
  assign n36000 = n688 | n35999 ;
  assign n36001 = n36000 ^ n13539 ^ n6355 ;
  assign n36002 = n34770 ^ n2148 ^ 1'b0 ;
  assign n36003 = n36001 & n36002 ;
  assign n36004 = n21142 ^ n8848 ^ 1'b0 ;
  assign n36005 = n23529 & n36004 ;
  assign n36006 = n36005 ^ n19821 ^ 1'b0 ;
  assign n36007 = n14858 ^ n5032 ^ 1'b0 ;
  assign n36008 = n14857 & n36007 ;
  assign n36009 = n9903 | n10254 ;
  assign n36010 = n13421 & ~n36009 ;
  assign n36011 = ~n36008 & n36010 ;
  assign n36012 = n551 | n36011 ;
  assign n36013 = n36012 ^ n2464 ^ 1'b0 ;
  assign n36014 = n36013 ^ n22048 ^ 1'b0 ;
  assign n36015 = n8018 ^ n1213 ^ 1'b0 ;
  assign n36016 = n4647 & ~n10093 ;
  assign n36017 = ~n3638 & n36016 ;
  assign n36018 = ~n14332 & n23779 ;
  assign n36019 = n36017 & n36018 ;
  assign n36020 = n36019 ^ n23397 ^ 1'b0 ;
  assign n36021 = n430 & n13677 ;
  assign n36022 = n11809 ^ n7414 ^ 1'b0 ;
  assign n36023 = ~n36021 & n36022 ;
  assign n36024 = ~n8319 & n21798 ;
  assign n36025 = n36024 ^ n2177 ^ 1'b0 ;
  assign n36026 = n18565 ^ n18451 ^ n4662 ;
  assign n36027 = ~n10164 & n36026 ;
  assign n36028 = n2776 & ~n4543 ;
  assign n36030 = ( n8300 & ~n10960 ) | ( n8300 & n12253 ) | ( ~n10960 & n12253 ) ;
  assign n36029 = n9253 ^ n4637 ^ n713 ;
  assign n36031 = n36030 ^ n36029 ^ n33624 ;
  assign n36032 = n772 & ~n23707 ;
  assign n36033 = n36032 ^ n8453 ^ 1'b0 ;
  assign n36038 = n9615 & ~n21510 ;
  assign n36039 = ~n2798 & n36038 ;
  assign n36034 = n892 | n13243 ;
  assign n36035 = n8625 & n28868 ;
  assign n36036 = n35335 | n36035 ;
  assign n36037 = ( n9230 & ~n36034 ) | ( n9230 & n36036 ) | ( ~n36034 & n36036 ) ;
  assign n36040 = n36039 ^ n36037 ^ 1'b0 ;
  assign n36043 = n237 | n12239 ;
  assign n36041 = n25833 ^ n5070 ^ 1'b0 ;
  assign n36042 = n31401 & n36041 ;
  assign n36044 = n36043 ^ n36042 ^ 1'b0 ;
  assign n36045 = ~n7945 & n15670 ;
  assign n36046 = n7945 & n36045 ;
  assign n36047 = n9081 | n36046 ;
  assign n36048 = n7561 & n19723 ;
  assign n36049 = n36047 & n36048 ;
  assign n36050 = ~n6389 & n14492 ;
  assign n36051 = n4543 ^ n3457 ^ 1'b0 ;
  assign n36052 = n9308 & ~n36051 ;
  assign n36053 = ~n19974 & n36052 ;
  assign n36054 = ~n41 & n36053 ;
  assign n36055 = n36050 & ~n36054 ;
  assign n36056 = ( n15940 & n29855 ) | ( n15940 & ~n36055 ) | ( n29855 & ~n36055 ) ;
  assign n36057 = ~n6074 & n17441 ;
  assign n36058 = ~n10769 & n23012 ;
  assign n36059 = n36058 ^ n12758 ^ 1'b0 ;
  assign n36060 = n15772 | n36059 ;
  assign n36061 = n10453 & n17838 ;
  assign n36062 = n28165 & ~n32813 ;
  assign n36063 = n11423 | n12428 ;
  assign n36064 = n36063 ^ n1079 ^ 1'b0 ;
  assign n36065 = n36064 ^ n27550 ^ 1'b0 ;
  assign n36066 = ( n14712 & ~n14791 ) | ( n14712 & n36065 ) | ( ~n14791 & n36065 ) ;
  assign n36067 = ~n3343 & n10557 ;
  assign n36068 = n36067 ^ n12292 ^ 1'b0 ;
  assign n36069 = n3620 & ~n15074 ;
  assign n36070 = n36069 ^ n21041 ^ 1'b0 ;
  assign n36071 = n13577 | n18404 ;
  assign n36072 = n36071 ^ n22128 ^ 1'b0 ;
  assign n36073 = ~n645 & n4468 ;
  assign n36074 = n26243 ^ n18984 ^ 1'b0 ;
  assign n36075 = ~n11724 & n32915 ;
  assign n36076 = n91 & n4826 ;
  assign n36077 = n13359 & n30046 ;
  assign n36078 = n36077 ^ n12358 ^ 1'b0 ;
  assign n36079 = n30196 ^ n29944 ^ n26449 ;
  assign n36080 = ~n30 & n19277 ;
  assign n36081 = ~n1609 & n3682 ;
  assign n36082 = ~n34574 & n36081 ;
  assign n36083 = ~n238 & n15421 ;
  assign n36084 = n4052 & n36083 ;
  assign n36085 = n35880 ^ n48 ^ 1'b0 ;
  assign n36086 = n36084 | n36085 ;
  assign n36087 = n7498 & ~n11519 ;
  assign n36088 = n36086 & n36087 ;
  assign n36089 = n15072 & ~n16162 ;
  assign n36090 = n36089 ^ n11098 ^ 1'b0 ;
  assign n36091 = n36090 ^ n3588 ^ 1'b0 ;
  assign n36092 = ( n12808 & ~n21061 ) | ( n12808 & n36091 ) | ( ~n21061 & n36091 ) ;
  assign n36093 = n32796 ^ n28984 ^ 1'b0 ;
  assign n36094 = n17295 | n21972 ;
  assign n36095 = n36093 | n36094 ;
  assign n36096 = n36095 ^ n25397 ^ n13827 ;
  assign n36097 = n36096 ^ n9770 ^ 1'b0 ;
  assign n36098 = n5109 & ~n36097 ;
  assign n36099 = n2435 & n36098 ;
  assign n36100 = n27146 ^ n14619 ^ n13337 ;
  assign n36101 = n24994 ^ n1918 ^ 1'b0 ;
  assign n36102 = n33402 ^ n2352 ^ 1'b0 ;
  assign n36103 = ~n2982 & n23914 ;
  assign n36104 = x10 | n17484 ;
  assign n36105 = n6115 & ~n9734 ;
  assign n36107 = n7749 ^ n854 ^ n383 ;
  assign n36108 = n36107 ^ n23733 ^ 1'b0 ;
  assign n36106 = ~n6075 & n8206 ;
  assign n36109 = n36108 ^ n36106 ^ 1'b0 ;
  assign n36110 = n31933 ^ n8797 ^ 1'b0 ;
  assign n36111 = n36109 | n36110 ;
  assign n36112 = n523 | n35926 ;
  assign n36113 = n34175 & n36112 ;
  assign n36114 = n16127 ^ n6938 ^ 1'b0 ;
  assign n36115 = ~n36113 & n36114 ;
  assign n36116 = n30339 ^ n14797 ^ 1'b0 ;
  assign n36117 = n3420 & n13537 ;
  assign n36118 = n1889 | n26546 ;
  assign n36119 = n36109 & ~n36118 ;
  assign n36120 = n25658 ^ n15728 ^ n6481 ;
  assign n36121 = n36120 ^ n9275 ^ 1'b0 ;
  assign n36122 = n25531 & n34256 ;
  assign n36123 = n3067 & n36122 ;
  assign n36124 = ( n18835 & n23615 ) | ( n18835 & ~n36123 ) | ( n23615 & ~n36123 ) ;
  assign n36125 = ~n12241 & n16035 ;
  assign n36126 = n36125 ^ n5831 ^ 1'b0 ;
  assign n36127 = n14466 & ~n36126 ;
  assign n36128 = n10079 ^ n5628 ^ 1'b0 ;
  assign n36129 = n16303 & ~n36128 ;
  assign n36130 = n22564 & ~n24272 ;
  assign n36131 = n29729 & n36130 ;
  assign n36132 = ( n8824 & n23535 ) | ( n8824 & n27533 ) | ( n23535 & n27533 ) ;
  assign n36133 = n18317 | n35182 ;
  assign n36134 = n36133 ^ n8688 ^ 1'b0 ;
  assign n36135 = n3652 | n17245 ;
  assign n36136 = n5854 & n26088 ;
  assign n36137 = n36136 ^ n16575 ^ 1'b0 ;
  assign n36138 = n10650 & ~n15802 ;
  assign n36139 = n36138 ^ n22549 ^ 1'b0 ;
  assign n36140 = n12005 ^ n9285 ^ 1'b0 ;
  assign n36141 = n24049 & ~n36140 ;
  assign n36142 = ~n15972 & n36141 ;
  assign n36143 = ( n6431 & n15470 ) | ( n6431 & n28173 ) | ( n15470 & n28173 ) ;
  assign n36144 = n36143 ^ n12932 ^ 1'b0 ;
  assign n36145 = n36144 ^ n11922 ^ 1'b0 ;
  assign n36146 = ~n972 & n2563 ;
  assign n36147 = n36146 ^ n8799 ^ 1'b0 ;
  assign n36148 = n36 | n29109 ;
  assign n36149 = n27180 ^ n10695 ^ 1'b0 ;
  assign n36150 = n10617 & n36149 ;
  assign n36152 = n1058 & ~n2403 ;
  assign n36153 = ~n3932 & n36152 ;
  assign n36151 = n1825 & n8278 ;
  assign n36154 = n36153 ^ n36151 ^ 1'b0 ;
  assign n36155 = n34989 ^ n2597 ^ 1'b0 ;
  assign n36156 = n13291 & ~n36155 ;
  assign n36157 = n36156 ^ n4288 ^ 1'b0 ;
  assign n36158 = n1151 & ~n18973 ;
  assign n36159 = ~n11361 & n36158 ;
  assign n36160 = n4628 & n34014 ;
  assign n36161 = n21436 & n28014 ;
  assign n36164 = n5876 & n10349 ;
  assign n36165 = n5815 | n36164 ;
  assign n36162 = n11340 & n12220 ;
  assign n36163 = n36162 ^ n1303 ^ 1'b0 ;
  assign n36166 = n36165 ^ n36163 ^ 1'b0 ;
  assign n36167 = n36166 ^ n30347 ^ n27095 ;
  assign n36168 = ( ~n16224 & n27415 ) | ( ~n16224 & n32347 ) | ( n27415 & n32347 ) ;
  assign n36169 = n10484 & ~n27258 ;
  assign n36170 = n36169 ^ n13760 ^ 1'b0 ;
  assign n36171 = n20311 ^ n14354 ^ n10353 ;
  assign n36172 = n12396 & n36171 ;
  assign n36173 = n6039 & n36172 ;
  assign n36174 = n6804 | n36173 ;
  assign n36175 = n25627 & ~n36174 ;
  assign n36176 = n22127 & ~n29351 ;
  assign n36177 = ~n12963 & n36176 ;
  assign n36178 = n21220 & ~n27863 ;
  assign n36179 = n12281 | n36178 ;
  assign n36180 = ( n702 & n1010 ) | ( n702 & n25707 ) | ( n1010 & n25707 ) ;
  assign n36181 = ( ~n8722 & n30256 ) | ( ~n8722 & n36180 ) | ( n30256 & n36180 ) ;
  assign n36182 = n17384 ^ n16200 ^ 1'b0 ;
  assign n36183 = n8631 & ~n36182 ;
  assign n36184 = n29593 ^ n14962 ^ 1'b0 ;
  assign n36185 = n849 & ~n3393 ;
  assign n36186 = n29726 & n36185 ;
  assign n36187 = n14752 & n36186 ;
  assign n36188 = ~n6684 & n8356 ;
  assign n36189 = ( ~n2694 & n20137 ) | ( ~n2694 & n36188 ) | ( n20137 & n36188 ) ;
  assign n36190 = ~n9950 & n28748 ;
  assign n36191 = n16641 ^ n209 ^ 1'b0 ;
  assign n36192 = n25672 | n36191 ;
  assign n36193 = n8030 | n20173 ;
  assign n36194 = n32583 | n36193 ;
  assign n36195 = ~n7368 & n16575 ;
  assign n36196 = ~n36194 & n36195 ;
  assign n36197 = n33252 ^ n32691 ^ 1'b0 ;
  assign n36198 = ~n9095 & n9246 ;
  assign n36199 = n8655 & n36198 ;
  assign n36200 = n9948 ^ n7357 ^ 1'b0 ;
  assign n36201 = n36200 ^ n20361 ^ n9430 ;
  assign n36202 = n36201 ^ n14086 ^ 1'b0 ;
  assign n36203 = ( n10839 & n28291 ) | ( n10839 & n36202 ) | ( n28291 & n36202 ) ;
  assign n36204 = n35197 ^ n15193 ^ n1803 ;
  assign n36205 = n73 & n11443 ;
  assign n36206 = n15767 ^ n4545 ^ 1'b0 ;
  assign n36207 = ~n19509 & n36206 ;
  assign n36208 = n26470 & ~n36207 ;
  assign n36209 = n2616 ^ n982 ^ 1'b0 ;
  assign n36210 = n36209 ^ n6880 ^ 1'b0 ;
  assign n36211 = n11919 & n36210 ;
  assign n36212 = n28765 & n31277 ;
  assign n36213 = n11204 ^ n575 ^ 1'b0 ;
  assign n36214 = n26983 | n36213 ;
  assign n36215 = n18679 | n30322 ;
  assign n36216 = n15292 ^ n13891 ^ n1706 ;
  assign n36217 = n35491 & n36216 ;
  assign n36218 = n6080 & n18076 ;
  assign n36219 = n28039 & n36218 ;
  assign n36220 = n36219 ^ n33801 ^ n9664 ;
  assign n36221 = n368 & ~n28669 ;
  assign n36222 = n36221 ^ n11033 ^ 1'b0 ;
  assign n36223 = ~n3375 & n36222 ;
  assign n36225 = n28292 ^ n5768 ^ 1'b0 ;
  assign n36224 = n7287 & ~n20439 ;
  assign n36226 = n36225 ^ n36224 ^ 1'b0 ;
  assign n36227 = n17349 & n20924 ;
  assign n36228 = n36227 ^ n16786 ^ 1'b0 ;
  assign n36229 = n24714 & n36228 ;
  assign n36230 = n14522 & n36229 ;
  assign n36231 = ( n9823 & ~n21867 ) | ( n9823 & n36230 ) | ( ~n21867 & n36230 ) ;
  assign n36232 = n19961 ^ n9248 ^ 1'b0 ;
  assign n36233 = n31055 ^ n26574 ^ 1'b0 ;
  assign n36234 = n36232 | n36233 ;
  assign n36235 = n36231 & ~n36234 ;
  assign n36236 = n36235 ^ n20289 ^ 1'b0 ;
  assign n36237 = n9830 ^ n637 ^ 1'b0 ;
  assign n36238 = n11402 & ~n36237 ;
  assign n36239 = n36238 ^ n10690 ^ n5209 ;
  assign n36240 = n2646 & ~n13256 ;
  assign n36242 = n14838 ^ n5324 ^ 1'b0 ;
  assign n36243 = n16146 & n36242 ;
  assign n36241 = n25650 & ~n33162 ;
  assign n36244 = n36243 ^ n36241 ^ 1'b0 ;
  assign n36245 = n20715 | n36244 ;
  assign n36246 = n77 | n36245 ;
  assign n36247 = n8143 ^ n1585 ^ 1'b0 ;
  assign n36248 = ~n33861 & n36247 ;
  assign n36249 = n11341 & n17165 ;
  assign n36250 = ~n12264 & n36249 ;
  assign n36251 = ( ~n4072 & n28374 ) | ( ~n4072 & n36250 ) | ( n28374 & n36250 ) ;
  assign n36252 = n36251 ^ n27545 ^ 1'b0 ;
  assign n36253 = n21569 & n36252 ;
  assign n36254 = n1642 | n6430 ;
  assign n36255 = n1642 & ~n36254 ;
  assign n36256 = ( n661 & ~n7133 ) | ( n661 & n36255 ) | ( ~n7133 & n36255 ) ;
  assign n36257 = n36256 ^ n9760 ^ 1'b0 ;
  assign n36258 = ~n3866 & n36257 ;
  assign n36259 = n1815 | n10305 ;
  assign n36260 = n36259 ^ n5370 ^ 1'b0 ;
  assign n36261 = n8385 & n21571 ;
  assign n36262 = n36260 & n36261 ;
  assign n36263 = ~n15746 & n31285 ;
  assign n36264 = n34189 ^ n17419 ^ n9167 ;
  assign n36265 = n18355 & n36264 ;
  assign n36266 = n17244 & n33021 ;
  assign n36267 = n20772 ^ n9449 ^ 1'b0 ;
  assign n36268 = ~n10550 & n36267 ;
  assign n36269 = n36266 & ~n36268 ;
  assign n36270 = n36269 ^ n35510 ^ n11079 ;
  assign n36271 = ( n884 & ~n13438 ) | ( n884 & n14011 ) | ( ~n13438 & n14011 ) ;
  assign n36272 = n16873 ^ n10114 ^ 1'b0 ;
  assign n36273 = n27689 ^ n25504 ^ n12119 ;
  assign n36274 = n1024 | n4605 ;
  assign n36275 = n36274 ^ n9171 ^ 1'b0 ;
  assign n36276 = n21660 ^ n11430 ^ 1'b0 ;
  assign n36277 = n3824 | n36276 ;
  assign n36278 = n20073 ^ n15837 ^ 1'b0 ;
  assign n36279 = n6491 & n11326 ;
  assign n36281 = n3989 & n12931 ;
  assign n36282 = ~n3989 & n36281 ;
  assign n36283 = n2918 & n36282 ;
  assign n36284 = n7216 & ~n36283 ;
  assign n36285 = n36283 & n36284 ;
  assign n36280 = n10056 | n22205 ;
  assign n36286 = n36285 ^ n36280 ^ 1'b0 ;
  assign n36287 = n36286 ^ n9276 ^ 1'b0 ;
  assign n36288 = n2384 & ~n36287 ;
  assign n36289 = ( n13034 & ~n36279 ) | ( n13034 & n36288 ) | ( ~n36279 & n36288 ) ;
  assign n36290 = n3698 & ~n28968 ;
  assign n36291 = n14605 & n22520 ;
  assign n36292 = n1399 & n36291 ;
  assign n36293 = ( n10811 & ~n14980 ) | ( n10811 & n15411 ) | ( ~n14980 & n15411 ) ;
  assign n36294 = n36293 ^ n29162 ^ n15946 ;
  assign n36295 = n12500 ^ n536 ^ 1'b0 ;
  assign n36296 = n31644 ^ n20776 ^ 1'b0 ;
  assign n36297 = ( n11132 & n24226 ) | ( n11132 & ~n36296 ) | ( n24226 & ~n36296 ) ;
  assign n36298 = n25097 ^ n15588 ^ 1'b0 ;
  assign n36299 = n25338 ^ n15386 ^ 1'b0 ;
  assign n36300 = n10402 & ~n14294 ;
  assign n36301 = n36300 ^ n24305 ^ 1'b0 ;
  assign n36302 = n14007 | n36301 ;
  assign n36303 = ( n5844 & n36299 ) | ( n5844 & n36302 ) | ( n36299 & n36302 ) ;
  assign n36304 = n16940 ^ n8799 ^ n187 ;
  assign n36305 = n26975 | n36304 ;
  assign n36306 = n36303 & ~n36305 ;
  assign n36307 = ( n14505 & ~n16476 ) | ( n14505 & n31929 ) | ( ~n16476 & n31929 ) ;
  assign n36308 = n25396 ^ n9800 ^ 1'b0 ;
  assign n36309 = n2039 & ~n13983 ;
  assign n36310 = n15454 & n36309 ;
  assign n36311 = n7388 & n19510 ;
  assign n36312 = ( n1300 & n34624 ) | ( n1300 & n36311 ) | ( n34624 & n36311 ) ;
  assign n36313 = n6383 ^ n5112 ^ 1'b0 ;
  assign n36314 = n6523 & n36313 ;
  assign n36315 = n33690 & n36314 ;
  assign n36316 = n20812 ^ n8663 ^ 1'b0 ;
  assign n36317 = n36316 ^ n20355 ^ 1'b0 ;
  assign n36318 = n7630 & n36317 ;
  assign n36319 = ( n7965 & n17866 ) | ( n7965 & n36318 ) | ( n17866 & n36318 ) ;
  assign n36320 = ~n10779 & n28311 ;
  assign n36321 = n33 & ~n6552 ;
  assign n36322 = ~n27100 & n36321 ;
  assign n36323 = n11769 ^ n9240 ^ 1'b0 ;
  assign n36324 = n36322 | n36323 ;
  assign n36325 = n30420 & ~n32667 ;
  assign n36326 = n459 & ~n7987 ;
  assign n36327 = n36326 ^ n8001 ^ 1'b0 ;
  assign n36328 = n30597 | n32998 ;
  assign n36329 = n36328 ^ n15037 ^ 1'b0 ;
  assign n36330 = ( ~n21181 & n36327 ) | ( ~n21181 & n36329 ) | ( n36327 & n36329 ) ;
  assign n36331 = n31708 ^ n6919 ^ 1'b0 ;
  assign n36332 = n3308 | n36331 ;
  assign n36333 = n36332 ^ n31348 ^ 1'b0 ;
  assign n36334 = n3243 & ~n8133 ;
  assign n36335 = n36334 ^ n13631 ^ 1'b0 ;
  assign n36336 = n10504 ^ n9127 ^ n2813 ;
  assign n36338 = n24890 ^ n13117 ^ n5377 ;
  assign n36337 = ( n3263 & n18374 ) | ( n3263 & ~n33178 ) | ( n18374 & ~n33178 ) ;
  assign n36339 = n36338 ^ n36337 ^ n13893 ;
  assign n36340 = n20309 & n26743 ;
  assign n36341 = n36339 & n36340 ;
  assign n36342 = n9397 ^ n3294 ^ 1'b0 ;
  assign n36343 = n11825 ^ n7137 ^ 1'b0 ;
  assign n36344 = n10830 | n15602 ;
  assign n36345 = n20161 | n36344 ;
  assign n36346 = ~n804 & n14985 ;
  assign n36347 = n1263 & ~n36346 ;
  assign n36348 = n5998 | n18895 ;
  assign n36349 = n18104 & ~n36348 ;
  assign n36350 = ~n36347 & n36349 ;
  assign n36351 = ~n3543 & n12126 ;
  assign n36352 = n20382 & n36351 ;
  assign n36353 = n36352 ^ n34044 ^ 1'b0 ;
  assign n36354 = ( n9358 & n13121 ) | ( n9358 & ~n35410 ) | ( n13121 & ~n35410 ) ;
  assign n36355 = n36354 ^ n1965 ^ 1'b0 ;
  assign n36356 = n6759 & n18845 ;
  assign n36357 = n36356 ^ n17784 ^ 1'b0 ;
  assign n36358 = n27183 & n36357 ;
  assign n36359 = n27941 ^ n16768 ^ 1'b0 ;
  assign n36360 = n19925 ^ n4345 ^ 1'b0 ;
  assign n36361 = n3303 | n36360 ;
  assign n36362 = n36361 ^ n874 ^ 1'b0 ;
  assign n36363 = ~n4289 & n36362 ;
  assign n36364 = ~n5277 & n36363 ;
  assign n36365 = n9079 & n36364 ;
  assign n36366 = n6126 & ~n9928 ;
  assign n36367 = n30934 & n36366 ;
  assign n36368 = n1515 | n36367 ;
  assign n36369 = n36368 ^ n1459 ^ 1'b0 ;
  assign n36370 = ~n25154 & n27305 ;
  assign n36371 = ~n36369 & n36370 ;
  assign n36372 = ~n1800 & n28507 ;
  assign n36373 = n25737 & ~n30373 ;
  assign n36374 = n36373 ^ n21561 ^ n5679 ;
  assign n36375 = ~n423 & n10644 ;
  assign n36376 = n36375 ^ n4803 ^ 1'b0 ;
  assign n36377 = n6956 & n36376 ;
  assign n36378 = n36377 ^ n63 ^ 1'b0 ;
  assign n36379 = n36378 ^ n316 ^ 1'b0 ;
  assign n36380 = n36379 ^ n19727 ^ 1'b0 ;
  assign n36389 = n15571 ^ n14152 ^ n54 ;
  assign n36386 = ~n12292 & n15958 ;
  assign n36387 = n12575 ^ n7260 ^ 1'b0 ;
  assign n36388 = n36386 & n36387 ;
  assign n36381 = n5603 | n8659 ;
  assign n36382 = n9347 & n20614 ;
  assign n36383 = n9172 & n36382 ;
  assign n36384 = ( n26465 & n36381 ) | ( n26465 & n36383 ) | ( n36381 & n36383 ) ;
  assign n36385 = n36384 ^ n4702 ^ 1'b0 ;
  assign n36390 = n36389 ^ n36388 ^ n36385 ;
  assign n36391 = ~n7272 & n27391 ;
  assign n36392 = n1220 & ~n11119 ;
  assign n36393 = n36392 ^ n2732 ^ 1'b0 ;
  assign n36394 = ~n31770 & n36393 ;
  assign n36395 = n4769 & n19487 ;
  assign n36396 = n36395 ^ n31794 ^ 1'b0 ;
  assign n36397 = n2497 & n24819 ;
  assign n36398 = ~n14392 & n36397 ;
  assign n36399 = n230 & ~n8526 ;
  assign n36400 = ~n12077 & n36399 ;
  assign n36401 = ~n19775 & n30072 ;
  assign n36402 = n26082 ^ n22472 ^ n17118 ;
  assign n36403 = n4092 & n18115 ;
  assign n36404 = n36403 ^ n25723 ^ 1'b0 ;
  assign n36405 = n17046 ^ n16572 ^ 1'b0 ;
  assign n36406 = n7031 ^ n6868 ^ 1'b0 ;
  assign n36407 = ~n10265 & n12165 ;
  assign n36408 = n36407 ^ n3125 ^ 1'b0 ;
  assign n36409 = n13276 & ~n36408 ;
  assign n36410 = ( ~n1387 & n5318 ) | ( ~n1387 & n17605 ) | ( n5318 & n17605 ) ;
  assign n36411 = n283 & ~n18675 ;
  assign n36412 = ~n4387 & n36411 ;
  assign n36413 = n15832 | n36412 ;
  assign n36414 = ~n13881 & n21363 ;
  assign n36415 = ~n36413 & n36414 ;
  assign n36416 = n11928 & ~n16070 ;
  assign n36417 = n36416 ^ n19600 ^ 1'b0 ;
  assign n36420 = n1348 | n17915 ;
  assign n36418 = ( n1000 & n4683 ) | ( n1000 & ~n16545 ) | ( n4683 & ~n16545 ) ;
  assign n36419 = n36418 ^ n24183 ^ n16963 ;
  assign n36421 = n36420 ^ n36419 ^ n35491 ;
  assign n36422 = n36032 ^ n3871 ^ 1'b0 ;
  assign n36423 = ~n25837 & n36422 ;
  assign n36424 = ~n242 & n16175 ;
  assign n36425 = ( n1261 & n10118 ) | ( n1261 & n14360 ) | ( n10118 & n14360 ) ;
  assign n36426 = n27663 & n36425 ;
  assign n36427 = n551 & n36426 ;
  assign n36428 = ( ~n8755 & n30105 ) | ( ~n8755 & n36427 ) | ( n30105 & n36427 ) ;
  assign n36429 = n18457 ^ n11229 ^ 1'b0 ;
  assign n36430 = n21087 & n36429 ;
  assign n36431 = n36428 & n36430 ;
  assign n36432 = ~n6748 & n11084 ;
  assign n36433 = n4975 & n36432 ;
  assign n36434 = n2258 & ~n3690 ;
  assign n36435 = n5576 & n36434 ;
  assign n36436 = n3322 & ~n36435 ;
  assign n36437 = n36436 ^ n1004 ^ 1'b0 ;
  assign n36438 = n36437 ^ n3832 ^ 1'b0 ;
  assign n36439 = ~n36433 & n36438 ;
  assign n36441 = n14204 ^ n1891 ^ 1'b0 ;
  assign n36442 = n9899 & n36441 ;
  assign n36440 = n20940 & ~n25163 ;
  assign n36443 = n36442 ^ n36440 ^ 1'b0 ;
  assign n36444 = n7017 | n21264 ;
  assign n36445 = n25792 | n36444 ;
  assign n36446 = ( n8418 & ~n27204 ) | ( n8418 & n36445 ) | ( ~n27204 & n36445 ) ;
  assign n36447 = n4968 & n36446 ;
  assign n36448 = n28564 & n36447 ;
  assign n36450 = n3650 & n11564 ;
  assign n36449 = n4124 | n6607 ;
  assign n36451 = n36450 ^ n36449 ^ 1'b0 ;
  assign n36452 = n28079 ^ n21467 ^ 1'b0 ;
  assign n36453 = n570 | n22403 ;
  assign n36454 = n10145 & ~n36453 ;
  assign n36455 = n36454 ^ n12847 ^ 1'b0 ;
  assign n36456 = n34408 ^ n26840 ^ 1'b0 ;
  assign n36457 = n16765 & n36456 ;
  assign n36458 = n21161 ^ n11249 ^ 1'b0 ;
  assign n36459 = n33093 & n36458 ;
  assign n36460 = ~n1410 & n36459 ;
  assign n36461 = n22843 & n36460 ;
  assign n36462 = n4670 & n36461 ;
  assign n36463 = n2670 & ~n6164 ;
  assign n36464 = n36463 ^ n9388 ^ n6514 ;
  assign n36465 = n10086 & n22575 ;
  assign n36466 = n15256 ^ n13402 ^ 1'b0 ;
  assign n36467 = n4719 & n10337 ;
  assign n36468 = n28582 ^ n4417 ^ 1'b0 ;
  assign n36469 = n704 | n2075 ;
  assign n36470 = n2075 & ~n36469 ;
  assign n36471 = n298 & ~n36470 ;
  assign n36472 = ~n298 & n36471 ;
  assign n36473 = n1263 & ~n12140 ;
  assign n36474 = n36472 & n36473 ;
  assign n36475 = n10679 & ~n36474 ;
  assign n36476 = n757 & n29175 ;
  assign n36477 = n4025 & n36476 ;
  assign n36478 = x3 & ~n10411 ;
  assign n36479 = ~x3 & n36478 ;
  assign n36480 = n36477 | n36479 ;
  assign n36481 = n36477 & ~n36480 ;
  assign n36482 = n36475 & ~n36481 ;
  assign n36483 = n36482 ^ n30416 ^ 1'b0 ;
  assign n36484 = n30242 ^ n16210 ^ 1'b0 ;
  assign n36485 = n8019 & ~n36484 ;
  assign n36486 = n10008 | n13705 ;
  assign n36487 = n22495 | n22804 ;
  assign n36488 = n36487 ^ n12400 ^ 1'b0 ;
  assign n36489 = ~n10572 & n36488 ;
  assign n36490 = n36489 ^ n8268 ^ 1'b0 ;
  assign n36491 = ( n5517 & ~n10792 ) | ( n5517 & n21518 ) | ( ~n10792 & n21518 ) ;
  assign n36492 = n36490 & ~n36491 ;
  assign n36493 = n23691 ^ n5122 ^ 1'b0 ;
  assign n36494 = n5261 & n36493 ;
  assign n36495 = n28550 & n36494 ;
  assign n36496 = n36495 ^ n34601 ^ 1'b0 ;
  assign n36497 = n1880 & n6176 ;
  assign n36498 = ~n23835 & n36497 ;
  assign n36499 = n8950 | n36498 ;
  assign n36500 = n3969 | n36499 ;
  assign n36501 = n4614 ^ n3307 ^ 1'b0 ;
  assign n36502 = n5599 | n36501 ;
  assign n36503 = n36502 ^ n18438 ^ 1'b0 ;
  assign n36504 = ~n31819 & n36503 ;
  assign n36505 = n9734 & ~n36504 ;
  assign n36506 = n24573 ^ n16500 ^ n9981 ;
  assign n36507 = n3183 & ~n20344 ;
  assign n36508 = n36507 ^ n11227 ^ 1'b0 ;
  assign n36509 = n10308 & n11238 ;
  assign n36510 = n36509 ^ n34812 ^ 1'b0 ;
  assign n36511 = n10323 | n25615 ;
  assign n36512 = n2660 & n23315 ;
  assign n36513 = ~n36511 & n36512 ;
  assign n36514 = n35054 ^ n23680 ^ 1'b0 ;
  assign n36515 = n1439 & ~n36514 ;
  assign n36516 = n13111 ^ n2986 ^ 1'b0 ;
  assign n36517 = n11238 ^ n9032 ^ 1'b0 ;
  assign n36518 = n8431 | n23646 ;
  assign n36519 = n6066 | n36518 ;
  assign n36520 = n31607 & n36519 ;
  assign n36521 = n16854 ^ n13092 ^ 1'b0 ;
  assign n36522 = n21640 ^ n1087 ^ 1'b0 ;
  assign n36523 = n17207 & n36522 ;
  assign n36524 = n31292 & n33690 ;
  assign n36525 = ( n32 & n3019 ) | ( n32 & n26169 ) | ( n3019 & n26169 ) ;
  assign n36526 = n13870 | n26514 ;
  assign n36527 = ~n10340 & n36526 ;
  assign n36528 = n7689 & ~n17576 ;
  assign n36533 = n5270 & n21632 ;
  assign n36534 = ~n28478 & n36533 ;
  assign n36532 = n2579 | n9994 ;
  assign n36535 = n36534 ^ n36532 ^ 1'b0 ;
  assign n36529 = n32944 ^ n22805 ^ 1'b0 ;
  assign n36530 = ~n27664 & n36529 ;
  assign n36531 = n30576 & n36530 ;
  assign n36536 = n36535 ^ n36531 ^ 1'b0 ;
  assign n36537 = n16210 ^ n10668 ^ 1'b0 ;
  assign n36538 = n14517 | n36537 ;
  assign n36539 = ( n13045 & n24422 ) | ( n13045 & ~n36538 ) | ( n24422 & ~n36538 ) ;
  assign n36540 = n36448 ^ n17206 ^ 1'b0 ;
  assign n36541 = ~n448 & n13056 ;
  assign n36542 = n24697 | n36541 ;
  assign n36545 = ~n756 & n984 ;
  assign n36546 = n36545 ^ n31046 ^ 1'b0 ;
  assign n36543 = ~n855 & n10265 ;
  assign n36544 = n3421 | n36543 ;
  assign n36547 = n36546 ^ n36544 ^ 1'b0 ;
  assign n36548 = ~n5113 & n20526 ;
  assign n36549 = n2261 | n36548 ;
  assign n36550 = n1500 | n18548 ;
  assign n36551 = n5620 | n36550 ;
  assign n36552 = n656 & n27595 ;
  assign n36553 = ~n36551 & n36552 ;
  assign n36554 = ( n8242 & n10023 ) | ( n8242 & ~n21387 ) | ( n10023 & ~n21387 ) ;
  assign n36555 = n6583 & n17976 ;
  assign n36556 = n2745 ^ n561 ^ 1'b0 ;
  assign n36557 = n4038 & ~n25031 ;
  assign n36558 = ( n10999 & n28285 ) | ( n10999 & ~n30989 ) | ( n28285 & ~n30989 ) ;
  assign n36559 = ~n24130 & n29593 ;
  assign n36560 = ~n5134 & n19991 ;
  assign n36561 = n36560 ^ n3642 ^ 1'b0 ;
  assign n36562 = n31809 | n33788 ;
  assign n36563 = n30233 & ~n36150 ;
  assign n36564 = n707 | n9317 ;
  assign n36566 = n20484 ^ n11777 ^ n3337 ;
  assign n36565 = n12018 | n22461 ;
  assign n36567 = n36566 ^ n36565 ^ 1'b0 ;
  assign n36568 = ~n15973 & n32801 ;
  assign n36569 = n36568 ^ n2139 ^ 1'b0 ;
  assign n36571 = n4838 ^ n316 ^ 1'b0 ;
  assign n36570 = n4324 & ~n9126 ;
  assign n36572 = n36571 ^ n36570 ^ 1'b0 ;
  assign n36573 = n14752 & n16177 ;
  assign n36574 = n36573 ^ n31650 ^ n4637 ;
  assign n36575 = n2451 | n5854 ;
  assign n36576 = n13282 | n36575 ;
  assign n36577 = n36576 ^ n12808 ^ 1'b0 ;
  assign n36578 = n32711 & ~n35092 ;
  assign n36579 = ( n2230 & n7989 ) | ( n2230 & ~n9449 ) | ( n7989 & ~n9449 ) ;
  assign n36580 = n22260 | n36579 ;
  assign n36581 = n33295 | n36580 ;
  assign n36582 = n25254 & ~n33101 ;
  assign n36583 = n2667 & ~n36582 ;
  assign n36584 = n2859 | n13974 ;
  assign n36586 = n14898 | n16096 ;
  assign n36585 = ( n10980 & n26773 ) | ( n10980 & n34150 ) | ( n26773 & n34150 ) ;
  assign n36587 = n36586 ^ n36585 ^ 1'b0 ;
  assign n36588 = n36584 & ~n36587 ;
  assign n36589 = ( n23531 & n33941 ) | ( n23531 & n36588 ) | ( n33941 & n36588 ) ;
  assign n36590 = n24666 ^ n18629 ^ n17740 ;
  assign n36591 = n21202 | n22766 ;
  assign n36592 = n36591 ^ n13481 ^ 1'b0 ;
  assign n36593 = n11603 & n36592 ;
  assign n36594 = ( n9757 & n32331 ) | ( n9757 & n33043 ) | ( n32331 & n33043 ) ;
  assign n36595 = ~n6571 & n36594 ;
  assign n36596 = n17525 & n36595 ;
  assign n36597 = n19190 | n36596 ;
  assign n36598 = n27522 | n36597 ;
  assign n36599 = n20443 ^ n10872 ^ 1'b0 ;
  assign n36600 = n6227 & n36599 ;
  assign n36601 = n36600 ^ n22272 ^ 1'b0 ;
  assign n36602 = ~n29831 & n36601 ;
  assign n36603 = n7365 ^ n5997 ^ 1'b0 ;
  assign n36604 = ~n4658 & n10400 ;
  assign n36605 = n33814 | n36604 ;
  assign n36606 = n36361 & ~n36605 ;
  assign n36608 = ~n16786 & n21703 ;
  assign n36609 = n36608 ^ n8896 ^ 1'b0 ;
  assign n36607 = n17656 & ~n29560 ;
  assign n36610 = n36609 ^ n36607 ^ 1'b0 ;
  assign n36611 = n36610 ^ n16321 ^ 1'b0 ;
  assign n36612 = n20355 ^ n3039 ^ 1'b0 ;
  assign n36613 = ~n12325 & n36612 ;
  assign n36614 = n29324 ^ n22303 ^ 1'b0 ;
  assign n36615 = ~n16883 & n36614 ;
  assign n36616 = n36615 ^ n22135 ^ 1'b0 ;
  assign n36617 = n25488 & n36616 ;
  assign n36618 = n30589 ^ n27216 ^ 1'b0 ;
  assign n36619 = n12421 ^ n10532 ^ 1'b0 ;
  assign n36620 = n4565 & ~n36619 ;
  assign n36621 = n36620 ^ n2791 ^ 1'b0 ;
  assign n36622 = ~n6316 & n25590 ;
  assign n36623 = ( n25737 & n36621 ) | ( n25737 & ~n36622 ) | ( n36621 & ~n36622 ) ;
  assign n36627 = n13145 ^ n3033 ^ 1'b0 ;
  assign n36628 = n19793 & ~n36627 ;
  assign n36629 = ~n4909 & n36628 ;
  assign n36624 = ~n7473 & n23309 ;
  assign n36625 = ~n2374 & n36624 ;
  assign n36626 = n9855 & n36625 ;
  assign n36630 = n36629 ^ n36626 ^ n30350 ;
  assign n36631 = n21019 | n36378 ;
  assign n36632 = n36631 ^ n7169 ^ 1'b0 ;
  assign n36633 = n36632 ^ n35419 ^ 1'b0 ;
  assign n36634 = n650 & n5537 ;
  assign n36635 = ( n13426 & n19456 ) | ( n13426 & ~n21680 ) | ( n19456 & ~n21680 ) ;
  assign n36636 = n36359 & ~n36635 ;
  assign n36637 = n923 ^ n209 ^ 1'b0 ;
  assign n36638 = n36637 ^ n18307 ^ 1'b0 ;
  assign n36639 = n32848 & ~n36638 ;
  assign n36640 = n11540 & n26685 ;
  assign n36641 = n1956 | n4830 ;
  assign n36642 = n36641 ^ n11974 ^ 1'b0 ;
  assign n36643 = n35661 | n36642 ;
  assign n36644 = n109 & n25010 ;
  assign n36645 = ~n22869 & n36644 ;
  assign n36646 = n36645 ^ n6850 ^ 1'b0 ;
  assign n36647 = n22429 & ~n36646 ;
  assign n36648 = n36647 ^ n25760 ^ 1'b0 ;
  assign n36649 = n14388 | n26283 ;
  assign n36650 = n5652 | n11123 ;
  assign n36651 = n36650 ^ n7550 ^ 1'b0 ;
  assign n36652 = n36651 ^ n29803 ^ n14057 ;
  assign n36653 = ~n31984 & n36652 ;
  assign n36654 = n28664 ^ n15706 ^ 1'b0 ;
  assign n36655 = n24193 ^ n17133 ^ n11546 ;
  assign n36656 = n9041 & ~n36655 ;
  assign n36657 = ( ~n12088 & n24866 ) | ( ~n12088 & n36656 ) | ( n24866 & n36656 ) ;
  assign n36658 = ( n1509 & ~n3696 ) | ( n1509 & n36657 ) | ( ~n3696 & n36657 ) ;
  assign n36659 = n25353 ^ n14246 ^ 1'b0 ;
  assign n36660 = n20188 | n36659 ;
  assign n36661 = n6139 & n11295 ;
  assign n36662 = ( n63 & n12371 ) | ( n63 & n16415 ) | ( n12371 & n16415 ) ;
  assign n36663 = n36661 & n36662 ;
  assign n36664 = n23042 ^ n13533 ^ n10808 ;
  assign n36665 = n36664 ^ n4186 ^ 1'b0 ;
  assign n36666 = n13037 | n36665 ;
  assign n36667 = ( ~n6558 & n36663 ) | ( ~n6558 & n36666 ) | ( n36663 & n36666 ) ;
  assign n36668 = ~n14763 & n36667 ;
  assign n36669 = n36668 ^ n7772 ^ 1'b0 ;
  assign n36670 = n30851 ^ n25445 ^ n15274 ;
  assign n36671 = n9651 & ~n31599 ;
  assign n36672 = n36671 ^ n34143 ^ n24262 ;
  assign n36673 = n18587 & n25610 ;
  assign n36674 = n27288 ^ n7734 ^ n3698 ;
  assign n36675 = ~n3926 & n4959 ;
  assign n36676 = n36675 ^ n31024 ^ 1'b0 ;
  assign n36677 = n3847 | n20374 ;
  assign n36678 = n36677 ^ n15052 ^ 1'b0 ;
  assign n36679 = n36678 ^ n411 ^ 1'b0 ;
  assign n36680 = ~n17945 & n27419 ;
  assign n36681 = n19323 & ~n36680 ;
  assign n36682 = ( n20436 & n26253 ) | ( n20436 & ~n36681 ) | ( n26253 & ~n36681 ) ;
  assign n36684 = n11171 ^ n7672 ^ n5970 ;
  assign n36685 = n17595 ^ n1181 ^ 1'b0 ;
  assign n36686 = n36684 & n36685 ;
  assign n36683 = n22398 ^ n20053 ^ 1'b0 ;
  assign n36687 = n36686 ^ n36683 ^ n27952 ;
  assign n36688 = ( n2544 & ~n4315 ) | ( n2544 & n17134 ) | ( ~n4315 & n17134 ) ;
  assign n36689 = ~n1653 & n17371 ;
  assign n36690 = n13873 & n36689 ;
  assign n36691 = n9013 & n13176 ;
  assign n36692 = n2045 & n7949 ;
  assign n36693 = n36692 ^ n12449 ^ 1'b0 ;
  assign n36694 = n36693 ^ n25427 ^ 1'b0 ;
  assign n36695 = n36691 | n36694 ;
  assign n36696 = n36690 | n36695 ;
  assign n36697 = n1166 & ~n36696 ;
  assign n36698 = ~n8554 & n8894 ;
  assign n36699 = ~n26064 & n36698 ;
  assign n36700 = n36699 ^ n24058 ^ n8683 ;
  assign n36701 = n36700 ^ n18132 ^ 1'b0 ;
  assign n36702 = n9111 & n36701 ;
  assign n36703 = n10956 ^ n2186 ^ 1'b0 ;
  assign n36704 = ~n654 & n36703 ;
  assign n36705 = n15645 | n24124 ;
  assign n36707 = n5612 ^ n2824 ^ 1'b0 ;
  assign n36706 = n6890 & n34118 ;
  assign n36708 = n36707 ^ n36706 ^ 1'b0 ;
  assign n36709 = n8665 & n17019 ;
  assign n36710 = n29558 | n36709 ;
  assign n36711 = n9081 | n36710 ;
  assign n36712 = n4083 & ~n8907 ;
  assign n36713 = n36712 ^ n11015 ^ 1'b0 ;
  assign n36714 = n36713 ^ n5986 ^ 1'b0 ;
  assign n36715 = n1784 & ~n36714 ;
  assign n36716 = ~n13011 & n16641 ;
  assign n36717 = ~n22230 & n36716 ;
  assign n36719 = n22791 ^ n448 ^ 1'b0 ;
  assign n36720 = n15265 | n36719 ;
  assign n36718 = n4241 | n33810 ;
  assign n36721 = n36720 ^ n36718 ^ 1'b0 ;
  assign n36722 = n3351 & ~n26149 ;
  assign n36723 = n8203 | n8522 ;
  assign n36724 = n36723 ^ n29022 ^ 1'b0 ;
  assign n36725 = ( n5312 & n6690 ) | ( n5312 & ~n27767 ) | ( n6690 & ~n27767 ) ;
  assign n36726 = ~n36724 & n36725 ;
  assign n36727 = n24153 & ~n25775 ;
  assign n36728 = n1109 & n36727 ;
  assign n36729 = n15315 & n20306 ;
  assign n36730 = n36729 ^ n4438 ^ 1'b0 ;
  assign n36731 = n28456 & n36730 ;
  assign n36732 = n3443 | n9816 ;
  assign n36733 = n32114 ^ n22761 ^ 1'b0 ;
  assign n36734 = n8996 | n19536 ;
  assign n36735 = n16838 & ~n36734 ;
  assign n36736 = n12241 & n36735 ;
  assign n36737 = n33235 ^ n15800 ^ 1'b0 ;
  assign n36738 = ~n5182 & n36737 ;
  assign n36739 = n9636 & n36738 ;
  assign n36740 = n30597 | n34189 ;
  assign n36741 = n11137 | n36740 ;
  assign n36742 = n3339 & ~n18268 ;
  assign n36743 = n14974 | n36742 ;
  assign n36744 = n36743 ^ n15608 ^ 1'b0 ;
  assign n36745 = n10870 & ~n36744 ;
  assign n36746 = n36745 ^ n20879 ^ 1'b0 ;
  assign n36747 = n1733 | n36746 ;
  assign n36748 = n36741 | n36747 ;
  assign n36749 = n9000 ^ n2597 ^ 1'b0 ;
  assign n36750 = ~n1822 & n2784 ;
  assign n36751 = n36750 ^ n22834 ^ 1'b0 ;
  assign n36752 = ( n548 & n3940 ) | ( n548 & n6679 ) | ( n3940 & n6679 ) ;
  assign n36753 = n36752 ^ n18692 ^ 1'b0 ;
  assign n36754 = ( n3879 & n4977 ) | ( n3879 & ~n36753 ) | ( n4977 & ~n36753 ) ;
  assign n36755 = ~n5844 & n26849 ;
  assign n36756 = n6276 & ~n17793 ;
  assign n36757 = n36756 ^ n13406 ^ 1'b0 ;
  assign n36758 = n12369 & n36757 ;
  assign n36759 = n36758 ^ n1589 ^ 1'b0 ;
  assign n36760 = n32919 ^ n26595 ^ 1'b0 ;
  assign n36761 = n24531 ^ n9696 ^ 1'b0 ;
  assign n36762 = n11150 & ~n14431 ;
  assign n36763 = n14578 ^ n2004 ^ 1'b0 ;
  assign n36764 = n369 & n4977 ;
  assign n36765 = n18432 & n36764 ;
  assign n36766 = n19518 ^ n18641 ^ 1'b0 ;
  assign n36767 = n31244 ^ n5639 ^ 1'b0 ;
  assign n36768 = n9899 & n36767 ;
  assign n36769 = ~n17266 & n36768 ;
  assign n36770 = n1822 & ~n4468 ;
  assign n36771 = n36770 ^ n5639 ^ 1'b0 ;
  assign n36772 = n25930 & ~n36771 ;
  assign n36773 = ~n4458 & n36772 ;
  assign n36774 = n36773 ^ n23743 ^ 1'b0 ;
  assign n36775 = n3299 & ~n7096 ;
  assign n36776 = n10915 ^ n5114 ^ 1'b0 ;
  assign n36777 = n36776 ^ n9517 ^ 1'b0 ;
  assign n36778 = ( n14033 & ~n36775 ) | ( n14033 & n36777 ) | ( ~n36775 & n36777 ) ;
  assign n36779 = n4171 & n28082 ;
  assign n36780 = n36779 ^ n9776 ^ 1'b0 ;
  assign n36781 = n12797 ^ n6284 ^ 1'b0 ;
  assign n36782 = n35267 & n36781 ;
  assign n36783 = n7686 | n12051 ;
  assign n36784 = n36783 ^ n14066 ^ 1'b0 ;
  assign n36785 = n36784 ^ n15925 ^ 1'b0 ;
  assign n36786 = n23628 & n36785 ;
  assign n36787 = ~n11262 & n36786 ;
  assign n36788 = n29816 ^ n18654 ^ 1'b0 ;
  assign n36789 = n21763 ^ n4309 ^ 1'b0 ;
  assign n36790 = n3159 | n36789 ;
  assign n36791 = n27191 | n36790 ;
  assign n36792 = n2505 & ~n36791 ;
  assign n36793 = n36792 ^ n1400 ^ 1'b0 ;
  assign n36794 = ( n11371 & n32155 ) | ( n11371 & ~n32715 ) | ( n32155 & ~n32715 ) ;
  assign n36795 = n20726 ^ n17136 ^ 1'b0 ;
  assign n36796 = n8575 | n36795 ;
  assign n36797 = n4274 & ~n29847 ;
  assign n36798 = ~n21628 & n33268 ;
  assign n36799 = ( n7987 & n8768 ) | ( n7987 & ~n12705 ) | ( n8768 & ~n12705 ) ;
  assign n36801 = ( n6915 & n8057 ) | ( n6915 & ~n14164 ) | ( n8057 & ~n14164 ) ;
  assign n36800 = ~n6220 & n7193 ;
  assign n36802 = n36801 ^ n36800 ^ 1'b0 ;
  assign n36803 = n1395 | n3412 ;
  assign n36804 = n3985 | n36803 ;
  assign n36805 = n20125 & ~n34412 ;
  assign n36806 = n30989 & n36805 ;
  assign n36807 = n36039 ^ n17088 ^ 1'b0 ;
  assign n36810 = ~n250 & n9509 ;
  assign n36811 = n21893 & ~n36810 ;
  assign n36812 = ~n29476 & n36811 ;
  assign n36808 = ( n12391 & n14236 ) | ( n12391 & n24996 ) | ( n14236 & n24996 ) ;
  assign n36809 = ~n5182 & n36808 ;
  assign n36813 = n36812 ^ n36809 ^ 1'b0 ;
  assign n36815 = n15767 & n30217 ;
  assign n36814 = n3429 | n10234 ;
  assign n36816 = n36815 ^ n36814 ^ 1'b0 ;
  assign n36817 = n25094 ^ n6696 ^ 1'b0 ;
  assign n36818 = n3981 ^ n223 ^ 1'b0 ;
  assign n36819 = n5210 & ~n7033 ;
  assign n36820 = ~n36818 & n36819 ;
  assign n36821 = ( n2064 & n13667 ) | ( n2064 & n13690 ) | ( n13667 & n13690 ) ;
  assign n36824 = n14617 | n15593 ;
  assign n36822 = n17561 ^ n7512 ^ 1'b0 ;
  assign n36823 = n14305 | n36822 ;
  assign n36825 = n36824 ^ n36823 ^ 1'b0 ;
  assign n36826 = ( n5300 & ~n29448 ) | ( n5300 & n36825 ) | ( ~n29448 & n36825 ) ;
  assign n36827 = n9197 | n28506 ;
  assign n36828 = ( n8470 & n13018 ) | ( n8470 & ~n13443 ) | ( n13018 & ~n13443 ) ;
  assign n36829 = n36828 ^ n21367 ^ 1'b0 ;
  assign n36830 = n10318 ^ n2475 ^ 1'b0 ;
  assign n36831 = n36829 & n36830 ;
  assign n36832 = n10164 & ~n21027 ;
  assign n36833 = n36832 ^ n9148 ^ 1'b0 ;
  assign n36834 = n16398 | n36833 ;
  assign n36835 = ~n36088 & n36834 ;
  assign n36836 = n36835 ^ n1078 ^ 1'b0 ;
  assign n36837 = n6930 & ~n9509 ;
  assign n36838 = n650 & n36837 ;
  assign n36839 = n11071 & ~n16038 ;
  assign n36840 = n9621 & n36839 ;
  assign n36841 = n24505 ^ n23549 ^ n22988 ;
  assign n36842 = n36841 ^ n34991 ^ 1'b0 ;
  assign n36843 = n10100 & ~n34368 ;
  assign n36844 = n36843 ^ n15839 ^ 1'b0 ;
  assign n36845 = n31092 ^ n25808 ^ n864 ;
  assign n36846 = n12836 & n12946 ;
  assign n36847 = n36846 ^ n1595 ^ 1'b0 ;
  assign n36848 = n8526 & ~n36847 ;
  assign n36849 = n33267 & ~n36848 ;
  assign n36850 = n10524 ^ n3420 ^ 1'b0 ;
  assign n36851 = ~n3663 & n36850 ;
  assign n36852 = ~n1127 & n4752 ;
  assign n36853 = n24169 & n36852 ;
  assign n36854 = n25598 | n27916 ;
  assign n36855 = n36854 ^ n33290 ^ 1'b0 ;
  assign n36856 = n7646 & n8197 ;
  assign n36857 = ~n7808 & n36856 ;
  assign n36858 = n36857 ^ n16045 ^ 1'b0 ;
  assign n36859 = n29721 ^ n11135 ^ n3038 ;
  assign n36860 = n36858 | n36859 ;
  assign n36861 = n8868 & ~n36860 ;
  assign n36862 = n36861 ^ n15042 ^ 1'b0 ;
  assign n36863 = n27152 ^ n1083 ^ 1'b0 ;
  assign n36864 = ~n4847 & n36863 ;
  assign n36865 = ( n2176 & n15569 ) | ( n2176 & ~n36864 ) | ( n15569 & ~n36864 ) ;
  assign n36866 = ~n7779 & n15154 ;
  assign n36867 = n6595 & n20969 ;
  assign n36868 = ~n36866 & n36867 ;
  assign n36869 = n7267 & ~n34450 ;
  assign n36870 = n36869 ^ n23 ^ 1'b0 ;
  assign n36871 = n3879 | n11818 ;
  assign n36872 = ~n2256 & n12377 ;
  assign n36873 = n36872 ^ n4252 ^ 1'b0 ;
  assign n36874 = n1122 & n15246 ;
  assign n36875 = n36874 ^ n16372 ^ 1'b0 ;
  assign n36876 = n20352 | n36875 ;
  assign n36877 = n6509 | n36876 ;
  assign n36878 = n36873 & ~n36877 ;
  assign n36879 = n32434 ^ n12589 ^ n5311 ;
  assign n36880 = n3551 ^ n408 ^ 1'b0 ;
  assign n36881 = n35592 & ~n36880 ;
  assign n36882 = n36881 ^ n25253 ^ 1'b0 ;
  assign n36888 = n6736 ^ n1907 ^ 1'b0 ;
  assign n36889 = n7755 | n11500 ;
  assign n36890 = n36889 ^ n13703 ^ 1'b0 ;
  assign n36891 = n36888 | n36890 ;
  assign n36883 = ~n8400 & n24065 ;
  assign n36884 = n34640 & n36883 ;
  assign n36885 = n36884 ^ n19091 ^ 1'b0 ;
  assign n36886 = n20671 & ~n22408 ;
  assign n36887 = n36885 | n36886 ;
  assign n36892 = n36891 ^ n36887 ^ 1'b0 ;
  assign n36893 = ~n18090 & n27906 ;
  assign n36894 = ~n2886 & n36893 ;
  assign n36895 = n28743 | n36894 ;
  assign n36899 = ( ~n115 & n1412 ) | ( ~n115 & n7599 ) | ( n1412 & n7599 ) ;
  assign n36896 = n11037 & n33347 ;
  assign n36897 = n36896 ^ n19356 ^ 1'b0 ;
  assign n36898 = n3313 & n36897 ;
  assign n36900 = n36899 ^ n36898 ^ n35254 ;
  assign n36901 = n112 | n33328 ;
  assign n36902 = n1716 & ~n36901 ;
  assign n36903 = n702 & ~n36902 ;
  assign n36904 = n36903 ^ n22508 ^ 1'b0 ;
  assign n36905 = n1401 & n1590 ;
  assign n36906 = n316 & n36905 ;
  assign n36907 = n1827 & ~n36906 ;
  assign n36908 = ~n13089 & n36907 ;
  assign n36909 = n26603 | n36908 ;
  assign n36910 = n36909 ^ n32697 ^ 1'b0 ;
  assign n36911 = n12484 ^ n8667 ^ 1'b0 ;
  assign n36912 = n19549 & ~n36911 ;
  assign n36913 = n1781 & n6804 ;
  assign n36916 = ( ~n5242 & n9692 ) | ( ~n5242 & n17352 ) | ( n9692 & n17352 ) ;
  assign n36914 = n29551 ^ n22974 ^ 1'b0 ;
  assign n36915 = n8497 & n36914 ;
  assign n36917 = n36916 ^ n36915 ^ n3133 ;
  assign n36918 = n8701 & ~n12945 ;
  assign n36919 = n36918 ^ n13876 ^ 1'b0 ;
  assign n36920 = n16051 & ~n16766 ;
  assign n36922 = n17274 & n20949 ;
  assign n36923 = ~n16478 & n36922 ;
  assign n36921 = ~n867 & n34806 ;
  assign n36924 = n36923 ^ n36921 ^ 1'b0 ;
  assign n36925 = n7035 & n36924 ;
  assign n36926 = n15080 | n15341 ;
  assign n36927 = ( ~n11536 & n27937 ) | ( ~n11536 & n36926 ) | ( n27937 & n36926 ) ;
  assign n36929 = n28120 ^ n25320 ^ 1'b0 ;
  assign n36930 = ~n5778 & n36929 ;
  assign n36928 = ( ~n532 & n18409 ) | ( ~n532 & n34345 ) | ( n18409 & n34345 ) ;
  assign n36931 = n36930 ^ n36928 ^ n34346 ;
  assign n36932 = n16073 ^ n14750 ^ 1'b0 ;
  assign n36933 = ~n8962 & n10752 ;
  assign n36934 = n36933 ^ n35231 ^ 1'b0 ;
  assign n36935 = n20968 | n30231 ;
  assign n36936 = ~n6050 & n12548 ;
  assign n36937 = n36936 ^ n8720 ^ 1'b0 ;
  assign n36938 = n13511 | n32871 ;
  assign n36939 = ( n390 & ~n14112 ) | ( n390 & n36938 ) | ( ~n14112 & n36938 ) ;
  assign n36940 = n6457 & n11302 ;
  assign n36941 = n12713 & ~n15597 ;
  assign n36942 = n6289 ^ n2152 ^ 1'b0 ;
  assign n36943 = n30474 ^ n16223 ^ 1'b0 ;
  assign n36944 = n13283 | n36943 ;
  assign n36946 = n8380 & n21552 ;
  assign n36947 = ~n41 & n36946 ;
  assign n36945 = n1969 & n17632 ;
  assign n36948 = n36947 ^ n36945 ^ 1'b0 ;
  assign n36949 = n6704 & n9244 ;
  assign n36950 = n36949 ^ n4044 ^ 1'b0 ;
  assign n36951 = n36950 ^ n32453 ^ 1'b0 ;
  assign n36953 = ~n11466 & n22516 ;
  assign n36954 = n36953 ^ n10968 ^ 1'b0 ;
  assign n36952 = ( ~n1279 & n2217 ) | ( ~n1279 & n3285 ) | ( n2217 & n3285 ) ;
  assign n36955 = n36954 ^ n36952 ^ n28025 ;
  assign n36956 = n607 | n19816 ;
  assign n36957 = n5384 ^ n2071 ^ 1'b0 ;
  assign n36958 = ~n18626 & n36957 ;
  assign n36959 = n36958 ^ n7584 ^ 1'b0 ;
  assign n36960 = n35750 | n36959 ;
  assign n36961 = n36960 ^ n14524 ^ 1'b0 ;
  assign n36963 = n9788 & ~n15437 ;
  assign n36962 = n10238 | n11567 ;
  assign n36964 = n36963 ^ n36962 ^ 1'b0 ;
  assign n36965 = n22687 ^ n17283 ^ 1'b0 ;
  assign n36966 = n102 | n32743 ;
  assign n36967 = n14597 ^ n375 ^ n304 ;
  assign n36972 = n12668 | n27278 ;
  assign n36973 = n12586 & ~n36972 ;
  assign n36968 = ~n4549 & n18247 ;
  assign n36969 = n4549 & n36968 ;
  assign n36970 = n36969 ^ n3333 ^ 1'b0 ;
  assign n36971 = n4102 | n36970 ;
  assign n36974 = n36973 ^ n36971 ^ 1'b0 ;
  assign n36975 = n22976 | n26563 ;
  assign n36976 = n15528 & ~n36975 ;
  assign n36977 = n29895 & ~n36976 ;
  assign n36978 = n29088 ^ n8257 ^ n4344 ;
  assign n36979 = ~n37 & n31001 ;
  assign n36980 = n32245 & n36979 ;
  assign n36981 = n10446 | n12235 ;
  assign n36982 = n36981 ^ n32006 ^ 1'b0 ;
  assign n36983 = n11488 & n18247 ;
  assign n36984 = n3432 & n5716 ;
  assign n36985 = n36983 & n36984 ;
  assign n36986 = n36985 ^ n18177 ^ 1'b0 ;
  assign n36987 = ~n36982 & n36986 ;
  assign n36988 = n36987 ^ n33567 ^ 1'b0 ;
  assign n36989 = n16651 ^ n13479 ^ 1'b0 ;
  assign n36990 = ~n24616 & n36989 ;
  assign n36991 = n10040 & n25764 ;
  assign n36992 = n36991 ^ n1064 ^ 1'b0 ;
  assign n36993 = n36992 ^ n17436 ^ 1'b0 ;
  assign n36994 = ~n19482 & n32621 ;
  assign n36995 = n6902 ^ n754 ^ 1'b0 ;
  assign n36996 = n345 & ~n20619 ;
  assign n36997 = n36995 & ~n36996 ;
  assign n36998 = n4569 | n8774 ;
  assign n36999 = n1813 & n36998 ;
  assign n37000 = n22290 & n36999 ;
  assign n37001 = ( ~n6833 & n27656 ) | ( ~n6833 & n37000 ) | ( n27656 & n37000 ) ;
  assign n37002 = ~n8885 & n28843 ;
  assign n37003 = n37002 ^ n13030 ^ 1'b0 ;
  assign n37004 = n7989 ^ n5534 ^ n962 ;
  assign n37005 = n15940 & ~n37004 ;
  assign n37006 = ~n11736 & n37005 ;
  assign n37007 = n16232 & n29119 ;
  assign n37009 = ~n4761 & n23428 ;
  assign n37008 = n21429 ^ n16660 ^ 1'b0 ;
  assign n37010 = n37009 ^ n37008 ^ n11536 ;
  assign n37011 = n37010 ^ n33038 ^ n11059 ;
  assign n37012 = n2461 & n36757 ;
  assign n37013 = n33641 ^ n20662 ^ 1'b0 ;
  assign n37014 = n963 | n37013 ;
  assign n37015 = n2350 | n7997 ;
  assign n37016 = n37015 ^ n18268 ^ 1'b0 ;
  assign n37017 = n37016 ^ n11129 ^ 1'b0 ;
  assign n37018 = ( n10441 & ~n17274 ) | ( n10441 & n34563 ) | ( ~n17274 & n34563 ) ;
  assign n37019 = n21401 & ~n37018 ;
  assign n37020 = n21997 & n37019 ;
  assign n37021 = n965 ^ n135 ^ 1'b0 ;
  assign n37022 = n37021 ^ n1664 ^ 1'b0 ;
  assign n37023 = n37022 ^ n30188 ^ n965 ;
  assign n37024 = ~n21350 & n25620 ;
  assign n37025 = ( ~n8551 & n13745 ) | ( ~n8551 & n37024 ) | ( n13745 & n37024 ) ;
  assign n37026 = ~n23763 & n32094 ;
  assign n37027 = n37026 ^ n6614 ^ 1'b0 ;
  assign n37028 = n637 | n11610 ;
  assign n37029 = n37028 ^ n3393 ^ 1'b0 ;
  assign n37030 = n28733 & n37029 ;
  assign n37031 = n5189 ^ n4626 ^ 1'b0 ;
  assign n37032 = n17643 & n20588 ;
  assign n37033 = ~n1542 & n16648 ;
  assign n37034 = n14510 ^ n7438 ^ 1'b0 ;
  assign n37035 = n37033 & ~n37034 ;
  assign n37036 = n3597 | n29218 ;
  assign n37037 = n18765 | n37036 ;
  assign n37038 = n37035 & n37037 ;
  assign n37039 = n37038 ^ n3098 ^ 1'b0 ;
  assign n37040 = n37039 ^ n29465 ^ 1'b0 ;
  assign n37041 = n22726 | n37040 ;
  assign n37042 = n30726 ^ n14409 ^ 1'b0 ;
  assign n37043 = n24121 ^ n23722 ^ n19426 ;
  assign n37044 = n6392 & n26936 ;
  assign n37045 = n5700 & ~n11000 ;
  assign n37046 = n34560 & n37045 ;
  assign n37047 = n37046 ^ n4113 ^ 1'b0 ;
  assign n37048 = n26449 & ~n37047 ;
  assign n37049 = n7550 & n13784 ;
  assign n37050 = ~n21546 & n36802 ;
  assign n37051 = ~n1767 & n37050 ;
  assign n37052 = n596 & ~n10462 ;
  assign n37053 = n14614 & n37052 ;
  assign n37054 = n27906 & ~n37053 ;
  assign n37055 = n37054 ^ n31356 ^ 1'b0 ;
  assign n37056 = ~n4128 & n8389 ;
  assign n37057 = n2228 & n37056 ;
  assign n37058 = n7557 & ~n21775 ;
  assign n37059 = n13015 & ~n14587 ;
  assign n37060 = n21570 & n37059 ;
  assign n37064 = n1010 | n10829 ;
  assign n37061 = n32 & ~n3469 ;
  assign n37062 = n23156 & n37061 ;
  assign n37063 = n37062 ^ n5281 ^ 1'b0 ;
  assign n37065 = n37064 ^ n37063 ^ 1'b0 ;
  assign n37066 = n37060 | n37065 ;
  assign n37067 = n8644 ^ n1064 ^ 1'b0 ;
  assign n37068 = ~n33667 & n37067 ;
  assign n37069 = n2884 & n27595 ;
  assign n37070 = n37069 ^ n318 ^ 1'b0 ;
  assign n37074 = n5538 & ~n36880 ;
  assign n37071 = n2674 & n12111 ;
  assign n37072 = n37071 ^ n2251 ^ 1'b0 ;
  assign n37073 = n25464 | n37072 ;
  assign n37075 = n37074 ^ n37073 ^ 1'b0 ;
  assign n37076 = n24907 & ~n37075 ;
  assign n37077 = n29298 ^ n5101 ^ 1'b0 ;
  assign n37078 = n6921 ^ n3209 ^ 1'b0 ;
  assign n37079 = n37077 | n37078 ;
  assign n37080 = n18428 ^ n3597 ^ 1'b0 ;
  assign n37081 = ~n13371 & n37080 ;
  assign n37082 = ~n33250 & n37081 ;
  assign n37083 = ( ~n4235 & n14593 ) | ( ~n4235 & n26013 ) | ( n14593 & n26013 ) ;
  assign n37084 = n31989 ^ n12127 ^ n7706 ;
  assign n37085 = n17852 ^ n9814 ^ n2955 ;
  assign n37086 = ( n5874 & n12632 ) | ( n5874 & ~n22804 ) | ( n12632 & ~n22804 ) ;
  assign n37087 = n37086 ^ n22576 ^ 1'b0 ;
  assign n37088 = n19171 | n37087 ;
  assign n37089 = n11403 & n13594 ;
  assign n37090 = n8945 & n37089 ;
  assign n37091 = ~n20218 & n37090 ;
  assign n37092 = n736 | n23171 ;
  assign n37093 = n37092 ^ n19360 ^ 1'b0 ;
  assign n37094 = n5185 ^ n2569 ^ 1'b0 ;
  assign n37095 = n4620 & ~n37094 ;
  assign n37096 = ~n37093 & n37095 ;
  assign n37099 = n2338 & ~n12270 ;
  assign n37100 = n13018 & ~n37099 ;
  assign n37101 = n37100 ^ n9436 ^ 1'b0 ;
  assign n37102 = n18568 & n37101 ;
  assign n37097 = n9388 & n20306 ;
  assign n37098 = n37097 ^ n1734 ^ 1'b0 ;
  assign n37103 = n37102 ^ n37098 ^ n31171 ;
  assign n37104 = n7261 & ~n37103 ;
  assign n37105 = n37104 ^ n4796 ^ 1'b0 ;
  assign n37106 = n1006 | n6615 ;
  assign n37107 = n37106 ^ n16540 ^ 1'b0 ;
  assign n37108 = n30251 & ~n37107 ;
  assign n37109 = n19863 ^ n1623 ^ 1'b0 ;
  assign n37110 = n27979 ^ n12366 ^ n1877 ;
  assign n37111 = n37110 ^ n11782 ^ 1'b0 ;
  assign n37112 = n33328 ^ n21762 ^ 1'b0 ;
  assign n37113 = n37112 ^ n7245 ^ 1'b0 ;
  assign n37114 = ( ~n4511 & n37111 ) | ( ~n4511 & n37113 ) | ( n37111 & n37113 ) ;
  assign n37115 = ( ~n9024 & n10025 ) | ( ~n9024 & n37114 ) | ( n10025 & n37114 ) ;
  assign n37116 = n2194 | n31177 ;
  assign n37117 = n9146 ^ n3991 ^ 1'b0 ;
  assign n37118 = n11806 & n23311 ;
  assign n37119 = n37118 ^ n3016 ^ 1'b0 ;
  assign n37120 = n12988 ^ n6032 ^ 1'b0 ;
  assign n37121 = n26434 ^ n5353 ^ n70 ;
  assign n37122 = n25760 ^ n10374 ^ 1'b0 ;
  assign n37123 = ( n8329 & ~n25419 ) | ( n8329 & n37122 ) | ( ~n25419 & n37122 ) ;
  assign n37126 = n35633 ^ n1096 ^ n41 ;
  assign n37124 = ( n14864 & ~n26204 ) | ( n14864 & n27982 ) | ( ~n26204 & n27982 ) ;
  assign n37125 = n16965 & n37124 ;
  assign n37127 = n37126 ^ n37125 ^ 1'b0 ;
  assign n37128 = n11934 ^ n8424 ^ 1'b0 ;
  assign n37129 = n3988 ^ n3312 ^ 1'b0 ;
  assign n37130 = n37129 ^ n6336 ^ n3571 ;
  assign n37131 = ~n37128 & n37130 ;
  assign n37132 = n37131 ^ n12260 ^ 1'b0 ;
  assign n37133 = ~n28751 & n37132 ;
  assign n37134 = n37133 ^ n32040 ^ 1'b0 ;
  assign n37135 = n26217 ^ n20781 ^ 1'b0 ;
  assign n37136 = ~n27974 & n37135 ;
  assign n37137 = ~n7805 & n16110 ;
  assign n37138 = n10277 & ~n37137 ;
  assign n37140 = n6097 & n21861 ;
  assign n37141 = ~n8950 & n37140 ;
  assign n37139 = n30776 ^ n29635 ^ 1'b0 ;
  assign n37142 = n37141 ^ n37139 ^ 1'b0 ;
  assign n37143 = n5394 & ~n24661 ;
  assign n37144 = n37143 ^ n26224 ^ 1'b0 ;
  assign n37145 = ~n14953 & n27178 ;
  assign n37146 = n37145 ^ n14485 ^ 1'b0 ;
  assign n37147 = n37146 ^ n18709 ^ 1'b0 ;
  assign n37148 = n15189 ^ n6762 ^ 1'b0 ;
  assign n37149 = ( n17788 & n23113 ) | ( n17788 & ~n25704 ) | ( n23113 & ~n25704 ) ;
  assign n37150 = n18521 & n37149 ;
  assign n37151 = ~n9905 & n31259 ;
  assign n37152 = n37151 ^ n9020 ^ 1'b0 ;
  assign n37153 = n7594 & n37152 ;
  assign n37154 = n37150 & n37153 ;
  assign n37155 = n15838 ^ n6595 ^ 1'b0 ;
  assign n37156 = ~n12460 & n37155 ;
  assign n37157 = ~n16703 & n37156 ;
  assign n37158 = n18573 ^ n3125 ^ 1'b0 ;
  assign n37159 = n13574 & ~n37158 ;
  assign n37160 = n24547 & n37159 ;
  assign n37161 = n338 & ~n3122 ;
  assign n37162 = ~n126 & n37161 ;
  assign n37163 = n8445 & n37162 ;
  assign n37164 = n36266 ^ n27846 ^ 1'b0 ;
  assign n37165 = n17432 | n37164 ;
  assign n37166 = n37163 & ~n37165 ;
  assign n37167 = n33043 ^ n20607 ^ 1'b0 ;
  assign n37168 = n7907 & n37167 ;
  assign n37169 = n7147 & n32331 ;
  assign n37170 = n37169 ^ n16096 ^ 1'b0 ;
  assign n37171 = ( n5616 & n37168 ) | ( n5616 & n37170 ) | ( n37168 & n37170 ) ;
  assign n37172 = ( n1697 & n9240 ) | ( n1697 & n21853 ) | ( n9240 & n21853 ) ;
  assign n37173 = n15347 & ~n25564 ;
  assign n37174 = n16007 ^ n14952 ^ 1'b0 ;
  assign n37175 = n37173 & ~n37174 ;
  assign n37176 = ~n24300 & n37175 ;
  assign n37177 = n37172 & n37176 ;
  assign n37178 = x0 & n236 ;
  assign n37184 = n1171 | n2239 ;
  assign n37185 = n22597 | n37184 ;
  assign n37179 = n5582 & ~n30664 ;
  assign n37180 = n14493 & n37179 ;
  assign n37181 = ~n23902 & n33679 ;
  assign n37182 = n37181 ^ n10631 ^ 1'b0 ;
  assign n37183 = n37180 | n37182 ;
  assign n37186 = n37185 ^ n37183 ^ 1'b0 ;
  assign n37187 = n11147 ^ n666 ^ 1'b0 ;
  assign n37188 = ~n6060 & n16082 ;
  assign n37189 = n37188 ^ n21904 ^ 1'b0 ;
  assign n37190 = n803 & ~n14707 ;
  assign n37191 = n37189 & n37190 ;
  assign n37192 = n37191 ^ n1397 ^ 1'b0 ;
  assign n37193 = n30182 ^ n22381 ^ n6771 ;
  assign n37194 = n37193 ^ n16331 ^ n11753 ;
  assign n37195 = n29847 ^ n25620 ^ 1'b0 ;
  assign n37196 = n17762 ^ n15739 ^ n953 ;
  assign n37197 = n28202 ^ n6927 ^ 1'b0 ;
  assign n37198 = n37196 & ~n37197 ;
  assign n37199 = n30122 ^ n13426 ^ 1'b0 ;
  assign n37200 = ~n32058 & n37199 ;
  assign n37201 = n6914 & n27647 ;
  assign n37202 = ~n13823 & n37201 ;
  assign n37203 = n37202 ^ n5142 ^ 1'b0 ;
  assign n37204 = ~n17621 & n32442 ;
  assign n37205 = n32686 | n37204 ;
  assign n37206 = n19714 ^ n3856 ^ 1'b0 ;
  assign n37207 = n19255 & ~n28019 ;
  assign n37208 = ~n11276 & n17870 ;
  assign n37209 = n28197 | n37208 ;
  assign n37210 = n32287 ^ n14076 ^ 1'b0 ;
  assign n37211 = n8766 & n37210 ;
  assign n37212 = ( x5 & n1457 ) | ( x5 & ~n8586 ) | ( n1457 & ~n8586 ) ;
  assign n37213 = n26859 ^ n11244 ^ 1'b0 ;
  assign n37214 = n37212 & ~n37213 ;
  assign n37215 = ( n17472 & n27341 ) | ( n17472 & ~n37214 ) | ( n27341 & ~n37214 ) ;
  assign n37216 = ~n15449 & n27673 ;
  assign n37217 = n37216 ^ n28857 ^ 1'b0 ;
  assign n37218 = ~n7925 & n37217 ;
  assign n37219 = n12355 | n16008 ;
  assign n37220 = n14452 & n33648 ;
  assign n37224 = ( n816 & n7165 ) | ( n816 & n8624 ) | ( n7165 & n8624 ) ;
  assign n37221 = ~n252 & n3957 ;
  assign n37222 = n252 & n37221 ;
  assign n37223 = n24356 | n37222 ;
  assign n37225 = n37224 ^ n37223 ^ 1'b0 ;
  assign n37226 = n21886 ^ n4422 ^ 1'b0 ;
  assign n37227 = n5612 & ~n13094 ;
  assign n37228 = n32127 & n37227 ;
  assign n37229 = n6453 | n19323 ;
  assign n37230 = n10402 | n14482 ;
  assign n37231 = n14371 ^ n11673 ^ 1'b0 ;
  assign n37232 = n24092 & n37231 ;
  assign n37233 = n3540 | n35974 ;
  assign n37234 = n37233 ^ n3491 ^ 1'b0 ;
  assign n37235 = n13785 | n37234 ;
  assign n37236 = n37235 ^ n13046 ^ 1'b0 ;
  assign n37237 = ~n15476 & n37236 ;
  assign n37238 = n37237 ^ n28184 ^ 1'b0 ;
  assign n37239 = n221 | n37238 ;
  assign n37240 = ~n27974 & n37239 ;
  assign n37241 = n30226 & ~n31608 ;
  assign n37242 = n8775 & ~n18104 ;
  assign n37243 = ~n4440 & n37242 ;
  assign n37244 = n35285 & ~n37243 ;
  assign n37245 = n29387 ^ n28831 ^ n2987 ;
  assign n37246 = n5727 | n8414 ;
  assign n37247 = n22562 ^ n14926 ^ 1'b0 ;
  assign n37248 = n6475 ^ n3362 ^ 1'b0 ;
  assign n37249 = n30846 & n37248 ;
  assign n37250 = ~n31415 & n37249 ;
  assign n37251 = n37250 ^ n4628 ^ 1'b0 ;
  assign n37252 = ~n19681 & n31613 ;
  assign n37253 = n31257 & ~n37252 ;
  assign n37254 = n37251 & n37253 ;
  assign n37255 = ~n28171 & n33685 ;
  assign n37256 = n37255 ^ n13107 ^ 1'b0 ;
  assign n37257 = n925 & ~n9986 ;
  assign n37258 = n37257 ^ n18155 ^ 1'b0 ;
  assign n37259 = n15077 & ~n18107 ;
  assign n37260 = n37258 & n37259 ;
  assign n37261 = ~n14694 & n34558 ;
  assign n37262 = n21570 ^ n9887 ^ 1'b0 ;
  assign n37263 = n734 & ~n37262 ;
  assign n37264 = n342 & n37263 ;
  assign n37265 = n14316 | n23662 ;
  assign n37266 = n37265 ^ n20835 ^ 1'b0 ;
  assign n37267 = n22107 & ~n37266 ;
  assign n37268 = n37267 ^ n1680 ^ 1'b0 ;
  assign n37269 = n28177 ^ n18215 ^ n9358 ;
  assign n37270 = n7958 ^ n2514 ^ 1'b0 ;
  assign n37271 = ( n12443 & n13700 ) | ( n12443 & ~n37270 ) | ( n13700 & ~n37270 ) ;
  assign n37272 = n26 & n1155 ;
  assign n37273 = ~n10551 & n37272 ;
  assign n37274 = ( n8345 & n23035 ) | ( n8345 & ~n37273 ) | ( n23035 & ~n37273 ) ;
  assign n37275 = n9059 & ~n37274 ;
  assign n37276 = n37275 ^ n6590 ^ 1'b0 ;
  assign n37277 = n4914 | n8885 ;
  assign n37281 = n13077 & n16625 ;
  assign n37282 = n37281 ^ n24093 ^ 1'b0 ;
  assign n37278 = n5902 & n7810 ;
  assign n37279 = n8886 & ~n37278 ;
  assign n37280 = n717 & n37279 ;
  assign n37283 = n37282 ^ n37280 ^ 1'b0 ;
  assign n37284 = n1054 & ~n30756 ;
  assign n37285 = n16796 ^ n9206 ^ 1'b0 ;
  assign n37286 = n37285 ^ n3222 ^ 1'b0 ;
  assign n37287 = n16126 ^ n6230 ^ 1'b0 ;
  assign n37288 = ~n14974 & n37287 ;
  assign n37289 = n12411 | n32070 ;
  assign n37290 = n37289 ^ n34563 ^ 1'b0 ;
  assign n37291 = n11965 | n16089 ;
  assign n37292 = n37291 ^ n10520 ^ 1'b0 ;
  assign n37293 = n24615 ^ n14748 ^ 1'b0 ;
  assign n37294 = n37292 | n37293 ;
  assign n37295 = n33096 ^ n20272 ^ 1'b0 ;
  assign n37296 = ~n11657 & n37295 ;
  assign n37297 = n28028 ^ n24022 ^ 1'b0 ;
  assign n37298 = n20764 ^ n15059 ^ 1'b0 ;
  assign n37299 = n9858 & n37298 ;
  assign n37300 = ( n4127 & n26815 ) | ( n4127 & n35451 ) | ( n26815 & n35451 ) ;
  assign n37301 = n8428 ^ n398 ^ 1'b0 ;
  assign n37302 = n37301 ^ n16329 ^ 1'b0 ;
  assign n37303 = n12921 ^ n2943 ^ 1'b0 ;
  assign n37304 = n13958 & n37303 ;
  assign n37305 = n10563 & ~n22461 ;
  assign n37306 = n37305 ^ n25539 ^ 1'b0 ;
  assign n37307 = ~n10929 & n13157 ;
  assign n37308 = n37307 ^ n1549 ^ 1'b0 ;
  assign n37309 = n2790 & ~n37234 ;
  assign n37310 = n3443 | n19987 ;
  assign n37311 = n870 | n37310 ;
  assign n37312 = n27975 ^ n14246 ^ n12604 ;
  assign n37313 = n37311 & n37312 ;
  assign n37314 = n37309 & n37313 ;
  assign n37315 = n37314 ^ n13286 ^ 1'b0 ;
  assign n37316 = n34273 ^ n5147 ^ 1'b0 ;
  assign n37317 = ~n4500 & n5264 ;
  assign n37318 = n17233 & n37317 ;
  assign n37319 = n8527 | n37318 ;
  assign n37320 = ~n18758 & n21204 ;
  assign n37321 = ~n15839 & n37320 ;
  assign n37322 = n37321 ^ n20255 ^ 1'b0 ;
  assign n37323 = ~n3918 & n35097 ;
  assign n37324 = ~n5654 & n11956 ;
  assign n37325 = n28872 & n37324 ;
  assign n37326 = ( n22514 & n24475 ) | ( n22514 & ~n37325 ) | ( n24475 & ~n37325 ) ;
  assign n37327 = ~n2687 & n2980 ;
  assign n37328 = n37327 ^ n12391 ^ 1'b0 ;
  assign n37329 = n18829 & ~n37328 ;
  assign n37330 = n37329 ^ n16722 ^ 1'b0 ;
  assign n37331 = n12927 | n16839 ;
  assign n37332 = n7115 & ~n37331 ;
  assign n37333 = n37332 ^ n34516 ^ 1'b0 ;
  assign n37334 = n3387 | n37333 ;
  assign n37335 = ( n1616 & ~n5724 ) | ( n1616 & n15414 ) | ( ~n5724 & n15414 ) ;
  assign n37336 = n37335 ^ n5502 ^ 1'b0 ;
  assign n37337 = n19443 & ~n30160 ;
  assign n37338 = n1848 | n10952 ;
  assign n37339 = n37338 ^ n9596 ^ 1'b0 ;
  assign n37340 = n8435 ^ n3158 ^ 1'b0 ;
  assign n37341 = n360 & ~n37340 ;
  assign n37342 = n37341 ^ x6 ^ 1'b0 ;
  assign n37343 = ~n9509 & n37342 ;
  assign n37344 = ~n37339 & n37343 ;
  assign n37345 = n33585 ^ n5361 ^ 1'b0 ;
  assign n37346 = n3918 & ~n37345 ;
  assign n37347 = n3898 & ~n13689 ;
  assign n37348 = ~n21183 & n37347 ;
  assign n37349 = n13608 | n37348 ;
  assign n37350 = n17543 | n37349 ;
  assign n37351 = n37350 ^ n1110 ^ 1'b0 ;
  assign n37352 = n448 & ~n37351 ;
  assign n37353 = n10229 & n37352 ;
  assign n37354 = n25627 ^ n10806 ^ 1'b0 ;
  assign n37355 = n13975 | n37354 ;
  assign n37356 = n5396 & ~n37355 ;
  assign n37357 = n16531 ^ n14718 ^ 1'b0 ;
  assign n37358 = n6524 & n8203 ;
  assign n37359 = n37358 ^ n29335 ^ 1'b0 ;
  assign n37360 = n5493 & n37359 ;
  assign n37361 = n3146 & n17946 ;
  assign n37362 = ~n37360 & n37361 ;
  assign n37363 = n10998 & ~n29900 ;
  assign n37364 = n31616 ^ n7903 ^ 1'b0 ;
  assign n37365 = n6925 & n10054 ;
  assign n37366 = n1912 & n37365 ;
  assign n37367 = n8414 & n14045 ;
  assign n37368 = n37367 ^ n11876 ^ 1'b0 ;
  assign n37369 = n37368 ^ n24463 ^ 1'b0 ;
  assign n37370 = n15289 & ~n37369 ;
  assign n37371 = n1549 & n37370 ;
  assign n37372 = n37371 ^ n13315 ^ 1'b0 ;
  assign n37373 = ( ~n28077 & n37366 ) | ( ~n28077 & n37372 ) | ( n37366 & n37372 ) ;
  assign n37374 = n22314 ^ n19895 ^ 1'b0 ;
  assign n37375 = n9837 | n23610 ;
  assign n37376 = n37374 & ~n37375 ;
  assign n37377 = n2041 & ~n10597 ;
  assign n37378 = ~n36268 & n37377 ;
  assign n37379 = n6379 & n29208 ;
  assign n37380 = ~n16771 & n24300 ;
  assign n37381 = n37380 ^ n5831 ^ 1'b0 ;
  assign n37382 = n30239 ^ n21134 ^ 1'b0 ;
  assign n37383 = n17991 & ~n24072 ;
  assign n37384 = n37383 ^ n19898 ^ 1'b0 ;
  assign n37385 = n1247 | n37384 ;
  assign n37386 = x10 & ~n18699 ;
  assign n37387 = n3564 & n6703 ;
  assign n37388 = n37387 ^ n34143 ^ n8414 ;
  assign n37389 = n21171 | n25726 ;
  assign n37390 = n37388 | n37389 ;
  assign n37391 = n31157 ^ n17030 ^ 1'b0 ;
  assign n37392 = n10656 & n37391 ;
  assign n37393 = n5418 ^ n637 ^ n41 ;
  assign n37394 = n11704 & n12787 ;
  assign n37395 = n7067 & n37394 ;
  assign n37396 = n22176 | n37395 ;
  assign n37397 = n37393 & ~n37396 ;
  assign n37399 = n17258 & n32703 ;
  assign n37398 = n13745 ^ n10295 ^ 1'b0 ;
  assign n37400 = n37399 ^ n37398 ^ 1'b0 ;
  assign n37402 = n4406 | n33128 ;
  assign n37403 = n37402 ^ n2542 ^ 1'b0 ;
  assign n37401 = n35010 & ~n35834 ;
  assign n37404 = n37403 ^ n37401 ^ 1'b0 ;
  assign n37405 = ~n9928 & n20030 ;
  assign n37406 = ~n37404 & n37405 ;
  assign n37407 = n5692 & n9613 ;
  assign n37408 = ~n15142 & n37407 ;
  assign n37409 = n32115 & ~n37408 ;
  assign n37410 = n35355 & n37409 ;
  assign n37411 = n22918 ^ n17895 ^ 1'b0 ;
  assign n37412 = ~n37323 & n37411 ;
  assign n37413 = ( n8978 & ~n19645 ) | ( n8978 & n23113 ) | ( ~n19645 & n23113 ) ;
  assign n37414 = n21482 ^ n9716 ^ 1'b0 ;
  assign n37415 = n4877 & ~n6099 ;
  assign n37416 = n37415 ^ n4173 ^ 1'b0 ;
  assign n37417 = n10414 & ~n37416 ;
  assign n37418 = n11988 | n13778 ;
  assign n37419 = n5878 & n32882 ;
  assign n37420 = ~n5354 & n37419 ;
  assign n37421 = n19865 ^ n9246 ^ 1'b0 ;
  assign n37422 = n6322 & ~n37421 ;
  assign n37423 = n9923 & n22815 ;
  assign n37424 = n37423 ^ n29185 ^ n14131 ;
  assign n37425 = n24640 ^ n23238 ^ n16756 ;
  assign n37426 = n18401 & n36669 ;
  assign n37427 = n37395 ^ n353 ^ 1'b0 ;
  assign n37428 = n26367 ^ n21660 ^ 1'b0 ;
  assign n37429 = n32801 & n37428 ;
  assign n37430 = n15871 ^ n7785 ^ 1'b0 ;
  assign n37431 = n24335 & n37430 ;
  assign n37432 = n37431 ^ n34929 ^ 1'b0 ;
  assign n37434 = ( n3580 & n8800 ) | ( n3580 & n19575 ) | ( n8800 & n19575 ) ;
  assign n37435 = n3698 | n37434 ;
  assign n37436 = n18488 & ~n37435 ;
  assign n37433 = n993 & ~n1046 ;
  assign n37437 = n37436 ^ n37433 ^ 1'b0 ;
  assign n37438 = n3994 & n18611 ;
  assign n37439 = n37438 ^ n37368 ^ 1'b0 ;
  assign n37440 = n1178 & n5738 ;
  assign n37441 = n37440 ^ n31769 ^ 1'b0 ;
  assign n37442 = n10827 ^ n4443 ^ 1'b0 ;
  assign n37443 = ~n10348 & n37442 ;
  assign n37444 = n37443 ^ n10492 ^ 1'b0 ;
  assign n37445 = ( n525 & n1423 ) | ( n525 & ~n2555 ) | ( n1423 & ~n2555 ) ;
  assign n37446 = n16510 ^ n2344 ^ 1'b0 ;
  assign n37447 = ~n37445 & n37446 ;
  assign n37448 = n11426 | n18052 ;
  assign n37449 = n36039 ^ n261 ^ 1'b0 ;
  assign n37450 = n14020 | n37449 ;
  assign n37451 = n31232 & n37450 ;
  assign n37453 = n2969 & ~n19871 ;
  assign n37454 = n37453 ^ n10865 ^ 1'b0 ;
  assign n37452 = n6874 & n34131 ;
  assign n37455 = n37454 ^ n37452 ^ n35952 ;
  assign n37456 = n17034 ^ n13021 ^ 1'b0 ;
  assign n37457 = n7996 & ~n15560 ;
  assign n37458 = n18758 & n37457 ;
  assign n37459 = n27572 ^ n13752 ^ n9907 ;
  assign n37460 = ~n37458 & n37459 ;
  assign n37461 = n31984 ^ n7943 ^ 1'b0 ;
  assign n37462 = n15249 ^ n13282 ^ n3528 ;
  assign n37463 = n3364 & ~n37462 ;
  assign n37464 = n18542 & ~n27925 ;
  assign n37465 = n37464 ^ n20334 ^ 1'b0 ;
  assign n37466 = ~n25171 & n25187 ;
  assign n37467 = n5831 | n37466 ;
  assign n37468 = n3609 | n37467 ;
  assign n37469 = n9362 ^ n1938 ^ 1'b0 ;
  assign n37470 = n2864 & ~n31615 ;
  assign n37471 = n34544 ^ n14772 ^ 1'b0 ;
  assign n37472 = n37471 ^ n8490 ^ 1'b0 ;
  assign n37473 = n16741 ^ n5311 ^ 1'b0 ;
  assign n37474 = n5353 | n21218 ;
  assign n37475 = n12490 & ~n37474 ;
  assign n37476 = n514 & n19539 ;
  assign n37477 = n28898 | n31694 ;
  assign n37478 = n33461 ^ n3127 ^ 1'b0 ;
  assign n37479 = n16304 & n27583 ;
  assign n37480 = n37479 ^ n10422 ^ 1'b0 ;
  assign n37481 = n28564 ^ n4899 ^ 1'b0 ;
  assign n37482 = ~n29138 & n37481 ;
  assign n37483 = n12310 & ~n16099 ;
  assign n37484 = ~n14273 & n21063 ;
  assign n37485 = n7694 & n37484 ;
  assign n37486 = n37483 | n37485 ;
  assign n37487 = n37486 ^ n31882 ^ 1'b0 ;
  assign n37488 = n9586 | n35349 ;
  assign n37489 = n32231 ^ n28699 ^ 1'b0 ;
  assign n37490 = n16205 & ~n25421 ;
  assign n37494 = n5990 & n13147 ;
  assign n37495 = n37494 ^ n22227 ^ 1'b0 ;
  assign n37496 = n13542 & n37495 ;
  assign n37497 = n37496 ^ n28988 ^ 1'b0 ;
  assign n37491 = ( n6978 & n13706 ) | ( n6978 & n19602 ) | ( n13706 & n19602 ) ;
  assign n37492 = n37491 ^ n8271 ^ 1'b0 ;
  assign n37493 = ~n13905 & n37492 ;
  assign n37498 = n37497 ^ n37493 ^ 1'b0 ;
  assign n37499 = n31073 ^ n31006 ^ 1'b0 ;
  assign n37500 = n774 & n37499 ;
  assign n37501 = n2335 & n6848 ;
  assign n37502 = ~n5350 & n37501 ;
  assign n37503 = n30419 ^ n17468 ^ 1'b0 ;
  assign n37504 = n37503 ^ n2447 ^ 1'b0 ;
  assign n37505 = ( n35313 & n37502 ) | ( n35313 & ~n37504 ) | ( n37502 & ~n37504 ) ;
  assign n37506 = n10528 & ~n16055 ;
  assign n37507 = n29490 & ~n32490 ;
  assign n37510 = ~n2084 & n8037 ;
  assign n37511 = n37510 ^ n11872 ^ 1'b0 ;
  assign n37508 = n10767 & n27064 ;
  assign n37509 = n6576 | n37508 ;
  assign n37512 = n37511 ^ n37509 ^ n3408 ;
  assign n37513 = n15177 & ~n37512 ;
  assign n37514 = n8745 & ~n32969 ;
  assign n37515 = n4066 & n37514 ;
  assign n37516 = n15926 & ~n28090 ;
  assign n37517 = n37516 ^ n7216 ^ 1'b0 ;
  assign n37518 = n12606 & n36995 ;
  assign n37519 = n17380 ^ n15651 ^ 1'b0 ;
  assign n37520 = ( n11861 & n12512 ) | ( n11861 & n37519 ) | ( n12512 & n37519 ) ;
  assign n37521 = n10899 ^ n10788 ^ 1'b0 ;
  assign n37522 = ( n7544 & n37520 ) | ( n7544 & n37521 ) | ( n37520 & n37521 ) ;
  assign n37523 = ( n20733 & n22151 ) | ( n20733 & ~n26940 ) | ( n22151 & ~n26940 ) ;
  assign n37524 = n37523 ^ n19320 ^ 1'b0 ;
  assign n37525 = n4520 & ~n37524 ;
  assign n37526 = n19041 ^ n13629 ^ 1'b0 ;
  assign n37527 = n3009 & ~n37526 ;
  assign n37528 = n778 & n8682 ;
  assign n37529 = n37528 ^ n32630 ^ n25604 ;
  assign n37530 = n37527 & n37529 ;
  assign n37531 = n4710 & n35380 ;
  assign n37532 = n15896 & n37531 ;
  assign n37533 = ~n2097 & n37532 ;
  assign n37534 = n30515 ^ n19461 ^ 1'b0 ;
  assign n37535 = n37534 ^ n16622 ^ n13670 ;
  assign n37537 = ~n2805 & n6299 ;
  assign n37538 = ~n10479 & n37537 ;
  assign n37536 = n8840 | n10648 ;
  assign n37539 = n37538 ^ n37536 ^ 1'b0 ;
  assign n37540 = n3761 ^ n427 ^ 1'b0 ;
  assign n37541 = n37540 ^ n6458 ^ n2418 ;
  assign n37542 = n13013 | n37541 ;
  assign n37543 = n6929 | n28841 ;
  assign n37544 = n32294 & n36973 ;
  assign n37545 = n37544 ^ n19833 ^ 1'b0 ;
  assign n37546 = n2910 | n9078 ;
  assign n37547 = n13396 | n37546 ;
  assign n37548 = n37547 ^ n27269 ^ 1'b0 ;
  assign n37549 = n22593 | n37548 ;
  assign n37550 = n4021 ^ n3308 ^ 1'b0 ;
  assign n37551 = n2596 & ~n14137 ;
  assign n37552 = n30514 & n37551 ;
  assign n37553 = n7096 ^ n5485 ^ 1'b0 ;
  assign n37554 = n19106 & n37553 ;
  assign n37555 = n18638 | n37554 ;
  assign n37556 = n864 | n32989 ;
  assign n37557 = n37556 ^ n2097 ^ 1'b0 ;
  assign n37558 = n6727 | n37557 ;
  assign n37559 = n8975 ^ n4434 ^ 1'b0 ;
  assign n37560 = n31815 | n37559 ;
  assign n37561 = n37560 ^ n5374 ^ 1'b0 ;
  assign n37562 = n12574 & ~n13314 ;
  assign n37563 = n27392 & n30760 ;
  assign n37564 = n37562 & n37563 ;
  assign n37565 = n33677 ^ n10046 ^ n10016 ;
  assign n37566 = n25421 & n37565 ;
  assign n37567 = n960 & ~n6524 ;
  assign n37568 = n37567 ^ n36569 ^ 1'b0 ;
  assign n37569 = ( n9154 & ~n12204 ) | ( n9154 & n14115 ) | ( ~n12204 & n14115 ) ;
  assign n37570 = n2514 ^ n1249 ^ 1'b0 ;
  assign n37571 = n21904 & n37570 ;
  assign n37572 = n2917 | n9072 ;
  assign n37573 = ( ~n16108 & n37571 ) | ( ~n16108 & n37572 ) | ( n37571 & n37572 ) ;
  assign n37574 = n24869 ^ n20417 ^ 1'b0 ;
  assign n37575 = n31720 ^ n23674 ^ n20674 ;
  assign n37576 = n18015 | n37575 ;
  assign n37577 = n26440 | n37576 ;
  assign n37578 = n37577 ^ n34846 ^ 1'b0 ;
  assign n37579 = ~n7818 & n37578 ;
  assign n37580 = n1427 & n6188 ;
  assign n37581 = n18164 ^ n11366 ^ n7596 ;
  assign n37582 = ( n15909 & n37507 ) | ( n15909 & ~n37581 ) | ( n37507 & ~n37581 ) ;
  assign n37583 = ( n2020 & ~n18325 ) | ( n2020 & n23744 ) | ( ~n18325 & n23744 ) ;
  assign n37584 = n14646 ^ n4269 ^ 1'b0 ;
  assign n37585 = n25349 ^ n22985 ^ 1'b0 ;
  assign n37586 = n3730 | n37585 ;
  assign n37587 = ~n1849 & n10579 ;
  assign n37588 = n27066 & n37587 ;
  assign n37589 = n11045 & ~n37588 ;
  assign n37590 = n5891 ^ n1658 ^ 1'b0 ;
  assign n37591 = n37589 & n37590 ;
  assign n37592 = n3988 & n37591 ;
  assign n37593 = n6622 | n36420 ;
  assign n37594 = n37592 & ~n37593 ;
  assign n37595 = n6603 ^ n2389 ^ 1'b0 ;
  assign n37596 = n24194 & ~n37595 ;
  assign n37597 = n37596 ^ n11458 ^ 1'b0 ;
  assign n37598 = n6317 & n19041 ;
  assign n37599 = n18969 & n37598 ;
  assign n37600 = n2135 & ~n11048 ;
  assign n37601 = n37600 ^ n25239 ^ 1'b0 ;
  assign n37602 = n614 & ~n37601 ;
  assign n37603 = ~n25960 & n37602 ;
  assign n37605 = n17838 | n32742 ;
  assign n37604 = n7243 & ~n29109 ;
  assign n37606 = n37605 ^ n37604 ^ 1'b0 ;
  assign n37607 = n7043 ^ n4813 ^ 1'b0 ;
  assign n37608 = n5944 & ~n6016 ;
  assign n37609 = ~n37607 & n37608 ;
  assign n37610 = n18657 ^ n10795 ^ 1'b0 ;
  assign n37611 = n25919 | n37610 ;
  assign n37612 = n30276 | n37611 ;
  assign n37613 = n1050 | n7761 ;
  assign n37614 = n27673 & ~n37613 ;
  assign n37615 = n8683 & ~n24071 ;
  assign n37616 = n37615 ^ n20498 ^ 1'b0 ;
  assign n37617 = n37616 ^ n20246 ^ 1'b0 ;
  assign n37618 = n35841 & ~n37617 ;
  assign n37619 = ~n11345 & n26446 ;
  assign n37620 = n8842 ^ n2918 ^ 1'b0 ;
  assign n37621 = n6381 & ~n28148 ;
  assign n37622 = ~n21550 & n37621 ;
  assign n37623 = n37622 ^ n28054 ^ 1'b0 ;
  assign n37624 = ~n8547 & n37623 ;
  assign n37625 = ( n386 & n1378 ) | ( n386 & n4207 ) | ( n1378 & n4207 ) ;
  assign n37626 = n37625 ^ n14401 ^ 1'b0 ;
  assign n37627 = n37626 ^ n25811 ^ n2005 ;
  assign n37628 = n16321 ^ n4183 ^ 1'b0 ;
  assign n37629 = n203 & ~n12311 ;
  assign n37630 = n12755 | n37629 ;
  assign n37631 = n37630 ^ n13726 ^ 1'b0 ;
  assign n37632 = n27607 ^ n21736 ^ 1'b0 ;
  assign n37633 = ( ~n8226 & n27566 ) | ( ~n8226 & n37632 ) | ( n27566 & n37632 ) ;
  assign n37634 = ( n16794 & n22319 ) | ( n16794 & n37633 ) | ( n22319 & n37633 ) ;
  assign n37635 = ~n12241 & n18204 ;
  assign n37636 = n14750 | n15811 ;
  assign n37637 = n37635 | n37636 ;
  assign n37638 = ( n3076 & n9753 ) | ( n3076 & ~n27915 ) | ( n9753 & ~n27915 ) ;
  assign n37639 = n1962 | n22724 ;
  assign n37640 = n37639 ^ n9785 ^ 1'b0 ;
  assign n37641 = ~n37638 & n37640 ;
  assign n37642 = n26408 ^ n15441 ^ 1'b0 ;
  assign n37643 = n17240 & ~n27511 ;
  assign n37644 = n3991 ^ n1167 ^ 1'b0 ;
  assign n37646 = ~n6009 & n29563 ;
  assign n37647 = ( n2628 & n17552 ) | ( n2628 & ~n37646 ) | ( n17552 & ~n37646 ) ;
  assign n37645 = n6052 | n24121 ;
  assign n37648 = n37647 ^ n37645 ^ 1'b0 ;
  assign n37649 = n13423 | n37648 ;
  assign n37650 = n9342 & ~n12277 ;
  assign n37651 = ~n24553 & n27688 ;
  assign n37652 = n29192 ^ n17895 ^ n7330 ;
  assign n37653 = n37652 ^ n10197 ^ 1'b0 ;
  assign n37654 = n2230 & ~n10035 ;
  assign n37655 = n9446 & n37654 ;
  assign n37656 = ( n9250 & ~n20707 ) | ( n9250 & n30273 ) | ( ~n20707 & n30273 ) ;
  assign n37657 = n33211 & n37656 ;
  assign n37658 = n37655 & n37657 ;
  assign n37659 = ~n5955 & n25887 ;
  assign n37660 = n18737 ^ n11454 ^ n2348 ;
  assign n37661 = n22733 ^ n14533 ^ n691 ;
  assign n37662 = ~n517 & n14548 ;
  assign n37663 = ~n15943 & n37662 ;
  assign n37664 = n37663 ^ n19505 ^ n14712 ;
  assign n37665 = ( n14964 & n37661 ) | ( n14964 & n37664 ) | ( n37661 & n37664 ) ;
  assign n37666 = ( n32211 & n37660 ) | ( n32211 & ~n37665 ) | ( n37660 & ~n37665 ) ;
  assign n37667 = n2760 & n22980 ;
  assign n37668 = n36 | n217 ;
  assign n37669 = n37668 ^ n17789 ^ 1'b0 ;
  assign n37670 = n37669 ^ n6091 ^ n3447 ;
  assign n37671 = n37670 ^ n21262 ^ n5761 ;
  assign n37672 = n21155 ^ n2431 ^ 1'b0 ;
  assign n37673 = ~n37671 & n37672 ;
  assign n37674 = n5531 & ~n8767 ;
  assign n37675 = n7208 & n22284 ;
  assign n37676 = n16082 & ~n23268 ;
  assign n37677 = ~n5167 & n37676 ;
  assign n37678 = n37677 ^ n8150 ^ 1'b0 ;
  assign n37679 = ~n10145 & n37678 ;
  assign n37680 = ~n9045 & n35884 ;
  assign n37681 = n1273 | n12779 ;
  assign n37682 = n18794 ^ n7817 ^ n5229 ;
  assign n37683 = ~n360 & n1105 ;
  assign n37684 = ~n5240 & n37683 ;
  assign n37685 = n17134 & n21649 ;
  assign n37686 = ( ~n82 & n37684 ) | ( ~n82 & n37685 ) | ( n37684 & n37685 ) ;
  assign n37687 = n12645 ^ n8359 ^ 1'b0 ;
  assign n37688 = n16171 ^ n1281 ^ 1'b0 ;
  assign n37689 = ~n5836 & n37688 ;
  assign n37690 = n5535 & ~n37689 ;
  assign n37691 = n34757 ^ n30210 ^ n19172 ;
  assign n37692 = n37691 ^ n15928 ^ 1'b0 ;
  assign n37693 = n19981 | n27253 ;
  assign n37694 = ~n9912 & n37033 ;
  assign n37695 = n37694 ^ n10665 ^ 1'b0 ;
  assign n37696 = n10376 & n16346 ;
  assign n37697 = n17369 ^ n11459 ^ n7269 ;
  assign n37698 = ~n7672 & n18749 ;
  assign n37699 = n37698 ^ n10313 ^ 1'b0 ;
  assign n37700 = n37697 & ~n37699 ;
  assign n37701 = ~n3235 & n7203 ;
  assign n37702 = ~n7203 & n37701 ;
  assign n37703 = n37702 ^ n245 ^ 1'b0 ;
  assign n37704 = n8128 | n37703 ;
  assign n37705 = n2745 | n37704 ;
  assign n37706 = n32052 & ~n37705 ;
  assign n37707 = n9527 & ~n37706 ;
  assign n37708 = ~n37700 & n37707 ;
  assign n37709 = n33128 ^ n6453 ^ 1'b0 ;
  assign n37710 = ~n6016 & n37709 ;
  assign n37711 = n37710 ^ n4827 ^ 1'b0 ;
  assign n37712 = n25740 ^ n14073 ^ 1'b0 ;
  assign n37713 = n8427 & ~n18638 ;
  assign n37714 = ~n37712 & n37713 ;
  assign n37716 = n14582 ^ n6603 ^ 1'b0 ;
  assign n37717 = n20294 & ~n37716 ;
  assign n37718 = n37717 ^ n8740 ^ 1'b0 ;
  assign n37715 = n23028 | n24852 ;
  assign n37719 = n37718 ^ n37715 ^ 1'b0 ;
  assign n37720 = n27671 ^ n12401 ^ 1'b0 ;
  assign n37721 = n13882 | n15608 ;
  assign n37722 = n37721 ^ n7645 ^ 1'b0 ;
  assign n37723 = n31271 ^ n12327 ^ 1'b0 ;
  assign n37724 = n29342 | n31514 ;
  assign n37725 = n33685 ^ n21848 ^ 1'b0 ;
  assign n37726 = n19084 ^ n7692 ^ 1'b0 ;
  assign n37727 = n10968 & n30787 ;
  assign n37728 = n8014 | n37727 ;
  assign n37729 = n4431 | n37728 ;
  assign n37731 = n1578 & n13110 ;
  assign n37732 = ~n5183 & n37731 ;
  assign n37730 = n6466 & n14313 ;
  assign n37733 = n37732 ^ n37730 ^ 1'b0 ;
  assign n37734 = n406 & n37733 ;
  assign n37735 = ~n21941 & n37734 ;
  assign n37736 = ~n4140 & n14440 ;
  assign n37737 = n21565 & n37736 ;
  assign n37738 = n7183 ^ n726 ^ 1'b0 ;
  assign n37739 = n19693 & ~n37738 ;
  assign n37740 = n14864 & n30068 ;
  assign n37741 = ~n23110 & n33445 ;
  assign n37742 = n9385 ^ n1891 ^ 1'b0 ;
  assign n37743 = ~n6998 & n37742 ;
  assign n37744 = n7850 | n37743 ;
  assign n37745 = n37744 ^ n15398 ^ 1'b0 ;
  assign n37746 = n3905 & n37745 ;
  assign n37747 = ~n21658 & n37746 ;
  assign n37749 = ~n11824 & n23774 ;
  assign n37748 = n3460 & n3677 ;
  assign n37750 = n37749 ^ n37748 ^ 1'b0 ;
  assign n37751 = n33079 ^ n11010 ^ 1'b0 ;
  assign n37752 = ( ~n3568 & n5098 ) | ( ~n3568 & n12985 ) | ( n5098 & n12985 ) ;
  assign n37753 = n5990 ^ n3214 ^ 1'b0 ;
  assign n37754 = n33736 | n37753 ;
  assign n37755 = n23375 ^ n21728 ^ 1'b0 ;
  assign n37756 = ~n240 & n37755 ;
  assign n37757 = n13331 ^ n6511 ^ 1'b0 ;
  assign n37758 = n10623 ^ n6273 ^ 1'b0 ;
  assign n37759 = n37757 | n37758 ;
  assign n37760 = n7380 | n14386 ;
  assign n37761 = n545 & ~n5370 ;
  assign n37762 = n14048 & n37761 ;
  assign n37763 = n11103 | n37762 ;
  assign n37764 = n30107 | n37763 ;
  assign n37765 = n37764 ^ n11118 ^ 1'b0 ;
  assign n37766 = n28014 ^ n2114 ^ 1'b0 ;
  assign n37767 = ~n8852 & n37766 ;
  assign n37768 = n26772 ^ n12687 ^ 1'b0 ;
  assign n37769 = n17832 & ~n37768 ;
  assign n37770 = n3864 & n5554 ;
  assign n37774 = n1250 | n2766 ;
  assign n37775 = n37774 ^ n6733 ^ 1'b0 ;
  assign n37776 = n37775 ^ n29426 ^ n3470 ;
  assign n37777 = n13031 & ~n16369 ;
  assign n37778 = n37776 & n37777 ;
  assign n37771 = n7350 & n25239 ;
  assign n37772 = ~n31449 & n37771 ;
  assign n37773 = n37772 ^ n7992 ^ 1'b0 ;
  assign n37779 = n37778 ^ n37773 ^ n8989 ;
  assign n37780 = n27405 ^ n25171 ^ n19140 ;
  assign n37781 = n23000 ^ n17407 ^ 1'b0 ;
  assign n37782 = n26833 | n37781 ;
  assign n37783 = ( n9494 & ~n32259 ) | ( n9494 & n37782 ) | ( ~n32259 & n37782 ) ;
  assign n37784 = ( n19985 & ~n33849 ) | ( n19985 & n37783 ) | ( ~n33849 & n37783 ) ;
  assign n37785 = ~n4889 & n6040 ;
  assign n37786 = n37785 ^ n23203 ^ 1'b0 ;
  assign n37787 = n21555 ^ n13881 ^ 1'b0 ;
  assign n37788 = n37786 | n37787 ;
  assign n37789 = n12133 & n12730 ;
  assign n37790 = n18857 ^ n1169 ^ 1'b0 ;
  assign n37791 = n30068 ^ n25402 ^ n8026 ;
  assign n37792 = n3130 & ~n16049 ;
  assign n37793 = n6752 & n37792 ;
  assign n37794 = n11470 | n37793 ;
  assign n37795 = n37794 ^ n27085 ^ 1'b0 ;
  assign n37796 = n10063 | n19986 ;
  assign n37797 = n2196 & ~n36858 ;
  assign n37798 = n24063 ^ n12789 ^ 1'b0 ;
  assign n37799 = ~n8291 & n37798 ;
  assign n37800 = n37799 ^ n3673 ^ 1'b0 ;
  assign n37801 = n23075 ^ n8913 ^ n7216 ;
  assign n37802 = n3491 & ~n9408 ;
  assign n37803 = ~n37801 & n37802 ;
  assign n37804 = ~n25081 & n37803 ;
  assign n37805 = n36839 ^ n2733 ^ 1'b0 ;
  assign n37806 = n36132 ^ n1166 ^ 1'b0 ;
  assign n37807 = ~n28957 & n37806 ;
  assign n37808 = n5557 | n7199 ;
  assign n37809 = ~n1958 & n2699 ;
  assign n37810 = n37809 ^ n32773 ^ 1'b0 ;
  assign n37811 = n23593 ^ n10328 ^ 1'b0 ;
  assign n37812 = n13555 & ~n37811 ;
  assign n37813 = n2857 | n9785 ;
  assign n37814 = n37813 ^ n26184 ^ 1'b0 ;
  assign n37815 = n7289 | n7702 ;
  assign n37816 = n19364 | n21813 ;
  assign n37817 = n22362 | n37816 ;
  assign n37818 = n11573 & n37817 ;
  assign n37819 = n12849 & n37818 ;
  assign n37820 = n1421 | n16780 ;
  assign n37821 = n13440 ^ n5316 ^ 1'b0 ;
  assign n37822 = n26941 ^ n6420 ^ 1'b0 ;
  assign n37823 = n28283 & n37822 ;
  assign n37824 = n16913 & n37823 ;
  assign n37825 = ~n32 & n37824 ;
  assign n37826 = n15849 ^ n401 ^ 1'b0 ;
  assign n37827 = n5582 ^ n881 ^ 1'b0 ;
  assign n37828 = n7252 & n37827 ;
  assign n37829 = n37828 ^ n35609 ^ 1'b0 ;
  assign n37830 = n25171 & n37829 ;
  assign n37831 = ~n6966 & n17890 ;
  assign n37832 = n19443 ^ n18124 ^ 1'b0 ;
  assign n37833 = n37831 & ~n37832 ;
  assign n37834 = n254 & n37833 ;
  assign n37835 = n8395 | n37106 ;
  assign n37836 = n37835 ^ n246 ^ 1'b0 ;
  assign n37837 = n11630 & n37836 ;
  assign n37838 = ( n15514 & ~n27818 ) | ( n15514 & n33433 ) | ( ~n27818 & n33433 ) ;
  assign n37839 = ~n18723 & n19560 ;
  assign n37840 = n6126 & ~n37839 ;
  assign n37841 = ~n15235 & n37840 ;
  assign n37842 = n21449 ^ n6291 ^ 1'b0 ;
  assign n37843 = ~n2568 & n37671 ;
  assign n37844 = n37843 ^ n26440 ^ 1'b0 ;
  assign n37845 = n691 | n9460 ;
  assign n37846 = n12793 | n37845 ;
  assign n37847 = n7312 ^ n37 ^ 1'b0 ;
  assign n37848 = ( n342 & n35503 ) | ( n342 & ~n37847 ) | ( n35503 & ~n37847 ) ;
  assign n37849 = n26453 & ~n30845 ;
  assign n37850 = n28400 & n37849 ;
  assign n37853 = ~n7032 & n24918 ;
  assign n37851 = n18863 & n19785 ;
  assign n37852 = n37851 ^ n18862 ^ 1'b0 ;
  assign n37854 = n37853 ^ n37852 ^ 1'b0 ;
  assign n37855 = n15805 & n18332 ;
  assign n37856 = n9395 & n37855 ;
  assign n37857 = n492 | n17610 ;
  assign n37858 = n37857 ^ n2787 ^ 1'b0 ;
  assign n37859 = n26145 ^ n25417 ^ n14749 ;
  assign n37860 = n24399 & ~n37859 ;
  assign n37861 = n22294 ^ n19856 ^ 1'b0 ;
  assign n37862 = n5312 & n37861 ;
  assign n37863 = ~n61 & n37862 ;
  assign n37864 = n16643 & n37863 ;
  assign n37865 = n31128 & ~n37864 ;
  assign n37866 = n22996 ^ n691 ^ 1'b0 ;
  assign n37867 = n37866 ^ n17804 ^ 1'b0 ;
  assign n37868 = n3558 | n24394 ;
  assign n37869 = n13224 ^ n3644 ^ 1'b0 ;
  assign n37870 = n1412 | n37869 ;
  assign n37871 = n2176 | n37870 ;
  assign n37872 = ( ~n16126 & n18139 ) | ( ~n16126 & n27402 ) | ( n18139 & n27402 ) ;
  assign n37873 = n37872 ^ n33938 ^ n5753 ;
  assign n37874 = n13823 | n17118 ;
  assign n37875 = ~n234 & n2289 ;
  assign n37876 = n2397 & ~n6737 ;
  assign n37877 = ( n16801 & ~n37875 ) | ( n16801 & n37876 ) | ( ~n37875 & n37876 ) ;
  assign n37878 = n5137 | n37877 ;
  assign n37880 = n11852 & n28299 ;
  assign n37881 = n37880 ^ n26178 ^ 1'b0 ;
  assign n37879 = n14638 & ~n25202 ;
  assign n37882 = n37881 ^ n37879 ^ n3376 ;
  assign n37883 = n13766 | n22157 ;
  assign n37884 = n3745 & ~n37883 ;
  assign n37885 = n14821 & ~n37884 ;
  assign n37886 = n12142 & n12184 ;
  assign n37887 = ~n36388 & n37886 ;
  assign n37888 = n29691 ^ n3950 ^ 1'b0 ;
  assign n37889 = n11593 & n29982 ;
  assign n37890 = n36090 & n37889 ;
  assign n37891 = n5261 & n10117 ;
  assign n37892 = ~n8555 & n37891 ;
  assign n37893 = ~n1553 & n9519 ;
  assign n37894 = n15302 | n23024 ;
  assign n37896 = ~n247 & n15470 ;
  assign n37895 = n6457 | n7286 ;
  assign n37897 = n37896 ^ n37895 ^ 1'b0 ;
  assign n37898 = ( ~n13420 & n20237 ) | ( ~n13420 & n37897 ) | ( n20237 & n37897 ) ;
  assign n37899 = n1827 & n16651 ;
  assign n37900 = ~n9631 & n37899 ;
  assign n37903 = n684 | n20596 ;
  assign n37904 = n19397 | n37903 ;
  assign n37901 = ( ~n4548 & n7253 ) | ( ~n4548 & n11795 ) | ( n7253 & n11795 ) ;
  assign n37902 = n26987 | n37901 ;
  assign n37905 = n37904 ^ n37902 ^ 1'b0 ;
  assign n37906 = n11642 | n15246 ;
  assign n37907 = n4348 & ~n37906 ;
  assign n37908 = ~n4549 & n37907 ;
  assign n37909 = ( n12658 & n29342 ) | ( n12658 & n30953 ) | ( n29342 & n30953 ) ;
  assign n37911 = n29778 ^ n1726 ^ 1'b0 ;
  assign n37910 = n32 & ~n10986 ;
  assign n37912 = n37911 ^ n37910 ^ 1'b0 ;
  assign n37916 = n9111 | n19180 ;
  assign n37917 = n25279 ^ n17849 ^ 1'b0 ;
  assign n37918 = n37916 & ~n37917 ;
  assign n37913 = n1411 & ~n31881 ;
  assign n37914 = ~n4779 & n37913 ;
  assign n37915 = n37914 ^ n29486 ^ 1'b0 ;
  assign n37919 = n37918 ^ n37915 ^ n31006 ;
  assign n37920 = n24374 ^ n6115 ^ 1'b0 ;
  assign n37921 = n26690 ^ n2177 ^ 1'b0 ;
  assign n37922 = n37921 ^ n5391 ^ 1'b0 ;
  assign n37923 = n31562 | n37922 ;
  assign n37924 = ~n2107 & n5070 ;
  assign n37925 = n23734 & n37924 ;
  assign n37926 = n4693 & ~n23419 ;
  assign n37927 = ~n5786 & n37926 ;
  assign n37928 = n37925 & n37927 ;
  assign n37929 = ~n2759 & n15660 ;
  assign n37930 = n17652 & ~n37929 ;
  assign n37931 = ~n35542 & n37930 ;
  assign n37932 = n37931 ^ n10598 ^ 1'b0 ;
  assign n37933 = n32118 ^ n3681 ^ 1'b0 ;
  assign n37934 = n17285 & n37933 ;
  assign n37935 = n22651 | n26099 ;
  assign n37936 = n1030 & ~n8357 ;
  assign n37937 = n37936 ^ n10358 ^ n9142 ;
  assign n37938 = ( ~n331 & n11120 ) | ( ~n331 & n20719 ) | ( n11120 & n20719 ) ;
  assign n37939 = n8815 | n14310 ;
  assign n37940 = n37938 | n37939 ;
  assign n37941 = n21929 ^ n4151 ^ 1'b0 ;
  assign n37942 = ( n8197 & n20042 ) | ( n8197 & n21332 ) | ( n20042 & n21332 ) ;
  assign n37943 = n29863 ^ n14172 ^ 1'b0 ;
  assign n37944 = ~n15053 & n37943 ;
  assign n37945 = n37077 ^ n813 ^ 1'b0 ;
  assign n37946 = n5287 | n37945 ;
  assign n37947 = n37944 | n37946 ;
  assign n37948 = n19588 & n23997 ;
  assign n37949 = n37948 ^ n19520 ^ 1'b0 ;
  assign n37950 = n890 | n10973 ;
  assign n37951 = ( n4830 & n34693 ) | ( n4830 & ~n37950 ) | ( n34693 & ~n37950 ) ;
  assign n37952 = n37951 ^ n26146 ^ n22891 ;
  assign n37953 = n5710 & n37952 ;
  assign n37954 = ~n811 & n16755 ;
  assign n37955 = n37953 & n37954 ;
  assign n37956 = ~n3925 & n15070 ;
  assign n37957 = n12100 & n37956 ;
  assign n37958 = n37957 ^ n10123 ^ 1'b0 ;
  assign n37959 = n9520 & ~n37958 ;
  assign n37962 = n6785 & n30122 ;
  assign n37963 = n37962 ^ n1457 ^ 1'b0 ;
  assign n37960 = n3825 & ~n22040 ;
  assign n37961 = n37960 ^ n11503 ^ 1'b0 ;
  assign n37964 = n37963 ^ n37961 ^ n4446 ;
  assign n37965 = n15306 ^ n4864 ^ 1'b0 ;
  assign n37966 = n26624 & ~n37965 ;
  assign n37967 = n32610 ^ n7848 ^ 1'b0 ;
  assign n37968 = n11030 & ~n37967 ;
  assign n37969 = n4977 & ~n10541 ;
  assign n37970 = n37969 ^ n33245 ^ n15498 ;
  assign n37971 = n14373 ^ n2868 ^ 1'b0 ;
  assign n37972 = n16499 | n37971 ;
  assign n37973 = n3805 | n37972 ;
  assign n37974 = n37973 ^ n25610 ^ n11652 ;
  assign n37975 = ( n18616 & ~n25283 ) | ( n18616 & n33732 ) | ( ~n25283 & n33732 ) ;
  assign n37976 = ( n10534 & n26446 ) | ( n10534 & n37975 ) | ( n26446 & n37975 ) ;
  assign n37977 = n5036 | n26795 ;
  assign n37978 = n24070 ^ n16124 ^ n156 ;
  assign n37979 = n15953 ^ n13754 ^ 1'b0 ;
  assign n37980 = n17447 & ~n37979 ;
  assign n37981 = ( n9972 & n37978 ) | ( n9972 & ~n37980 ) | ( n37978 & ~n37980 ) ;
  assign n37982 = n37977 | n37981 ;
  assign n37983 = n30377 & ~n37982 ;
  assign n37984 = n7040 | n13514 ;
  assign n37985 = n17131 & n35612 ;
  assign n37986 = ~n33653 & n37985 ;
  assign n37987 = ~n3189 & n4647 ;
  assign n37988 = ~n1237 & n37987 ;
  assign n37989 = n32036 & ~n37988 ;
  assign n37990 = n37989 ^ n18945 ^ 1'b0 ;
  assign n37991 = ~n4624 & n31708 ;
  assign n37992 = n3024 & ~n11656 ;
  assign n37993 = ~n5776 & n37992 ;
  assign n37994 = n21552 | n26873 ;
  assign n37995 = n22085 ^ n5165 ^ 1'b0 ;
  assign n37996 = n37995 ^ n5702 ^ 1'b0 ;
  assign n37997 = ~n9973 & n35198 ;
  assign n37998 = n18157 | n37997 ;
  assign n37999 = n15323 & ~n37998 ;
  assign n38000 = n19805 & ~n37999 ;
  assign n38001 = n10971 | n19985 ;
  assign n38002 = n38000 | n38001 ;
  assign n38003 = ~n5880 & n13923 ;
  assign n38004 = n38003 ^ n33021 ^ 1'b0 ;
  assign n38005 = n38004 ^ n21518 ^ n12255 ;
  assign n38006 = n1276 & ~n26820 ;
  assign n38007 = n38006 ^ n10347 ^ 1'b0 ;
  assign n38008 = n4096 | n38007 ;
  assign n38009 = n38008 ^ n10420 ^ 1'b0 ;
  assign n38010 = n4048 & ~n9801 ;
  assign n38011 = n38010 ^ n32975 ^ 1'b0 ;
  assign n38012 = n2357 & n7508 ;
  assign n38013 = n38012 ^ n20788 ^ 1'b0 ;
  assign n38014 = n18132 ^ n10769 ^ 1'b0 ;
  assign n38015 = n5725 | n38014 ;
  assign n38016 = n36425 ^ n4223 ^ 1'b0 ;
  assign n38017 = n13193 & ~n38016 ;
  assign n38018 = n38017 ^ n18600 ^ 1'b0 ;
  assign n38019 = ( n16207 & n16568 ) | ( n16207 & n38018 ) | ( n16568 & n38018 ) ;
  assign n38020 = n5817 ^ n4966 ^ 1'b0 ;
  assign n38021 = n15601 | n38020 ;
  assign n38022 = n38019 | n38021 ;
  assign n38023 = n16325 | n17251 ;
  assign n38024 = n38023 ^ n20306 ^ 1'b0 ;
  assign n38025 = n14272 ^ n5673 ^ 1'b0 ;
  assign n38026 = ~n3821 & n38025 ;
  assign n38027 = n38026 ^ n31259 ^ n8350 ;
  assign n38031 = n1882 & ~n28525 ;
  assign n38028 = n4860 | n10140 ;
  assign n38029 = n24482 | n38028 ;
  assign n38030 = n38029 ^ n15009 ^ 1'b0 ;
  assign n38032 = n38031 ^ n38030 ^ 1'b0 ;
  assign n38033 = n19875 ^ n498 ^ 1'b0 ;
  assign n38034 = n38033 ^ n21683 ^ 1'b0 ;
  assign n38035 = n1582 & ~n35510 ;
  assign n38036 = ~n10254 & n38035 ;
  assign n38037 = ~n15761 & n22469 ;
  assign n38038 = n469 | n38037 ;
  assign n38039 = n38038 ^ n11575 ^ 1'b0 ;
  assign n38040 = n4906 & n35609 ;
  assign n38041 = ~n6044 & n27821 ;
  assign n38042 = n20213 & n23221 ;
  assign n38043 = n38042 ^ n22493 ^ 1'b0 ;
  assign n38044 = n11642 & n24316 ;
  assign n38045 = n20576 ^ n9687 ^ 1'b0 ;
  assign n38046 = n411 | n38045 ;
  assign n38047 = n38046 ^ n676 ^ 1'b0 ;
  assign n38048 = n22464 | n29788 ;
  assign n38049 = ( n19815 & n34266 ) | ( n19815 & ~n38048 ) | ( n34266 & ~n38048 ) ;
  assign n38050 = n9968 ^ n6157 ^ 1'b0 ;
  assign n38051 = n16510 | n22027 ;
  assign n38052 = ~n11229 & n38051 ;
  assign n38053 = n38050 & n38052 ;
  assign n38054 = n21550 & ~n38053 ;
  assign n38055 = n38054 ^ n6879 ^ 1'b0 ;
  assign n38057 = ( n2667 & n3130 ) | ( n2667 & n3263 ) | ( n3130 & n3263 ) ;
  assign n38058 = n38057 ^ n36713 ^ n27493 ;
  assign n38056 = n836 & n13396 ;
  assign n38059 = n38058 ^ n38056 ^ 1'b0 ;
  assign n38060 = n21489 ^ n3460 ^ 1'b0 ;
  assign n38061 = ~n1849 & n24998 ;
  assign n38062 = ~n7188 & n38061 ;
  assign n38063 = ~n26495 & n38062 ;
  assign n38064 = n38060 & n38063 ;
  assign n38065 = ~n4578 & n14849 ;
  assign n38066 = n15394 | n38065 ;
  assign n38067 = n10600 ^ n6704 ^ 1'b0 ;
  assign n38068 = n22068 & ~n38067 ;
  assign n38069 = n9999 & ~n12925 ;
  assign n38070 = ~n18036 & n38069 ;
  assign n38071 = n16171 ^ n8493 ^ 1'b0 ;
  assign n38077 = n3737 | n16471 ;
  assign n38078 = n38077 ^ n18919 ^ 1'b0 ;
  assign n38079 = ~n2068 & n38078 ;
  assign n38080 = n987 & ~n38079 ;
  assign n38072 = n1564 & ~n15953 ;
  assign n38073 = n38072 ^ n1502 ^ 1'b0 ;
  assign n38074 = n38073 ^ n13642 ^ 1'b0 ;
  assign n38075 = n22411 & n38074 ;
  assign n38076 = n14002 & n38075 ;
  assign n38081 = n38080 ^ n38076 ^ n9457 ;
  assign n38082 = n19170 ^ n1095 ^ 1'b0 ;
  assign n38083 = ~n20426 & n38082 ;
  assign n38084 = n3867 & ~n12949 ;
  assign n38085 = ~n15386 & n38084 ;
  assign n38086 = n2933 | n7583 ;
  assign n38087 = n38085 & ~n38086 ;
  assign n38088 = n2524 ^ n712 ^ 1'b0 ;
  assign n38089 = n27041 ^ n12606 ^ n2915 ;
  assign n38090 = n19857 & ~n30608 ;
  assign n38091 = ( n999 & n38089 ) | ( n999 & n38090 ) | ( n38089 & n38090 ) ;
  assign n38092 = n24976 & ~n38091 ;
  assign n38093 = n5244 & n5979 ;
  assign n38094 = n38093 ^ n6745 ^ 1'b0 ;
  assign n38095 = n2695 & ~n21946 ;
  assign n38096 = n38094 | n38095 ;
  assign n38097 = n26363 ^ n20859 ^ n10016 ;
  assign n38098 = ( n7106 & ~n26805 ) | ( n7106 & n38097 ) | ( ~n26805 & n38097 ) ;
  assign n38099 = n28245 ^ n7380 ^ 1'b0 ;
  assign n38100 = ( ~n8046 & n8205 ) | ( ~n8046 & n9814 ) | ( n8205 & n9814 ) ;
  assign n38101 = n38100 ^ n7820 ^ 1'b0 ;
  assign n38102 = n1903 | n11222 ;
  assign n38103 = n19150 & ~n38102 ;
  assign n38104 = n8526 & ~n17094 ;
  assign n38105 = n38104 ^ n4729 ^ 1'b0 ;
  assign n38106 = n17488 & ~n38105 ;
  assign n38107 = ~n5486 & n38106 ;
  assign n38108 = n10722 ^ n1744 ^ 1'b0 ;
  assign n38109 = n29930 ^ n23091 ^ n3020 ;
  assign n38110 = ~n12403 & n30310 ;
  assign n38111 = n38110 ^ n834 ^ 1'b0 ;
  assign n38112 = n8813 | n33343 ;
  assign n38113 = n26823 ^ n21271 ^ 1'b0 ;
  assign n38114 = n16321 ^ n473 ^ 1'b0 ;
  assign n38115 = n8794 | n38114 ;
  assign n38116 = n8955 | n38115 ;
  assign n38117 = n1318 & ~n38116 ;
  assign n38118 = n38117 ^ n32109 ^ n29029 ;
  assign n38119 = n5638 & n34404 ;
  assign n38120 = ~n18756 & n25582 ;
  assign n38121 = n16661 | n19968 ;
  assign n38122 = n16605 & ~n38121 ;
  assign n38123 = n933 ^ n216 ^ 1'b0 ;
  assign n38124 = n23094 & n38123 ;
  assign n38125 = n13467 | n17451 ;
  assign n38126 = n13684 & ~n38125 ;
  assign n38127 = n38124 | n38126 ;
  assign n38128 = n26476 & n28540 ;
  assign n38129 = n38128 ^ n36027 ^ 1'b0 ;
  assign n38130 = n6304 | n31329 ;
  assign n38131 = n38130 ^ n15316 ^ 1'b0 ;
  assign n38132 = ~n4141 & n29657 ;
  assign n38133 = n38132 ^ n624 ^ 1'b0 ;
  assign n38134 = n38133 ^ n23825 ^ 1'b0 ;
  assign n38135 = n20654 | n38134 ;
  assign n38136 = ( n1489 & ~n15208 ) | ( n1489 & n16632 ) | ( ~n15208 & n16632 ) ;
  assign n38137 = n20919 & n38136 ;
  assign n38138 = n5268 & n6533 ;
  assign n38139 = ( n14187 & ~n24665 ) | ( n14187 & n30156 ) | ( ~n24665 & n30156 ) ;
  assign n38140 = n8761 ^ n5180 ^ n1882 ;
  assign n38141 = ( n4738 & n13889 ) | ( n4738 & n23283 ) | ( n13889 & n23283 ) ;
  assign n38142 = n38141 ^ n26378 ^ 1'b0 ;
  assign n38143 = n38142 ^ n6743 ^ 1'b0 ;
  assign n38144 = ~n16896 & n38143 ;
  assign n38145 = ( n38139 & n38140 ) | ( n38139 & ~n38144 ) | ( n38140 & ~n38144 ) ;
  assign n38146 = n15297 ^ n14204 ^ 1'b0 ;
  assign n38147 = n4665 & n15579 ;
  assign n38148 = n7271 | n38147 ;
  assign n38149 = n38148 ^ n34320 ^ 1'b0 ;
  assign n38150 = n27910 & ~n38045 ;
  assign n38151 = n27525 ^ n2466 ^ 1'b0 ;
  assign n38152 = n14755 & n38151 ;
  assign n38153 = ~n4866 & n38152 ;
  assign n38154 = n21057 & ~n32946 ;
  assign n38155 = n38154 ^ n10718 ^ 1'b0 ;
  assign n38156 = n38155 ^ n32256 ^ 1'b0 ;
  assign n38157 = n11121 | n38156 ;
  assign n38158 = ~n4447 & n8383 ;
  assign n38159 = ( n6261 & n18510 ) | ( n6261 & ~n27340 ) | ( n18510 & ~n27340 ) ;
  assign n38160 = n22947 ^ n1049 ^ 1'b0 ;
  assign n38161 = n1272 & ~n38160 ;
  assign n38162 = n16153 & n18096 ;
  assign n38163 = n38162 ^ n5348 ^ 1'b0 ;
  assign n38164 = n38163 ^ n36374 ^ 1'b0 ;
  assign n38165 = n6098 & ~n24140 ;
  assign n38166 = n24647 ^ n408 ^ 1'b0 ;
  assign n38167 = n24096 & n38166 ;
  assign n38168 = n9713 & n38167 ;
  assign n38169 = n16468 & n38168 ;
  assign n38175 = n10721 | n14740 ;
  assign n38170 = n23847 ^ n4285 ^ 1'b0 ;
  assign n38171 = n18847 ^ n16382 ^ n12503 ;
  assign n38172 = n10467 | n38171 ;
  assign n38173 = n38172 ^ n24670 ^ 1'b0 ;
  assign n38174 = n38170 | n38173 ;
  assign n38176 = n38175 ^ n38174 ^ n20662 ;
  assign n38177 = n11171 | n14949 ;
  assign n38178 = n15730 & ~n36695 ;
  assign n38179 = ~n16284 & n38178 ;
  assign n38180 = n18378 & n25149 ;
  assign n38181 = n10240 | n21139 ;
  assign n38182 = n38181 ^ n29932 ^ 1'b0 ;
  assign n38183 = n35612 ^ n29952 ^ 1'b0 ;
  assign n38184 = n32540 & ~n38183 ;
  assign n38185 = n25660 ^ n5565 ^ 1'b0 ;
  assign n38186 = n33311 | n38185 ;
  assign n38191 = n7565 ^ n47 ^ 1'b0 ;
  assign n38190 = n4740 | n27781 ;
  assign n38187 = n21953 | n32034 ;
  assign n38188 = n2667 & ~n38187 ;
  assign n38189 = n38188 ^ n14332 ^ n12459 ;
  assign n38192 = n38191 ^ n38190 ^ n38189 ;
  assign n38193 = n25625 ^ n7862 ^ 1'b0 ;
  assign n38194 = ~n1996 & n17664 ;
  assign n38195 = n38194 ^ n865 ^ 1'b0 ;
  assign n38196 = n38195 ^ n33820 ^ 1'b0 ;
  assign n38197 = n13541 | n37323 ;
  assign n38198 = n8856 & ~n38197 ;
  assign n38206 = n8527 ^ n7124 ^ 1'b0 ;
  assign n38203 = n11764 ^ n4548 ^ 1'b0 ;
  assign n38199 = n22917 ^ n3868 ^ 1'b0 ;
  assign n38200 = ~n25623 & n38199 ;
  assign n38201 = ~n8298 & n38200 ;
  assign n38202 = n3918 & ~n38201 ;
  assign n38204 = n38203 ^ n38202 ^ 1'b0 ;
  assign n38205 = n38204 ^ n3706 ^ 1'b0 ;
  assign n38207 = n38206 ^ n38205 ^ 1'b0 ;
  assign n38208 = n29401 ^ n5418 ^ n2294 ;
  assign n38209 = n863 & ~n7362 ;
  assign n38210 = n7639 & n38209 ;
  assign n38211 = ~n13862 & n18542 ;
  assign n38212 = ~n38210 & n38211 ;
  assign n38213 = n27411 ^ n17637 ^ 1'b0 ;
  assign n38214 = n8722 | n38213 ;
  assign n38215 = n10949 | n11478 ;
  assign n38216 = n38215 ^ n12830 ^ 1'b0 ;
  assign n38217 = n17447 & ~n38216 ;
  assign n38218 = n38217 ^ n5329 ^ 1'b0 ;
  assign n38219 = n38158 ^ n6128 ^ 1'b0 ;
  assign n38220 = n38218 & n38219 ;
  assign n38221 = ~n2525 & n16407 ;
  assign n38222 = ( ~n19725 & n20726 ) | ( ~n19725 & n38221 ) | ( n20726 & n38221 ) ;
  assign n38223 = n36446 ^ n19744 ^ 1'b0 ;
  assign n38224 = n18888 ^ n1552 ^ 1'b0 ;
  assign n38225 = ~n3755 & n14042 ;
  assign n38226 = n38224 | n38225 ;
  assign n38227 = n9063 & ~n22239 ;
  assign n38228 = n38227 ^ n23858 ^ 1'b0 ;
  assign n38229 = n38228 ^ n1786 ^ 1'b0 ;
  assign n38230 = n2370 & ~n28742 ;
  assign n38231 = n38230 ^ n23095 ^ n12285 ;
  assign n38232 = ( n29685 & n35961 ) | ( n29685 & n38231 ) | ( n35961 & n38231 ) ;
  assign n38233 = ~n1149 & n5372 ;
  assign n38234 = n1064 & ~n38233 ;
  assign n38235 = n5292 & n38234 ;
  assign n38236 = n4729 ^ n3608 ^ 1'b0 ;
  assign n38237 = ~n24639 & n38236 ;
  assign n38238 = n17535 ^ n8234 ^ n3919 ;
  assign n38240 = n33162 ^ n11583 ^ n1179 ;
  assign n38239 = n36321 ^ n9996 ^ n2597 ;
  assign n38241 = n38240 ^ n38239 ^ 1'b0 ;
  assign n38242 = n928 & ~n10408 ;
  assign n38243 = n8655 & n38242 ;
  assign n38244 = ( n341 & ~n1296 ) | ( n341 & n1662 ) | ( ~n1296 & n1662 ) ;
  assign n38245 = n14886 & ~n38244 ;
  assign n38246 = n38245 ^ n5038 ^ 1'b0 ;
  assign n38247 = ~n6288 & n9004 ;
  assign n38248 = ( n5298 & n25518 ) | ( n5298 & n38247 ) | ( n25518 & n38247 ) ;
  assign n38250 = n7893 & n11243 ;
  assign n38251 = ( ~n5568 & n8927 ) | ( ~n5568 & n38250 ) | ( n8927 & n38250 ) ;
  assign n38249 = ~n5630 & n13649 ;
  assign n38252 = n38251 ^ n38249 ^ 1'b0 ;
  assign n38254 = n16363 & ~n35878 ;
  assign n38253 = n8143 | n31242 ;
  assign n38255 = n38254 ^ n38253 ^ 1'b0 ;
  assign n38256 = ~n332 & n6320 ;
  assign n38257 = n8177 ^ n4579 ^ n2390 ;
  assign n38258 = n38257 ^ n14802 ^ n9696 ;
  assign n38259 = n7427 & ~n38258 ;
  assign n38266 = ~n1327 & n8847 ;
  assign n38263 = ~n12536 & n12600 ;
  assign n38264 = n3784 & n38263 ;
  assign n38260 = ~n890 & n1071 ;
  assign n38261 = ~n21671 & n38260 ;
  assign n38262 = n12055 | n38261 ;
  assign n38265 = n38264 ^ n38262 ^ 1'b0 ;
  assign n38267 = n38266 ^ n38265 ^ 1'b0 ;
  assign n38268 = n31429 ^ n14805 ^ 1'b0 ;
  assign n38269 = n9186 & ~n9440 ;
  assign n38271 = n9222 & n22859 ;
  assign n38270 = n8743 & n33263 ;
  assign n38272 = n38271 ^ n38270 ^ 1'b0 ;
  assign n38277 = n4599 ^ n604 ^ 1'b0 ;
  assign n38278 = n11781 & ~n38277 ;
  assign n38273 = n7393 ^ n2440 ^ 1'b0 ;
  assign n38274 = n38273 ^ n14447 ^ 1'b0 ;
  assign n38275 = n6388 & ~n38274 ;
  assign n38276 = n38275 ^ n10657 ^ n5843 ;
  assign n38279 = n38278 ^ n38276 ^ n10034 ;
  assign n38280 = n5595 | n23787 ;
  assign n38281 = n2246 & ~n38280 ;
  assign n38282 = ( ~n30179 & n38279 ) | ( ~n30179 & n38281 ) | ( n38279 & n38281 ) ;
  assign n38283 = n7661 | n10859 ;
  assign n38284 = n3882 ^ n962 ^ 1'b0 ;
  assign n38285 = ~n5783 & n38284 ;
  assign n38286 = n6357 & ~n7556 ;
  assign n38287 = ~n7994 & n38286 ;
  assign n38288 = n13410 & ~n38287 ;
  assign n38289 = ( ~n6466 & n38285 ) | ( ~n6466 & n38288 ) | ( n38285 & n38288 ) ;
  assign n38290 = n4102 | n13537 ;
  assign n38291 = n38290 ^ n26474 ^ 1'b0 ;
  assign n38292 = n38289 & ~n38291 ;
  assign n38293 = n11898 & ~n38292 ;
  assign n38294 = n38293 ^ n31282 ^ 1'b0 ;
  assign n38295 = n1810 & n33236 ;
  assign n38296 = n38295 ^ n14375 ^ 1'b0 ;
  assign n38297 = n38296 ^ n10305 ^ 1'b0 ;
  assign n38298 = n20885 ^ n6702 ^ 1'b0 ;
  assign n38299 = ( n28833 & n28847 ) | ( n28833 & ~n38298 ) | ( n28847 & ~n38298 ) ;
  assign n38300 = n19696 & n21375 ;
  assign n38301 = n38300 ^ n21730 ^ 1'b0 ;
  assign n38302 = n8979 | n38301 ;
  assign n38303 = ~n19306 & n19749 ;
  assign n38304 = n38303 ^ n24264 ^ 1'b0 ;
  assign n38305 = n406 & ~n38304 ;
  assign n38306 = n38305 ^ n27689 ^ 1'b0 ;
  assign n38307 = n960 ^ n230 ^ 1'b0 ;
  assign n38308 = n3530 & n4297 ;
  assign n38309 = n8452 & n38308 ;
  assign n38310 = ( n3277 & ~n7584 ) | ( n3277 & n38309 ) | ( ~n7584 & n38309 ) ;
  assign n38311 = n38310 ^ n9004 ^ 1'b0 ;
  assign n38312 = n15753 | n38311 ;
  assign n38313 = n38307 & ~n38312 ;
  assign n38315 = n3007 ^ n2130 ^ 1'b0 ;
  assign n38316 = n9507 | n38315 ;
  assign n38317 = n7228 & ~n11825 ;
  assign n38318 = ~n38316 & n38317 ;
  assign n38319 = n13383 & n38318 ;
  assign n38314 = n455 & n8575 ;
  assign n38320 = n38319 ^ n38314 ^ 1'b0 ;
  assign n38321 = n38320 ^ n37577 ^ 1'b0 ;
  assign n38324 = n16551 ^ n8745 ^ n2466 ;
  assign n38322 = n18240 & n26464 ;
  assign n38323 = n13678 & n38322 ;
  assign n38325 = n38324 ^ n38323 ^ n11423 ;
  assign n38328 = n16143 ^ n10333 ^ 1'b0 ;
  assign n38326 = n13169 | n29838 ;
  assign n38327 = n31576 & n38326 ;
  assign n38329 = n38328 ^ n38327 ^ 1'b0 ;
  assign n38330 = n25668 ^ n24399 ^ 1'b0 ;
  assign n38331 = n10703 & n15820 ;
  assign n38333 = ~n44 & n8347 ;
  assign n38334 = n38333 ^ n1838 ^ 1'b0 ;
  assign n38332 = n5713 & n24854 ;
  assign n38335 = n38334 ^ n38332 ^ 1'b0 ;
  assign n38336 = n26149 | n29657 ;
  assign n38337 = n25503 ^ n12266 ^ 1'b0 ;
  assign n38338 = n38336 & n38337 ;
  assign n38339 = n7300 | n25900 ;
  assign n38340 = ~n4560 & n38339 ;
  assign n38341 = ~n2605 & n15912 ;
  assign n38342 = ~n35796 & n38341 ;
  assign n38343 = ~n7290 & n25480 ;
  assign n38344 = n4578 ^ n3389 ^ n46 ;
  assign n38345 = ( ~n33619 & n38343 ) | ( ~n33619 & n38344 ) | ( n38343 & n38344 ) ;
  assign n38347 = n5781 | n11891 ;
  assign n38348 = ~n27425 & n38347 ;
  assign n38346 = n36651 ^ n18712 ^ 1'b0 ;
  assign n38349 = n38348 ^ n38346 ^ 1'b0 ;
  assign n38350 = ~n27525 & n29426 ;
  assign n38356 = n5753 & n13522 ;
  assign n38357 = n1397 & n38356 ;
  assign n38352 = n8080 | n13040 ;
  assign n38351 = n2282 & n27982 ;
  assign n38353 = n38352 ^ n38351 ^ 1'b0 ;
  assign n38354 = n10333 & ~n38353 ;
  assign n38355 = ~n28853 & n38354 ;
  assign n38358 = n38357 ^ n38355 ^ 1'b0 ;
  assign n38359 = n14421 | n20995 ;
  assign n38360 = n13866 & ~n38359 ;
  assign n38361 = ( ~n1760 & n2734 ) | ( ~n1760 & n10201 ) | ( n2734 & n10201 ) ;
  assign n38362 = n17411 & n37431 ;
  assign n38363 = ~n9760 & n38362 ;
  assign n38364 = n12596 | n24820 ;
  assign n38365 = n6180 ^ n3762 ^ 1'b0 ;
  assign n38366 = n35564 & ~n37520 ;
  assign n38367 = ~n25103 & n38366 ;
  assign n38368 = n38367 ^ n35781 ^ n12481 ;
  assign n38369 = n5963 | n7520 ;
  assign n38370 = n17055 & ~n38369 ;
  assign n38371 = n969 | n13984 ;
  assign n38372 = ( n1815 & ~n7019 ) | ( n1815 & n38371 ) | ( ~n7019 & n38371 ) ;
  assign n38373 = n8778 & ~n38372 ;
  assign n38374 = n36219 ^ n4781 ^ 1'b0 ;
  assign n38375 = ~n11667 & n38374 ;
  assign n38376 = n32554 & ~n38044 ;
  assign n38377 = ~n33083 & n38376 ;
  assign n38380 = ( n4280 & n20089 ) | ( n4280 & n33931 ) | ( n20089 & n33931 ) ;
  assign n38378 = n28425 ^ n2001 ^ 1'b0 ;
  assign n38379 = n2115 & n38378 ;
  assign n38381 = n38380 ^ n38379 ^ 1'b0 ;
  assign n38382 = n18049 ^ n10313 ^ 1'b0 ;
  assign n38383 = ~n10850 & n38382 ;
  assign n38384 = ~n17039 & n38383 ;
  assign n38385 = ~n1511 & n19564 ;
  assign n38386 = n25564 & n38385 ;
  assign n38387 = n38386 ^ n17734 ^ 1'b0 ;
  assign n38388 = ~n538 & n12249 ;
  assign n38389 = n2879 | n4296 ;
  assign n38390 = n17445 | n38389 ;
  assign n38391 = ( n13500 & n38388 ) | ( n13500 & n38390 ) | ( n38388 & n38390 ) ;
  assign n38392 = ( ~n2082 & n2305 ) | ( ~n2082 & n4917 ) | ( n2305 & n4917 ) ;
  assign n38393 = n14443 | n20718 ;
  assign n38394 = n38393 ^ n24193 ^ 1'b0 ;
  assign n38395 = n38392 & ~n38394 ;
  assign n38396 = n3606 | n32293 ;
  assign n38399 = n26680 | n37189 ;
  assign n38400 = n38399 ^ n35 ^ 1'b0 ;
  assign n38401 = n1444 & ~n38400 ;
  assign n38397 = n34273 ^ n27040 ^ 1'b0 ;
  assign n38398 = n9564 & n38397 ;
  assign n38402 = n38401 ^ n38398 ^ n11400 ;
  assign n38403 = n14876 ^ n7159 ^ 1'b0 ;
  assign n38404 = n10488 ^ n1917 ^ 1'b0 ;
  assign n38405 = n22660 ^ n7920 ^ 1'b0 ;
  assign n38406 = n3153 & n38405 ;
  assign n38407 = n38406 ^ n17652 ^ 1'b0 ;
  assign n38408 = n23676 & n24285 ;
  assign n38409 = n38408 ^ n24051 ^ 1'b0 ;
  assign n38410 = ~n32201 & n38409 ;
  assign n38411 = n6205 & n22700 ;
  assign n38412 = n15804 & n18859 ;
  assign n38413 = n9238 & n9696 ;
  assign n38414 = n8486 & ~n38413 ;
  assign n38415 = n38414 ^ n3466 ^ 1'b0 ;
  assign n38416 = n38415 ^ n3531 ^ 1'b0 ;
  assign n38417 = ~n8365 & n33874 ;
  assign n38418 = n19478 ^ n9260 ^ 1'b0 ;
  assign n38419 = ~n26642 & n35429 ;
  assign n38420 = n38419 ^ n19170 ^ 1'b0 ;
  assign n38422 = n12080 & n14083 ;
  assign n38421 = ~n4904 & n31461 ;
  assign n38423 = n38422 ^ n38421 ^ 1'b0 ;
  assign n38424 = n29524 & n32147 ;
  assign n38425 = n21210 & n38424 ;
  assign n38427 = n17974 ^ n3273 ^ 1'b0 ;
  assign n38428 = ( ~n7687 & n23093 ) | ( ~n7687 & n38427 ) | ( n23093 & n38427 ) ;
  assign n38426 = n2644 & n22267 ;
  assign n38429 = n38428 ^ n38426 ^ 1'b0 ;
  assign n38430 = n18246 ^ n18188 ^ 1'b0 ;
  assign n38431 = n21131 ^ n7357 ^ n289 ;
  assign n38432 = n18945 | n38431 ;
  assign n38433 = n2790 | n38432 ;
  assign n38434 = n26257 ^ n13608 ^ 1'b0 ;
  assign n38435 = ~n6723 & n38434 ;
  assign n38436 = n13770 & n38435 ;
  assign n38437 = n206 & n38436 ;
  assign n38438 = n7692 & n38437 ;
  assign n38439 = n15198 & ~n33393 ;
  assign n38440 = n38439 ^ n10072 ^ 1'b0 ;
  assign n38441 = n19463 ^ n15467 ^ n1596 ;
  assign n38442 = n31299 ^ n4668 ^ 1'b0 ;
  assign n38443 = n6045 | n38442 ;
  assign n38445 = n20521 ^ n12826 ^ n11873 ;
  assign n38446 = n38445 ^ n13133 ^ n8376 ;
  assign n38444 = n7599 & ~n21448 ;
  assign n38447 = n38446 ^ n38444 ^ 1'b0 ;
  assign n38448 = n9321 | n38092 ;
  assign n38449 = n38447 & ~n38448 ;
  assign n38450 = n25640 ^ n17125 ^ 1'b0 ;
  assign n38451 = n2568 | n24472 ;
  assign n38452 = n38451 ^ n15166 ^ 1'b0 ;
  assign n38453 = n5856 | n19198 ;
  assign n38454 = n36314 ^ n18893 ^ 1'b0 ;
  assign n38455 = n10976 & n38435 ;
  assign n38456 = n38455 ^ n1927 ^ 1'b0 ;
  assign n38457 = ~n3069 & n5735 ;
  assign n38458 = n38457 ^ n1206 ^ 1'b0 ;
  assign n38459 = n1891 & ~n30219 ;
  assign n38460 = ~n38458 & n38459 ;
  assign n38461 = n22843 ^ x11 ^ 1'b0 ;
  assign n38462 = n38460 | n38461 ;
  assign n38463 = n7176 & n38462 ;
  assign n38464 = n2686 & n18553 ;
  assign n38465 = n38464 ^ n23068 ^ 1'b0 ;
  assign n38466 = ( n2722 & ~n11202 ) | ( n2722 & n23961 ) | ( ~n11202 & n23961 ) ;
  assign n38467 = n10875 ^ n5412 ^ 1'b0 ;
  assign n38468 = n2084 | n30057 ;
  assign n38469 = n37267 ^ n19618 ^ n8119 ;
  assign n38470 = n22601 ^ n3175 ^ 1'b0 ;
  assign n38471 = n28063 & n38470 ;
  assign n38472 = n12794 | n36379 ;
  assign n38473 = n38472 ^ n36060 ^ 1'b0 ;
  assign n38474 = n12677 ^ n5504 ^ 1'b0 ;
  assign n38475 = ~n16759 & n38474 ;
  assign n38476 = ~n37013 & n38475 ;
  assign n38477 = ~n3582 & n6326 ;
  assign n38478 = n38477 ^ n34134 ^ 1'b0 ;
  assign n38479 = ( n2567 & ~n12617 ) | ( n2567 & n18977 ) | ( ~n12617 & n18977 ) ;
  assign n38480 = n17765 | n38479 ;
  assign n38481 = n38480 ^ n8588 ^ 1'b0 ;
  assign n38482 = ( ~n411 & n1791 ) | ( ~n411 & n36009 ) | ( n1791 & n36009 ) ;
  assign n38483 = ~n8260 & n38482 ;
  assign n38484 = n37379 ^ n4789 ^ 1'b0 ;
  assign n38485 = n12801 | n38484 ;
  assign n38486 = n29344 ^ n12075 ^ 1'b0 ;
  assign n38487 = n19549 & n29513 ;
  assign n38496 = n7914 ^ n4480 ^ n4115 ;
  assign n38494 = n640 | n18504 ;
  assign n38495 = n863 | n38494 ;
  assign n38497 = n38496 ^ n38495 ^ 1'b0 ;
  assign n38498 = n38497 ^ n4738 ^ 1'b0 ;
  assign n38491 = n7287 & n7630 ;
  assign n38488 = ~n6076 & n22233 ;
  assign n38489 = n38488 ^ n11355 ^ n7888 ;
  assign n38490 = n38489 ^ n15537 ^ n14943 ;
  assign n38492 = n38491 ^ n38490 ^ n32537 ;
  assign n38493 = ~n36359 & n38492 ;
  assign n38499 = n38498 ^ n38493 ^ 1'b0 ;
  assign n38503 = n1069 & ~n19947 ;
  assign n38504 = n9968 & n38503 ;
  assign n38500 = n9061 ^ n2871 ^ 1'b0 ;
  assign n38501 = n10709 | n11123 ;
  assign n38502 = n38500 | n38501 ;
  assign n38505 = n38504 ^ n38502 ^ 1'b0 ;
  assign n38506 = n9794 | n37852 ;
  assign n38507 = n38505 & ~n38506 ;
  assign n38508 = ~n8801 & n14760 ;
  assign n38509 = n38508 ^ n15493 ^ 1'b0 ;
  assign n38510 = ( n9162 & ~n10946 ) | ( n9162 & n38509 ) | ( ~n10946 & n38509 ) ;
  assign n38511 = n37429 & ~n37621 ;
  assign n38513 = n13558 & n14938 ;
  assign n38512 = ~n4646 & n6869 ;
  assign n38514 = n38513 ^ n38512 ^ 1'b0 ;
  assign n38515 = n30127 | n38514 ;
  assign n38516 = n23739 ^ n11059 ^ n7583 ;
  assign n38517 = n25244 | n38516 ;
  assign n38518 = n38517 ^ n15972 ^ 1'b0 ;
  assign n38519 = n1766 | n30621 ;
  assign n38520 = n16492 & ~n38519 ;
  assign n38521 = ( n11378 & n20911 ) | ( n11378 & n36331 ) | ( n20911 & n36331 ) ;
  assign n38522 = n38521 ^ n9357 ^ 1'b0 ;
  assign n38523 = n2083 | n28164 ;
  assign n38524 = ( n1893 & n5254 ) | ( n1893 & ~n10718 ) | ( n5254 & ~n10718 ) ;
  assign n38525 = n7126 | n24745 ;
  assign n38526 = n38524 & ~n38525 ;
  assign n38527 = n38526 ^ n9183 ^ 1'b0 ;
  assign n38528 = n7650 & n23428 ;
  assign n38529 = ~n26681 & n38528 ;
  assign n38530 = n12537 | n26179 ;
  assign n38531 = n20788 | n38530 ;
  assign n38532 = n25591 ^ n3045 ^ 1'b0 ;
  assign n38533 = n38532 ^ n25128 ^ 1'b0 ;
  assign n38534 = n26540 ^ n23077 ^ 1'b0 ;
  assign n38535 = n34116 ^ n15772 ^ 1'b0 ;
  assign n38536 = n1050 | n6457 ;
  assign n38537 = n27178 | n38536 ;
  assign n38538 = n2864 | n19285 ;
  assign n38539 = n38538 ^ n11724 ^ 1'b0 ;
  assign n38540 = n38539 ^ n36594 ^ 1'b0 ;
  assign n38541 = n11899 ^ n7138 ^ 1'b0 ;
  assign n38542 = n2126 & n38541 ;
  assign n38543 = n8897 ^ n714 ^ 1'b0 ;
  assign n38544 = n85 & ~n38543 ;
  assign n38545 = n36535 | n38544 ;
  assign n38546 = n16693 & ~n28664 ;
  assign n38547 = n26450 & n38546 ;
  assign n38548 = n4721 & n9393 ;
  assign n38549 = n26918 | n38548 ;
  assign n38550 = n3696 & n38549 ;
  assign n38551 = n1312 | n2601 ;
  assign n38552 = ~n19034 & n38551 ;
  assign n38553 = n38552 ^ n27922 ^ 1'b0 ;
  assign n38554 = ~n1022 & n29310 ;
  assign n38555 = ~n1828 & n38554 ;
  assign n38556 = n9076 ^ n3146 ^ 1'b0 ;
  assign n38557 = n36139 & ~n38556 ;
  assign n38558 = n38555 & n38557 ;
  assign n38559 = n38431 ^ n4368 ^ 1'b0 ;
  assign n38560 = n17991 ^ n2378 ^ n2341 ;
  assign n38561 = n9909 & ~n15801 ;
  assign n38562 = n915 & ~n38561 ;
  assign n38563 = n38562 ^ n5667 ^ 1'b0 ;
  assign n38564 = n6673 & ~n9341 ;
  assign n38565 = ~n38563 & n38564 ;
  assign n38566 = ( n2421 & n9070 ) | ( n2421 & n15900 ) | ( n9070 & n15900 ) ;
  assign n38567 = n7399 ^ n1402 ^ 1'b0 ;
  assign n38568 = n16316 & ~n38567 ;
  assign n38569 = n38568 ^ n20704 ^ 1'b0 ;
  assign n38570 = n33944 & n38569 ;
  assign n38571 = ~n38566 & n38570 ;
  assign n38572 = n7929 & n18712 ;
  assign n38573 = n38572 ^ n10062 ^ 1'b0 ;
  assign n38574 = n27845 ^ n10267 ^ 1'b0 ;
  assign n38575 = n38574 ^ n2778 ^ n1633 ;
  assign n38576 = n3609 & n13821 ;
  assign n38577 = n38576 ^ n29567 ^ 1'b0 ;
  assign n38578 = n17194 & n31128 ;
  assign n38579 = ~n15965 & n38578 ;
  assign n38580 = n23838 | n23980 ;
  assign n38581 = n15254 ^ n6951 ^ 1'b0 ;
  assign n38582 = n38265 | n38581 ;
  assign n38583 = n38580 & ~n38582 ;
  assign n38584 = n4925 & n14829 ;
  assign n38585 = n38584 ^ n2423 ^ 1'b0 ;
  assign n38586 = n38585 ^ n4180 ^ 1'b0 ;
  assign n38587 = n9395 | n38586 ;
  assign n38588 = n32352 & n38587 ;
  assign n38589 = n19748 ^ n16003 ^ 1'b0 ;
  assign n38590 = n38588 | n38589 ;
  assign n38591 = n25747 ^ n23963 ^ n12857 ;
  assign n38593 = n14331 ^ n5811 ^ 1'b0 ;
  assign n38592 = n30915 & n37503 ;
  assign n38594 = n38593 ^ n38592 ^ 1'b0 ;
  assign n38595 = n5979 ^ n1915 ^ 1'b0 ;
  assign n38596 = ( ~n6478 & n9623 ) | ( ~n6478 & n38595 ) | ( n9623 & n38595 ) ;
  assign n38597 = n14285 ^ n283 ^ 1'b0 ;
  assign n38598 = n7467 | n38597 ;
  assign n38599 = n38598 ^ n17378 ^ 1'b0 ;
  assign n38600 = n18453 & ~n38599 ;
  assign n38601 = ~n33008 & n38600 ;
  assign n38602 = ~n38596 & n38601 ;
  assign n38603 = ~n2992 & n27759 ;
  assign n38604 = n33326 & n38603 ;
  assign n38605 = ~n68 & n35860 ;
  assign n38606 = n16871 & ~n25550 ;
  assign n38607 = n38606 ^ n14916 ^ 1'b0 ;
  assign n38608 = ( n8748 & n27353 ) | ( n8748 & ~n38607 ) | ( n27353 & ~n38607 ) ;
  assign n38609 = n38608 ^ n19727 ^ 1'b0 ;
  assign n38610 = n36664 ^ n26664 ^ 1'b0 ;
  assign n38611 = ( ~n84 & n29563 ) | ( ~n84 & n38610 ) | ( n29563 & n38610 ) ;
  assign n38613 = n926 & n2328 ;
  assign n38614 = ~n33736 & n34001 ;
  assign n38615 = ( n1563 & n38613 ) | ( n1563 & n38614 ) | ( n38613 & n38614 ) ;
  assign n38612 = n4120 & ~n16536 ;
  assign n38616 = n38615 ^ n38612 ^ 1'b0 ;
  assign n38617 = ( n5088 & ~n11100 ) | ( n5088 & n38616 ) | ( ~n11100 & n38616 ) ;
  assign n38618 = n38617 ^ n16785 ^ 1'b0 ;
  assign n38619 = ~n1267 & n25334 ;
  assign n38620 = ( n30832 & n32045 ) | ( n30832 & n38619 ) | ( n32045 & n38619 ) ;
  assign n38621 = n16955 & n28993 ;
  assign n38622 = n25181 & ~n38621 ;
  assign n38623 = n26783 ^ n6128 ^ 1'b0 ;
  assign n38624 = n2124 & n38623 ;
  assign n38625 = n5790 ^ n1303 ^ 1'b0 ;
  assign n38626 = n38624 & ~n38625 ;
  assign n38627 = n18074 ^ n5120 ^ 1'b0 ;
  assign n38628 = n963 & ~n38627 ;
  assign n38629 = ~n2721 & n13440 ;
  assign n38630 = ~n1614 & n2613 ;
  assign n38631 = n12134 ^ n11819 ^ 1'b0 ;
  assign n38632 = ( ~n645 & n16082 ) | ( ~n645 & n38631 ) | ( n16082 & n38631 ) ;
  assign n38633 = n10773 & ~n38632 ;
  assign n38634 = ( n1487 & n5114 ) | ( n1487 & n16540 ) | ( n5114 & n16540 ) ;
  assign n38635 = n38634 ^ n36380 ^ n20355 ;
  assign n38637 = n22930 ^ n2149 ^ 1'b0 ;
  assign n38638 = n14912 ^ n10350 ^ 1'b0 ;
  assign n38639 = ~n38637 & n38638 ;
  assign n38636 = n2270 & ~n7678 ;
  assign n38640 = n38639 ^ n38636 ^ 1'b0 ;
  assign n38641 = n2413 & ~n19983 ;
  assign n38642 = n7383 & n38641 ;
  assign n38643 = ~n26405 & n29840 ;
  assign n38644 = n38642 & n38643 ;
  assign n38645 = n7918 & ~n14639 ;
  assign n38646 = n38645 ^ n12139 ^ 1'b0 ;
  assign n38647 = n38646 ^ n30441 ^ n1043 ;
  assign n38648 = n2732 ^ n43 ^ 1'b0 ;
  assign n38649 = ~n21895 & n38648 ;
  assign n38650 = n38649 ^ n25335 ^ 1'b0 ;
  assign n38651 = n11378 ^ n11290 ^ n7807 ;
  assign n38652 = n7240 | n38651 ;
  assign n38653 = n16576 ^ n5239 ^ 1'b0 ;
  assign n38654 = n11072 & n38653 ;
  assign n38655 = n35182 ^ n14112 ^ 1'b0 ;
  assign n38656 = n38654 & n38655 ;
  assign n38657 = n28199 ^ n23469 ^ n9483 ;
  assign n38658 = ( n14016 & ~n34194 ) | ( n14016 & n38657 ) | ( ~n34194 & n38657 ) ;
  assign n38659 = n3195 | n12106 ;
  assign n38660 = n7207 ^ n2734 ^ 1'b0 ;
  assign n38661 = n38660 ^ n22981 ^ 1'b0 ;
  assign n38662 = ( n1596 & n7477 ) | ( n1596 & ~n13331 ) | ( n7477 & ~n13331 ) ;
  assign n38663 = ( n19780 & ~n29341 ) | ( n19780 & n38662 ) | ( ~n29341 & n38662 ) ;
  assign n38664 = n23529 ^ n14188 ^ n961 ;
  assign n38668 = ( n9837 & n13580 ) | ( n9837 & ~n13860 ) | ( n13580 & ~n13860 ) ;
  assign n38665 = n7228 & n13921 ;
  assign n38666 = n9615 & n38665 ;
  assign n38667 = n10568 & ~n38666 ;
  assign n38669 = n38668 ^ n38667 ^ 1'b0 ;
  assign n38670 = n13464 | n38669 ;
  assign n38671 = n31788 ^ n9284 ^ 1'b0 ;
  assign n38672 = ~n1766 & n38671 ;
  assign n38673 = n38672 ^ n14201 ^ 1'b0 ;
  assign n38674 = n13202 ^ n4044 ^ n2778 ;
  assign n38675 = n35552 & n38674 ;
  assign n38676 = n2836 ^ n2059 ^ 1'b0 ;
  assign n38677 = n8455 | n38676 ;
  assign n38678 = n20526 | n38677 ;
  assign n38679 = n8768 & n28316 ;
  assign n38680 = n38679 ^ n5311 ^ 1'b0 ;
  assign n38681 = n15260 | n23546 ;
  assign n38682 = ~n1442 & n9434 ;
  assign n38683 = n38682 ^ n6474 ^ 1'b0 ;
  assign n38684 = ~n8480 & n38683 ;
  assign n38685 = n38684 ^ n7516 ^ 1'b0 ;
  assign n38686 = n15376 ^ n4936 ^ 1'b0 ;
  assign n38687 = n15879 | n38686 ;
  assign n38688 = n38687 ^ n21347 ^ 1'b0 ;
  assign n38689 = n23937 & ~n38688 ;
  assign n38690 = n8197 & n38689 ;
  assign n38691 = n22961 & ~n33944 ;
  assign n38692 = n37396 & ~n38691 ;
  assign n38693 = n22241 & ~n38692 ;
  assign n38694 = n38690 & n38693 ;
  assign n38695 = n2831 & ~n6368 ;
  assign n38696 = n38695 ^ n3461 ^ 1'b0 ;
  assign n38697 = n4713 | n10649 ;
  assign n38698 = ~n10727 & n38697 ;
  assign n38699 = ~n26821 & n33468 ;
  assign n38700 = n25 & n38699 ;
  assign n38701 = n13881 & ~n27146 ;
  assign n38702 = n38701 ^ n36112 ^ 1'b0 ;
  assign n38703 = ~n16903 & n23743 ;
  assign n38704 = n6877 ^ n3255 ^ 1'b0 ;
  assign n38705 = n38703 & ~n38704 ;
  assign n38706 = n21556 ^ n296 ^ 1'b0 ;
  assign n38707 = n8205 | n31864 ;
  assign n38708 = n34076 ^ n228 ^ 1'b0 ;
  assign n38709 = n9459 ^ n2674 ^ 1'b0 ;
  assign n38710 = ~n1041 & n38709 ;
  assign n38711 = n1312 & n38710 ;
  assign n38712 = n34733 & n38711 ;
  assign n38713 = n3934 & n9304 ;
  assign n38714 = n16033 | n38713 ;
  assign n38715 = n38712 & ~n38714 ;
  assign n38716 = ( n6889 & ~n27940 ) | ( n6889 & n38715 ) | ( ~n27940 & n38715 ) ;
  assign n38717 = n18164 ^ n4006 ^ n3803 ;
  assign n38718 = n38717 ^ n5822 ^ 1'b0 ;
  assign n38719 = n334 & ~n18848 ;
  assign n38720 = n38719 ^ n2008 ^ 1'b0 ;
  assign n38721 = n38720 ^ n30966 ^ 1'b0 ;
  assign n38722 = ~n9921 & n38721 ;
  assign n38724 = n3495 & n3898 ;
  assign n38725 = n32689 & n38724 ;
  assign n38723 = n22865 & ~n23718 ;
  assign n38726 = n38725 ^ n38723 ^ 1'b0 ;
  assign n38727 = n25630 ^ n3866 ^ 1'b0 ;
  assign n38728 = n11788 | n38727 ;
  assign n38729 = n38726 | n38728 ;
  assign n38730 = n12468 | n36682 ;
  assign n38731 = ~n3959 & n23290 ;
  assign n38732 = n8177 ^ n8094 ^ 1'b0 ;
  assign n38733 = n38731 & ~n38732 ;
  assign n38735 = n3040 & ~n16324 ;
  assign n38734 = n36529 ^ n28789 ^ n4708 ;
  assign n38736 = n38735 ^ n38734 ^ 1'b0 ;
  assign n38737 = ~n2082 & n35669 ;
  assign n38738 = n18100 ^ n11382 ^ n2469 ;
  assign n38739 = n24051 & ~n38738 ;
  assign n38740 = n38739 ^ n26924 ^ 1'b0 ;
  assign n38741 = n26293 ^ n5391 ^ 1'b0 ;
  assign n38742 = n556 & n3505 ;
  assign n38743 = n38742 ^ n10195 ^ 1'b0 ;
  assign n38744 = n38743 ^ n19468 ^ n14864 ;
  assign n38745 = ( ~n15356 & n20078 ) | ( ~n15356 & n38744 ) | ( n20078 & n38744 ) ;
  assign n38746 = n10498 & n15146 ;
  assign n38747 = n25460 ^ n11695 ^ 1'b0 ;
  assign n38748 = n9452 | n18226 ;
  assign n38749 = n4350 & n24739 ;
  assign n38753 = n2165 & n3818 ;
  assign n38750 = n17166 ^ n7076 ^ 1'b0 ;
  assign n38751 = n1977 & n38750 ;
  assign n38752 = ~n9074 & n38751 ;
  assign n38754 = n38753 ^ n38752 ^ 1'b0 ;
  assign n38755 = n33664 ^ n762 ^ 1'b0 ;
  assign n38756 = n9111 & ~n38755 ;
  assign n38757 = n2170 & n16304 ;
  assign n38758 = ~n38756 & n38757 ;
  assign n38759 = n27950 ^ n11301 ^ n201 ;
  assign n38760 = n3938 | n18014 ;
  assign n38761 = n38760 ^ n10151 ^ 1'b0 ;
  assign n38762 = n25074 ^ n18921 ^ 1'b0 ;
  assign n38763 = n14514 & ~n38762 ;
  assign n38764 = n26404 ^ n17755 ^ 1'b0 ;
  assign n38765 = n38763 & n38764 ;
  assign n38766 = n22472 ^ n17687 ^ 1'b0 ;
  assign n38767 = ( n10217 & n13946 ) | ( n10217 & ~n14798 ) | ( n13946 & ~n14798 ) ;
  assign n38768 = n38767 ^ n7690 ^ 1'b0 ;
  assign n38769 = ~n21029 & n38768 ;
  assign n38770 = ~n694 & n38769 ;
  assign n38771 = n14428 & ~n38770 ;
  assign n38772 = n33884 & ~n38771 ;
  assign n38773 = n38766 & n38772 ;
  assign n38776 = n10274 ^ n3386 ^ 1'b0 ;
  assign n38774 = ~n3580 & n35308 ;
  assign n38775 = n38774 ^ n20696 ^ 1'b0 ;
  assign n38777 = n38776 ^ n38775 ^ n12838 ;
  assign n38778 = ( ~n14030 & n15638 ) | ( ~n14030 & n28798 ) | ( n15638 & n28798 ) ;
  assign n38779 = n35456 ^ n15321 ^ 1'b0 ;
  assign n38780 = n4060 | n24662 ;
  assign n38781 = n19971 ^ n2100 ^ 1'b0 ;
  assign n38782 = n36102 & n38781 ;
  assign n38783 = n19894 & ~n23987 ;
  assign n38784 = n7932 & n11019 ;
  assign n38785 = n38784 ^ n36258 ^ 1'b0 ;
  assign n38786 = n5576 | n38785 ;
  assign n38787 = n1031 | n38786 ;
  assign n38788 = n38787 ^ n8285 ^ 1'b0 ;
  assign n38789 = ( ~n2504 & n12626 ) | ( ~n2504 & n20120 ) | ( n12626 & n20120 ) ;
  assign n38790 = n38789 ^ n13082 ^ 1'b0 ;
  assign n38793 = n10163 & ~n29072 ;
  assign n38791 = ~n1937 & n12248 ;
  assign n38792 = n38791 ^ n25088 ^ 1'b0 ;
  assign n38794 = n38793 ^ n38792 ^ n30062 ;
  assign n38796 = n2413 & ~n3906 ;
  assign n38797 = n38796 ^ n3914 ^ 1'b0 ;
  assign n38795 = ~n16711 & n36556 ;
  assign n38798 = n38797 ^ n38795 ^ 1'b0 ;
  assign n38799 = n2354 ^ n1455 ^ 1'b0 ;
  assign n38800 = ~n4502 & n38799 ;
  assign n38801 = n14547 ^ n2825 ^ 1'b0 ;
  assign n38802 = n28303 | n38801 ;
  assign n38803 = n2620 | n38802 ;
  assign n38804 = n28874 ^ n5654 ^ 1'b0 ;
  assign n38805 = n38803 & ~n38804 ;
  assign n38806 = n25760 & ~n28472 ;
  assign n38807 = ( n7019 & ~n38805 ) | ( n7019 & n38806 ) | ( ~n38805 & n38806 ) ;
  assign n38808 = n26404 ^ n8847 ^ 1'b0 ;
  assign n38809 = n33597 & ~n38808 ;
  assign n38810 = n3135 | n27000 ;
  assign n38811 = n38810 ^ n21977 ^ n4021 ;
  assign n38812 = n16639 ^ n15953 ^ n8047 ;
  assign n38813 = n21222 ^ n645 ^ 1'b0 ;
  assign n38814 = ~n38812 & n38813 ;
  assign n38815 = n10594 ^ n4364 ^ n1060 ;
  assign n38816 = n38815 ^ n5256 ^ 1'b0 ;
  assign n38817 = n38816 ^ n3309 ^ 1'b0 ;
  assign n38818 = n26790 & n38817 ;
  assign n38819 = n3679 ^ n978 ^ 1'b0 ;
  assign n38820 = ~n25218 & n38819 ;
  assign n38821 = ~n587 & n4683 ;
  assign n38822 = n38821 ^ n14379 ^ n6916 ;
  assign n38823 = n230 & n3376 ;
  assign n38824 = n38823 ^ n28 ^ 1'b0 ;
  assign n38825 = n15934 ^ n320 ^ 1'b0 ;
  assign n38826 = n38825 ^ n3579 ^ 1'b0 ;
  assign n38827 = n21520 & ~n38826 ;
  assign n38828 = ( n20954 & ~n37649 ) | ( n20954 & n38827 ) | ( ~n37649 & n38827 ) ;
  assign n38829 = n26499 & n38828 ;
  assign n38830 = n1959 & ~n16944 ;
  assign n38831 = n17825 ^ n17171 ^ 1'b0 ;
  assign n38832 = n8490 & n38831 ;
  assign n38833 = n8330 ^ n326 ^ 1'b0 ;
  assign n38834 = n8729 & ~n38833 ;
  assign n38835 = n14179 ^ n12445 ^ 1'b0 ;
  assign n38836 = n17372 & n38835 ;
  assign n38837 = n12302 & n29511 ;
  assign n38838 = n13796 & n38837 ;
  assign n38839 = n9530 ^ n6625 ^ 1'b0 ;
  assign n38840 = n38838 | n38839 ;
  assign n38841 = n28641 ^ n8941 ^ 1'b0 ;
  assign n38842 = ( n19927 & n38840 ) | ( n19927 & n38841 ) | ( n38840 & n38841 ) ;
  assign n38843 = ( ~n7332 & n18240 ) | ( ~n7332 & n38842 ) | ( n18240 & n38842 ) ;
  assign n38844 = n36185 ^ n31520 ^ n12796 ;
  assign n38845 = ~n1416 & n10578 ;
  assign n38846 = n38428 ^ n25120 ^ 1'b0 ;
  assign n38847 = n9309 & n38846 ;
  assign n38848 = n32777 ^ n690 ^ 1'b0 ;
  assign n38849 = ~n21752 & n38848 ;
  assign n38850 = n33028 ^ n27992 ^ 1'b0 ;
  assign n38851 = n38849 | n38850 ;
  assign n38852 = n2686 & ~n4221 ;
  assign n38853 = ( ~n2886 & n5585 ) | ( ~n2886 & n11673 ) | ( n5585 & n11673 ) ;
  assign n38854 = n5135 & n38853 ;
  assign n38855 = n38852 & n38854 ;
  assign n38856 = n38855 ^ n14611 ^ 1'b0 ;
  assign n38857 = ( n5878 & ~n26938 ) | ( n5878 & n38856 ) | ( ~n26938 & n38856 ) ;
  assign n38860 = n21312 ^ n4543 ^ 1'b0 ;
  assign n38859 = ~n6657 & n28532 ;
  assign n38858 = n2832 & ~n24270 ;
  assign n38861 = n38860 ^ n38859 ^ n38858 ;
  assign n38862 = n17666 ^ n2793 ^ 1'b0 ;
  assign n38863 = n20386 & ~n38862 ;
  assign n38864 = n38863 ^ n398 ^ 1'b0 ;
  assign n38865 = n9479 ^ n7133 ^ 1'b0 ;
  assign n38866 = n3273 | n38865 ;
  assign n38867 = n14829 & ~n16406 ;
  assign n38868 = n38866 & n38867 ;
  assign n38869 = n38868 ^ n32372 ^ 1'b0 ;
  assign n38870 = n27376 ^ n19212 ^ n16248 ;
  assign n38871 = n38870 ^ n27187 ^ 1'b0 ;
  assign n38872 = ~n23978 & n38871 ;
  assign n38873 = n32173 & n38872 ;
  assign n38874 = n4842 & n14731 ;
  assign n38875 = n38874 ^ n9288 ^ 1'b0 ;
  assign n38876 = n38875 ^ n22818 ^ 1'b0 ;
  assign n38877 = n33459 | n33482 ;
  assign n38878 = n38877 ^ n6948 ^ 1'b0 ;
  assign n38879 = ~n9441 & n17033 ;
  assign n38880 = n38879 ^ n35242 ^ 1'b0 ;
  assign n38881 = ~n11646 & n22477 ;
  assign n38882 = n38881 ^ n15184 ^ 1'b0 ;
  assign n38883 = n8372 ^ n1273 ^ 1'b0 ;
  assign n38884 = n14671 & n38883 ;
  assign n38885 = n38884 ^ n23917 ^ 1'b0 ;
  assign n38886 = ~n2832 & n36623 ;
  assign n38887 = n38886 ^ n17976 ^ 1'b0 ;
  assign n38888 = n4975 ^ n3011 ^ n822 ;
  assign n38889 = ~n249 & n34793 ;
  assign n38890 = n28323 & n38889 ;
  assign n38891 = n38890 ^ n8542 ^ 1'b0 ;
  assign n38892 = n38888 & n38891 ;
  assign n38893 = n27897 & ~n38247 ;
  assign n38894 = n28939 & n38893 ;
  assign n38895 = n38894 ^ n23563 ^ 1'b0 ;
  assign n38896 = ( n436 & ~n6625 ) | ( n436 & n12060 ) | ( ~n6625 & n12060 ) ;
  assign n38897 = n38895 | n38896 ;
  assign n38898 = n8641 & n15789 ;
  assign n38899 = n27788 & n38898 ;
  assign n38901 = ( n5580 & n11111 ) | ( n5580 & n15382 ) | ( n11111 & n15382 ) ;
  assign n38902 = n38901 ^ n23392 ^ 1'b0 ;
  assign n38903 = n10910 & ~n38902 ;
  assign n38900 = n8474 & n17925 ;
  assign n38904 = n38903 ^ n38900 ^ 1'b0 ;
  assign n38905 = n19180 ^ n6206 ^ 1'b0 ;
  assign n38906 = n87 | n11750 ;
  assign n38907 = n38906 ^ n2077 ^ 1'b0 ;
  assign n38908 = n5533 & n18130 ;
  assign n38909 = n26034 & ~n38908 ;
  assign n38910 = ( ~n10990 & n14443 ) | ( ~n10990 & n27405 ) | ( n14443 & n27405 ) ;
  assign n38911 = n37236 & n38910 ;
  assign n38912 = n25039 & n38911 ;
  assign n38913 = n26913 ^ n21952 ^ 1'b0 ;
  assign n38914 = n26540 & n35074 ;
  assign n38918 = n15112 ^ n9117 ^ n2579 ;
  assign n38916 = ( ~x10 & n563 ) | ( ~x10 & n5359 ) | ( n563 & n5359 ) ;
  assign n38915 = n7150 & n22466 ;
  assign n38917 = n38916 ^ n38915 ^ 1'b0 ;
  assign n38919 = n38918 ^ n38917 ^ 1'b0 ;
  assign n38920 = n38919 ^ n35719 ^ n34999 ;
  assign n38921 = n10123 & n13699 ;
  assign n38922 = n38921 ^ n26159 ^ 1'b0 ;
  assign n38923 = n12100 ^ n3925 ^ 1'b0 ;
  assign n38924 = n1107 & ~n20627 ;
  assign n38925 = n38923 & n38924 ;
  assign n38926 = n24822 ^ n12752 ^ 1'b0 ;
  assign n38927 = n24555 ^ n15950 ^ 1'b0 ;
  assign n38928 = n13798 ^ n6571 ^ 1'b0 ;
  assign n38929 = n34589 ^ n17455 ^ 1'b0 ;
  assign n38930 = n16269 ^ n594 ^ 1'b0 ;
  assign n38931 = n24249 | n38930 ;
  assign n38932 = n7572 | n30189 ;
  assign n38933 = n5342 | n35571 ;
  assign n38934 = n38933 ^ n15490 ^ 1'b0 ;
  assign n38935 = n7929 & ~n26770 ;
  assign n38936 = n5099 & ~n5740 ;
  assign n38937 = ~n38935 & n38936 ;
  assign n38938 = ~n740 & n11129 ;
  assign n38939 = n38938 ^ n24332 ^ n11038 ;
  assign n38940 = n9705 | n38939 ;
  assign n38941 = n1407 | n38940 ;
  assign n38943 = n14101 | n30638 ;
  assign n38942 = n10118 | n13969 ;
  assign n38944 = n38943 ^ n38942 ^ 1'b0 ;
  assign n38945 = n10212 & n38944 ;
  assign n38946 = n10875 & ~n15317 ;
  assign n38947 = n3313 & ~n5309 ;
  assign n38948 = ~n4743 & n38947 ;
  assign n38949 = n7414 & n9621 ;
  assign n38950 = n38949 ^ n5756 ^ 1'b0 ;
  assign n38951 = n38950 ^ n22941 ^ 1'b0 ;
  assign n38952 = n9014 ^ n6835 ^ n611 ;
  assign n38953 = n10304 ^ n2236 ^ 1'b0 ;
  assign n38954 = n806 & n38953 ;
  assign n38955 = ( n2745 & n38952 ) | ( n2745 & n38954 ) | ( n38952 & n38954 ) ;
  assign n38956 = n4380 & n38955 ;
  assign n38957 = n38956 ^ n8122 ^ 1'b0 ;
  assign n38958 = n8520 & ~n38957 ;
  assign n38961 = n5333 & n5692 ;
  assign n38962 = n38961 ^ n4126 ^ 1'b0 ;
  assign n38959 = n17287 & ~n18996 ;
  assign n38960 = n38959 ^ n30371 ^ 1'b0 ;
  assign n38963 = n38962 ^ n38960 ^ 1'b0 ;
  assign n38970 = n13418 ^ n6639 ^ 1'b0 ;
  assign n38971 = ~n448 & n38970 ;
  assign n38964 = n30235 ^ n2594 ^ 1'b0 ;
  assign n38965 = n7035 & ~n38964 ;
  assign n38966 = n11902 ^ n11731 ^ 1'b0 ;
  assign n38967 = n209 | n38966 ;
  assign n38968 = n38967 ^ n4614 ^ n1250 ;
  assign n38969 = n38965 & ~n38968 ;
  assign n38972 = n38971 ^ n38969 ^ 1'b0 ;
  assign n38973 = n31420 ^ n9118 ^ 1'b0 ;
  assign n38974 = n36099 & n38973 ;
  assign n38975 = n9339 & ~n19560 ;
  assign n38976 = n38975 ^ n9120 ^ 1'b0 ;
  assign n38977 = n36419 ^ n5965 ^ 1'b0 ;
  assign n38978 = n12111 | n38977 ;
  assign n38979 = ~n14687 & n21245 ;
  assign n38980 = ( n2228 & n7268 ) | ( n2228 & ~n10449 ) | ( n7268 & ~n10449 ) ;
  assign n38981 = n37356 ^ n18690 ^ 1'b0 ;
  assign n38982 = ~n10490 & n16706 ;
  assign n38985 = n3923 & ~n23958 ;
  assign n38983 = n22850 ^ n8443 ^ 1'b0 ;
  assign n38984 = ~n8355 & n38983 ;
  assign n38986 = n38985 ^ n38984 ^ 1'b0 ;
  assign n38987 = ~n7128 & n38986 ;
  assign n38988 = n34122 ^ n1213 ^ 1'b0 ;
  assign n38989 = n38987 & ~n38988 ;
  assign n38990 = ~n7607 & n29457 ;
  assign n38991 = n14213 & n38990 ;
  assign n38992 = n15907 ^ n10715 ^ 1'b0 ;
  assign n38993 = n15803 ^ n9050 ^ 1'b0 ;
  assign n38995 = n3736 | n8126 ;
  assign n38996 = n38995 ^ n8086 ^ 1'b0 ;
  assign n38994 = ~n5312 & n30301 ;
  assign n38997 = n38996 ^ n38994 ^ 1'b0 ;
  assign n38998 = n18097 & n32762 ;
  assign n38999 = n8249 & n11301 ;
  assign n39000 = ~n442 & n469 ;
  assign n39001 = ~n3301 & n39000 ;
  assign n39002 = n475 & n17787 ;
  assign n39003 = n5329 | n16419 ;
  assign n39004 = n39003 ^ n3779 ^ 1'b0 ;
  assign n39005 = n21683 ^ n18926 ^ 1'b0 ;
  assign n39006 = ( n39002 & ~n39004 ) | ( n39002 & n39005 ) | ( ~n39004 & n39005 ) ;
  assign n39007 = ( n31130 & ~n39001 ) | ( n31130 & n39006 ) | ( ~n39001 & n39006 ) ;
  assign n39008 = ~n9616 & n15334 ;
  assign n39009 = n1088 & ~n39008 ;
  assign n39010 = ~n11464 & n27027 ;
  assign n39011 = n39010 ^ n15359 ^ 1'b0 ;
  assign n39012 = n17933 & n38917 ;
  assign n39013 = n8355 | n28277 ;
  assign n39014 = n39013 ^ n6635 ^ 1'b0 ;
  assign n39015 = n624 & ~n19995 ;
  assign n39016 = n39014 & n39015 ;
  assign n39017 = n35491 ^ n27766 ^ 1'b0 ;
  assign n39018 = n4340 | n39017 ;
  assign n39019 = n1362 | n39018 ;
  assign n39020 = n9887 | n39019 ;
  assign n39021 = n39020 ^ n15885 ^ n13051 ;
  assign n39022 = n37128 ^ n20453 ^ 1'b0 ;
  assign n39023 = n19527 ^ n6189 ^ 1'b0 ;
  assign n39024 = n17641 ^ n16820 ^ 1'b0 ;
  assign n39025 = n2060 | n18695 ;
  assign n39026 = n39025 ^ n25485 ^ 1'b0 ;
  assign n39027 = n18638 ^ n10170 ^ 1'b0 ;
  assign n39028 = n3767 | n39027 ;
  assign n39029 = n16218 ^ n11063 ^ 1'b0 ;
  assign n39030 = n15925 | n39029 ;
  assign n39031 = n39030 ^ n30927 ^ 1'b0 ;
  assign n39032 = n21318 | n31292 ;
  assign n39033 = n17280 ^ n6292 ^ 1'b0 ;
  assign n39034 = n39033 ^ n3257 ^ n371 ;
  assign n39035 = n13054 ^ n6917 ^ 1'b0 ;
  assign n39036 = n39035 ^ n37175 ^ 1'b0 ;
  assign n39037 = n20311 ^ n10938 ^ 1'b0 ;
  assign n39038 = ~n15150 & n39037 ;
  assign n39039 = ~n32109 & n39038 ;
  assign n39040 = n39039 ^ n16532 ^ 1'b0 ;
  assign n39041 = n7078 & n24509 ;
  assign n39042 = n39040 & n39041 ;
  assign n39043 = n39042 ^ n36163 ^ n31696 ;
  assign n39044 = n32689 ^ n15250 ^ 1'b0 ;
  assign n39045 = n32262 ^ n28338 ^ 1'b0 ;
  assign n39046 = n35951 | n39045 ;
  assign n39047 = n39046 ^ n250 ^ 1'b0 ;
  assign n39048 = ~n5583 & n18325 ;
  assign n39052 = n2778 | n25115 ;
  assign n39053 = n39052 ^ n8577 ^ 1'b0 ;
  assign n39050 = n1376 | n5469 ;
  assign n39051 = n28843 | n39050 ;
  assign n39049 = ( n9261 & n29660 ) | ( n9261 & ~n30808 ) | ( n29660 & ~n30808 ) ;
  assign n39054 = n39053 ^ n39051 ^ n39049 ;
  assign n39055 = n5205 & ~n11344 ;
  assign n39056 = n39055 ^ n7841 ^ 1'b0 ;
  assign n39057 = ~n26571 & n39056 ;
  assign n39058 = n21578 & ~n25590 ;
  assign n39059 = ( ~n3762 & n6447 ) | ( ~n3762 & n39058 ) | ( n6447 & n39058 ) ;
  assign n39060 = n11964 & ~n35036 ;
  assign n39061 = n37655 & n39060 ;
  assign n39062 = n9638 ^ n3686 ^ 1'b0 ;
  assign n39063 = n11307 | n36041 ;
  assign n39066 = ( n4068 & n7518 ) | ( n4068 & ~n9634 ) | ( n7518 & ~n9634 ) ;
  assign n39067 = n39066 ^ n18218 ^ n10307 ;
  assign n39068 = n39067 ^ n753 ^ 1'b0 ;
  assign n39064 = n19228 ^ n7808 ^ n3534 ;
  assign n39065 = n15684 | n39064 ;
  assign n39069 = n39068 ^ n39065 ^ 1'b0 ;
  assign n39071 = n24532 ^ n6847 ^ n6644 ;
  assign n39070 = ~n13379 & n15197 ;
  assign n39072 = n39071 ^ n39070 ^ 1'b0 ;
  assign n39073 = n5932 & ~n32501 ;
  assign n39074 = n39073 ^ n2276 ^ 1'b0 ;
  assign n39075 = n15277 ^ n2631 ^ 1'b0 ;
  assign n39076 = ( ~n7569 & n38275 ) | ( ~n7569 & n39075 ) | ( n38275 & n39075 ) ;
  assign n39077 = ~n2186 & n33445 ;
  assign n39078 = n17551 & n39077 ;
  assign n39079 = n20136 & n39078 ;
  assign n39080 = ~n25073 & n39079 ;
  assign n39081 = n48 & n39080 ;
  assign n39082 = n514 & ~n1193 ;
  assign n39083 = n33526 ^ n473 ^ 1'b0 ;
  assign n39084 = n28188 ^ n20559 ^ 1'b0 ;
  assign n39085 = ~n473 & n39084 ;
  assign n39087 = ( n12408 & n21603 ) | ( n12408 & ~n26565 ) | ( n21603 & ~n26565 ) ;
  assign n39086 = ~n5420 & n16851 ;
  assign n39088 = n39087 ^ n39086 ^ 1'b0 ;
  assign n39089 = n9415 & ~n18231 ;
  assign n39090 = n39089 ^ n10199 ^ 1'b0 ;
  assign n39091 = n23666 | n39090 ;
  assign n39092 = n39091 ^ n9317 ^ 1'b0 ;
  assign n39096 = n750 & ~n10224 ;
  assign n39097 = n21054 & n39096 ;
  assign n39093 = n3659 & n5572 ;
  assign n39094 = n39093 ^ n3939 ^ 1'b0 ;
  assign n39095 = n11314 | n39094 ;
  assign n39098 = n39097 ^ n39095 ^ 1'b0 ;
  assign n39099 = n7862 & ~n9537 ;
  assign n39100 = n9537 & n39099 ;
  assign n39101 = n23040 | n39100 ;
  assign n39102 = n39101 ^ n19600 ^ 1'b0 ;
  assign n39103 = n39102 ^ n22545 ^ 1'b0 ;
  assign n39104 = n953 & ~n22194 ;
  assign n39105 = n39104 ^ n7081 ^ 1'b0 ;
  assign n39106 = n39105 ^ n33722 ^ n10556 ;
  assign n39107 = n7108 | n17712 ;
  assign n39108 = n39106 & ~n39107 ;
  assign n39109 = n9227 & ~n28302 ;
  assign n39110 = n19197 & n39109 ;
  assign n39111 = n9078 ^ n5978 ^ 1'b0 ;
  assign n39112 = n1807 & ~n39111 ;
  assign n39113 = n7020 & n21912 ;
  assign n39114 = n15309 ^ n4345 ^ 1'b0 ;
  assign n39115 = ~n39113 & n39114 ;
  assign n39116 = n36321 ^ n17649 ^ 1'b0 ;
  assign n39117 = n30703 | n39116 ;
  assign n39118 = n39117 ^ n1167 ^ 1'b0 ;
  assign n39119 = n2089 ^ n396 ^ 1'b0 ;
  assign n39120 = n14206 & n39119 ;
  assign n39121 = ~n2610 & n18565 ;
  assign n39122 = n39121 ^ n10068 ^ 1'b0 ;
  assign n39123 = n39122 ^ n21387 ^ 1'b0 ;
  assign n39124 = n12116 | n39123 ;
  assign n39127 = n34212 ^ n3824 ^ 1'b0 ;
  assign n39128 = n39127 ^ n16021 ^ n1269 ;
  assign n39125 = n4918 | n5044 ;
  assign n39126 = n32944 & ~n39125 ;
  assign n39129 = n39128 ^ n39126 ^ n16715 ;
  assign n39130 = n3435 | n24296 ;
  assign n39131 = n39130 ^ n27122 ^ 1'b0 ;
  assign n39132 = ~n10537 & n34486 ;
  assign n39133 = n39131 & n39132 ;
  assign n39134 = n2083 | n11589 ;
  assign n39135 = n5688 | n39134 ;
  assign n39136 = n39135 ^ n7284 ^ 1'b0 ;
  assign n39137 = n3161 & n6313 ;
  assign n39138 = n39137 ^ n6689 ^ 1'b0 ;
  assign n39139 = n39138 ^ n153 ^ 1'b0 ;
  assign n39140 = n1415 ^ n147 ^ 1'b0 ;
  assign n39141 = ( n6639 & ~n8120 ) | ( n6639 & n39140 ) | ( ~n8120 & n39140 ) ;
  assign n39142 = n39141 ^ n7112 ^ 1'b0 ;
  assign n39143 = n10473 ^ n187 ^ 1'b0 ;
  assign n39144 = n18302 ^ n3650 ^ n777 ;
  assign n39145 = n22881 & n39144 ;
  assign n39146 = n4072 & n39145 ;
  assign n39147 = n6851 & n23686 ;
  assign n39148 = n1032 & n34173 ;
  assign n39150 = ( n448 & n2463 ) | ( n448 & n5937 ) | ( n2463 & n5937 ) ;
  assign n39151 = n39150 ^ n31906 ^ n20872 ;
  assign n39149 = n21056 ^ n17943 ^ n7944 ;
  assign n39152 = n39151 ^ n39149 ^ 1'b0 ;
  assign n39153 = n33003 ^ n2094 ^ 1'b0 ;
  assign n39154 = n3286 | n8936 ;
  assign n39155 = n27605 ^ n4038 ^ 1'b0 ;
  assign n39156 = n6943 & ~n39155 ;
  assign n39157 = ( ~n11225 & n17838 ) | ( ~n11225 & n28749 ) | ( n17838 & n28749 ) ;
  assign n39158 = n13316 ^ n5722 ^ 1'b0 ;
  assign n39159 = n32339 & ~n39158 ;
  assign n39160 = n7031 ^ n1378 ^ 1'b0 ;
  assign n39161 = n39160 ^ n5867 ^ 1'b0 ;
  assign n39162 = ~n11743 & n39161 ;
  assign n39163 = n1182 & n11652 ;
  assign n39164 = n12070 | n17199 ;
  assign n39165 = n20351 & ~n39164 ;
  assign n39166 = ~n13040 & n39165 ;
  assign n39167 = n14047 ^ n3581 ^ 1'b0 ;
  assign n39168 = n39166 & n39167 ;
  assign n39169 = ( n26126 & n39163 ) | ( n26126 & ~n39168 ) | ( n39163 & ~n39168 ) ;
  assign n39170 = n1841 | n12696 ;
  assign n39171 = n39170 ^ n762 ^ 1'b0 ;
  assign n39172 = ( n10026 & n12641 ) | ( n10026 & n39171 ) | ( n12641 & n39171 ) ;
  assign n39173 = n39172 ^ n20962 ^ 1'b0 ;
  assign n39175 = ( ~n1988 & n20890 ) | ( ~n1988 & n21262 ) | ( n20890 & n21262 ) ;
  assign n39174 = ~n8967 & n10679 ;
  assign n39176 = n39175 ^ n39174 ^ 1'b0 ;
  assign n39177 = n39176 ^ n70 ^ 1'b0 ;
  assign n39178 = n15389 & ~n39177 ;
  assign n39179 = n39178 ^ n12136 ^ 1'b0 ;
  assign n39184 = n22624 ^ n18031 ^ n8313 ;
  assign n39185 = ~n2718 & n39184 ;
  assign n39186 = n39185 ^ n22094 ^ n21895 ;
  assign n39180 = n6890 & n26430 ;
  assign n39181 = n38166 ^ n20460 ^ 1'b0 ;
  assign n39182 = n39180 & ~n39181 ;
  assign n39183 = n17838 & n39182 ;
  assign n39187 = n39186 ^ n39183 ^ 1'b0 ;
  assign n39188 = ~n147 & n4563 ;
  assign n39189 = n29257 ^ n18929 ^ 1'b0 ;
  assign n39191 = n3993 | n6931 ;
  assign n39192 = n29863 | n39191 ;
  assign n39190 = ~n10509 & n34677 ;
  assign n39193 = n39192 ^ n39190 ^ 1'b0 ;
  assign n39194 = n9065 | n14543 ;
  assign n39195 = n39194 ^ n9438 ^ 1'b0 ;
  assign n39196 = n39195 ^ n4218 ^ 1'b0 ;
  assign n39197 = n26307 & ~n39196 ;
  assign n39198 = n13795 & ~n15214 ;
  assign n39199 = x3 | n2486 ;
  assign n39207 = n34912 ^ n6948 ^ 1'b0 ;
  assign n39208 = n5862 | n39207 ;
  assign n39204 = ~n2208 & n17825 ;
  assign n39205 = n39204 ^ n5455 ^ 1'b0 ;
  assign n39206 = n21663 & ~n39205 ;
  assign n39209 = n39208 ^ n39206 ^ 1'b0 ;
  assign n39200 = n20608 & n22008 ;
  assign n39201 = n39200 ^ n16531 ^ 1'b0 ;
  assign n39202 = n39201 ^ n37901 ^ n11054 ;
  assign n39203 = n39202 ^ n22918 ^ 1'b0 ;
  assign n39210 = n39209 ^ n39203 ^ 1'b0 ;
  assign n39211 = n453 | n3578 ;
  assign n39212 = n3989 | n39211 ;
  assign n39213 = ( n2569 & ~n4678 ) | ( n2569 & n39212 ) | ( ~n4678 & n39212 ) ;
  assign n39214 = n38985 ^ n34000 ^ 1'b0 ;
  assign n39215 = n22883 | n39214 ;
  assign n39216 = n11873 & ~n23137 ;
  assign n39217 = n12252 & n39216 ;
  assign n39218 = n12670 & n39217 ;
  assign n39219 = n1137 | n23089 ;
  assign n39220 = n20134 | n39219 ;
  assign n39221 = n19312 | n26172 ;
  assign n39222 = n7645 & n39221 ;
  assign n39223 = ~n11195 & n39222 ;
  assign n39224 = ( n3442 & n3906 ) | ( n3442 & n4681 ) | ( n3906 & n4681 ) ;
  assign n39225 = n7470 ^ n1439 ^ 1'b0 ;
  assign n39226 = n21409 | n39225 ;
  assign n39227 = n9987 & n10635 ;
  assign n39228 = n39226 | n39227 ;
  assign n39229 = n39228 ^ n21184 ^ 1'b0 ;
  assign n39230 = n4615 ^ n1073 ^ 1'b0 ;
  assign n39231 = ~n4045 & n39230 ;
  assign n39232 = n39231 ^ n12332 ^ n7295 ;
  assign n39233 = n10373 & n17443 ;
  assign n39234 = n39233 ^ n9504 ^ 1'b0 ;
  assign n39235 = ( n2221 & n15326 ) | ( n2221 & n39234 ) | ( n15326 & n39234 ) ;
  assign n39236 = n34431 ^ n16086 ^ n2062 ;
  assign n39237 = n16454 ^ n3630 ^ 1'b0 ;
  assign n39238 = n3040 & ~n39237 ;
  assign n39239 = n39238 ^ n15641 ^ 1'b0 ;
  assign n39240 = n39239 ^ n28297 ^ n7681 ;
  assign n39241 = n12856 & n20612 ;
  assign n39242 = n39241 ^ n8979 ^ 1'b0 ;
  assign n39243 = ~n2815 & n6666 ;
  assign n39244 = ~n39242 & n39243 ;
  assign n39245 = n39244 ^ n20387 ^ n1621 ;
  assign n39246 = ~n2899 & n15012 ;
  assign n39248 = ( n4147 & n5535 ) | ( n4147 & ~n9796 ) | ( n5535 & ~n9796 ) ;
  assign n39249 = n39248 ^ n23459 ^ 1'b0 ;
  assign n39247 = ~n10093 & n28516 ;
  assign n39250 = n39249 ^ n39247 ^ 1'b0 ;
  assign n39254 = n16477 & n31407 ;
  assign n39251 = n10263 & ~n22098 ;
  assign n39252 = n39251 ^ n13207 ^ 1'b0 ;
  assign n39253 = n12906 & ~n39252 ;
  assign n39255 = n39254 ^ n39253 ^ 1'b0 ;
  assign n39256 = ( n39246 & n39250 ) | ( n39246 & ~n39255 ) | ( n39250 & ~n39255 ) ;
  assign n39257 = n16372 & n39256 ;
  assign n39258 = n8334 | n30671 ;
  assign n39259 = n39258 ^ n11276 ^ 1'b0 ;
  assign n39260 = n39259 ^ n26239 ^ 1'b0 ;
  assign n39261 = n13136 & ~n15114 ;
  assign n39262 = n39260 & n39261 ;
  assign n39263 = n17993 | n39262 ;
  assign n39264 = n39263 ^ n36424 ^ 1'b0 ;
  assign n39265 = n5493 & ~n26408 ;
  assign n39266 = n34666 & n39265 ;
  assign n39267 = n35601 ^ n34824 ^ n11554 ;
  assign n39268 = ~n14029 & n39267 ;
  assign n39269 = n18928 ^ n18143 ^ 1'b0 ;
  assign n39270 = n16771 ^ n4334 ^ 1'b0 ;
  assign n39271 = n14912 & n39270 ;
  assign n39272 = n32192 & ~n39271 ;
  assign n39273 = n6657 & n28451 ;
  assign n39274 = n39273 ^ n7912 ^ 1'b0 ;
  assign n39275 = ~n525 & n39274 ;
  assign n39276 = n17243 ^ n3844 ^ 1'b0 ;
  assign n39277 = ~n12958 & n37102 ;
  assign n39278 = n23364 & n32112 ;
  assign n39279 = n39278 ^ n2966 ^ 1'b0 ;
  assign n39280 = n17579 ^ n523 ^ 1'b0 ;
  assign n39281 = n22223 & ~n39280 ;
  assign n39282 = n39279 & n39281 ;
  assign n39283 = ~n39277 & n39282 ;
  assign n39284 = n6731 & ~n8881 ;
  assign n39285 = n36393 ^ n20501 ^ 1'b0 ;
  assign n39286 = n1800 & ~n30090 ;
  assign n39287 = ~n1800 & n39286 ;
  assign n39288 = n4487 & n39287 ;
  assign n39289 = n39288 ^ n12858 ^ n1709 ;
  assign n39290 = n969 | n24815 ;
  assign n39291 = n39290 ^ n7147 ^ 1'b0 ;
  assign n39292 = n1858 & ~n9197 ;
  assign n39293 = n39292 ^ n14661 ^ 1'b0 ;
  assign n39294 = n19653 ^ n6553 ^ 1'b0 ;
  assign n39295 = n33209 & n39294 ;
  assign n39296 = n9676 | n24251 ;
  assign n39297 = n39296 ^ n13577 ^ 1'b0 ;
  assign n39298 = n7067 ^ n6000 ^ 1'b0 ;
  assign n39299 = n1880 & ~n39298 ;
  assign n39300 = ~n1426 & n37672 ;
  assign n39301 = ~n39299 & n39300 ;
  assign n39302 = n28884 ^ n13511 ^ 1'b0 ;
  assign n39303 = n22693 & ~n39302 ;
  assign n39304 = n5936 | n37942 ;
  assign n39305 = n39303 | n39304 ;
  assign n39306 = n5584 | n18109 ;
  assign n39307 = n39306 ^ n1083 ^ 1'b0 ;
  assign n39308 = n39307 ^ n14864 ^ 1'b0 ;
  assign n39309 = n39308 ^ n18085 ^ n14961 ;
  assign n39310 = n21262 ^ n12863 ^ n6139 ;
  assign n39311 = n39309 & ~n39310 ;
  assign n39315 = n10935 | n38460 ;
  assign n39316 = n29903 | n39315 ;
  assign n39312 = n2062 & ~n4889 ;
  assign n39313 = n31527 & n39312 ;
  assign n39314 = ( n6142 & n10260 ) | ( n6142 & n39313 ) | ( n10260 & n39313 ) ;
  assign n39317 = n39316 ^ n39314 ^ 1'b0 ;
  assign n39318 = n32264 ^ n21828 ^ n11361 ;
  assign n39319 = n36229 ^ n10457 ^ 1'b0 ;
  assign n39320 = n2545 & n26573 ;
  assign n39321 = n39320 ^ n11345 ^ 1'b0 ;
  assign n39322 = ( ~n3234 & n4966 ) | ( ~n3234 & n16112 ) | ( n4966 & n16112 ) ;
  assign n39323 = ( n1549 & n11999 ) | ( n1549 & ~n38336 ) | ( n11999 & ~n38336 ) ;
  assign n39324 = ~n17146 & n39323 ;
  assign n39325 = n39324 ^ n4044 ^ 1'b0 ;
  assign n39326 = ( ~n7457 & n31882 ) | ( ~n7457 & n39325 ) | ( n31882 & n39325 ) ;
  assign n39327 = ~n20311 & n31795 ;
  assign n39328 = n39327 ^ n18454 ^ 1'b0 ;
  assign n39329 = n25103 ^ n16136 ^ 1'b0 ;
  assign n39330 = ~n4308 & n36194 ;
  assign n39331 = ~n39329 & n39330 ;
  assign n39332 = ( n5229 & n8782 ) | ( n5229 & n10623 ) | ( n8782 & n10623 ) ;
  assign n39333 = n15355 | n39332 ;
  assign n39334 = ~n32794 & n39333 ;
  assign n39335 = n22866 & n39334 ;
  assign n39336 = n27466 ^ n5650 ^ 1'b0 ;
  assign n39337 = n39336 ^ n28153 ^ 1'b0 ;
  assign n39338 = n35526 | n39150 ;
  assign n39339 = n39337 & ~n39338 ;
  assign n39340 = n3943 & ~n13550 ;
  assign n39341 = n39340 ^ n1332 ^ 1'b0 ;
  assign n39342 = n34055 & n39341 ;
  assign n39343 = n39342 ^ n24537 ^ n2495 ;
  assign n39344 = n11873 ^ n4584 ^ 1'b0 ;
  assign n39345 = n9140 & n33253 ;
  assign n39346 = ~n3565 & n25918 ;
  assign n39347 = n31964 & n39346 ;
  assign n39348 = n11690 | n39347 ;
  assign n39349 = n39348 ^ n1487 ^ 1'b0 ;
  assign n39350 = ~n40 & n10531 ;
  assign n39351 = n5832 | n20931 ;
  assign n39352 = ~n30374 & n39351 ;
  assign n39353 = n39350 & n39352 ;
  assign n39354 = n6737 | n39353 ;
  assign n39355 = n39354 ^ n4214 ^ 1'b0 ;
  assign n39359 = n26355 ^ n25372 ^ n361 ;
  assign n39356 = ~n3501 & n12658 ;
  assign n39357 = n39356 ^ n19917 ^ n11301 ;
  assign n39358 = n14246 & ~n39357 ;
  assign n39360 = n39359 ^ n39358 ^ 1'b0 ;
  assign n39361 = n5214 ^ n3389 ^ 1'b0 ;
  assign n39362 = n14112 ^ n1359 ^ 1'b0 ;
  assign n39363 = ~n6431 & n9299 ;
  assign n39364 = ( n6128 & n22235 ) | ( n6128 & n39363 ) | ( n22235 & n39363 ) ;
  assign n39365 = ~n12969 & n14297 ;
  assign n39366 = n39365 ^ n12741 ^ 1'b0 ;
  assign n39367 = n7376 & n11244 ;
  assign n39368 = n39367 ^ n36538 ^ 1'b0 ;
  assign n39369 = ~n17186 & n39368 ;
  assign n39370 = n36064 ^ n22185 ^ 1'b0 ;
  assign n39371 = n21564 | n30634 ;
  assign n39372 = n39371 ^ n21331 ^ 1'b0 ;
  assign n39373 = n27737 ^ n24553 ^ 1'b0 ;
  assign n39374 = ~n5584 & n39373 ;
  assign n39375 = ~n4252 & n15726 ;
  assign n39376 = n39375 ^ n9769 ^ 1'b0 ;
  assign n39377 = ~n6343 & n17815 ;
  assign n39378 = ~n22193 & n39377 ;
  assign n39379 = ~n543 & n39378 ;
  assign n39380 = n38175 ^ n135 ^ 1'b0 ;
  assign n39381 = n17487 & ~n39380 ;
  assign n39382 = n4231 & n26852 ;
  assign n39383 = n39382 ^ n26179 ^ 1'b0 ;
  assign n39384 = n6903 & ~n11285 ;
  assign n39385 = ( n11427 & n39383 ) | ( n11427 & n39384 ) | ( n39383 & n39384 ) ;
  assign n39386 = n10881 & ~n32540 ;
  assign n39387 = n11306 | n20627 ;
  assign n39388 = n1231 & n26521 ;
  assign n39389 = n39388 ^ n4310 ^ 1'b0 ;
  assign n39390 = n39389 ^ n20439 ^ 1'b0 ;
  assign n39391 = ~n39387 & n39390 ;
  assign n39392 = n15537 & n39391 ;
  assign n39393 = n39392 ^ n16368 ^ 1'b0 ;
  assign n39394 = n34761 ^ n1472 ^ 1'b0 ;
  assign n39395 = n10211 & ~n39394 ;
  assign n39396 = ~n3824 & n11994 ;
  assign n39397 = ( n14949 & ~n16351 ) | ( n14949 & n39396 ) | ( ~n16351 & n39396 ) ;
  assign n39398 = n39397 ^ n6560 ^ 1'b0 ;
  assign n39399 = n2296 & n20871 ;
  assign n39400 = n39399 ^ n30850 ^ n1082 ;
  assign n39401 = n26453 ^ n12211 ^ 1'b0 ;
  assign n39402 = n8826 | n39401 ;
  assign n39403 = n4461 | n27608 ;
  assign n39404 = n39403 ^ n38863 ^ 1'b0 ;
  assign n39405 = n33 & ~n32150 ;
  assign n39406 = n2098 | n39405 ;
  assign n39407 = ( ~n1875 & n14110 ) | ( ~n1875 & n36038 ) | ( n14110 & n36038 ) ;
  assign n39408 = n15274 ^ n11035 ^ 1'b0 ;
  assign n39409 = n39407 & n39408 ;
  assign n39413 = ( n682 & n2250 ) | ( n682 & n28885 ) | ( n2250 & n28885 ) ;
  assign n39410 = n28786 | n36810 ;
  assign n39411 = n10348 & ~n39410 ;
  assign n39412 = n39411 ^ n2882 ^ 1'b0 ;
  assign n39414 = n39413 ^ n39412 ^ n17457 ;
  assign n39415 = n8185 & ~n27247 ;
  assign n39416 = n7724 & n12415 ;
  assign n39417 = n39416 ^ n38392 ^ 1'b0 ;
  assign n39418 = ~n16500 & n39417 ;
  assign n39419 = n39418 ^ n2755 ^ 1'b0 ;
  assign n39420 = n538 | n11978 ;
  assign n39421 = n11978 & ~n39420 ;
  assign n39422 = ~n955 & n18622 ;
  assign n39423 = n955 & n39422 ;
  assign n39424 = n39421 | n39423 ;
  assign n39425 = n39424 ^ n630 ^ 1'b0 ;
  assign n39426 = n17504 | n39425 ;
  assign n39427 = n10894 | n32911 ;
  assign n39428 = n9858 | n18613 ;
  assign n39429 = n9858 & ~n39428 ;
  assign n39430 = n10649 ^ n3750 ^ 1'b0 ;
  assign n39431 = n39430 ^ n9228 ^ n6087 ;
  assign n39432 = n72 | n4521 ;
  assign n39433 = n27623 ^ n24197 ^ 1'b0 ;
  assign n39434 = n4877 | n39433 ;
  assign n39435 = n19813 ^ n1145 ^ 1'b0 ;
  assign n39436 = n5996 | n13028 ;
  assign n39437 = n37450 & ~n39436 ;
  assign n39438 = n18975 ^ n18613 ^ 1'b0 ;
  assign n39439 = ~n11656 & n39438 ;
  assign n39440 = n21905 & n39439 ;
  assign n39441 = n26960 ^ n12017 ^ 1'b0 ;
  assign n39442 = ~n2806 & n39441 ;
  assign n39443 = ( n9666 & n11150 ) | ( n9666 & ~n38172 ) | ( n11150 & ~n38172 ) ;
  assign n39444 = n39443 ^ n22615 ^ 1'b0 ;
  assign n39445 = ~n423 & n11271 ;
  assign n39446 = n18837 ^ n12946 ^ 1'b0 ;
  assign n39447 = n13901 & n14207 ;
  assign n39448 = n20312 & n39447 ;
  assign n39449 = ( n6729 & n39446 ) | ( n6729 & n39448 ) | ( n39446 & n39448 ) ;
  assign n39450 = n39445 | n39449 ;
  assign n39451 = n39450 ^ n30915 ^ 1'b0 ;
  assign n39452 = n21165 ^ n11941 ^ 1'b0 ;
  assign n39453 = n31733 & n39452 ;
  assign n39454 = ~n11947 & n39453 ;
  assign n39455 = n878 ^ n263 ^ 1'b0 ;
  assign n39456 = n39455 ^ n10408 ^ 1'b0 ;
  assign n39457 = n32606 & ~n39456 ;
  assign n39458 = n35534 ^ n34756 ^ 1'b0 ;
  assign n39459 = n17881 & ~n39396 ;
  assign n39460 = ( n1918 & n39458 ) | ( n1918 & ~n39459 ) | ( n39458 & ~n39459 ) ;
  assign n39461 = n26697 ^ n408 ^ 1'b0 ;
  assign n39462 = ~n4393 & n36437 ;
  assign n39463 = n39462 ^ n36906 ^ 1'b0 ;
  assign n39464 = n30935 ^ n16707 ^ 1'b0 ;
  assign n39465 = n8615 & n39464 ;
  assign n39466 = n39465 ^ n16028 ^ 1'b0 ;
  assign n39467 = ~n2621 & n39466 ;
  assign n39468 = n24032 & n39467 ;
  assign n39469 = n2022 & ~n6657 ;
  assign n39470 = n39469 ^ n8421 ^ 1'b0 ;
  assign n39471 = n18225 ^ n18074 ^ 1'b0 ;
  assign n39472 = n33644 | n39471 ;
  assign n39473 = n39472 ^ n1962 ^ 1'b0 ;
  assign n39474 = ( n2405 & ~n34398 ) | ( n2405 & n39473 ) | ( ~n34398 & n39473 ) ;
  assign n39475 = n39470 & n39474 ;
  assign n39476 = n20206 & n39475 ;
  assign n39477 = n8941 ^ n543 ^ 1'b0 ;
  assign n39478 = n29010 & ~n39477 ;
  assign n39479 = ( n3702 & n16038 ) | ( n3702 & n39478 ) | ( n16038 & n39478 ) ;
  assign n39480 = n10123 & n23143 ;
  assign n39481 = n30551 & ~n39480 ;
  assign n39482 = n39479 & n39481 ;
  assign n39484 = n23335 & ~n25611 ;
  assign n39485 = n39484 ^ n31158 ^ 1'b0 ;
  assign n39486 = n39485 ^ n2358 ^ 1'b0 ;
  assign n39483 = ~n5987 & n34035 ;
  assign n39487 = n39486 ^ n39483 ^ 1'b0 ;
  assign n39488 = n10263 ^ n8807 ^ n8310 ;
  assign n39489 = n39488 ^ n13798 ^ 1'b0 ;
  assign n39490 = n39489 ^ n8085 ^ 1'b0 ;
  assign n39491 = ~n13256 & n39490 ;
  assign n39492 = n18712 ^ n6320 ^ 1'b0 ;
  assign n39493 = ~n21043 & n39492 ;
  assign n39494 = n19923 ^ n3385 ^ n2348 ;
  assign n39495 = ~n1670 & n27860 ;
  assign n39496 = n39495 ^ n18510 ^ 1'b0 ;
  assign n39497 = n6756 & n39496 ;
  assign n39498 = n16731 | n20047 ;
  assign n39499 = n26821 ^ n76 ^ 1'b0 ;
  assign n39500 = n18748 ^ n7925 ^ 1'b0 ;
  assign n39501 = ~n13817 & n39500 ;
  assign n39502 = ~n39499 & n39501 ;
  assign n39503 = n39502 ^ n20217 ^ 1'b0 ;
  assign n39504 = ~n7772 & n12340 ;
  assign n39505 = n22936 ^ n13049 ^ 1'b0 ;
  assign n39506 = n8163 & n39505 ;
  assign n39510 = n2146 & ~n23941 ;
  assign n39511 = n39510 ^ n2431 ^ 1'b0 ;
  assign n39507 = n11137 & n26184 ;
  assign n39508 = ~n11137 & n39507 ;
  assign n39509 = n18596 | n39508 ;
  assign n39512 = n39511 ^ n39509 ^ 1'b0 ;
  assign n39513 = n17130 | n37544 ;
  assign n39514 = ~n8848 & n33154 ;
  assign n39515 = n30416 ^ n21186 ^ n18923 ;
  assign n39516 = ~n7813 & n32449 ;
  assign n39517 = n26195 & n39516 ;
  assign n39518 = n12166 ^ n74 ^ 1'b0 ;
  assign n39519 = n18652 ^ n16447 ^ 1'b0 ;
  assign n39520 = n4562 & n39519 ;
  assign n39521 = n8034 & n26566 ;
  assign n39522 = n39521 ^ n9251 ^ 1'b0 ;
  assign n39523 = n39520 & ~n39522 ;
  assign n39524 = ~n34793 & n39523 ;
  assign n39528 = n3967 | n20250 ;
  assign n39525 = n192 | n38509 ;
  assign n39526 = n8282 & ~n39525 ;
  assign n39527 = n39526 ^ n31476 ^ n12760 ;
  assign n39529 = n39528 ^ n39527 ^ n37335 ;
  assign n39530 = n39529 ^ n32748 ^ 1'b0 ;
  assign n39531 = n27788 | n39530 ;
  assign n39532 = ~n4511 & n18495 ;
  assign n39533 = n39532 ^ n22672 ^ 1'b0 ;
  assign n39534 = ( ~n13004 & n24444 ) | ( ~n13004 & n24972 ) | ( n24444 & n24972 ) ;
  assign n39535 = n36185 & ~n39534 ;
  assign n39536 = n19190 ^ n13710 ^ 1'b0 ;
  assign n39537 = n485 | n863 ;
  assign n39538 = n38100 ^ n22232 ^ 1'b0 ;
  assign n39539 = n39537 & n39538 ;
  assign n39540 = n22592 | n39539 ;
  assign n39541 = n2338 & ~n37559 ;
  assign n39542 = ~n22768 & n39541 ;
  assign n39543 = n567 & ~n9588 ;
  assign n39544 = n39543 ^ n12442 ^ 1'b0 ;
  assign n39545 = n35069 ^ n4132 ^ 1'b0 ;
  assign n39546 = ( ~n33275 & n39544 ) | ( ~n33275 & n39545 ) | ( n39544 & n39545 ) ;
  assign n39547 = ~n39542 & n39546 ;
  assign n39548 = ~n29441 & n39547 ;
  assign n39549 = ~n2785 & n26104 ;
  assign n39550 = n3390 & ~n12323 ;
  assign n39551 = n39550 ^ n26794 ^ 1'b0 ;
  assign n39552 = n18408 | n39551 ;
  assign n39553 = n13284 & n25556 ;
  assign n39554 = ~n27534 & n39553 ;
  assign n39555 = n3428 & ~n5657 ;
  assign n39556 = n19848 ^ n7699 ^ 1'b0 ;
  assign n39557 = ~n39555 & n39556 ;
  assign n39558 = ~n7672 & n14163 ;
  assign n39559 = n39558 ^ n11495 ^ 1'b0 ;
  assign n39560 = n13181 ^ n113 ^ 1'b0 ;
  assign n39561 = n21733 | n39560 ;
  assign n39562 = n11290 | n16502 ;
  assign n39563 = n39562 ^ n13789 ^ 1'b0 ;
  assign n39564 = ~n5311 & n27046 ;
  assign n39565 = n39564 ^ n29478 ^ n2887 ;
  assign n39566 = n16417 | n17402 ;
  assign n39567 = n39566 ^ n19568 ^ 1'b0 ;
  assign n39568 = n39567 ^ n17100 ^ n12373 ;
  assign n39569 = n39071 | n39568 ;
  assign n39570 = n3252 ^ n2489 ^ 1'b0 ;
  assign n39571 = n21751 | n39570 ;
  assign n39572 = n6743 ^ n1346 ^ 1'b0 ;
  assign n39573 = n11490 & ~n21607 ;
  assign n39574 = ~n39572 & n39573 ;
  assign n39575 = ~n4363 & n26308 ;
  assign n39576 = n2795 ^ n2340 ^ 1'b0 ;
  assign n39577 = n39576 ^ n23276 ^ n15636 ;
  assign n39578 = n16897 ^ n3892 ^ 1'b0 ;
  assign n39579 = n17803 | n39578 ;
  assign n39580 = n29517 | n39579 ;
  assign n39581 = n34935 & ~n39580 ;
  assign n39582 = n39581 ^ n4330 ^ 1'b0 ;
  assign n39583 = n39577 & ~n39582 ;
  assign n39584 = n18321 ^ n1706 ^ 1'b0 ;
  assign n39585 = n2363 & n19833 ;
  assign n39586 = n39585 ^ n1069 ^ 1'b0 ;
  assign n39587 = n28789 & ~n39586 ;
  assign n39588 = n39584 & n39587 ;
  assign n39589 = n14711 ^ n9855 ^ 1'b0 ;
  assign n39590 = n32112 ^ n4294 ^ 1'b0 ;
  assign n39591 = ( n21436 & n39589 ) | ( n21436 & n39590 ) | ( n39589 & n39590 ) ;
  assign n39593 = n35457 ^ n10739 ^ 1'b0 ;
  assign n39594 = ~n2330 & n39593 ;
  assign n39595 = n39594 ^ n395 ^ 1'b0 ;
  assign n39596 = n14583 & n39595 ;
  assign n39597 = n11359 & n39596 ;
  assign n39598 = n20056 | n39597 ;
  assign n39592 = n14769 ^ n6407 ^ 1'b0 ;
  assign n39599 = n39598 ^ n39592 ^ 1'b0 ;
  assign n39600 = n15646 & n39599 ;
  assign n39601 = n315 & ~n39600 ;
  assign n39602 = n6384 | n18820 ;
  assign n39603 = n8960 & ~n39602 ;
  assign n39604 = n17050 & n28203 ;
  assign n39605 = n11772 & n39604 ;
  assign n39606 = n2630 | n5219 ;
  assign n39607 = n25031 & ~n39606 ;
  assign n39608 = n39605 & n39607 ;
  assign n39609 = n29117 ^ n27538 ^ 1'b0 ;
  assign n39610 = ~n39608 & n39609 ;
  assign n39611 = n151 | n21565 ;
  assign n39612 = n14623 & ~n39611 ;
  assign n39613 = n39612 ^ n15036 ^ 1'b0 ;
  assign n39614 = n20092 & ~n39613 ;
  assign n39615 = n38367 ^ n17951 ^ n4292 ;
  assign n39616 = n10319 | n19304 ;
  assign n39617 = n39616 ^ n5963 ^ 1'b0 ;
  assign n39618 = n7265 ^ n7187 ^ 1'b0 ;
  assign n39619 = ( n10253 & n39617 ) | ( n10253 & n39618 ) | ( n39617 & n39618 ) ;
  assign n39620 = ~n177 & n738 ;
  assign n39621 = n2836 & n39620 ;
  assign n39622 = n3897 | n39621 ;
  assign n39623 = n27000 | n39622 ;
  assign n39624 = n15868 | n39623 ;
  assign n39625 = n26561 | n32238 ;
  assign n39626 = n20282 ^ n17282 ^ 1'b0 ;
  assign n39627 = n17875 ^ n8260 ^ 1'b0 ;
  assign n39628 = n14506 | n39627 ;
  assign n39629 = n39628 ^ n4740 ^ 1'b0 ;
  assign n39630 = ( n7354 & n16910 ) | ( n7354 & n37799 ) | ( n16910 & n37799 ) ;
  assign n39631 = n7481 | n21264 ;
  assign n39632 = ( n4977 & n6269 ) | ( n4977 & ~n39631 ) | ( n6269 & ~n39631 ) ;
  assign n39633 = n5202 & n18811 ;
  assign n39634 = ( n7086 & ~n25933 ) | ( n7086 & n39633 ) | ( ~n25933 & n39633 ) ;
  assign n39635 = n19074 & n20812 ;
  assign n39636 = n4685 & ~n12436 ;
  assign n39637 = ~n17197 & n39636 ;
  assign n39638 = n36504 ^ n26791 ^ 1'b0 ;
  assign n39639 = ~n12225 & n39638 ;
  assign n39640 = n14831 ^ n13032 ^ 1'b0 ;
  assign n39641 = ( ~n8367 & n10790 ) | ( ~n8367 & n39640 ) | ( n10790 & n39640 ) ;
  assign n39643 = n4897 & ~n11487 ;
  assign n39644 = n21683 & n39643 ;
  assign n39642 = n16705 ^ n2008 ^ n1204 ;
  assign n39645 = n39644 ^ n39642 ^ 1'b0 ;
  assign n39646 = ~n39641 & n39645 ;
  assign n39647 = n27022 ^ n13343 ^ 1'b0 ;
  assign n39648 = n26450 | n39647 ;
  assign n39649 = n39646 & ~n39648 ;
  assign n39650 = n11386 | n12442 ;
  assign n39651 = n39650 ^ n3844 ^ 1'b0 ;
  assign n39652 = n9785 | n23983 ;
  assign n39653 = n28543 & n32801 ;
  assign n39654 = n39653 ^ n5044 ^ 1'b0 ;
  assign n39655 = ( n9955 & n18484 ) | ( n9955 & n39654 ) | ( n18484 & n39654 ) ;
  assign n39656 = ~n8449 & n39655 ;
  assign n39657 = n39656 ^ n5301 ^ 1'b0 ;
  assign n39658 = ~n10129 & n31718 ;
  assign n39659 = n39658 ^ n18268 ^ 1'b0 ;
  assign n39660 = ~n9005 & n22515 ;
  assign n39661 = n39660 ^ n31507 ^ 1'b0 ;
  assign n39662 = n5047 & n32540 ;
  assign n39663 = n39662 ^ n30227 ^ 1'b0 ;
  assign n39664 = ~n27921 & n36594 ;
  assign n39665 = n39663 & n39664 ;
  assign n39666 = n33638 ^ n8942 ^ 1'b0 ;
  assign n39667 = n3737 | n6590 ;
  assign n39668 = ( n481 & n5978 ) | ( n481 & n39667 ) | ( n5978 & n39667 ) ;
  assign n39669 = n16149 ^ n1532 ^ 1'b0 ;
  assign n39670 = n19883 & n39669 ;
  assign n39671 = n12311 & ~n36753 ;
  assign n39672 = n39670 | n39671 ;
  assign n39673 = n29634 ^ n28410 ^ 1'b0 ;
  assign n39674 = n36886 | n39673 ;
  assign n39675 = n12963 ^ n8010 ^ 1'b0 ;
  assign n39676 = n39675 ^ n18619 ^ n13443 ;
  assign n39677 = n39676 ^ n25611 ^ n17951 ;
  assign n39678 = n16500 & ~n21424 ;
  assign n39679 = n13021 & n39678 ;
  assign n39680 = n28394 ^ n15823 ^ n14748 ;
  assign n39681 = n18719 ^ n13752 ^ 1'b0 ;
  assign n39682 = n28511 | n39681 ;
  assign n39683 = ( n22016 & n39680 ) | ( n22016 & n39682 ) | ( n39680 & n39682 ) ;
  assign n39684 = n28462 | n32358 ;
  assign n39685 = n39684 ^ n24041 ^ 1'b0 ;
  assign n39686 = n14585 & ~n39685 ;
  assign n39687 = ~n10743 & n39686 ;
  assign n39688 = ~n11058 & n12708 ;
  assign n39689 = n15341 & n39688 ;
  assign n39690 = n39689 ^ n1888 ^ 1'b0 ;
  assign n39691 = n35355 ^ n20612 ^ 1'b0 ;
  assign n39692 = n39690 & ~n39691 ;
  assign n39693 = n9438 & ~n35312 ;
  assign n39694 = n15672 | n26837 ;
  assign n39695 = n39694 ^ n7906 ^ 1'b0 ;
  assign n39696 = n39695 ^ n14752 ^ 1'b0 ;
  assign n39697 = n46 & n39696 ;
  assign n39698 = ~n12053 & n26167 ;
  assign n39699 = n7545 & ~n39698 ;
  assign n39700 = ~n9039 & n20971 ;
  assign n39701 = ~n32649 & n35521 ;
  assign n39702 = n39701 ^ n1988 ^ 1'b0 ;
  assign n39703 = n31065 & n39702 ;
  assign n39704 = ~n3732 & n39703 ;
  assign n39705 = ( n8655 & n16756 ) | ( n8655 & ~n25268 ) | ( n16756 & ~n25268 ) ;
  assign n39706 = n34371 & ~n39705 ;
  assign n39707 = n39706 ^ n572 ^ 1'b0 ;
  assign n39708 = n9061 ^ n2859 ^ 1'b0 ;
  assign n39710 = n23521 ^ n5751 ^ 1'b0 ;
  assign n39709 = n4652 ^ n3408 ^ 1'b0 ;
  assign n39711 = n39710 ^ n39709 ^ n30182 ;
  assign n39712 = n6676 ^ n4977 ^ 1'b0 ;
  assign n39713 = ~n408 & n39712 ;
  assign n39714 = n5021 & ~n39713 ;
  assign n39715 = n39714 ^ n20849 ^ 1'b0 ;
  assign n39716 = ~n39711 & n39715 ;
  assign n39717 = n7650 & n21414 ;
  assign n39719 = n442 & n35057 ;
  assign n39718 = n1442 | n18479 ;
  assign n39720 = n39719 ^ n39718 ^ 1'b0 ;
  assign n39721 = n39720 ^ n8816 ^ n7898 ;
  assign n39725 = n28480 ^ n18927 ^ n177 ;
  assign n39722 = ~n2004 & n29447 ;
  assign n39723 = n39722 ^ n13451 ^ 1'b0 ;
  assign n39724 = n26437 & n39723 ;
  assign n39726 = n39725 ^ n39724 ^ n15359 ;
  assign n39727 = n9399 ^ n63 ^ 1'b0 ;
  assign n39728 = n39727 ^ n16739 ^ 1'b0 ;
  assign n39730 = n5935 & ~n16643 ;
  assign n39731 = n39730 ^ n14148 ^ 1'b0 ;
  assign n39729 = n856 & ~n16934 ;
  assign n39732 = n39731 ^ n39729 ^ 1'b0 ;
  assign n39733 = n14047 ^ n63 ^ 1'b0 ;
  assign n39734 = ~n5557 & n11090 ;
  assign n39735 = ~n9372 & n39734 ;
  assign n39736 = n39735 ^ n4605 ^ 1'b0 ;
  assign n39737 = n39733 & n39736 ;
  assign n39738 = n19509 ^ n12261 ^ n7768 ;
  assign n39739 = n39738 ^ n4345 ^ n2835 ;
  assign n39740 = n2251 & n2289 ;
  assign n39741 = n39740 ^ n12327 ^ 1'b0 ;
  assign n39742 = n4685 & n39741 ;
  assign n39743 = n34693 ^ n5392 ^ 1'b0 ;
  assign n39744 = n15788 ^ n4878 ^ 1'b0 ;
  assign n39745 = n39743 & n39744 ;
  assign n39746 = n13538 & ~n16176 ;
  assign n39747 = n9827 ^ n5840 ^ 1'b0 ;
  assign n39748 = ~n17413 & n39747 ;
  assign n39749 = n1962 & ~n4627 ;
  assign n39750 = n39749 ^ n38831 ^ 1'b0 ;
  assign n39751 = n16106 & ~n26458 ;
  assign n39752 = n39751 ^ n14916 ^ n10094 ;
  assign n39753 = n39752 ^ n10643 ^ 1'b0 ;
  assign n39754 = ~n28290 & n39753 ;
  assign n39755 = ~n3769 & n22626 ;
  assign n39756 = n9141 & n39755 ;
  assign n39757 = n6487 & n23443 ;
  assign n39758 = n39757 ^ n39237 ^ n37342 ;
  assign n39759 = n16513 | n39758 ;
  assign n39760 = n39759 ^ n3274 ^ 1'b0 ;
  assign n39761 = n39760 ^ n22052 ^ n7317 ;
  assign n39762 = n21691 & n39761 ;
  assign n39763 = ( n321 & ~n11593 ) | ( n321 & n32580 ) | ( ~n11593 & n32580 ) ;
  assign n39764 = n35202 ^ n12164 ^ 1'b0 ;
  assign n39765 = ( n18662 & n26712 ) | ( n18662 & n39764 ) | ( n26712 & n39764 ) ;
  assign n39766 = n963 & n10784 ;
  assign n39767 = ~n963 & n39766 ;
  assign n39768 = n8490 & n10784 ;
  assign n39769 = ~n8490 & n39768 ;
  assign n39770 = n4869 & n39769 ;
  assign n39771 = n39770 ^ n10091 ^ 1'b0 ;
  assign n39772 = n691 | n39771 ;
  assign n39773 = n39767 & ~n39772 ;
  assign n39774 = n11830 & ~n39773 ;
  assign n39775 = n39773 & n39774 ;
  assign n39776 = n3308 & ~n7490 ;
  assign n39777 = n15876 | n34647 ;
  assign n39778 = n28177 | n39777 ;
  assign n39779 = n4729 | n13251 ;
  assign n39780 = ~n9539 & n14755 ;
  assign n39781 = n12698 ^ n6021 ^ 1'b0 ;
  assign n39782 = n15805 & ~n39781 ;
  assign n39783 = ~n1319 & n39782 ;
  assign n39784 = n1295 & n16643 ;
  assign n39785 = n26802 ^ n11925 ^ n3059 ;
  assign n39786 = n22790 | n32315 ;
  assign n39787 = n601 & ~n2883 ;
  assign n39788 = n39787 ^ n39708 ^ 1'b0 ;
  assign n39789 = n11656 ^ n1185 ^ 1'b0 ;
  assign n39790 = ( ~n15987 & n28080 ) | ( ~n15987 & n38311 ) | ( n28080 & n38311 ) ;
  assign n39791 = n36599 ^ n28592 ^ n17742 ;
  assign n39792 = n6853 & ~n18883 ;
  assign n39793 = n39792 ^ n25591 ^ 1'b0 ;
  assign n39794 = n5374 | n24392 ;
  assign n39795 = n39794 ^ n24356 ^ 1'b0 ;
  assign n39796 = n5272 & ~n5342 ;
  assign n39797 = ~n2039 & n39796 ;
  assign n39798 = n39797 ^ n34813 ^ n25446 ;
  assign n39799 = n25787 | n39798 ;
  assign n39800 = n11581 & ~n39799 ;
  assign n39801 = n31129 ^ n10105 ^ 1'b0 ;
  assign n39802 = ~n23392 & n39801 ;
  assign n39803 = ~n7510 & n9736 ;
  assign n39804 = n34485 ^ n13041 ^ 1'b0 ;
  assign n39805 = n32078 ^ n2919 ^ 1'b0 ;
  assign n39806 = n13642 & n39805 ;
  assign n39807 = ~n14188 & n36661 ;
  assign n39808 = n39807 ^ n35536 ^ 1'b0 ;
  assign n39809 = n10288 & ~n39808 ;
  assign n39810 = ~n17064 & n39809 ;
  assign n39811 = n32347 & n39810 ;
  assign n39812 = n4750 & ~n11093 ;
  assign n39813 = n38783 & ~n39812 ;
  assign n39814 = n2357 & n26286 ;
  assign n39815 = n39814 ^ n7494 ^ n771 ;
  assign n39816 = n6875 | n31315 ;
  assign n39817 = n23118 ^ n225 ^ 1'b0 ;
  assign n39818 = n12058 & ~n17338 ;
  assign n39819 = n39818 ^ n6275 ^ 1'b0 ;
  assign n39822 = n3201 ^ x10 ^ 1'b0 ;
  assign n39823 = n26888 & ~n39822 ;
  assign n39824 = n39823 ^ n36038 ^ 1'b0 ;
  assign n39825 = n39824 ^ n14204 ^ 1'b0 ;
  assign n39826 = n17173 & ~n39825 ;
  assign n39820 = ~n3501 & n11032 ;
  assign n39821 = n39820 ^ n27392 ^ 1'b0 ;
  assign n39827 = n39826 ^ n39821 ^ n1891 ;
  assign n39828 = n18929 ^ n12801 ^ n935 ;
  assign n39829 = n16637 ^ n3786 ^ 1'b0 ;
  assign n39830 = n7016 & n39829 ;
  assign n39831 = n18117 ^ n6970 ^ n2147 ;
  assign n39832 = n20659 & ~n39831 ;
  assign n39833 = n39832 ^ n14315 ^ n1188 ;
  assign n39834 = n3698 | n39833 ;
  assign n39835 = n39834 ^ n9658 ^ 1'b0 ;
  assign n39836 = n39432 ^ n12277 ^ 1'b0 ;
  assign n39837 = n39495 & ~n39836 ;
  assign n39838 = n2266 & n6801 ;
  assign n39839 = n39838 ^ n19170 ^ 1'b0 ;
  assign n39840 = ~n48 & n39839 ;
  assign n39845 = n31005 ^ n2476 ^ 1'b0 ;
  assign n39843 = n9700 ^ n8664 ^ 1'b0 ;
  assign n39844 = n37677 | n39843 ;
  assign n39846 = n39845 ^ n39844 ^ 1'b0 ;
  assign n39841 = n12348 & n31694 ;
  assign n39842 = ~n23501 & n39841 ;
  assign n39847 = n39846 ^ n39842 ^ 1'b0 ;
  assign n39848 = n25128 ^ n791 ^ 1'b0 ;
  assign n39849 = n36417 | n39848 ;
  assign n39850 = ~n4383 & n22013 ;
  assign n39851 = n37 & ~n7947 ;
  assign n39852 = ~n5359 & n39851 ;
  assign n39853 = n12461 & ~n39852 ;
  assign n39854 = n6020 & n39853 ;
  assign n39855 = n33409 ^ n20972 ^ n11009 ;
  assign n39858 = n3321 & ~n12036 ;
  assign n39856 = n8691 ^ n4281 ^ 1'b0 ;
  assign n39857 = n12076 & ~n39856 ;
  assign n39859 = n39858 ^ n39857 ^ 1'b0 ;
  assign n39860 = n1296 | n10587 ;
  assign n39861 = ( n30729 & n33416 ) | ( n30729 & n39860 ) | ( n33416 & n39860 ) ;
  assign n39862 = ~n9473 & n26740 ;
  assign n39863 = n39862 ^ n18683 ^ 1'b0 ;
  assign n39864 = n6569 | n9573 ;
  assign n39865 = n20070 & ~n39864 ;
  assign n39866 = ( ~n13051 & n14008 ) | ( ~n13051 & n39865 ) | ( n14008 & n39865 ) ;
  assign n39867 = ( n10883 & ~n24505 ) | ( n10883 & n35029 ) | ( ~n24505 & n35029 ) ;
  assign n39868 = n2995 & ~n18268 ;
  assign n39869 = ~n2320 & n13818 ;
  assign n39870 = n39869 ^ n36194 ^ 1'b0 ;
  assign n39871 = ( ~n3191 & n27143 ) | ( ~n3191 & n39870 ) | ( n27143 & n39870 ) ;
  assign n39872 = ~n10814 & n12409 ;
  assign n39873 = n3035 & n10422 ;
  assign n39874 = n20311 & n39873 ;
  assign n39875 = ~n21596 & n39874 ;
  assign n39876 = n23221 ^ n18132 ^ 1'b0 ;
  assign n39877 = n39876 ^ n3682 ^ n3377 ;
  assign n39878 = n9146 & n22641 ;
  assign n39879 = n39878 ^ n28593 ^ 1'b0 ;
  assign n39880 = ~n181 & n39879 ;
  assign n39881 = n4102 & ~n9020 ;
  assign n39882 = n19753 ^ n15744 ^ 1'b0 ;
  assign n39883 = n11374 & n39882 ;
  assign n39884 = n4685 & n39883 ;
  assign n39885 = ~n39881 & n39884 ;
  assign n39886 = n9416 ^ n6134 ^ 1'b0 ;
  assign n39887 = n21943 | n25995 ;
  assign n39888 = n39887 ^ n453 ^ 1'b0 ;
  assign n39889 = ~n7962 & n36359 ;
  assign n39890 = ( ~n13579 & n16102 ) | ( ~n13579 & n39889 ) | ( n16102 & n39889 ) ;
  assign n39891 = n18728 ^ n7225 ^ 1'b0 ;
  assign n39892 = n27391 ^ n8608 ^ 1'b0 ;
  assign n39893 = ( n18493 & n21967 ) | ( n18493 & n39892 ) | ( n21967 & n39892 ) ;
  assign n39899 = n24518 ^ n8720 ^ n4142 ;
  assign n39895 = n20200 | n20659 ;
  assign n39896 = n24900 | n39895 ;
  assign n39894 = n3059 | n13107 ;
  assign n39897 = n39896 ^ n39894 ^ 1'b0 ;
  assign n39898 = ~n13684 & n39897 ;
  assign n39900 = n39899 ^ n39898 ^ 1'b0 ;
  assign n39901 = ~n17748 & n39900 ;
  assign n39902 = n11668 & ~n14777 ;
  assign n39903 = n39902 ^ n2012 ^ 1'b0 ;
  assign n39904 = n25610 ^ n19429 ^ 1'b0 ;
  assign n39905 = n22583 ^ n18136 ^ 1'b0 ;
  assign n39906 = n34958 | n39905 ;
  assign n39907 = n592 | n12007 ;
  assign n39908 = n23188 ^ n10943 ^ 1'b0 ;
  assign n39909 = n33189 & ~n39908 ;
  assign n39910 = n3039 | n10440 ;
  assign n39911 = n39910 ^ n10507 ^ 1'b0 ;
  assign n39912 = n2044 | n39911 ;
  assign n39913 = n11870 & ~n39912 ;
  assign n39914 = n39913 ^ n15767 ^ 1'b0 ;
  assign n39915 = n37888 ^ n4072 ^ 1'b0 ;
  assign n39916 = n11120 & n39915 ;
  assign n39917 = n6731 & n27276 ;
  assign n39918 = ~n34972 & n39917 ;
  assign n39919 = ( n24202 & ~n34016 ) | ( n24202 & n39474 ) | ( ~n34016 & n39474 ) ;
  assign n39920 = n20801 ^ n14253 ^ 1'b0 ;
  assign n39921 = n39920 ^ n19657 ^ 1'b0 ;
  assign n39922 = n14570 ^ n9180 ^ n6010 ;
  assign n39923 = n39922 ^ n35505 ^ 1'b0 ;
  assign n39924 = n10368 | n29199 ;
  assign n39925 = n25095 ^ n13514 ^ 1'b0 ;
  assign n39926 = ~n30563 & n39925 ;
  assign n39927 = n9239 ^ n5657 ^ n1116 ;
  assign n39928 = n39927 ^ n2328 ^ n962 ;
  assign n39929 = n13710 ^ n3148 ^ 1'b0 ;
  assign n39930 = n39929 ^ n21532 ^ n18932 ;
  assign n39931 = n3922 & n23128 ;
  assign n39932 = n39931 ^ n9885 ^ 1'b0 ;
  assign n39933 = n31732 & n34089 ;
  assign n39934 = ~n12139 & n39933 ;
  assign n39942 = n11980 & n28749 ;
  assign n39940 = n5502 | n8195 ;
  assign n39937 = n8426 ^ n993 ^ 1'b0 ;
  assign n39935 = n17128 ^ n7133 ^ n2422 ;
  assign n39936 = n12300 | n39935 ;
  assign n39938 = n39937 ^ n39936 ^ 1'b0 ;
  assign n39939 = n23295 & ~n39938 ;
  assign n39941 = n39940 ^ n39939 ^ 1'b0 ;
  assign n39943 = n39942 ^ n39941 ^ 1'b0 ;
  assign n39944 = n26293 ^ n12782 ^ 1'b0 ;
  assign n39945 = n1223 & ~n32961 ;
  assign n39946 = n5199 | n19402 ;
  assign n39947 = ( n4189 & ~n5458 ) | ( n4189 & n39946 ) | ( ~n5458 & n39946 ) ;
  assign n39950 = ~n4915 & n36425 ;
  assign n39951 = ~n9392 & n39950 ;
  assign n39948 = n23787 ^ n22716 ^ 1'b0 ;
  assign n39949 = n26631 & ~n39948 ;
  assign n39952 = n39951 ^ n39949 ^ 1'b0 ;
  assign n39953 = n39952 ^ n15314 ^ 1'b0 ;
  assign n39954 = n24687 | n39953 ;
  assign n39955 = ~n2401 & n39105 ;
  assign n39956 = n35247 | n37616 ;
  assign n39957 = n13533 ^ n1092 ^ 1'b0 ;
  assign n39958 = ( n15353 & n39956 ) | ( n15353 & ~n39957 ) | ( n39956 & ~n39957 ) ;
  assign n39959 = ~n636 & n1300 ;
  assign n39960 = n13832 & n39959 ;
  assign n39961 = ( n6093 & n15801 ) | ( n6093 & n22869 ) | ( n15801 & n22869 ) ;
  assign n39962 = n39961 ^ n26567 ^ 1'b0 ;
  assign n39963 = n12097 & ~n39962 ;
  assign n39964 = ~n9902 & n36266 ;
  assign n39965 = ~n5806 & n24512 ;
  assign n39966 = n15195 ^ n9027 ^ 1'b0 ;
  assign n39967 = n4322 & ~n39966 ;
  assign n39968 = ~n3159 & n13707 ;
  assign n39969 = ~n2623 & n39968 ;
  assign n39970 = n39969 ^ n9015 ^ 1'b0 ;
  assign n39971 = n39970 ^ n18303 ^ 1'b0 ;
  assign n39972 = n7236 ^ n6118 ^ n4318 ;
  assign n39973 = n1761 | n39972 ;
  assign n39974 = ~n15367 & n39973 ;
  assign n39975 = n8913 ^ n6293 ^ 1'b0 ;
  assign n39976 = ~n521 & n39975 ;
  assign n39977 = n39976 ^ n37344 ^ 1'b0 ;
  assign n39978 = n8294 & ~n39977 ;
  assign n39979 = n31697 ^ n21347 ^ 1'b0 ;
  assign n39980 = n11839 & ~n39979 ;
  assign n39981 = n8598 & n39980 ;
  assign n39982 = n37376 ^ n11704 ^ 1'b0 ;
  assign n39983 = n13870 ^ n7558 ^ 1'b0 ;
  assign n39984 = ~n34612 & n37912 ;
  assign n39985 = n39984 ^ n23118 ^ 1'b0 ;
  assign n39986 = n3176 | n21528 ;
  assign n39987 = n39986 ^ n16476 ^ 1'b0 ;
  assign n39988 = ~x10 & n1803 ;
  assign n39989 = ( n6289 & ~n23111 ) | ( n6289 & n39988 ) | ( ~n23111 & n39988 ) ;
  assign n39990 = ~n27767 & n39989 ;
  assign n39991 = n39990 ^ n32448 ^ 1'b0 ;
  assign n39992 = n39987 & n39991 ;
  assign n39993 = n16771 | n28235 ;
  assign n39994 = n39993 ^ n19599 ^ 1'b0 ;
  assign n39995 = n4507 & n19848 ;
  assign n39996 = ~n39994 & n39995 ;
  assign n39997 = ( n2294 & ~n9290 ) | ( n2294 & n9503 ) | ( ~n9290 & n9503 ) ;
  assign n39998 = n2190 & n39997 ;
  assign n39999 = n24266 & ~n39998 ;
  assign n40000 = n10955 & n39999 ;
  assign n40001 = n24715 | n31401 ;
  assign n40002 = n29479 ^ n20902 ^ n5044 ;
  assign n40003 = n5153 | n5233 ;
  assign n40004 = n40003 ^ n401 ^ 1'b0 ;
  assign n40005 = n31052 | n40004 ;
  assign n40006 = ~n8806 & n14067 ;
  assign n40007 = ~n6682 & n40006 ;
  assign n40008 = n40007 ^ n32576 ^ 1'b0 ;
  assign n40009 = n40008 ^ n7056 ^ 1'b0 ;
  assign n40010 = x10 & n40009 ;
  assign n40011 = n6613 & n40010 ;
  assign n40012 = n11402 ^ n10108 ^ 1'b0 ;
  assign n40013 = ~n4341 & n40012 ;
  assign n40014 = n40013 ^ n25511 ^ 1'b0 ;
  assign n40015 = n40014 ^ n10292 ^ 1'b0 ;
  assign n40016 = n4674 | n28986 ;
  assign n40017 = n40016 ^ n14855 ^ 1'b0 ;
  assign n40018 = n10263 & ~n40017 ;
  assign n40019 = n32133 & ~n40018 ;
  assign n40020 = n9666 | n35202 ;
  assign n40021 = n20227 ^ n14951 ^ 1'b0 ;
  assign n40022 = ~n18855 & n40021 ;
  assign n40023 = n40022 ^ n34271 ^ 1'b0 ;
  assign n40024 = ~n40020 & n40023 ;
  assign n40025 = n2983 | n34966 ;
  assign n40026 = ~n2813 & n40025 ;
  assign n40027 = n40026 ^ n16556 ^ 1'b0 ;
  assign n40028 = n10731 & n40027 ;
  assign n40029 = n40028 ^ n17457 ^ 1'b0 ;
  assign n40030 = n40029 ^ n7363 ^ 1'b0 ;
  assign n40031 = n9599 & n40030 ;
  assign n40032 = n40031 ^ n4099 ^ 1'b0 ;
  assign n40033 = ~n4920 & n12810 ;
  assign n40034 = n31021 & n40033 ;
  assign n40035 = ~n21701 & n40034 ;
  assign n40036 = n1658 | n10907 ;
  assign n40037 = n40036 ^ n22532 ^ 1'b0 ;
  assign n40038 = n40037 ^ n22886 ^ 1'b0 ;
  assign n40039 = n16122 & ~n31096 ;
  assign n40040 = n12036 ^ n2233 ^ 1'b0 ;
  assign n40041 = n14790 ^ n6595 ^ 1'b0 ;
  assign n40042 = ~n40040 & n40041 ;
  assign n40043 = ~n40039 & n40042 ;
  assign n40044 = ( ~n4591 & n20756 ) | ( ~n4591 & n31621 ) | ( n20756 & n31621 ) ;
  assign n40045 = n6055 & n40044 ;
  assign n40046 = n3155 & ~n4446 ;
  assign n40047 = n875 & n40046 ;
  assign n40048 = n20137 & ~n40047 ;
  assign n40049 = ~n39780 & n40048 ;
  assign n40050 = n9049 & n29534 ;
  assign n40051 = n5156 & n40050 ;
  assign n40052 = ( n1400 & n6412 ) | ( n1400 & n9360 ) | ( n6412 & n9360 ) ;
  assign n40053 = ( n1962 & n2563 ) | ( n1962 & ~n23580 ) | ( n2563 & ~n23580 ) ;
  assign n40054 = n502 & n16820 ;
  assign n40055 = n36738 & n40054 ;
  assign n40056 = n40055 ^ n25313 ^ 1'b0 ;
  assign n40057 = n35727 ^ n16066 ^ 1'b0 ;
  assign n40058 = n32133 | n40057 ;
  assign n40059 = n475 & n36656 ;
  assign n40060 = n40059 ^ n36339 ^ 1'b0 ;
  assign n40061 = n4165 & n21663 ;
  assign n40062 = n22369 ^ n9373 ^ 1'b0 ;
  assign n40066 = n28090 ^ n14771 ^ 1'b0 ;
  assign n40067 = n15138 | n40066 ;
  assign n40065 = n35934 ^ n29940 ^ 1'b0 ;
  assign n40068 = n40067 ^ n40065 ^ n14421 ;
  assign n40063 = n2787 | n3961 ;
  assign n40064 = n27441 | n40063 ;
  assign n40069 = n40068 ^ n40064 ^ 1'b0 ;
  assign n40070 = ~n31953 & n40069 ;
  assign n40071 = n8135 & n12484 ;
  assign n40072 = n13064 | n31879 ;
  assign n40073 = n39962 ^ n729 ^ 1'b0 ;
  assign n40074 = n40073 ^ n32882 ^ 1'b0 ;
  assign n40075 = n7167 | n40074 ;
  assign n40076 = n6939 | n18736 ;
  assign n40077 = n40076 ^ n11723 ^ 1'b0 ;
  assign n40078 = n37021 & n40077 ;
  assign n40079 = ~n1290 & n35774 ;
  assign n40080 = n2485 & n8305 ;
  assign n40081 = n7393 & ~n19683 ;
  assign n40082 = n9687 | n40081 ;
  assign n40083 = ~n13266 & n14011 ;
  assign n40084 = n40083 ^ n35313 ^ 1'b0 ;
  assign n40085 = n10563 & n12212 ;
  assign n40086 = n38319 & n40085 ;
  assign n40087 = n17171 ^ n10578 ^ n4126 ;
  assign n40088 = ~n22562 & n25028 ;
  assign n40089 = ( n631 & ~n28017 ) | ( n631 & n40088 ) | ( ~n28017 & n40088 ) ;
  assign n40090 = n13261 & ~n36828 ;
  assign n40091 = ~n25604 & n40090 ;
  assign n40092 = n18950 & ~n40091 ;
  assign n40093 = n1602 | n5691 ;
  assign n40094 = n5691 & ~n40093 ;
  assign n40095 = n5892 & ~n40094 ;
  assign n40098 = ~n9956 & n11598 ;
  assign n40099 = ~n11598 & n40098 ;
  assign n40100 = n10223 | n13909 ;
  assign n40101 = n10223 & ~n40100 ;
  assign n40102 = ~n1315 & n40101 ;
  assign n40103 = n40099 | n40102 ;
  assign n40104 = n40099 & ~n40103 ;
  assign n40096 = n11500 & ~n25475 ;
  assign n40097 = n40096 ^ n36300 ^ n2552 ;
  assign n40105 = n40104 ^ n40097 ^ 1'b0 ;
  assign n40106 = n40095 | n40105 ;
  assign n40107 = n28643 | n40106 ;
  assign n40108 = ( n4724 & ~n9583 ) | ( n4724 & n10445 ) | ( ~n9583 & n10445 ) ;
  assign n40109 = ( n9889 & n27262 ) | ( n9889 & n40108 ) | ( n27262 & n40108 ) ;
  assign n40110 = ( n1148 & n3119 ) | ( n1148 & ~n35506 ) | ( n3119 & ~n35506 ) ;
  assign n40111 = n14815 ^ n2271 ^ 1'b0 ;
  assign n40112 = n8693 & ~n40111 ;
  assign n40113 = ~n6882 & n40112 ;
  assign n40114 = n8026 & n40113 ;
  assign n40115 = n7640 ^ n1886 ^ 1'b0 ;
  assign n40116 = n6442 & n40115 ;
  assign n40117 = n40116 ^ n33847 ^ n12931 ;
  assign n40118 = n20328 & ~n30456 ;
  assign n40119 = n40118 ^ n21840 ^ 1'b0 ;
  assign n40120 = n3876 ^ n2984 ^ 1'b0 ;
  assign n40121 = n40119 & ~n40120 ;
  assign n40122 = n14132 & ~n40121 ;
  assign n40123 = n28164 & ~n40122 ;
  assign n40124 = n20715 ^ n4417 ^ 1'b0 ;
  assign n40125 = ~n7062 & n16880 ;
  assign n40126 = n40125 ^ n19644 ^ 1'b0 ;
  assign n40127 = n2989 & ~n13520 ;
  assign n40128 = n12683 ^ n435 ^ 1'b0 ;
  assign n40129 = n21723 | n40128 ;
  assign n40130 = ~n2956 & n40129 ;
  assign n40131 = n7017 & ~n9790 ;
  assign n40132 = ~n40130 & n40131 ;
  assign n40133 = n35417 ^ n17746 ^ n14030 ;
  assign n40134 = n33771 ^ n791 ^ n614 ;
  assign n40135 = n9060 | n10090 ;
  assign n40136 = ~n38999 & n40135 ;
  assign n40137 = n15849 ^ n1305 ^ 1'b0 ;
  assign n40138 = n32029 ^ n13650 ^ n7363 ;
  assign n40139 = n40137 & n40138 ;
  assign n40140 = n4817 | n29089 ;
  assign n40142 = n6611 | n13855 ;
  assign n40143 = n40142 ^ n30189 ^ 1'b0 ;
  assign n40141 = n33720 | n37189 ;
  assign n40144 = n40143 ^ n40141 ^ 1'b0 ;
  assign n40145 = ( n25303 & ~n35199 ) | ( n25303 & n40144 ) | ( ~n35199 & n40144 ) ;
  assign n40147 = n115 & n7260 ;
  assign n40148 = ~n10649 & n40147 ;
  assign n40149 = n36286 ^ n769 ^ 1'b0 ;
  assign n40150 = ~n40148 & n40149 ;
  assign n40146 = n11185 ^ n5920 ^ 1'b0 ;
  assign n40151 = n40150 ^ n40146 ^ 1'b0 ;
  assign n40153 = n7022 ^ n5298 ^ 1'b0 ;
  assign n40154 = n5160 & n40153 ;
  assign n40155 = ~n14628 & n40154 ;
  assign n40156 = n40155 ^ n9325 ^ 1'b0 ;
  assign n40157 = ( n6313 & n7859 ) | ( n6313 & n40156 ) | ( n7859 & n40156 ) ;
  assign n40152 = ~n19066 & n23666 ;
  assign n40158 = n40157 ^ n40152 ^ n37516 ;
  assign n40159 = n25232 ^ n22414 ^ 1'b0 ;
  assign n40160 = n35562 ^ n27072 ^ 1'b0 ;
  assign n40161 = n40159 & ~n40160 ;
  assign n40162 = ( n9620 & n12644 ) | ( n9620 & ~n27816 ) | ( n12644 & ~n27816 ) ;
  assign n40163 = ( n3426 & n11438 ) | ( n3426 & n18462 ) | ( n11438 & n18462 ) ;
  assign n40164 = ( n20269 & ~n40162 ) | ( n20269 & n40163 ) | ( ~n40162 & n40163 ) ;
  assign n40166 = n1492 & ~n29331 ;
  assign n40165 = n13267 ^ n5714 ^ 1'b0 ;
  assign n40167 = n40166 ^ n40165 ^ n2580 ;
  assign n40168 = n4436 ^ n791 ^ 1'b0 ;
  assign n40169 = n26519 ^ n12631 ^ 1'b0 ;
  assign n40170 = n10254 | n40169 ;
  assign n40171 = n6868 & ~n12421 ;
  assign n40172 = n4027 | n25291 ;
  assign n40173 = n40171 | n40172 ;
  assign n40174 = n37700 & n39658 ;
  assign n40175 = n40174 ^ n30472 ^ 1'b0 ;
  assign n40176 = n33753 ^ n4110 ^ 1'b0 ;
  assign n40177 = n31415 | n40176 ;
  assign n40178 = n1948 & ~n23869 ;
  assign n40179 = n40178 ^ n29927 ^ 1'b0 ;
  assign n40180 = n29927 ^ n17832 ^ 1'b0 ;
  assign n40181 = n31548 & n40180 ;
  assign n40182 = n33953 ^ n20062 ^ 1'b0 ;
  assign n40183 = n583 & ~n40182 ;
  assign n40184 = n40183 ^ n37972 ^ 1'b0 ;
  assign n40186 = ( n374 & ~n6516 ) | ( n374 & n20429 ) | ( ~n6516 & n20429 ) ;
  assign n40185 = n9275 & ~n11074 ;
  assign n40187 = n40186 ^ n40185 ^ 1'b0 ;
  assign n40188 = ( n5057 & n18730 ) | ( n5057 & n32819 ) | ( n18730 & n32819 ) ;
  assign n40189 = n16652 ^ n6942 ^ 1'b0 ;
  assign n40192 = n515 | n6353 ;
  assign n40193 = n40192 ^ n27439 ^ n17118 ;
  assign n40190 = ( n5324 & n22410 ) | ( n5324 & ~n24817 ) | ( n22410 & ~n24817 ) ;
  assign n40191 = n22198 & ~n40190 ;
  assign n40194 = n40193 ^ n40191 ^ 1'b0 ;
  assign n40195 = n10049 | n21010 ;
  assign n40196 = n40195 ^ n37353 ^ n14957 ;
  assign n40197 = n23697 ^ n15179 ^ 1'b0 ;
  assign n40198 = ( n1400 & ~n34252 ) | ( n1400 & n40197 ) | ( ~n34252 & n40197 ) ;
  assign n40199 = n1343 & n3838 ;
  assign n40200 = n14201 ^ n11410 ^ n10017 ;
  assign n40201 = n40200 ^ n3781 ^ 1'b0 ;
  assign n40202 = n1523 & ~n40201 ;
  assign n40203 = n3669 | n5007 ;
  assign n40204 = n40203 ^ n6516 ^ 1'b0 ;
  assign n40205 = n40124 ^ n19291 ^ 1'b0 ;
  assign n40206 = n11696 & ~n40205 ;
  assign n40207 = ( ~n3866 & n22090 ) | ( ~n3866 & n28079 ) | ( n22090 & n28079 ) ;
  assign n40208 = n5391 ^ n4134 ^ 1'b0 ;
  assign n40209 = n40208 ^ n9489 ^ 1'b0 ;
  assign n40210 = n19079 ^ n12874 ^ 1'b0 ;
  assign n40211 = n25022 & n40210 ;
  assign n40212 = ( ~n24444 & n27270 ) | ( ~n24444 & n40211 ) | ( n27270 & n40211 ) ;
  assign n40213 = n40209 | n40212 ;
  assign n40214 = n40213 ^ n30729 ^ 1'b0 ;
  assign n40215 = n101 & ~n4188 ;
  assign n40216 = ~n101 & n40215 ;
  assign n40217 = n5707 & ~n40216 ;
  assign n40218 = ~n5707 & n40217 ;
  assign n40219 = n40218 ^ n17094 ^ 1'b0 ;
  assign n40220 = n40219 ^ n22307 ^ 1'b0 ;
  assign n40221 = n12252 & ~n40220 ;
  assign n40222 = ~n15779 & n18741 ;
  assign n40223 = n12202 & n40222 ;
  assign n40224 = n1426 | n27583 ;
  assign n40231 = n6102 & ~n21770 ;
  assign n40230 = n30812 ^ n10849 ^ n2474 ;
  assign n40225 = n14168 ^ n4053 ^ 1'b0 ;
  assign n40226 = n572 & n40225 ;
  assign n40227 = n6074 ^ n2083 ^ 1'b0 ;
  assign n40228 = n3510 & ~n40227 ;
  assign n40229 = ~n40226 & n40228 ;
  assign n40232 = n40231 ^ n40230 ^ n40229 ;
  assign n40233 = n3874 ^ n1167 ^ 1'b0 ;
  assign n40234 = n40171 & n40233 ;
  assign n40235 = n11017 | n14864 ;
  assign n40236 = ~n1280 & n9218 ;
  assign n40238 = n28203 ^ n23042 ^ 1'b0 ;
  assign n40239 = n10258 | n40238 ;
  assign n40237 = n15912 ^ n7267 ^ 1'b0 ;
  assign n40240 = n40239 ^ n40237 ^ n3892 ;
  assign n40241 = n31328 ^ n21810 ^ 1'b0 ;
  assign n40244 = n22678 & ~n29650 ;
  assign n40242 = n32328 ^ n9704 ^ n5095 ;
  assign n40243 = n20078 & ~n40242 ;
  assign n40245 = n40244 ^ n40243 ^ 1'b0 ;
  assign n40246 = ~n24345 & n25987 ;
  assign n40247 = ~n6648 & n38593 ;
  assign n40248 = n40247 ^ n36762 ^ n26416 ;
  assign n40249 = n2519 & n40248 ;
  assign n40250 = n3365 | n7841 ;
  assign n40251 = n40250 ^ n3923 ^ 1'b0 ;
  assign n40252 = n40251 ^ n31556 ^ 1'b0 ;
  assign n40253 = n38073 ^ n20273 ^ 1'b0 ;
  assign n40254 = n27979 & n40253 ;
  assign n40255 = n5933 & ~n15856 ;
  assign n40256 = n40255 ^ n37977 ^ 1'b0 ;
  assign n40257 = ~n18140 & n29559 ;
  assign n40258 = n20518 ^ n20213 ^ n14766 ;
  assign n40259 = n1393 & ~n40258 ;
  assign n40260 = n40259 ^ n38502 ^ n24123 ;
  assign n40261 = ~n5740 & n10385 ;
  assign n40262 = n40261 ^ n6353 ^ 1'b0 ;
  assign n40263 = n4450 ^ n108 ^ 1'b0 ;
  assign n40264 = n6888 & ~n40263 ;
  assign n40265 = ~n16030 & n40264 ;
  assign n40266 = ~n40262 & n40265 ;
  assign n40267 = ~n122 & n10178 ;
  assign n40268 = ( ~n1948 & n40266 ) | ( ~n1948 & n40267 ) | ( n40266 & n40267 ) ;
  assign n40269 = n40268 ^ n8566 ^ 1'b0 ;
  assign n40270 = n25460 ^ n17465 ^ n13312 ;
  assign n40271 = n37198 & ~n40270 ;
  assign n40272 = n12925 & n40271 ;
  assign n40273 = ( n4769 & n22695 ) | ( n4769 & ~n27540 ) | ( n22695 & ~n27540 ) ;
  assign n40274 = n23481 | n38561 ;
  assign n40275 = n6374 | n40274 ;
  assign n40276 = n15704 | n27032 ;
  assign n40277 = n40275 | n40276 ;
  assign n40278 = n41 & n26500 ;
  assign n40301 = n21140 ^ n23 ^ 1'b0 ;
  assign n40279 = ~n287 & n1674 ;
  assign n40280 = n287 & n40279 ;
  assign n40281 = n121 & ~n3925 ;
  assign n40282 = n40280 & n40281 ;
  assign n40283 = n695 & n1801 ;
  assign n40284 = n40282 & n40283 ;
  assign n40285 = n771 & n1881 ;
  assign n40286 = ~n771 & n40285 ;
  assign n40287 = n6537 & n7279 ;
  assign n40288 = n40286 & n40287 ;
  assign n40289 = n11241 | n40288 ;
  assign n40290 = n40288 & ~n40289 ;
  assign n40291 = n40284 & ~n40290 ;
  assign n40292 = ~n139 & n40291 ;
  assign n40295 = n2412 & n10038 ;
  assign n40296 = ~n2412 & n40295 ;
  assign n40297 = n2094 & n40296 ;
  assign n40293 = n850 & ~n2587 ;
  assign n40294 = n2587 & n40293 ;
  assign n40298 = n40297 ^ n40294 ^ 1'b0 ;
  assign n40299 = ~n40292 & n40298 ;
  assign n40300 = n30977 & n40299 ;
  assign n40302 = n40301 ^ n40300 ^ 1'b0 ;
  assign n40303 = n145 & ~n33488 ;
  assign n40304 = n16739 & n40303 ;
  assign n40305 = ~n31962 & n40304 ;
  assign n40307 = n10253 & ~n19363 ;
  assign n40306 = ~n14307 & n24806 ;
  assign n40308 = n40307 ^ n40306 ^ 1'b0 ;
  assign n40309 = n34467 & ~n40308 ;
  assign n40310 = n6807 & n40309 ;
  assign n40311 = n11126 ^ n8359 ^ 1'b0 ;
  assign n40313 = n22678 ^ n15197 ^ 1'b0 ;
  assign n40312 = n91 & n18095 ;
  assign n40314 = n40313 ^ n40312 ^ 1'b0 ;
  assign n40315 = n35188 & n40314 ;
  assign n40316 = n40315 ^ n7702 ^ 1'b0 ;
  assign n40317 = n1533 | n11495 ;
  assign n40318 = n32963 & n40317 ;
  assign n40319 = n9631 & n12281 ;
  assign n40320 = n13960 ^ n10267 ^ n411 ;
  assign n40321 = ( ~n12413 & n18039 ) | ( ~n12413 & n40320 ) | ( n18039 & n40320 ) ;
  assign n40322 = n40321 ^ n19978 ^ n7133 ;
  assign n40323 = ( n23920 & n25888 ) | ( n23920 & n40322 ) | ( n25888 & n40322 ) ;
  assign n40324 = n24970 | n25934 ;
  assign n40325 = n9565 | n18025 ;
  assign n40326 = n13125 & ~n19420 ;
  assign n40327 = ~n40325 & n40326 ;
  assign n40329 = n12373 ^ n3642 ^ 1'b0 ;
  assign n40328 = ~n23573 & n31455 ;
  assign n40330 = n40329 ^ n40328 ^ 1'b0 ;
  assign n40331 = ~n13362 & n40330 ;
  assign n40332 = n32473 ^ n14440 ^ 1'b0 ;
  assign n40333 = n6576 & n40332 ;
  assign n40334 = n5373 & n40333 ;
  assign n40338 = n17860 & ~n26447 ;
  assign n40339 = n40338 ^ n575 ^ 1'b0 ;
  assign n40335 = n4183 & n34424 ;
  assign n40336 = ~n6458 & n40335 ;
  assign n40337 = n1318 | n40336 ;
  assign n40340 = n40339 ^ n40337 ^ 1'b0 ;
  assign n40341 = ~n8365 & n25706 ;
  assign n40342 = ~n23514 & n40341 ;
  assign n40343 = n20529 & ~n32245 ;
  assign n40344 = n17494 ^ n1120 ^ 1'b0 ;
  assign n40345 = ~n17828 & n40344 ;
  assign n40346 = n40345 ^ n24340 ^ 1'b0 ;
  assign n40347 = n3234 ^ n141 ^ n113 ;
  assign n40348 = n4351 | n40347 ;
  assign n40353 = n11500 | n13023 ;
  assign n40354 = n18886 | n40353 ;
  assign n40349 = n15197 ^ n401 ^ 1'b0 ;
  assign n40350 = n10579 ^ n7400 ^ 1'b0 ;
  assign n40351 = n40349 & ~n40350 ;
  assign n40352 = n40351 ^ n17749 ^ n412 ;
  assign n40355 = n40354 ^ n40352 ^ 1'b0 ;
  assign n40356 = n23338 ^ n14360 ^ n11292 ;
  assign n40357 = n40356 ^ n4214 ^ 1'b0 ;
  assign n40358 = ~n29216 & n40357 ;
  assign n40359 = n9238 | n27242 ;
  assign n40360 = n40359 ^ n29693 ^ 1'b0 ;
  assign n40361 = n17795 ^ n8160 ^ 1'b0 ;
  assign n40362 = n10326 & ~n40361 ;
  assign n40363 = ~n8603 & n25994 ;
  assign n40364 = n16231 ^ n15476 ^ n12112 ;
  assign n40365 = n40363 & ~n40364 ;
  assign n40367 = n792 ^ n733 ^ 1'b0 ;
  assign n40368 = n5867 ^ n4305 ^ 1'b0 ;
  assign n40369 = n40367 | n40368 ;
  assign n40366 = n20671 & ~n33944 ;
  assign n40370 = n40369 ^ n40366 ^ 1'b0 ;
  assign n40371 = ~n11420 & n19070 ;
  assign n40372 = n40371 ^ n5549 ^ 1'b0 ;
  assign n40373 = n40372 ^ n21512 ^ 1'b0 ;
  assign n40375 = n11680 | n20628 ;
  assign n40376 = n40375 ^ n7053 ^ 1'b0 ;
  assign n40374 = n2287 & ~n14578 ;
  assign n40377 = n40376 ^ n40374 ^ n35969 ;
  assign n40378 = n9264 ^ n8490 ^ n2097 ;
  assign n40379 = n14177 & n40378 ;
  assign n40380 = n13817 & n40379 ;
  assign n40381 = n40380 ^ n10234 ^ 1'b0 ;
  assign n40382 = n9962 & ~n15569 ;
  assign n40383 = n24268 & ~n29084 ;
  assign n40384 = ( n4301 & n17840 ) | ( n4301 & n36752 ) | ( n17840 & n36752 ) ;
  assign n40385 = n19987 ^ n17974 ^ n5924 ;
  assign n40386 = n9118 | n32919 ;
  assign n40387 = n4185 | n40386 ;
  assign n40388 = n14745 ^ n5521 ^ n308 ;
  assign n40389 = n40388 ^ n3252 ^ 1'b0 ;
  assign n40390 = n11601 ^ n1734 ^ 1'b0 ;
  assign n40391 = ~n7779 & n40390 ;
  assign n40392 = ( n5930 & n16259 ) | ( n5930 & ~n40391 ) | ( n16259 & ~n40391 ) ;
  assign n40394 = n14547 ^ n13133 ^ 1'b0 ;
  assign n40393 = n6657 & ~n8465 ;
  assign n40395 = n40394 ^ n40393 ^ 1'b0 ;
  assign n40396 = ~n24834 & n29769 ;
  assign n40397 = n16485 ^ n7970 ^ 1'b0 ;
  assign n40398 = ~n14048 & n40397 ;
  assign n40399 = n23539 ^ n10219 ^ n2667 ;
  assign n40400 = n40399 ^ n11713 ^ 1'b0 ;
  assign n40401 = n37387 & n40400 ;
  assign n40402 = n7115 ^ n684 ^ 1'b0 ;
  assign n40403 = n11925 ^ n2362 ^ 1'b0 ;
  assign n40404 = n2246 | n40403 ;
  assign n40405 = n15029 ^ n13507 ^ n7925 ;
  assign n40406 = n37523 ^ n31935 ^ n19320 ;
  assign n40407 = n31617 ^ n14960 ^ 1'b0 ;
  assign n40408 = n24237 | n40407 ;
  assign n40409 = n19478 ^ n9959 ^ 1'b0 ;
  assign n40410 = n23835 & ~n40409 ;
  assign n40411 = n12987 ^ n3034 ^ 1'b0 ;
  assign n40412 = n40410 & n40411 ;
  assign n40413 = ~n14363 & n40412 ;
  assign n40414 = n7594 & n8523 ;
  assign n40415 = n13363 ^ n6149 ^ 1'b0 ;
  assign n40416 = n7267 & ~n10223 ;
  assign n40417 = n40415 & n40416 ;
  assign n40418 = n8356 & ~n40417 ;
  assign n40419 = ~n7448 & n10012 ;
  assign n40420 = n12541 & n34542 ;
  assign n40421 = n32809 ^ n18876 ^ n15461 ;
  assign n40422 = n15892 | n38061 ;
  assign n40423 = ( n18514 & ~n26581 ) | ( n18514 & n26589 ) | ( ~n26581 & n26589 ) ;
  assign n40424 = n5135 & n40423 ;
  assign n40425 = n37884 ^ n28044 ^ 1'b0 ;
  assign n40426 = n12603 | n18513 ;
  assign n40427 = ~n14292 & n16159 ;
  assign n40428 = n527 & ~n40427 ;
  assign n40429 = ~n5102 & n40428 ;
  assign n40430 = ~n9055 & n40277 ;
  assign n40431 = n40430 ^ n680 ^ 1'b0 ;
  assign n40432 = n34825 ^ n17245 ^ 1'b0 ;
  assign n40433 = n1842 ^ n588 ^ 1'b0 ;
  assign n40434 = n4701 & n40433 ;
  assign n40435 = n1993 | n17037 ;
  assign n40436 = n24785 | n40435 ;
  assign n40437 = n3085 | n23962 ;
  assign n40438 = n8550 & ~n40437 ;
  assign n40439 = n40436 & ~n40438 ;
  assign n40440 = n23204 & n40439 ;
  assign n40441 = ( n7363 & ~n21817 ) | ( n7363 & n40440 ) | ( ~n21817 & n40440 ) ;
  assign n40442 = ~n2992 & n18509 ;
  assign n40443 = n29476 ^ n27668 ^ 1'b0 ;
  assign n40444 = n25633 & n40443 ;
  assign n40445 = n15626 & n25482 ;
  assign n40446 = n40445 ^ n3647 ^ 1'b0 ;
  assign n40447 = ( n12202 & n14886 ) | ( n12202 & n40446 ) | ( n14886 & n40446 ) ;
  assign n40448 = n10103 | n38588 ;
  assign n40449 = n40448 ^ n14414 ^ n8811 ;
  assign n40450 = n15051 ^ n4930 ^ 1'b0 ;
  assign n40451 = ( n11264 & n12622 ) | ( n11264 & ~n33466 ) | ( n12622 & ~n33466 ) ;
  assign n40452 = n3644 & ~n3911 ;
  assign n40453 = ~n40451 & n40452 ;
  assign n40454 = n5342 ^ n411 ^ 1'b0 ;
  assign n40455 = ~n23942 & n40454 ;
  assign n40456 = ~n18036 & n40455 ;
  assign n40457 = n28765 & ~n40456 ;
  assign n40459 = ( ~n7565 & n8597 ) | ( ~n7565 & n9565 ) | ( n8597 & n9565 ) ;
  assign n40458 = n19087 ^ n7940 ^ 1'b0 ;
  assign n40460 = n40459 ^ n40458 ^ n13993 ;
  assign n40461 = ~n18528 & n22556 ;
  assign n40462 = n40461 ^ n10321 ^ 1'b0 ;
  assign n40463 = n22741 & n40462 ;
  assign n40464 = ~n35261 & n40463 ;
  assign n40465 = n24411 ^ n15250 ^ n10553 ;
  assign n40466 = n890 | n19536 ;
  assign n40467 = n19207 | n40466 ;
  assign n40468 = n11159 & n40467 ;
  assign n40469 = n40465 & n40468 ;
  assign n40470 = n8524 & n25755 ;
  assign n40471 = n24978 & n40470 ;
  assign n40472 = n3433 & ~n40471 ;
  assign n40473 = n40472 ^ n10123 ^ 1'b0 ;
  assign n40477 = ~n228 & n22052 ;
  assign n40474 = n17963 ^ n17801 ^ n9863 ;
  assign n40475 = ( n22736 & n25146 ) | ( n22736 & ~n40474 ) | ( n25146 & ~n40474 ) ;
  assign n40476 = n6938 & ~n40475 ;
  assign n40478 = n40477 ^ n40476 ^ 1'b0 ;
  assign n40479 = ~n22495 & n32937 ;
  assign n40480 = n40479 ^ n39090 ^ 1'b0 ;
  assign n40482 = n326 & n13626 ;
  assign n40481 = n6713 & ~n13554 ;
  assign n40483 = n40482 ^ n40481 ^ 1'b0 ;
  assign n40484 = n5279 & n32995 ;
  assign n40485 = n40484 ^ n4540 ^ 1'b0 ;
  assign n40486 = n1922 & ~n11674 ;
  assign n40487 = n8334 | n40486 ;
  assign n40488 = n35592 ^ n17302 ^ 1'b0 ;
  assign n40489 = ~n7284 & n20817 ;
  assign n40490 = n3542 & n40489 ;
  assign n40491 = n38216 & ~n40490 ;
  assign n40492 = n8516 ^ n1000 ^ n319 ;
  assign n40493 = ~n15130 & n40492 ;
  assign n40494 = n20473 ^ n15987 ^ 1'b0 ;
  assign n40495 = ~n3168 & n40494 ;
  assign n40496 = n8365 | n17019 ;
  assign n40497 = n40496 ^ n6135 ^ 1'b0 ;
  assign n40498 = ( n21027 & n28047 ) | ( n21027 & ~n40497 ) | ( n28047 & ~n40497 ) ;
  assign n40499 = n21624 ^ n16793 ^ n7786 ;
  assign n40500 = n6010 | n14881 ;
  assign n40501 = n9227 | n40500 ;
  assign n40502 = n11915 ^ n11063 ^ 1'b0 ;
  assign n40503 = n20099 ^ n14690 ^ n9506 ;
  assign n40504 = n19510 ^ n7163 ^ n1339 ;
  assign n40505 = n8782 & ~n16489 ;
  assign n40506 = n40505 ^ n213 ^ 1'b0 ;
  assign n40507 = n40504 & n40506 ;
  assign n40508 = n40507 ^ n3214 ^ 1'b0 ;
  assign n40509 = n27350 ^ n16647 ^ 1'b0 ;
  assign n40510 = ~n5570 & n40509 ;
  assign n40511 = n40155 ^ n26332 ^ 1'b0 ;
  assign n40512 = n31055 ^ n18709 ^ 1'b0 ;
  assign n40513 = n17559 ^ n2991 ^ 1'b0 ;
  assign n40514 = n6353 | n40513 ;
  assign n40515 = ~n7977 & n19235 ;
  assign n40519 = n4189 | n12209 ;
  assign n40516 = n519 & ~n26143 ;
  assign n40517 = n18669 ^ n8220 ^ n7251 ;
  assign n40518 = n40516 & n40517 ;
  assign n40520 = n40519 ^ n40518 ^ 1'b0 ;
  assign n40521 = n25672 | n36890 ;
  assign n40522 = n4207 | n4232 ;
  assign n40523 = n40522 ^ n28805 ^ 1'b0 ;
  assign n40524 = n27064 ^ n15799 ^ 1'b0 ;
  assign n40525 = n40523 & ~n40524 ;
  assign n40526 = n18896 & n29685 ;
  assign n40527 = ~n40525 & n40526 ;
  assign n40528 = n2754 & ~n21492 ;
  assign n40529 = n40528 ^ n2560 ^ 1'b0 ;
  assign n40530 = ~n4079 & n33677 ;
  assign n40531 = n40530 ^ n12635 ^ 1'b0 ;
  assign n40532 = n7690 & n19354 ;
  assign n40533 = n29663 & n40532 ;
  assign n40535 = n38141 ^ n26426 ^ n867 ;
  assign n40534 = ~n5710 & n9108 ;
  assign n40536 = n40535 ^ n40534 ^ 1'b0 ;
  assign n40537 = n23747 ^ x3 ^ 1'b0 ;
  assign n40538 = n21299 | n40537 ;
  assign n40539 = n25680 & n38051 ;
  assign n40540 = ( n2529 & n19325 ) | ( n2529 & n27024 ) | ( n19325 & n27024 ) ;
  assign n40541 = n35526 & n40540 ;
  assign n40542 = n40541 ^ n5554 ^ 1'b0 ;
  assign n40543 = n27009 & ~n37710 ;
  assign n40544 = n24421 ^ n16454 ^ 1'b0 ;
  assign n40545 = n3076 & n40544 ;
  assign n40546 = n25995 ^ n1553 ^ 1'b0 ;
  assign n40547 = n10470 | n12541 ;
  assign n40548 = n16319 ^ n6753 ^ n6564 ;
  assign n40549 = n40548 ^ n13376 ^ n3330 ;
  assign n40550 = ( ~n15607 & n35426 ) | ( ~n15607 & n35635 ) | ( n35426 & n35635 ) ;
  assign n40551 = n3959 & n7021 ;
  assign n40552 = n18620 & ~n40551 ;
  assign n40553 = n27882 ^ n16124 ^ n2397 ;
  assign n40554 = n3912 & ~n40553 ;
  assign n40555 = n16264 | n21723 ;
  assign n40556 = n40555 ^ n22818 ^ 1'b0 ;
  assign n40557 = n34944 & n40556 ;
  assign n40558 = n18124 & n40557 ;
  assign n40559 = n10977 & ~n15324 ;
  assign n40560 = n40559 ^ n17564 ^ 1'b0 ;
  assign n40561 = n33760 ^ n25539 ^ 1'b0 ;
  assign n40562 = n38528 & n40561 ;
  assign n40563 = ~n40560 & n40562 ;
  assign n40564 = n2374 & ~n2657 ;
  assign n40565 = n40564 ^ n4769 ^ 1'b0 ;
  assign n40566 = n10646 & ~n19850 ;
  assign n40567 = ~n8242 & n40566 ;
  assign n40568 = n816 & ~n11611 ;
  assign n40569 = n39150 & n40568 ;
  assign n40570 = n26820 ^ n7852 ^ 1'b0 ;
  assign n40571 = n5420 ^ n1592 ^ 1'b0 ;
  assign n40572 = n6016 | n40571 ;
  assign n40573 = n40572 ^ n31516 ^ 1'b0 ;
  assign n40574 = n40570 & n40573 ;
  assign n40575 = n9737 | n10044 ;
  assign n40576 = n40575 ^ n1326 ^ 1'b0 ;
  assign n40577 = ~n27066 & n40576 ;
  assign n40578 = ( n2476 & n5520 ) | ( n2476 & n9533 ) | ( n5520 & n9533 ) ;
  assign n40579 = n40578 ^ n24779 ^ n3082 ;
  assign n40580 = n25813 & n40579 ;
  assign n40581 = n40580 ^ n9768 ^ 1'b0 ;
  assign n40582 = n2115 & ~n40581 ;
  assign n40583 = ~n11594 & n40582 ;
  assign n40584 = n40583 ^ n16319 ^ 1'b0 ;
  assign n40585 = ~n11929 & n23335 ;
  assign n40586 = n14409 | n29650 ;
  assign n40587 = n38802 | n40586 ;
  assign n40588 = ~n18539 & n40587 ;
  assign n40589 = n20173 | n25227 ;
  assign n40590 = n11538 | n18986 ;
  assign n40591 = n40590 ^ n28334 ^ 1'b0 ;
  assign n40592 = n1481 & n39275 ;
  assign n40593 = ~n8712 & n21935 ;
  assign n40594 = n2280 & n40593 ;
  assign n40595 = ~n4339 & n40594 ;
  assign n40596 = n607 & n26165 ;
  assign n40601 = n1290 & ~n6638 ;
  assign n40602 = n15979 | n40601 ;
  assign n40597 = n8952 ^ n543 ^ 1'b0 ;
  assign n40598 = n24361 & ~n40597 ;
  assign n40599 = ~n39874 & n40598 ;
  assign n40600 = n40599 ^ n24984 ^ 1'b0 ;
  assign n40603 = n40602 ^ n40600 ^ n31288 ;
  assign n40604 = n24676 ^ n23459 ^ 1'b0 ;
  assign n40605 = n22312 | n24991 ;
  assign n40606 = n40604 & ~n40605 ;
  assign n40607 = ( ~n4426 & n11135 ) | ( ~n4426 & n21171 ) | ( n11135 & n21171 ) ;
  assign n40608 = n10079 | n19316 ;
  assign n40609 = n17780 | n40608 ;
  assign n40610 = ~n40607 & n40609 ;
  assign n40611 = ~n3772 & n40610 ;
  assign n40612 = n379 & n8440 ;
  assign n40613 = n33760 | n36683 ;
  assign n40616 = n10171 & ~n12166 ;
  assign n40614 = ~n21679 & n24200 ;
  assign n40615 = n13013 & n40614 ;
  assign n40617 = n40616 ^ n40615 ^ 1'b0 ;
  assign n40618 = ~n3346 & n12355 ;
  assign n40619 = ~n1220 & n40618 ;
  assign n40620 = ( ~n2403 & n21010 ) | ( ~n2403 & n40619 ) | ( n21010 & n40619 ) ;
  assign n40621 = n12901 | n13660 ;
  assign n40622 = n21548 | n40621 ;
  assign n40623 = ~n10005 & n40622 ;
  assign n40624 = ~n6733 & n40623 ;
  assign n40625 = n19927 & ~n40624 ;
  assign n40626 = n40625 ^ n18130 ^ 1'b0 ;
  assign n40627 = ~n18735 & n24841 ;
  assign n40628 = n6278 & n40627 ;
  assign n40629 = n17493 ^ n3891 ^ 1'b0 ;
  assign n40630 = n40628 & ~n40629 ;
  assign n40631 = n6743 & ~n23893 ;
  assign n40632 = n10223 & n40631 ;
  assign n40633 = n4105 | n40632 ;
  assign n40634 = ( n22925 & n26085 ) | ( n22925 & n37258 ) | ( n26085 & n37258 ) ;
  assign n40635 = n9504 ^ n8210 ^ 1'b0 ;
  assign n40636 = n37766 ^ n14035 ^ 1'b0 ;
  assign n40637 = n23427 & ~n40636 ;
  assign n40638 = n35224 | n37106 ;
  assign n40639 = ~n31819 & n38330 ;
  assign n40640 = n40639 ^ n11267 ^ 1'b0 ;
  assign n40641 = ( n23 & n9425 ) | ( n23 & ~n13585 ) | ( n9425 & ~n13585 ) ;
  assign n40642 = n40641 ^ n17692 ^ 1'b0 ;
  assign n40643 = n29438 ^ n13382 ^ 1'b0 ;
  assign n40644 = n20954 | n30079 ;
  assign n40645 = n29187 | n40644 ;
  assign n40646 = n15956 | n16488 ;
  assign n40647 = n6530 | n40646 ;
  assign n40648 = n2250 & n3833 ;
  assign n40653 = n8421 | n30029 ;
  assign n40654 = n40653 ^ n11490 ^ 1'b0 ;
  assign n40649 = n39869 ^ n6541 ^ 1'b0 ;
  assign n40650 = n40649 ^ n23256 ^ n9236 ;
  assign n40651 = n40650 ^ n12722 ^ 1'b0 ;
  assign n40652 = n25964 | n40651 ;
  assign n40655 = n40654 ^ n40652 ^ n7067 ;
  assign n40656 = n11766 & ~n28986 ;
  assign n40657 = n5882 & n40656 ;
  assign n40658 = n8794 ^ n6873 ^ 1'b0 ;
  assign n40659 = n29229 & n40658 ;
  assign n40660 = ~n22452 & n30262 ;
  assign n40661 = n9734 & n12931 ;
  assign n40662 = n6877 & n40661 ;
  assign n40663 = n1540 & ~n40662 ;
  assign n40665 = n26081 ^ n22139 ^ n20891 ;
  assign n40664 = ~n10907 & n20290 ;
  assign n40666 = n40665 ^ n40664 ^ 1'b0 ;
  assign n40667 = n11929 ^ n9571 ^ n3237 ;
  assign n40668 = ~n24687 & n40667 ;
  assign n40676 = ( n16005 & n20079 ) | ( n16005 & n29813 ) | ( n20079 & n29813 ) ;
  assign n40670 = n34345 ^ n30392 ^ 1'b0 ;
  assign n40671 = n13699 & n40670 ;
  assign n40672 = ~n2832 & n40671 ;
  assign n40673 = n40672 ^ n10745 ^ 1'b0 ;
  assign n40669 = n16212 & ~n28111 ;
  assign n40674 = n40673 ^ n40669 ^ 1'b0 ;
  assign n40675 = n40674 ^ n15534 ^ 1'b0 ;
  assign n40677 = n40676 ^ n40675 ^ 1'b0 ;
  assign n40678 = n15579 & n27307 ;
  assign n40679 = n40581 & n40678 ;
  assign n40680 = n27811 & ~n40679 ;
  assign n40681 = n40680 ^ n8063 ^ n7553 ;
  assign n40682 = ~n11219 & n16398 ;
  assign n40685 = n5350 & ~n36534 ;
  assign n40686 = n40685 ^ n23565 ^ 1'b0 ;
  assign n40683 = n25604 & n37847 ;
  assign n40684 = n40683 ^ n18368 ^ 1'b0 ;
  assign n40687 = n40686 ^ n40684 ^ 1'b0 ;
  assign n40688 = n8775 & n17272 ;
  assign n40691 = ~n823 & n10399 ;
  assign n40689 = n20022 & n24805 ;
  assign n40690 = ~n14345 & n40689 ;
  assign n40692 = n40691 ^ n40690 ^ n17273 ;
  assign n40693 = n10935 ^ n2946 ^ 1'b0 ;
  assign n40696 = n18499 ^ n100 ^ 1'b0 ;
  assign n40697 = n5484 & ~n40696 ;
  assign n40694 = ( n3844 & n4996 ) | ( n3844 & ~n7580 ) | ( n4996 & ~n7580 ) ;
  assign n40695 = n16065 & ~n40694 ;
  assign n40698 = n40697 ^ n40695 ^ 1'b0 ;
  assign n40699 = ( n12119 & n15047 ) | ( n12119 & n40698 ) | ( n15047 & n40698 ) ;
  assign n40700 = ~n2819 & n25885 ;
  assign n40701 = n27012 | n33137 ;
  assign n40702 = n4280 | n10379 ;
  assign n40703 = n4724 & ~n40702 ;
  assign n40704 = ( n5484 & ~n25313 ) | ( n5484 & n40703 ) | ( ~n25313 & n40703 ) ;
  assign n40705 = n33032 ^ n14516 ^ 1'b0 ;
  assign n40706 = n31292 | n34564 ;
  assign n40707 = n16616 & ~n22669 ;
  assign n40708 = n24670 ^ n6361 ^ n722 ;
  assign n40709 = n25941 & ~n40708 ;
  assign n40714 = n10212 ^ n4011 ^ 1'b0 ;
  assign n40710 = n4826 | n4923 ;
  assign n40711 = n15912 & ~n40710 ;
  assign n40712 = n40711 ^ n16131 ^ 1'b0 ;
  assign n40713 = n40712 ^ n6372 ^ n2182 ;
  assign n40715 = n40714 ^ n40713 ^ n4604 ;
  assign n40716 = ( ~n23164 & n27739 ) | ( ~n23164 & n39640 ) | ( n27739 & n39640 ) ;
  assign n40717 = ~n9712 & n22235 ;
  assign n40718 = ( n5301 & ~n40716 ) | ( n5301 & n40717 ) | ( ~n40716 & n40717 ) ;
  assign n40719 = n21741 ^ n12247 ^ 1'b0 ;
  assign n40720 = n6995 & n12921 ;
  assign n40721 = n7626 & ~n40720 ;
  assign n40722 = n40721 ^ n1846 ^ 1'b0 ;
  assign n40723 = n20716 ^ n2729 ^ 1'b0 ;
  assign n40724 = n40723 ^ n29479 ^ 1'b0 ;
  assign n40725 = ~n30279 & n39075 ;
  assign n40726 = n40724 & n40725 ;
  assign n40729 = n9448 & ~n24705 ;
  assign n40727 = n30726 & ~n33713 ;
  assign n40728 = n40727 ^ n6874 ^ 1'b0 ;
  assign n40730 = n40729 ^ n40728 ^ n5160 ;
  assign n40731 = n29088 ^ n431 ^ 1'b0 ;
  assign n40732 = n40731 ^ n13725 ^ 1'b0 ;
  assign n40733 = n29115 | n32475 ;
  assign n40734 = n26926 & n30544 ;
  assign n40736 = n20688 & n27996 ;
  assign n40735 = n1125 & n15989 ;
  assign n40737 = n40736 ^ n40735 ^ 1'b0 ;
  assign n40738 = ~n1965 & n3877 ;
  assign n40739 = n40738 ^ n13643 ^ n676 ;
  assign n40740 = n40739 ^ n38239 ^ 1'b0 ;
  assign n40741 = n7358 & n25067 ;
  assign n40742 = ~x0 & n40741 ;
  assign n40743 = n40742 ^ n11678 ^ 1'b0 ;
  assign n40744 = n11850 & n40743 ;
  assign n40745 = n8323 & ~n40744 ;
  assign n40746 = ( n9026 & n18510 ) | ( n9026 & ~n40745 ) | ( n18510 & ~n40745 ) ;
  assign n40747 = n37403 ^ n13025 ^ 1'b0 ;
  assign n40748 = n332 | n40747 ;
  assign n40749 = n40748 ^ n1800 ^ 1'b0 ;
  assign n40750 = n40749 ^ n31283 ^ n4813 ;
  assign n40751 = n9326 ^ n776 ^ 1'b0 ;
  assign n40752 = n14564 & n40751 ;
  assign n40753 = n15340 & n38553 ;
  assign n40754 = ~n40752 & n40753 ;
  assign n40758 = n12211 ^ n12119 ^ 1'b0 ;
  assign n40759 = n16268 & ~n40758 ;
  assign n40755 = n15020 & ~n27097 ;
  assign n40756 = ~n26802 & n40755 ;
  assign n40757 = n6474 | n40756 ;
  assign n40760 = n40759 ^ n40757 ^ 1'b0 ;
  assign n40761 = ( n717 & ~n3390 ) | ( n717 & n38009 ) | ( ~n3390 & n38009 ) ;
  assign n40762 = n18697 ^ n1172 ^ 1'b0 ;
  assign n40763 = n9138 & n40762 ;
  assign n40764 = ~n9638 & n32621 ;
  assign n40765 = ~n40763 & n40764 ;
  assign n40766 = n5011 & ~n40765 ;
  assign n40767 = n27416 & n40766 ;
  assign n40768 = n108 & ~n12695 ;
  assign n40769 = n2987 & n40768 ;
  assign n40771 = n11074 ^ n5627 ^ n2798 ;
  assign n40770 = n18387 ^ n91 ^ 1'b0 ;
  assign n40772 = n40771 ^ n40770 ^ n8927 ;
  assign n40773 = n17531 ^ n11701 ^ 1'b0 ;
  assign n40774 = n10968 & n14827 ;
  assign n40775 = n37159 ^ n13626 ^ 1'b0 ;
  assign n40776 = n11640 & ~n40775 ;
  assign n40777 = ( n34443 & n40774 ) | ( n34443 & ~n40776 ) | ( n40774 & ~n40776 ) ;
  assign n40778 = n9399 ^ n1159 ^ 1'b0 ;
  assign n40779 = n40777 | n40778 ;
  assign n40780 = ~n15310 & n19258 ;
  assign n40781 = n40780 ^ n14605 ^ 1'b0 ;
  assign n40782 = n1704 | n40781 ;
  assign n40783 = n40782 ^ n35091 ^ 1'b0 ;
  assign n40784 = n27673 & n40438 ;
  assign n40785 = ( n21862 & n32159 ) | ( n21862 & n40784 ) | ( n32159 & n40784 ) ;
  assign n40786 = n10718 & n15198 ;
  assign n40787 = ~n8614 & n40786 ;
  assign n40788 = n16145 ^ n6068 ^ n4785 ;
  assign n40789 = n40787 & n40788 ;
  assign n40790 = n33255 ^ n30598 ^ 1'b0 ;
  assign n40791 = n14698 | n40790 ;
  assign n40792 = n12499 | n24676 ;
  assign n40793 = n40792 ^ n20943 ^ 1'b0 ;
  assign n40794 = n4005 & n4988 ;
  assign n40795 = n25247 ^ n5563 ^ 1'b0 ;
  assign n40796 = ( ~n2569 & n40794 ) | ( ~n2569 & n40795 ) | ( n40794 & n40795 ) ;
  assign n40797 = n36098 ^ n10209 ^ 1'b0 ;
  assign n40798 = n33217 ^ n7144 ^ 1'b0 ;
  assign n40799 = n9996 ^ n6606 ^ 1'b0 ;
  assign n40800 = n37332 ^ n6711 ^ 1'b0 ;
  assign n40801 = n6990 & ~n40800 ;
  assign n40802 = n40801 ^ n17075 ^ 1'b0 ;
  assign n40803 = n10477 | n14587 ;
  assign n40804 = n8210 & ~n36078 ;
  assign n40805 = n36078 & n40804 ;
  assign n40806 = ~n18964 & n40805 ;
  assign n40807 = n1403 | n5515 ;
  assign n40808 = n5515 & ~n40807 ;
  assign n40809 = n4487 & ~n40808 ;
  assign n40810 = ~n4487 & n40809 ;
  assign n40811 = n10769 & ~n40810 ;
  assign n40812 = n40811 ^ n1465 ^ 1'b0 ;
  assign n40813 = n40806 | n40812 ;
  assign n40814 = n19402 | n23376 ;
  assign n40815 = n2805 | n29970 ;
  assign n40816 = n12206 & ~n40815 ;
  assign n40817 = n40816 ^ n35410 ^ 1'b0 ;
  assign n40818 = n24856 ^ n4485 ^ 1'b0 ;
  assign n40819 = n11897 | n19807 ;
  assign n40820 = ~n36861 & n40819 ;
  assign n40821 = n40820 ^ n17123 ^ 1'b0 ;
  assign n40822 = n24414 ^ n17349 ^ n16602 ;
  assign n40823 = n40822 ^ n23375 ^ 1'b0 ;
  assign n40824 = ~n34120 & n40823 ;
  assign n40825 = n33043 & n40824 ;
  assign n40826 = n10361 | n13965 ;
  assign n40827 = n40826 ^ n25813 ^ 1'b0 ;
  assign n40828 = n10186 ^ n6067 ^ n1846 ;
  assign n40829 = ~n12879 & n21198 ;
  assign n40830 = ~n40828 & n40829 ;
  assign n40831 = n16786 ^ n11572 ^ 1'b0 ;
  assign n40832 = ~n35074 & n40831 ;
  assign n40833 = n40832 ^ n10060 ^ 1'b0 ;
  assign n40834 = ~n16594 & n23153 ;
  assign n40835 = n29973 & ~n40834 ;
  assign n40836 = n12301 ^ n11204 ^ n7104 ;
  assign n40837 = n23971 & n28480 ;
  assign n40838 = n40837 ^ n18541 ^ 1'b0 ;
  assign n40839 = n7860 | n11634 ;
  assign n40840 = n40839 ^ n4708 ^ 1'b0 ;
  assign n40841 = n7434 & n16182 ;
  assign n40842 = n17208 ^ n5813 ^ 1'b0 ;
  assign n40843 = n5333 | n19985 ;
  assign n40844 = ( n16650 & ~n40842 ) | ( n16650 & n40843 ) | ( ~n40842 & n40843 ) ;
  assign n40845 = n3720 & ~n13743 ;
  assign n40846 = n23304 ^ n10902 ^ 1'b0 ;
  assign n40847 = ~n2846 & n40846 ;
  assign n40848 = n17671 | n26395 ;
  assign n40849 = n34983 ^ n15195 ^ 1'b0 ;
  assign n40850 = n8759 | n40849 ;
  assign n40851 = n3584 ^ n601 ^ 1'b0 ;
  assign n40852 = ~n28360 & n40851 ;
  assign n40853 = n12600 & n28216 ;
  assign n40854 = ~n15617 & n40853 ;
  assign n40855 = n30662 ^ n19145 ^ 1'b0 ;
  assign n40856 = ~n40854 & n40855 ;
  assign n40857 = n10411 ^ n2618 ^ 1'b0 ;
  assign n40858 = n25829 | n40857 ;
  assign n40859 = n4985 ^ n2678 ^ 1'b0 ;
  assign n40860 = n40859 ^ n13007 ^ 1'b0 ;
  assign n40861 = ( n575 & ~n5197 ) | ( n575 & n38955 ) | ( ~n5197 & n38955 ) ;
  assign n40862 = n4985 | n12951 ;
  assign n40863 = n17897 | n40862 ;
  assign n40864 = n3027 & ~n40863 ;
  assign n40865 = n28188 ^ n2779 ^ 1'b0 ;
  assign n40866 = n27222 | n40865 ;
  assign n40867 = n7856 & ~n40866 ;
  assign n40868 = n2312 | n3198 ;
  assign n40869 = n40868 ^ n24307 ^ 1'b0 ;
  assign n40870 = n40867 & n40869 ;
  assign n40871 = ( n1974 & ~n20383 ) | ( n1974 & n36713 ) | ( ~n20383 & n36713 ) ;
  assign n40872 = n13979 & n20993 ;
  assign n40873 = n40872 ^ n57 ^ 1'b0 ;
  assign n40874 = n40873 ^ n12697 ^ 1'b0 ;
  assign n40875 = n28742 | n40874 ;
  assign n40876 = n17499 & ~n40875 ;
  assign n40877 = n28246 ^ n15590 ^ 1'b0 ;
  assign n40878 = n40876 | n40877 ;
  assign n40879 = n16990 & ~n21677 ;
  assign n40880 = n40879 ^ n3763 ^ 1'b0 ;
  assign n40882 = n23841 ^ n18631 ^ 1'b0 ;
  assign n40881 = n7686 | n10677 ;
  assign n40883 = n40882 ^ n40881 ^ 1'b0 ;
  assign n40884 = ~n401 & n40883 ;
  assign n40885 = n13933 ^ n3131 ^ 1'b0 ;
  assign n40886 = n13946 ^ n6595 ^ 1'b0 ;
  assign n40887 = n11167 & ~n40886 ;
  assign n40888 = n36695 & n39419 ;
  assign n40889 = n27072 ^ n20679 ^ 1'b0 ;
  assign n40890 = n19091 ^ n8032 ^ n143 ;
  assign n40891 = n3736 | n40890 ;
  assign n40892 = n40891 ^ n16603 ^ 1'b0 ;
  assign n40893 = n35927 & n40892 ;
  assign n40894 = n40893 ^ n7389 ^ 1'b0 ;
  assign n40895 = n29650 & ~n40894 ;
  assign n40896 = n4543 & n6455 ;
  assign n40897 = n8591 ^ n5147 ^ 1'b0 ;
  assign n40898 = n13192 ^ n3382 ^ 1'b0 ;
  assign n40899 = n7213 & ~n15940 ;
  assign n40900 = n40899 ^ n14597 ^ 1'b0 ;
  assign n40903 = n25260 | n27159 ;
  assign n40901 = n34345 ^ n5657 ^ n2952 ;
  assign n40902 = n15916 | n40901 ;
  assign n40904 = n40903 ^ n40902 ^ 1'b0 ;
  assign n40905 = n30926 & n40904 ;
  assign n40906 = n40446 ^ n13238 ^ 1'b0 ;
  assign n40907 = ~n1964 & n40906 ;
  assign n40913 = n6356 & ~n6402 ;
  assign n40914 = ~n18337 & n40913 ;
  assign n40910 = n5032 ^ n2815 ^ 1'b0 ;
  assign n40908 = n10452 | n34753 ;
  assign n40909 = n16218 & n40908 ;
  assign n40911 = n40910 ^ n40909 ^ 1'b0 ;
  assign n40912 = n23779 & n40911 ;
  assign n40915 = n40914 ^ n40912 ^ 1'b0 ;
  assign n40916 = n30085 ^ n11860 ^ 1'b0 ;
  assign n40917 = n6342 & ~n12928 ;
  assign n40918 = n9081 & ~n40917 ;
  assign n40919 = ~n24569 & n30158 ;
  assign n40920 = n40919 ^ n29395 ^ n21587 ;
  assign n40921 = n5595 & ~n31164 ;
  assign n40922 = n9036 & n15977 ;
  assign n40923 = n40921 & n40922 ;
  assign n40924 = n22466 & ~n36321 ;
  assign n40925 = n473 & n40924 ;
  assign n40926 = n31935 | n40925 ;
  assign n40927 = n26772 | n35572 ;
  assign n40929 = ( ~n2352 & n7113 ) | ( ~n2352 & n18638 ) | ( n7113 & n18638 ) ;
  assign n40930 = n40929 ^ n24939 ^ n18412 ;
  assign n40928 = ~n8117 & n17556 ;
  assign n40931 = n40930 ^ n40928 ^ 1'b0 ;
  assign n40932 = n12323 ^ n7020 ^ 1'b0 ;
  assign n40933 = n40932 ^ n17565 ^ 1'b0 ;
  assign n40934 = n2747 | n40933 ;
  assign n40935 = n17754 & ~n24260 ;
  assign n40936 = n40935 ^ n24183 ^ 1'b0 ;
  assign n40937 = n40934 & ~n40936 ;
  assign n40938 = n29185 ^ n23152 ^ 1'b0 ;
  assign n40939 = n40938 ^ n990 ^ 1'b0 ;
  assign n40940 = n17247 ^ n462 ^ 1'b0 ;
  assign n40941 = n3915 ^ n1104 ^ 1'b0 ;
  assign n40942 = ( n882 & n40940 ) | ( n882 & ~n40941 ) | ( n40940 & ~n40941 ) ;
  assign n40944 = ( ~n2563 & n12438 ) | ( ~n2563 & n28866 ) | ( n12438 & n28866 ) ;
  assign n40943 = n8728 & n10799 ;
  assign n40945 = n40944 ^ n40943 ^ 1'b0 ;
  assign n40946 = n21725 & ~n40774 ;
  assign n40947 = n30725 & ~n40946 ;
  assign n40948 = ~n23727 & n40947 ;
  assign n40949 = n2113 & ~n40948 ;
  assign n40950 = n17062 & n40949 ;
  assign n40951 = n960 & ~n12290 ;
  assign n40952 = ( ~n11385 & n18526 ) | ( ~n11385 & n40951 ) | ( n18526 & n40951 ) ;
  assign n40953 = n3060 & n11195 ;
  assign n40954 = ~n23514 & n40953 ;
  assign n40955 = n40954 ^ n13404 ^ n532 ;
  assign n40956 = ( n11393 & n36187 ) | ( n11393 & n40955 ) | ( n36187 & n40955 ) ;
  assign n40957 = n31359 & n35796 ;
  assign n40958 = n21315 & n40957 ;
  assign n40959 = n40958 ^ n24484 ^ n13101 ;
  assign n40960 = n37051 ^ n12086 ^ n8228 ;
  assign n40961 = n7122 & n40960 ;
  assign n40962 = n7771 & ~n9716 ;
  assign n40963 = n40962 ^ n9139 ^ 1'b0 ;
  assign n40964 = ~n10699 & n18702 ;
  assign n40965 = n27167 ^ n13965 ^ 1'b0 ;
  assign n40966 = n12734 & n40965 ;
  assign n40967 = ~n20385 & n40966 ;
  assign n40968 = n40967 ^ n349 ^ 1'b0 ;
  assign n40969 = n2985 & ~n38020 ;
  assign n40970 = ~n2345 & n40969 ;
  assign n40971 = n31530 & ~n38870 ;
  assign n40972 = n33340 ^ n11210 ^ 1'b0 ;
  assign n40973 = n12083 | n21035 ;
  assign n40974 = n40973 ^ n18530 ^ 1'b0 ;
  assign n40975 = n1888 & ~n9938 ;
  assign n40976 = n14393 | n24296 ;
  assign n40977 = ~n7081 & n14102 ;
  assign n40978 = n40977 ^ n9003 ^ 1'b0 ;
  assign n40979 = n18699 & n40978 ;
  assign n40980 = ( n5249 & n26474 ) | ( n5249 & n32113 ) | ( n26474 & n32113 ) ;
  assign n40981 = n33784 | n40938 ;
  assign n40982 = n15949 & n24922 ;
  assign n40983 = n40982 ^ n12013 ^ 1'b0 ;
  assign n40984 = n108 & n8882 ;
  assign n40985 = n1071 & n40984 ;
  assign n40986 = n37289 ^ n25687 ^ 1'b0 ;
  assign n40991 = ~n4216 & n6408 ;
  assign n40987 = n12436 ^ n8938 ^ 1'b0 ;
  assign n40988 = n40987 ^ n2216 ^ 1'b0 ;
  assign n40989 = n40988 ^ n27278 ^ 1'b0 ;
  assign n40990 = n18876 & ~n40989 ;
  assign n40992 = n40991 ^ n40990 ^ n21200 ;
  assign n40993 = n6114 & ~n12409 ;
  assign n40994 = n29781 ^ n11090 ^ 1'b0 ;
  assign n40995 = n40993 & ~n40994 ;
  assign n40996 = n8798 & n12898 ;
  assign n40997 = n11245 | n18911 ;
  assign n40998 = n40996 & ~n40997 ;
  assign n40999 = ~n22483 & n40998 ;
  assign n41000 = n11519 ^ n2889 ^ 1'b0 ;
  assign n41001 = n26467 & n41000 ;
  assign n41002 = n1234 | n12658 ;
  assign n41003 = n10659 ^ n6841 ^ n5450 ;
  assign n41004 = n17523 & n41003 ;
  assign n41005 = n41004 ^ n1276 ^ 1'b0 ;
  assign n41006 = ( n1037 & ~n41002 ) | ( n1037 & n41005 ) | ( ~n41002 & n41005 ) ;
  assign n41007 = ( n14783 & ~n18950 ) | ( n14783 & n19169 ) | ( ~n18950 & n19169 ) ;
  assign n41008 = n41007 ^ n1007 ^ 1'b0 ;
  assign n41009 = n9723 | n17295 ;
  assign n41010 = n20751 ^ n6128 ^ 1'b0 ;
  assign n41011 = n7425 | n41010 ;
  assign n41012 = n20078 & ~n35496 ;
  assign n41013 = n2552 & n35079 ;
  assign n41014 = n488 & n41013 ;
  assign n41015 = n39158 ^ n34471 ^ n19653 ;
  assign n41016 = n3694 & ~n17493 ;
  assign n41017 = ~n9578 & n41016 ;
  assign n41018 = ( n4489 & n16389 ) | ( n4489 & ~n41017 ) | ( n16389 & ~n41017 ) ;
  assign n41022 = n26427 ^ n4765 ^ n3479 ;
  assign n41021 = n1622 & ~n10391 ;
  assign n41023 = n41022 ^ n41021 ^ 1'b0 ;
  assign n41019 = n11330 & ~n15091 ;
  assign n41020 = n25221 & n41019 ;
  assign n41024 = n41023 ^ n41020 ^ 1'b0 ;
  assign n41025 = ~n7161 & n20638 ;
  assign n41026 = n41025 ^ n28761 ^ 1'b0 ;
  assign n41027 = ~n13778 & n29650 ;
  assign n41028 = ~n23469 & n38662 ;
  assign n41029 = n4593 ^ n1476 ^ n115 ;
  assign n41030 = n10596 | n41029 ;
  assign n41031 = n6785 | n41030 ;
  assign n41032 = n16329 | n21429 ;
  assign n41033 = n41032 ^ n35112 ^ 1'b0 ;
  assign n41034 = ~n4792 & n41033 ;
  assign n41035 = n39913 ^ n2499 ^ 1'b0 ;
  assign n41036 = ( n15421 & ~n33045 ) | ( n15421 & n38596 ) | ( ~n33045 & n38596 ) ;
  assign n41037 = n31241 ^ n7506 ^ 1'b0 ;
  assign n41038 = n29970 | n41037 ;
  assign n41039 = ~n12371 & n23851 ;
  assign n41040 = n38785 & n41039 ;
  assign n41041 = n7520 ^ n7122 ^ 1'b0 ;
  assign n41042 = ~n17084 & n41041 ;
  assign n41043 = n41042 ^ n33402 ^ 1'b0 ;
  assign n41044 = n14653 & ~n41043 ;
  assign n41045 = ~n22127 & n41044 ;
  assign n41046 = n11547 ^ n1129 ^ 1'b0 ;
  assign n41047 = n5370 | n14965 ;
  assign n41048 = n41047 ^ n28086 ^ 1'b0 ;
  assign n41049 = n41046 & n41048 ;
  assign n41050 = ( n2391 & n30703 ) | ( n2391 & n41049 ) | ( n30703 & n41049 ) ;
  assign n41051 = n18100 ^ n11893 ^ 1'b0 ;
  assign n41052 = ~n29193 & n41051 ;
  assign n41053 = ( n3579 & ~n6490 ) | ( n3579 & n41052 ) | ( ~n6490 & n41052 ) ;
  assign n41054 = n22127 ^ n12711 ^ 1'b0 ;
  assign n41055 = n12053 & ~n25591 ;
  assign n41056 = n250 & n41055 ;
  assign n41057 = n29371 & n41056 ;
  assign n41058 = n25407 ^ n1293 ^ 1'b0 ;
  assign n41059 = ~n850 & n41058 ;
  assign n41060 = n40323 ^ n2314 ^ 1'b0 ;
  assign n41061 = n41059 | n41060 ;
  assign n41062 = n6433 & n10202 ;
  assign n41063 = n41062 ^ n21955 ^ 1'b0 ;
  assign n41064 = n26733 & ~n41063 ;
  assign n41065 = n7101 | n24681 ;
  assign n41066 = n38821 & ~n41065 ;
  assign n41067 = n31634 ^ n5080 ^ 1'b0 ;
  assign n41068 = n7360 & n41067 ;
  assign n41069 = n41068 ^ n1579 ^ 1'b0 ;
  assign n41070 = n13256 ^ n8720 ^ n7102 ;
  assign n41071 = n652 & ~n41070 ;
  assign n41072 = n41071 ^ n9898 ^ 1'b0 ;
  assign n41073 = n41072 ^ n29671 ^ 1'b0 ;
  assign n41074 = n5180 ^ n2108 ^ 1'b0 ;
  assign n41075 = n3057 & n41074 ;
  assign n41076 = n1587 | n35116 ;
  assign n41077 = n13004 ^ n1506 ^ 1'b0 ;
  assign n41078 = n41077 ^ n18556 ^ 1'b0 ;
  assign n41079 = n35998 ^ n33896 ^ 1'b0 ;
  assign n41080 = n2563 ^ n1746 ^ 1'b0 ;
  assign n41081 = n41079 | n41080 ;
  assign n41082 = n145 & ~n11568 ;
  assign n41083 = n41082 ^ n44 ^ 1'b0 ;
  assign n41084 = n27532 & ~n41083 ;
  assign n41085 = n41084 ^ n26794 ^ 1'b0 ;
  assign n41086 = n20407 | n41085 ;
  assign n41087 = ~n11218 & n11243 ;
  assign n41088 = n41087 ^ n22473 ^ 1'b0 ;
  assign n41089 = ( n2661 & n26912 ) | ( n2661 & ~n41088 ) | ( n26912 & ~n41088 ) ;
  assign n41090 = n4313 & ~n38065 ;
  assign n41091 = n41089 | n41090 ;
  assign n41092 = ~n5171 & n16580 ;
  assign n41093 = n13298 ^ n11554 ^ 1'b0 ;
  assign n41094 = n57 & n41093 ;
  assign n41095 = n23588 ^ n18080 ^ 1'b0 ;
  assign n41098 = n1537 | n3853 ;
  assign n41099 = n41098 ^ n132 ^ 1'b0 ;
  assign n41096 = n11753 ^ n2157 ^ 1'b0 ;
  assign n41097 = n13930 | n41096 ;
  assign n41100 = n41099 ^ n41097 ^ 1'b0 ;
  assign n41101 = n15131 | n41100 ;
  assign n41102 = n41101 ^ n23675 ^ 1'b0 ;
  assign n41103 = ~n15086 & n23302 ;
  assign n41104 = n28831 & n31964 ;
  assign n41105 = n17377 & n30455 ;
  assign n41106 = n9278 ^ n1888 ^ 1'b0 ;
  assign n41107 = n40001 & n41106 ;
  assign n41108 = ~n41105 & n41107 ;
  assign n41109 = ~n8964 & n20745 ;
  assign n41110 = n5329 | n30002 ;
  assign n41111 = n3588 & ~n41110 ;
  assign n41112 = n41111 ^ n14107 ^ n5570 ;
  assign n41113 = n9806 | n29054 ;
  assign n41114 = n5490 | n41113 ;
  assign n41115 = n41114 ^ n39095 ^ 1'b0 ;
  assign n41116 = n8804 & ~n41115 ;
  assign n41117 = n41116 ^ n9692 ^ 1'b0 ;
  assign n41118 = ( n1204 & n10290 ) | ( n1204 & n22334 ) | ( n10290 & n22334 ) ;
  assign n41119 = ~n25914 & n41118 ;
  assign n41120 = ~n12779 & n23913 ;
  assign n41121 = n41120 ^ n607 ^ 1'b0 ;
  assign n41122 = n560 & n14715 ;
  assign n41123 = n41122 ^ n13208 ^ 1'b0 ;
  assign n41124 = n24761 & n26218 ;
  assign n41125 = n10578 & n14695 ;
  assign n41126 = ~n1815 & n26994 ;
  assign n41127 = n41126 ^ n6128 ^ 1'b0 ;
  assign n41128 = n1810 & ~n41127 ;
  assign n41129 = n11761 & n41128 ;
  assign n41130 = ~n1004 & n4772 ;
  assign n41131 = n10339 & n41130 ;
  assign n41132 = ~n11916 & n12178 ;
  assign n41133 = ~n398 & n33207 ;
  assign n41134 = n41133 ^ n40108 ^ 1'b0 ;
  assign n41135 = n458 & ~n41134 ;
  assign n41136 = n16841 & ~n41135 ;
  assign n41137 = n13151 | n33423 ;
  assign n41138 = n41137 ^ n40313 ^ 1'b0 ;
  assign n41139 = n1942 | n24044 ;
  assign n41140 = ( n6024 & n39292 ) | ( n6024 & n41139 ) | ( n39292 & n41139 ) ;
  assign n41141 = n4674 | n23261 ;
  assign n41142 = n38445 & ~n41141 ;
  assign n41143 = n14395 & n28063 ;
  assign n41144 = n41142 & n41143 ;
  assign n41145 = n10430 | n25995 ;
  assign n41146 = n126 & ~n41145 ;
  assign n41147 = ~n22090 & n40840 ;
  assign n41148 = n91 & n41147 ;
  assign n41149 = n20847 ^ n8043 ^ 1'b0 ;
  assign n41150 = n34299 & n41149 ;
  assign n41151 = n41150 ^ n7065 ^ 1'b0 ;
  assign n41152 = n41151 ^ n14979 ^ 1'b0 ;
  assign n41153 = ~n2581 & n32382 ;
  assign n41154 = n1419 & n41153 ;
  assign n41155 = ~n10815 & n24715 ;
  assign n41156 = n3793 & n41155 ;
  assign n41157 = n12989 | n28618 ;
  assign n41158 = n41157 ^ n109 ^ 1'b0 ;
  assign n41159 = ~n41156 & n41158 ;
  assign n41160 = n40 & ~n2667 ;
  assign n41161 = n7974 & n8656 ;
  assign n41162 = n41161 ^ n9895 ^ 1'b0 ;
  assign n41163 = n9764 & ~n19596 ;
  assign n41164 = n3466 & n41163 ;
  assign n41165 = n3810 & ~n18416 ;
  assign n41166 = ~n1055 & n36126 ;
  assign n41167 = ( n15452 & ~n21474 ) | ( n15452 & n29774 ) | ( ~n21474 & n29774 ) ;
  assign n41168 = ~n1327 & n3637 ;
  assign n41169 = n41168 ^ n19974 ^ 1'b0 ;
  assign n41170 = n41169 ^ n23500 ^ n4892 ;
  assign n41171 = n18577 ^ n9105 ^ n3345 ;
  assign n41172 = n21134 & ~n41171 ;
  assign n41173 = n41172 ^ n5809 ^ 1'b0 ;
  assign n41174 = n11101 ^ n10348 ^ n2374 ;
  assign n41175 = n35369 ^ n20545 ^ 1'b0 ;
  assign n41176 = ~n41174 & n41175 ;
  assign n41177 = n1933 | n22134 ;
  assign n41178 = n41177 ^ n281 ^ 1'b0 ;
  assign n41179 = n2216 & n41178 ;
  assign n41180 = n41179 ^ n34191 ^ 1'b0 ;
  assign n41183 = n4116 | n6574 ;
  assign n41181 = n28453 ^ n2284 ^ 1'b0 ;
  assign n41182 = n7759 & ~n41181 ;
  assign n41184 = n41183 ^ n41182 ^ n16622 ;
  assign n41185 = n19238 ^ n13081 ^ 1'b0 ;
  assign n41186 = n6121 ^ n622 ^ 1'b0 ;
  assign n41187 = n3811 | n22312 ;
  assign n41188 = n41186 | n41187 ;
  assign n41189 = n2070 ^ n885 ^ 1'b0 ;
  assign n41190 = n9721 | n41189 ;
  assign n41191 = ( n3387 & n18221 ) | ( n3387 & n31334 ) | ( n18221 & n31334 ) ;
  assign n41192 = n11925 ^ n5302 ^ n2517 ;
  assign n41193 = n23658 ^ n7490 ^ 1'b0 ;
  assign n41197 = n39489 ^ n1319 ^ 1'b0 ;
  assign n41194 = ( n1126 & n14649 ) | ( n1126 & n20356 ) | ( n14649 & n20356 ) ;
  assign n41195 = n5939 | n41194 ;
  assign n41196 = n1668 | n41195 ;
  assign n41198 = n41197 ^ n41196 ^ 1'b0 ;
  assign n41199 = n32343 & ~n39067 ;
  assign n41200 = n6589 & n41199 ;
  assign n41201 = n11213 & ~n12171 ;
  assign n41202 = n581 & ~n6618 ;
  assign n41205 = n5667 & ~n8452 ;
  assign n41206 = ~n4997 & n41205 ;
  assign n41204 = n17604 | n31639 ;
  assign n41207 = n41206 ^ n41204 ^ 1'b0 ;
  assign n41203 = n3781 & ~n6353 ;
  assign n41208 = n41207 ^ n41203 ^ 1'b0 ;
  assign n41209 = n32619 ^ n27657 ^ n9658 ;
  assign n41210 = n41209 ^ n30110 ^ n63 ;
  assign n41211 = n41210 ^ n4622 ^ n342 ;
  assign n41212 = ( n15068 & n29029 ) | ( n15068 & n41211 ) | ( n29029 & n41211 ) ;
  assign n41213 = n35569 & ~n36400 ;
  assign n41214 = n41213 ^ n20943 ^ 1'b0 ;
  assign n41215 = n41214 ^ n6254 ^ 1'b0 ;
  assign n41216 = n22605 ^ n17932 ^ n1662 ;
  assign n41217 = ( n8594 & n13819 ) | ( n8594 & ~n41216 ) | ( n13819 & ~n41216 ) ;
  assign n41218 = n32777 ^ n30338 ^ n20602 ;
  assign n41219 = n41218 ^ n23763 ^ 1'b0 ;
  assign n41220 = ~n4490 & n28651 ;
  assign n41221 = n40490 ^ n14835 ^ 1'b0 ;
  assign n41222 = n31085 ^ n19383 ^ n2294 ;
  assign n41223 = n23739 ^ n19270 ^ 1'b0 ;
  assign n41224 = n41223 ^ n6266 ^ 1'b0 ;
  assign n41226 = n20793 & ~n39841 ;
  assign n41225 = n12321 & n14386 ;
  assign n41227 = n41226 ^ n41225 ^ 1'b0 ;
  assign n41228 = ~n15870 & n23535 ;
  assign n41230 = n179 | n1979 ;
  assign n41231 = n21781 & ~n41230 ;
  assign n41229 = ~n13923 & n27133 ;
  assign n41232 = n41231 ^ n41229 ^ 1'b0 ;
  assign n41235 = n8624 ^ n1391 ^ 1'b0 ;
  assign n41233 = ~n9793 & n15586 ;
  assign n41234 = n32761 & n41233 ;
  assign n41236 = n41235 ^ n41234 ^ n35883 ;
  assign n41237 = ~n15926 & n23903 ;
  assign n41238 = n5639 & ~n26257 ;
  assign n41239 = n41238 ^ n23795 ^ 1'b0 ;
  assign n41240 = n28898 & ~n41239 ;
  assign n41241 = n41240 ^ n26971 ^ 1'b0 ;
  assign n41242 = n28816 ^ n23449 ^ 1'b0 ;
  assign n41243 = n41241 & ~n41242 ;
  assign n41244 = n35099 ^ n949 ^ 1'b0 ;
  assign n41245 = n33648 ^ n26178 ^ 1'b0 ;
  assign n41246 = n29813 ^ n6221 ^ 1'b0 ;
  assign n41247 = n34468 & n41246 ;
  assign n41249 = n16871 ^ n4319 ^ 1'b0 ;
  assign n41248 = n958 & ~n24745 ;
  assign n41250 = n41249 ^ n41248 ^ 1'b0 ;
  assign n41251 = ~n16030 & n41250 ;
  assign n41253 = n4482 | n28805 ;
  assign n41254 = n37775 | n41253 ;
  assign n41252 = n213 & n7516 ;
  assign n41255 = n41254 ^ n41252 ^ 1'b0 ;
  assign n41256 = n40774 ^ n17133 ^ 1'b0 ;
  assign n41257 = n41255 & n41256 ;
  assign n41258 = n17438 ^ n10420 ^ 1'b0 ;
  assign n41259 = n12840 | n41258 ;
  assign n41260 = n38912 & ~n41259 ;
  assign n41263 = ~n3307 & n22261 ;
  assign n41261 = n10375 & n24527 ;
  assign n41262 = n41261 ^ n16822 ^ 1'b0 ;
  assign n41264 = n41263 ^ n41262 ^ n9128 ;
  assign n41265 = n25933 | n27867 ;
  assign n41266 = n41265 ^ n32398 ^ 1'b0 ;
  assign n41267 = n14507 ^ n2986 ^ 1'b0 ;
  assign n41268 = n6533 & ~n11066 ;
  assign n41269 = ~n11582 & n41268 ;
  assign n41270 = n29664 | n32770 ;
  assign n41271 = n11718 & ~n41270 ;
  assign n41272 = ~n7505 & n14798 ;
  assign n41273 = n41271 & ~n41272 ;
  assign n41274 = n41269 | n41273 ;
  assign n41275 = n5335 ^ n3818 ^ 1'b0 ;
  assign n41276 = n5888 & ~n12275 ;
  assign n41277 = n10391 & n41276 ;
  assign n41278 = n25573 ^ n21784 ^ 1'b0 ;
  assign n41279 = n22286 | n41278 ;
  assign n41280 = ( n289 & n24749 ) | ( n289 & ~n36212 ) | ( n24749 & ~n36212 ) ;
  assign n41281 = n23615 ^ n3969 ^ 1'b0 ;
  assign n41282 = n33093 & ~n41281 ;
  assign n41283 = ~n2759 & n3351 ;
  assign n41284 = n41283 ^ n4491 ^ 1'b0 ;
  assign n41285 = ~n3546 & n9560 ;
  assign n41286 = ~n7618 & n41285 ;
  assign n41287 = ~n33326 & n41286 ;
  assign n41288 = n21936 & ~n41287 ;
  assign n41289 = n36227 & n41288 ;
  assign n41290 = n33091 ^ n28922 ^ n26189 ;
  assign n41291 = n2104 | n30529 ;
  assign n41292 = n13199 & ~n41291 ;
  assign n41293 = n41292 ^ n8101 ^ 1'b0 ;
  assign n41294 = ( n16682 & n37348 ) | ( n16682 & ~n41293 ) | ( n37348 & ~n41293 ) ;
  assign n41295 = n604 | n15729 ;
  assign n41296 = n41295 ^ n17603 ^ 1'b0 ;
  assign n41297 = n34713 & n41296 ;
  assign n41298 = n17617 & n27489 ;
  assign n41299 = ~n41297 & n41298 ;
  assign n41300 = n32431 ^ n4084 ^ 1'b0 ;
  assign n41301 = n2281 & n41300 ;
  assign n41302 = n7265 | n10596 ;
  assign n41303 = n17042 | n41302 ;
  assign n41304 = ( n15720 & n31461 ) | ( n15720 & n41303 ) | ( n31461 & n41303 ) ;
  assign n41305 = n9086 & n41304 ;
  assign n41306 = n6264 & n41305 ;
  assign n41307 = n21138 ^ n13151 ^ 1'b0 ;
  assign n41308 = n11585 & ~n41307 ;
  assign n41309 = n15994 & n25924 ;
  assign n41310 = ( n8090 & n41308 ) | ( n8090 & n41309 ) | ( n41308 & n41309 ) ;
  assign n41311 = ~n18695 & n23108 ;
  assign n41312 = ~n32096 & n41311 ;
  assign n41313 = n41312 ^ n8480 ^ 1'b0 ;
  assign n41314 = n41313 ^ n12506 ^ 1'b0 ;
  assign n41316 = n20921 ^ n13808 ^ 1'b0 ;
  assign n41317 = n29112 & ~n36144 ;
  assign n41318 = ~n41316 & n41317 ;
  assign n41315 = ( n962 & ~n6553 ) | ( n962 & n20386 ) | ( ~n6553 & n20386 ) ;
  assign n41319 = n41318 ^ n41315 ^ 1'b0 ;
  assign n41320 = n5743 ^ n188 ^ 1'b0 ;
  assign n41321 = n16230 | n41320 ;
  assign n41322 = n41319 & ~n41321 ;
  assign n41323 = ~n11998 & n22411 ;
  assign n41324 = n2990 & n41323 ;
  assign n41325 = n556 & ~n15464 ;
  assign n41326 = n41325 ^ n4927 ^ 1'b0 ;
  assign n41327 = n16837 | n24431 ;
  assign n41328 = n21253 & ~n41327 ;
  assign n41329 = ~n5350 & n41328 ;
  assign n41330 = n1628 & ~n11465 ;
  assign n41331 = n11465 & n41330 ;
  assign n41332 = n14236 & ~n20443 ;
  assign n41333 = n20443 & n41332 ;
  assign n41334 = ( n3638 & ~n41331 ) | ( n3638 & n41333 ) | ( ~n41331 & n41333 ) ;
  assign n41335 = n24512 ^ n16468 ^ 1'b0 ;
  assign n41336 = n20529 | n41335 ;
  assign n41337 = n25157 | n32122 ;
  assign n41338 = n41337 ^ n18111 ^ 1'b0 ;
  assign n41339 = n2041 & ~n12880 ;
  assign n41340 = ~n2041 & n41339 ;
  assign n41341 = n41340 ^ n21913 ^ 1'b0 ;
  assign n41342 = n10517 & ~n41341 ;
  assign n41343 = ( ~n10106 & n12323 ) | ( ~n10106 & n19592 ) | ( n12323 & n19592 ) ;
  assign n41344 = n102 & ~n17793 ;
  assign n41346 = ~n7500 & n33274 ;
  assign n41347 = n41346 ^ n14711 ^ 1'b0 ;
  assign n41345 = n11743 ^ n7165 ^ x7 ;
  assign n41348 = n41347 ^ n41345 ^ n7699 ;
  assign n41349 = ~n41344 & n41348 ;
  assign n41350 = n17718 & n26503 ;
  assign n41351 = n41350 ^ n4851 ^ 1'b0 ;
  assign n41352 = ( ~n14256 & n40720 ) | ( ~n14256 & n41351 ) | ( n40720 & n41351 ) ;
  assign n41353 = n9658 ^ n6562 ^ 1'b0 ;
  assign n41354 = n41353 ^ n39224 ^ 1'b0 ;
  assign n41355 = n2257 & ~n41354 ;
  assign n41356 = n15859 ^ n15456 ^ 1'b0 ;
  assign n41357 = n20929 & n41356 ;
  assign n41358 = n40865 ^ n21552 ^ 1'b0 ;
  assign n41359 = n41357 & ~n41358 ;
  assign n41360 = n8866 & n41359 ;
  assign n41361 = n41360 ^ n38060 ^ 1'b0 ;
  assign n41362 = n5868 | n30948 ;
  assign n41363 = n41362 ^ n473 ^ 1'b0 ;
  assign n41364 = ~n3600 & n20525 ;
  assign n41365 = ~n570 & n41364 ;
  assign n41366 = n22586 & ~n41365 ;
  assign n41367 = n41363 & n41366 ;
  assign n41368 = ( ~n14758 & n41361 ) | ( ~n14758 & n41367 ) | ( n41361 & n41367 ) ;
  assign n41369 = n6511 & n41368 ;
  assign n41370 = n22488 & n41369 ;
  assign n41371 = ~n1256 & n8631 ;
  assign n41372 = ~n1177 & n14531 ;
  assign n41375 = n1389 & n11195 ;
  assign n41373 = n9079 | n15210 ;
  assign n41374 = n16959 & ~n41373 ;
  assign n41376 = n41375 ^ n41374 ^ n2507 ;
  assign n41377 = n30489 ^ n24311 ^ n22662 ;
  assign n41378 = n8906 | n40214 ;
  assign n41379 = ( n10586 & ~n13123 ) | ( n10586 & n37470 ) | ( ~n13123 & n37470 ) ;
  assign n41380 = n20824 ^ n8055 ^ 1'b0 ;
  assign n41381 = ~n14452 & n41380 ;
  assign n41382 = n41381 ^ n35405 ^ 1'b0 ;
  assign n41383 = n1751 & n6892 ;
  assign n41384 = n41383 ^ n14611 ^ 1'b0 ;
  assign n41385 = n41384 ^ n7694 ^ 1'b0 ;
  assign n41386 = ~n17373 & n41385 ;
  assign n41387 = n27673 & n40024 ;
  assign n41388 = n2497 & n41387 ;
  assign n41389 = n4575 & n19354 ;
  assign n41391 = n10094 ^ n2418 ^ 1'b0 ;
  assign n41392 = n6903 & ~n21732 ;
  assign n41393 = ~n41391 & n41392 ;
  assign n41394 = ( n3288 & ~n9274 ) | ( n3288 & n41393 ) | ( ~n9274 & n41393 ) ;
  assign n41395 = n41394 ^ n19267 ^ 1'b0 ;
  assign n41396 = n1940 & n41395 ;
  assign n41397 = n41396 ^ n27192 ^ 1'b0 ;
  assign n41398 = n25487 & n41397 ;
  assign n41390 = n21075 ^ n8591 ^ 1'b0 ;
  assign n41399 = n41398 ^ n41390 ^ n22070 ;
  assign n41400 = n744 | n21262 ;
  assign n41401 = n41400 ^ n7020 ^ 1'b0 ;
  assign n41402 = n13268 | n41401 ;
  assign n41403 = n40146 ^ n37540 ^ 1'b0 ;
  assign n41404 = n23131 | n32530 ;
  assign n41405 = n41404 ^ n17617 ^ 1'b0 ;
  assign n41406 = n10593 ^ n8575 ^ 1'b0 ;
  assign n41407 = n1940 & n3385 ;
  assign n41408 = n35516 & n41407 ;
  assign n41409 = ~n8043 & n29897 ;
  assign n41411 = n5848 & ~n9504 ;
  assign n41410 = n31177 | n33178 ;
  assign n41412 = n41411 ^ n41410 ^ 1'b0 ;
  assign n41413 = n4859 | n8082 ;
  assign n41414 = n4859 & ~n41413 ;
  assign n41415 = n41253 & ~n41414 ;
  assign n41416 = n41415 ^ n4467 ^ 1'b0 ;
  assign n41417 = n8574 | n14129 ;
  assign n41418 = n19898 | n41417 ;
  assign n41419 = n24053 ^ n7267 ^ 1'b0 ;
  assign n41420 = n3119 & ~n41419 ;
  assign n41421 = n25 | n20220 ;
  assign n41422 = n41421 ^ n19426 ^ 1'b0 ;
  assign n41423 = n3604 | n9303 ;
  assign n41426 = n6874 ^ n5990 ^ 1'b0 ;
  assign n41424 = ~n2466 & n15789 ;
  assign n41425 = n41424 ^ n29198 ^ 1'b0 ;
  assign n41427 = n41426 ^ n41425 ^ n40333 ;
  assign n41428 = n5939 | n11768 ;
  assign n41429 = n41428 ^ n7388 ^ 1'b0 ;
  assign n41430 = n37334 ^ n33368 ^ 1'b0 ;
  assign n41431 = n24909 & ~n41430 ;
  assign n41432 = n1891 | n6044 ;
  assign n41433 = n11216 & n20835 ;
  assign n41434 = n41432 | n41433 ;
  assign n41435 = n21918 & ~n41434 ;
  assign n41436 = n13832 & n41435 ;
  assign n41437 = n31394 ^ n15059 ^ 1'b0 ;
  assign n41438 = n17883 | n19186 ;
  assign n41439 = ~n15391 & n41438 ;
  assign n41440 = n40367 & n41439 ;
  assign n41441 = n22690 ^ n10494 ^ 1'b0 ;
  assign n41442 = n26963 & n41441 ;
  assign n41443 = n11535 ^ n5554 ^ 1'b0 ;
  assign n41444 = n7907 ^ n1345 ^ 1'b0 ;
  assign n41445 = n41444 ^ n37689 ^ n1450 ;
  assign n41446 = n19204 & n27068 ;
  assign n41447 = n12049 ^ n7121 ^ 1'b0 ;
  assign n41448 = n41447 ^ n26565 ^ 1'b0 ;
  assign n41449 = n22411 & n41448 ;
  assign n41450 = n3054 | n4847 ;
  assign n41451 = n41450 ^ n19052 ^ 1'b0 ;
  assign n41452 = n34086 ^ n19839 ^ 1'b0 ;
  assign n41453 = ~n41451 & n41452 ;
  assign n41454 = n16491 & n24347 ;
  assign n41455 = n41454 ^ n37185 ^ 1'b0 ;
  assign n41456 = n41455 ^ n1463 ^ 1'b0 ;
  assign n41465 = n9915 ^ n6428 ^ 1'b0 ;
  assign n41457 = ~n14017 & n21795 ;
  assign n41458 = n41457 ^ n6067 ^ 1'b0 ;
  assign n41459 = n35048 ^ n567 ^ 1'b0 ;
  assign n41460 = ~n26428 & n41459 ;
  assign n41461 = ~n13172 & n21905 ;
  assign n41462 = ~n41460 & n41461 ;
  assign n41463 = ( n7930 & n41458 ) | ( n7930 & n41462 ) | ( n41458 & n41462 ) ;
  assign n41464 = n7295 | n41463 ;
  assign n41466 = n41465 ^ n41464 ^ 1'b0 ;
  assign n41467 = n7694 & ~n41466 ;
  assign n41468 = n19810 ^ n4159 ^ n424 ;
  assign n41469 = n7707 & n12304 ;
  assign n41471 = ~n14069 & n23282 ;
  assign n41472 = n41471 ^ n23493 ^ n3216 ;
  assign n41470 = n17491 & ~n23718 ;
  assign n41473 = n41472 ^ n41470 ^ 1'b0 ;
  assign n41474 = ~n3575 & n23046 ;
  assign n41475 = ( n6066 & n9901 ) | ( n6066 & n13524 ) | ( n9901 & n13524 ) ;
  assign n41476 = n41475 ^ n37263 ^ 1'b0 ;
  assign n41477 = n20745 ^ n980 ^ 1'b0 ;
  assign n41478 = n41476 & n41477 ;
  assign n41479 = n27374 ^ n21148 ^ 1'b0 ;
  assign n41480 = ( ~n4815 & n34563 ) | ( ~n4815 & n38117 ) | ( n34563 & n38117 ) ;
  assign n41481 = n19935 ^ n15581 ^ 1'b0 ;
  assign n41482 = n41481 ^ n23802 ^ 1'b0 ;
  assign n41483 = ~n7836 & n41482 ;
  assign n41484 = ~n35139 & n41483 ;
  assign n41485 = n41484 ^ n40333 ^ 1'b0 ;
  assign n41486 = n11225 ^ n6356 ^ n4949 ;
  assign n41487 = ( n12482 & n20177 ) | ( n12482 & n41486 ) | ( n20177 & n41486 ) ;
  assign n41488 = n14533 | n41487 ;
  assign n41489 = n24216 | n41488 ;
  assign n41490 = n19710 ^ n3843 ^ n744 ;
  assign n41491 = n20048 ^ n1346 ^ 1'b0 ;
  assign n41492 = n41490 | n41491 ;
  assign n41493 = n29088 ^ n14131 ^ 1'b0 ;
  assign n41494 = n17413 | n41493 ;
  assign n41495 = n41494 ^ n37388 ^ 1'b0 ;
  assign n41496 = n18447 | n41495 ;
  assign n41497 = n41496 ^ n2582 ^ 1'b0 ;
  assign n41498 = n3313 & n41497 ;
  assign n41499 = n12445 ^ n1069 ^ 1'b0 ;
  assign n41500 = n24011 & ~n41499 ;
  assign n41501 = n4458 ^ n779 ^ 1'b0 ;
  assign n41502 = ~n1000 & n41501 ;
  assign n41503 = n8228 & n41502 ;
  assign n41504 = n39456 ^ n6016 ^ n1364 ;
  assign n41505 = n31383 ^ n22022 ^ 1'b0 ;
  assign n41506 = n7766 & ~n36596 ;
  assign n41507 = n41506 ^ n20665 ^ 1'b0 ;
  assign n41508 = ~n27954 & n37551 ;
  assign n41509 = n40720 ^ n15649 ^ 1'b0 ;
  assign n41510 = n32973 ^ n20288 ^ 1'b0 ;
  assign n41511 = n3313 & n23672 ;
  assign n41512 = n13603 & n23950 ;
  assign n41513 = ~n24274 & n41512 ;
  assign n41514 = n41513 ^ n9033 ^ 1'b0 ;
  assign n41515 = ( n6001 & n6941 ) | ( n6001 & n13040 ) | ( n6941 & n13040 ) ;
  assign n41516 = n12784 ^ n8071 ^ 1'b0 ;
  assign n41517 = n3295 ^ n649 ^ 1'b0 ;
  assign n41518 = ~n41516 & n41517 ;
  assign n41519 = n41518 ^ n14141 ^ n9630 ;
  assign n41520 = n41515 & ~n41519 ;
  assign n41521 = ~n32256 & n41520 ;
  assign n41522 = n29611 & n32096 ;
  assign n41523 = n41522 ^ n19630 ^ n3088 ;
  assign n41524 = ~n3790 & n20146 ;
  assign n41525 = ~n35190 & n41524 ;
  assign n41526 = n16787 ^ n131 ^ 1'b0 ;
  assign n41527 = ( n6866 & n6885 ) | ( n6866 & ~n41526 ) | ( n6885 & ~n41526 ) ;
  assign n41528 = n41527 ^ n10846 ^ n10405 ;
  assign n41529 = n41528 ^ n26007 ^ n8106 ;
  assign n41530 = n1832 & ~n41529 ;
  assign n41531 = n41525 & n41530 ;
  assign n41532 = ( n8738 & n12704 ) | ( n8738 & n40117 ) | ( n12704 & n40117 ) ;
  assign n41533 = ~n12596 & n41532 ;
  assign n41534 = n12402 ^ n3457 ^ 1'b0 ;
  assign n41535 = n9706 ^ n1768 ^ 1'b0 ;
  assign n41536 = n12261 ^ n249 ^ 1'b0 ;
  assign n41537 = ~n13371 & n41536 ;
  assign n41538 = n10106 & n15999 ;
  assign n41539 = n41538 ^ n17082 ^ 1'b0 ;
  assign n41540 = ~n411 & n17954 ;
  assign n41541 = n39868 | n40862 ;
  assign n41542 = n41541 ^ n9832 ^ 1'b0 ;
  assign n41543 = ~n183 & n6693 ;
  assign n41544 = n1665 & n41543 ;
  assign n41545 = n41544 ^ n3714 ^ 1'b0 ;
  assign n41546 = n16550 & n41545 ;
  assign n41547 = ~n6174 & n18926 ;
  assign n41548 = ~n11772 & n41547 ;
  assign n41549 = n626 & ~n38073 ;
  assign n41550 = ~n18172 & n41549 ;
  assign n41551 = ( n2139 & n21985 ) | ( n2139 & n23900 ) | ( n21985 & n23900 ) ;
  assign n41552 = n2418 | n17915 ;
  assign n41553 = ~n11456 & n26776 ;
  assign n41554 = n41552 & ~n41553 ;
  assign n41555 = n39883 ^ n21079 ^ 1'b0 ;
  assign n41556 = n27507 | n41555 ;
  assign n41557 = n41556 ^ n25755 ^ 1'b0 ;
  assign n41558 = n41557 ^ n13399 ^ 1'b0 ;
  assign n41559 = n5904 & n41558 ;
  assign n41560 = n1084 & n40425 ;
  assign n41561 = n15726 ^ n3731 ^ 1'b0 ;
  assign n41562 = ~n1866 & n36930 ;
  assign n41563 = ~n10551 & n41562 ;
  assign n41564 = ( n20212 & n24580 ) | ( n20212 & n41563 ) | ( n24580 & n41563 ) ;
  assign n41565 = n10289 & ~n41564 ;
  assign n41566 = n22117 ^ n14684 ^ 1'b0 ;
  assign n41567 = n24956 ^ n11416 ^ 1'b0 ;
  assign n41568 = n41567 ^ n4140 ^ 1'b0 ;
  assign n41569 = n8768 & ~n32133 ;
  assign n41570 = ~n7357 & n41569 ;
  assign n41571 = n6686 & ~n41570 ;
  assign n41572 = n39281 ^ n20676 ^ 1'b0 ;
  assign n41573 = n4844 & ~n22777 ;
  assign n41574 = ~n17155 & n28646 ;
  assign n41575 = n41574 ^ n756 ^ 1'b0 ;
  assign n41576 = n41575 ^ n15742 ^ 1'b0 ;
  assign n41577 = n17107 & ~n36722 ;
  assign n41578 = n41577 ^ n13496 ^ 1'b0 ;
  assign n41579 = ( n2142 & ~n4551 ) | ( n2142 & n28292 ) | ( ~n4551 & n28292 ) ;
  assign n41580 = n34556 ^ n15498 ^ 1'b0 ;
  assign n41581 = n5348 & n41580 ;
  assign n41582 = n7954 & ~n41581 ;
  assign n41583 = ~n2687 & n25877 ;
  assign n41584 = n23810 & n28841 ;
  assign n41585 = n10254 & n19529 ;
  assign n41586 = ~n5549 & n41585 ;
  assign n41587 = n41586 ^ n29617 ^ n5886 ;
  assign n41588 = ~n8851 & n14523 ;
  assign n41589 = n41588 ^ n32133 ^ n20199 ;
  assign n41590 = n5915 | n41589 ;
  assign n41591 = n13574 ^ n3790 ^ 1'b0 ;
  assign n41592 = n34589 & ~n41591 ;
  assign n41593 = n12844 & n17617 ;
  assign n41594 = ( ~n11227 & n28664 ) | ( ~n11227 & n30068 ) | ( n28664 & n30068 ) ;
  assign n41595 = n40044 ^ n4458 ^ 1'b0 ;
  assign n41596 = n25560 & ~n26793 ;
  assign n41597 = n10380 & ~n11510 ;
  assign n41598 = n41597 ^ n6050 ^ 1'b0 ;
  assign n41599 = n41598 ^ n2563 ^ 1'b0 ;
  assign n41600 = n15079 ^ n11356 ^ 1'b0 ;
  assign n41601 = n41599 & n41600 ;
  assign n41602 = n28892 & ~n32054 ;
  assign n41603 = ~n41601 & n41602 ;
  assign n41604 = n15266 & n21439 ;
  assign n41605 = n12014 | n29632 ;
  assign n41606 = n7510 & ~n41605 ;
  assign n41607 = n40702 ^ n31006 ^ n12366 ;
  assign n41608 = ( x10 & ~n1586 ) | ( x10 & n2576 ) | ( ~n1586 & n2576 ) ;
  assign n41610 = n25325 ^ n17099 ^ n7386 ;
  assign n41611 = n41610 ^ n17893 ^ 1'b0 ;
  assign n41609 = n23094 ^ n2089 ^ n43 ;
  assign n41612 = n41611 ^ n41609 ^ n25237 ;
  assign n41613 = n6804 ^ n1596 ^ 1'b0 ;
  assign n41614 = ~n21776 & n41613 ;
  assign n41615 = n7208 & ~n17712 ;
  assign n41616 = ~n41614 & n41615 ;
  assign n41617 = n25039 ^ n16691 ^ n12185 ;
  assign n41618 = n21182 & ~n41617 ;
  assign n41619 = n17783 & n41618 ;
  assign n41620 = n22778 & n41619 ;
  assign n41621 = n6024 & ~n11854 ;
  assign n41622 = n14422 | n41621 ;
  assign n41623 = n41622 ^ n25039 ^ 1'b0 ;
  assign n41624 = n4304 & n16736 ;
  assign n41625 = n41624 ^ n28825 ^ 1'b0 ;
  assign n41626 = n13345 & ~n41625 ;
  assign n41627 = n18859 ^ n2451 ^ 1'b0 ;
  assign n41628 = n32094 & ~n39113 ;
  assign n41629 = n41628 ^ n1970 ^ 1'b0 ;
  assign n41632 = n1381 | n1816 ;
  assign n41633 = ~n5176 & n41632 ;
  assign n41630 = n5751 | n28755 ;
  assign n41631 = n17292 | n41630 ;
  assign n41634 = n41633 ^ n41631 ^ n19198 ;
  assign n41635 = ( n8299 & n10826 ) | ( n8299 & ~n41634 ) | ( n10826 & ~n41634 ) ;
  assign n41636 = ( n2761 & n15383 ) | ( n2761 & n38562 ) | ( n15383 & n38562 ) ;
  assign n41637 = n41636 ^ n5219 ^ 1'b0 ;
  assign n41638 = n7124 & n41637 ;
  assign n41639 = n4121 & ~n29563 ;
  assign n41640 = ~n6544 & n41639 ;
  assign n41641 = n17920 & ~n41640 ;
  assign n41642 = n7753 & n41641 ;
  assign n41643 = n5285 | n7891 ;
  assign n41644 = n41643 ^ n4807 ^ 1'b0 ;
  assign n41645 = n41642 | n41644 ;
  assign n41646 = ~n22935 & n39264 ;
  assign n41647 = n41646 ^ n23933 ^ 1'b0 ;
  assign n41649 = n12986 | n13974 ;
  assign n41648 = n8143 | n39872 ;
  assign n41650 = n41649 ^ n41648 ^ 1'b0 ;
  assign n41651 = n5001 & n8163 ;
  assign n41652 = n17022 & ~n41651 ;
  assign n41653 = n41652 ^ n30062 ^ n25560 ;
  assign n41654 = ~n6647 & n41653 ;
  assign n41655 = n2687 | n14533 ;
  assign n41656 = n41655 ^ n32347 ^ 1'b0 ;
  assign n41657 = n10202 ^ n1371 ^ 1'b0 ;
  assign n41658 = n41657 ^ n6413 ^ 1'b0 ;
  assign n41659 = n36822 ^ n17980 ^ 1'b0 ;
  assign n41660 = n14570 & ~n41659 ;
  assign n41661 = n38907 ^ n166 ^ 1'b0 ;
  assign n41662 = n2570 & n41661 ;
  assign n41664 = n17280 & n24956 ;
  assign n41665 = n41664 ^ n12767 ^ n9120 ;
  assign n41666 = n13755 & ~n41665 ;
  assign n41663 = n4345 & n20166 ;
  assign n41667 = n41666 ^ n41663 ^ 1'b0 ;
  assign n41668 = n24143 | n27532 ;
  assign n41669 = n40017 ^ n14961 ^ 1'b0 ;
  assign n41670 = n13939 | n41669 ;
  assign n41671 = n1131 & ~n41670 ;
  assign n41672 = n41671 ^ n24169 ^ 1'b0 ;
  assign n41673 = ~n1787 & n3786 ;
  assign n41674 = n41673 ^ n23744 ^ 1'b0 ;
  assign n41675 = ~n15872 & n22610 ;
  assign n41676 = ~n6288 & n41675 ;
  assign n41677 = n23265 ^ n68 ^ 1'b0 ;
  assign n41678 = n41676 | n41677 ;
  assign n41679 = ~n9290 & n12111 ;
  assign n41680 = ~n16704 & n18785 ;
  assign n41681 = n41680 ^ n25427 ^ 1'b0 ;
  assign n41682 = n5033 & ~n41681 ;
  assign n41683 = n14049 | n39683 ;
  assign n41684 = n41683 ^ n24319 ^ 1'b0 ;
  assign n41685 = n7447 | n10411 ;
  assign n41686 = n8767 & ~n41685 ;
  assign n41687 = n14554 & ~n29259 ;
  assign n41688 = n41687 ^ n13921 ^ 1'b0 ;
  assign n41693 = n283 & n2326 ;
  assign n41694 = n41693 ^ n8498 ^ 1'b0 ;
  assign n41689 = n1704 ^ n607 ^ 1'b0 ;
  assign n41690 = n73 | n41689 ;
  assign n41691 = n31835 ^ n23520 ^ n3234 ;
  assign n41692 = n41690 | n41691 ;
  assign n41695 = n41694 ^ n41692 ^ 1'b0 ;
  assign n41696 = n41695 ^ n8206 ^ 1'b0 ;
  assign n41697 = n24758 ^ n6277 ^ 1'b0 ;
  assign n41698 = n18826 | n24130 ;
  assign n41699 = n41698 ^ n8943 ^ 1'b0 ;
  assign n41700 = ~n17956 & n41699 ;
  assign n41701 = n18240 & n41700 ;
  assign n41702 = n41701 ^ n19169 ^ 1'b0 ;
  assign n41703 = n38073 ^ n9384 ^ n6236 ;
  assign n41704 = n40895 ^ n4290 ^ 1'b0 ;
  assign n41705 = ~n41703 & n41704 ;
  assign n41706 = n34990 ^ n14611 ^ n4741 ;
  assign n41707 = n11346 ^ n2428 ^ 1'b0 ;
  assign n41708 = n32794 ^ n11137 ^ 1'b0 ;
  assign n41709 = n5949 | n41708 ;
  assign n41710 = n41709 ^ n10241 ^ 1'b0 ;
  assign n41711 = ~n13708 & n22095 ;
  assign n41712 = n39798 & n41711 ;
  assign n41713 = n1353 & n19345 ;
  assign n41714 = n41713 ^ n24543 ^ 1'b0 ;
  assign n41715 = n41714 ^ n34993 ^ n7520 ;
  assign n41716 = n41715 ^ n6699 ^ 1'b0 ;
  assign n41717 = n99 & ~n24063 ;
  assign n41718 = ( n13689 & n26798 ) | ( n13689 & n41717 ) | ( n26798 & n41717 ) ;
  assign n41719 = ~n8851 & n17807 ;
  assign n41720 = ~n1341 & n9989 ;
  assign n41721 = n41720 ^ n13010 ^ 1'b0 ;
  assign n41722 = n607 ^ n293 ^ 1'b0 ;
  assign n41723 = ~n8147 & n41722 ;
  assign n41724 = n21809 ^ n8977 ^ 1'b0 ;
  assign n41725 = n41723 & n41724 ;
  assign n41726 = n9485 & ~n38168 ;
  assign n41727 = n41726 ^ n26815 ^ 1'b0 ;
  assign n41728 = n18162 ^ n7771 ^ 1'b0 ;
  assign n41729 = n3508 & ~n10754 ;
  assign n41730 = n16006 ^ n9437 ^ 1'b0 ;
  assign n41731 = n37541 & ~n41730 ;
  assign n41732 = ~n11748 & n33072 ;
  assign n41733 = n41732 ^ n8397 ^ 1'b0 ;
  assign n41734 = n17909 ^ n13870 ^ 1'b0 ;
  assign n41735 = n41443 & ~n41734 ;
  assign n41736 = n41735 ^ n12209 ^ 1'b0 ;
  assign n41737 = ~n11868 & n23975 ;
  assign n41738 = n13752 & ~n27543 ;
  assign n41739 = n3551 & ~n5329 ;
  assign n41740 = n13275 ^ n9116 ^ 1'b0 ;
  assign n41741 = ( n346 & n31533 ) | ( n346 & ~n41740 ) | ( n31533 & ~n41740 ) ;
  assign n41742 = n7037 | n41741 ;
  assign n41743 = ~n9655 & n28792 ;
  assign n41744 = n41743 ^ n15080 ^ 1'b0 ;
  assign n41745 = n7020 | n30901 ;
  assign n41746 = n41745 ^ n19545 ^ 1'b0 ;
  assign n41747 = n3717 & n41746 ;
  assign n41748 = ~n38030 & n41747 ;
  assign n41749 = n32777 ^ n24980 ^ n2573 ;
  assign n41750 = n41749 ^ n24157 ^ 1'b0 ;
  assign n41751 = n5941 | n41750 ;
  assign n41752 = n41748 & ~n41751 ;
  assign n41753 = n13326 ^ n4914 ^ 1'b0 ;
  assign n41754 = n5562 & ~n17833 ;
  assign n41755 = ~n20332 & n41754 ;
  assign n41756 = ( n10780 & ~n13751 ) | ( n10780 & n26099 ) | ( ~n13751 & n26099 ) ;
  assign n41757 = n38717 ^ n32686 ^ 1'b0 ;
  assign n41758 = n18912 ^ n6550 ^ 1'b0 ;
  assign n41759 = n16321 | n41758 ;
  assign n41760 = n41759 ^ n41271 ^ 1'b0 ;
  assign n41762 = ( n14425 & n16480 ) | ( n14425 & ~n20662 ) | ( n16480 & ~n20662 ) ;
  assign n41761 = n4732 | n24288 ;
  assign n41763 = n41762 ^ n41761 ^ 1'b0 ;
  assign n41764 = n27340 & ~n31703 ;
  assign n41765 = ~n32376 & n41764 ;
  assign n41766 = n41765 ^ n10055 ^ 1'b0 ;
  assign n41767 = ~n6445 & n22964 ;
  assign n41769 = n25560 ^ n19246 ^ 1'b0 ;
  assign n41770 = n27995 ^ n10820 ^ n4093 ;
  assign n41771 = n41769 & n41770 ;
  assign n41772 = n41771 ^ n27452 ^ n4291 ;
  assign n41768 = n2023 | n40143 ;
  assign n41773 = n41772 ^ n41768 ^ 1'b0 ;
  assign n41774 = n17561 & n19982 ;
  assign n41775 = n30079 & n41774 ;
  assign n41776 = ( n3793 & n28185 ) | ( n3793 & n31863 ) | ( n28185 & n31863 ) ;
  assign n41777 = ~n41775 & n41776 ;
  assign n41778 = n41775 & n41777 ;
  assign n41779 = ~n14539 & n15610 ;
  assign n41780 = ~n31760 & n41779 ;
  assign n41781 = n30366 ^ n12527 ^ 1'b0 ;
  assign n41782 = ~n3634 & n41781 ;
  assign n41783 = n10084 | n15101 ;
  assign n41784 = n31070 | n41783 ;
  assign n41785 = n13636 & n41784 ;
  assign n41786 = n41785 ^ n2650 ^ 1'b0 ;
  assign n41787 = n960 & ~n1634 ;
  assign n41788 = n41787 ^ n38562 ^ 1'b0 ;
  assign n41789 = n17008 ^ n13977 ^ n59 ;
  assign n41790 = n41789 ^ n36986 ^ n12554 ;
  assign n41791 = n1995 & n16556 ;
  assign n41792 = n1628 | n41791 ;
  assign n41793 = n41792 ^ n30895 ^ 1'b0 ;
  assign n41794 = n10145 ^ n4830 ^ 1'b0 ;
  assign n41795 = n12358 & n41794 ;
  assign n41796 = n25155 ^ n1487 ^ 1'b0 ;
  assign n41797 = n41795 & ~n41796 ;
  assign n41798 = n10720 & n41797 ;
  assign n41799 = n41798 ^ n7941 ^ 1'b0 ;
  assign n41800 = ( ~n2225 & n9995 ) | ( ~n2225 & n18015 ) | ( n9995 & n18015 ) ;
  assign n41801 = n18458 | n41800 ;
  assign n41802 = n40800 & ~n41801 ;
  assign n41803 = ~n25242 & n26281 ;
  assign n41804 = n34649 & n41803 ;
  assign n41805 = n38528 ^ n3665 ^ n612 ;
  assign n41806 = ~n7804 & n10063 ;
  assign n41807 = n17643 & n25059 ;
  assign n41808 = n17402 & n22929 ;
  assign n41809 = n9269 ^ n8527 ^ 1'b0 ;
  assign n41810 = ~n41808 & n41809 ;
  assign n41811 = n36634 & n41810 ;
  assign n41812 = n12340 ^ n4760 ^ 1'b0 ;
  assign n41813 = n41812 ^ n26132 ^ 1'b0 ;
  assign n41814 = n26829 & ~n41813 ;
  assign n41815 = ~n7768 & n10983 ;
  assign n41816 = ~n4752 & n41815 ;
  assign n41817 = n33849 | n41816 ;
  assign n41818 = n4574 & ~n30339 ;
  assign n41819 = n1868 | n41818 ;
  assign n41820 = n1868 & ~n41819 ;
  assign n41821 = n21846 | n41820 ;
  assign n41822 = n41820 & ~n41821 ;
  assign n41823 = n34859 ^ n20695 ^ 1'b0 ;
  assign n41824 = n12349 & ~n30538 ;
  assign n41825 = n14409 & n41824 ;
  assign n41826 = n8175 & ~n11986 ;
  assign n41827 = n41825 & n41826 ;
  assign n41828 = n41827 ^ n1688 ^ 1'b0 ;
  assign n41829 = ~n5339 & n16342 ;
  assign n41830 = n41829 ^ n28014 ^ 1'b0 ;
  assign n41831 = n23942 ^ n3365 ^ 1'b0 ;
  assign n41832 = n31251 ^ n28498 ^ 1'b0 ;
  assign n41833 = n5265 & ~n41832 ;
  assign n41834 = n21728 & n41833 ;
  assign n41835 = n6817 ^ n4536 ^ 1'b0 ;
  assign n41836 = n24345 & ~n27024 ;
  assign n41837 = n5003 | n41836 ;
  assign n41838 = n8249 & n31664 ;
  assign n41839 = n41838 ^ n1800 ^ 1'b0 ;
  assign n41840 = n15378 ^ n621 ^ 1'b0 ;
  assign n41841 = n17308 & ~n41840 ;
  assign n41842 = ~n4584 & n23014 ;
  assign n41843 = n471 & ~n28872 ;
  assign n41844 = n265 | n5311 ;
  assign n41845 = n19433 & ~n41844 ;
  assign n41846 = n34228 ^ n1135 ^ 1'b0 ;
  assign n41847 = n3970 & n41846 ;
  assign n41848 = n23723 & n26979 ;
  assign n41849 = n1305 & ~n15459 ;
  assign n41850 = n41849 ^ n788 ^ 1'b0 ;
  assign n41852 = n8509 ^ n6041 ^ 1'b0 ;
  assign n41851 = n7882 | n27128 ;
  assign n41853 = n41852 ^ n41851 ^ 1'b0 ;
  assign n41854 = n6978 | n27984 ;
  assign n41855 = n32759 ^ n16261 ^ 1'b0 ;
  assign n41856 = n9490 | n41855 ;
  assign n41857 = n41856 ^ n32159 ^ 1'b0 ;
  assign n41858 = n41854 & ~n41857 ;
  assign n41859 = ~n14009 & n41858 ;
  assign n41860 = n15897 ^ n8636 ^ 1'b0 ;
  assign n41861 = n36311 & n41860 ;
  assign n41862 = n10118 & ~n12211 ;
  assign n41863 = n41862 ^ n19363 ^ 1'b0 ;
  assign n41864 = n21381 | n37648 ;
  assign n41865 = n7804 & ~n15109 ;
  assign n41866 = ~n1079 & n41865 ;
  assign n41867 = n18773 ^ n17906 ^ n301 ;
  assign n41868 = ( ~n2801 & n41866 ) | ( ~n2801 & n41867 ) | ( n41866 & n41867 ) ;
  assign n41869 = n542 & ~n19650 ;
  assign n41870 = n10467 ^ n2990 ^ 1'b0 ;
  assign n41871 = n16942 | n41870 ;
  assign n41872 = n2146 | n41871 ;
  assign n41878 = n5277 ^ n263 ^ 1'b0 ;
  assign n41873 = n15784 ^ n2745 ^ 1'b0 ;
  assign n41874 = n20845 | n41873 ;
  assign n41875 = ~n383 & n30082 ;
  assign n41876 = n41874 & n41875 ;
  assign n41877 = n1496 & ~n41876 ;
  assign n41879 = n41878 ^ n41877 ^ 1'b0 ;
  assign n41880 = ~n15886 & n30389 ;
  assign n41881 = n33917 & n41880 ;
  assign n41882 = n231 | n25919 ;
  assign n41883 = n41882 ^ n27816 ^ 1'b0 ;
  assign n41884 = n5003 & n41883 ;
  assign n41885 = n2152 | n4135 ;
  assign n41886 = ( n12695 & ~n20014 ) | ( n12695 & n41885 ) | ( ~n20014 & n41885 ) ;
  assign n41887 = n30924 ^ n16853 ^ 1'b0 ;
  assign n41888 = ~n4025 & n41887 ;
  assign n41889 = n12626 & n27293 ;
  assign n41890 = n36958 ^ n28795 ^ n8558 ;
  assign n41891 = ~n9630 & n17800 ;
  assign n41892 = n34144 ^ n17736 ^ 1'b0 ;
  assign n41893 = n4339 & ~n15138 ;
  assign n41894 = n4795 & n41893 ;
  assign n41895 = ~n19098 & n29474 ;
  assign n41896 = n38811 ^ n11226 ^ 1'b0 ;
  assign n41897 = n41895 & n41896 ;
  assign n41898 = n18571 ^ n6673 ^ n6289 ;
  assign n41899 = n41898 ^ n27104 ^ 1'b0 ;
  assign n41900 = ( n4877 & ~n29194 ) | ( n4877 & n41899 ) | ( ~n29194 & n41899 ) ;
  assign n41901 = n4378 & n5240 ;
  assign n41902 = n34153 & n39680 ;
  assign n41903 = ( n4105 & ~n12143 ) | ( n4105 & n41902 ) | ( ~n12143 & n41902 ) ;
  assign n41904 = n28817 | n41903 ;
  assign n41908 = n5815 ^ n4431 ^ 1'b0 ;
  assign n41905 = n2745 | n10329 ;
  assign n41906 = n7365 | n41905 ;
  assign n41907 = n41906 ^ n18466 ^ 1'b0 ;
  assign n41909 = n41908 ^ n41907 ^ 1'b0 ;
  assign n41910 = ~n4742 & n14240 ;
  assign n41911 = n41910 ^ n21705 ^ 1'b0 ;
  assign n41912 = n6570 & ~n35140 ;
  assign n41913 = n11194 ^ n2418 ^ 1'b0 ;
  assign n41914 = n10852 | n41913 ;
  assign n41915 = n7587 & ~n13354 ;
  assign n41916 = n12180 & n41915 ;
  assign n41917 = n3415 & n14503 ;
  assign n41918 = n20311 & n41917 ;
  assign n41919 = n29880 & ~n41918 ;
  assign n41920 = n16233 ^ n2606 ^ 1'b0 ;
  assign n41921 = n102 & ~n41920 ;
  assign n41922 = n20942 & ~n41921 ;
  assign n41923 = ( n13198 & n21861 ) | ( n13198 & ~n34174 ) | ( n21861 & ~n34174 ) ;
  assign n41924 = n780 | n41923 ;
  assign n41925 = n41924 ^ x6 ^ 1'b0 ;
  assign n41926 = ~n41922 & n41925 ;
  assign n41927 = n1368 | n12421 ;
  assign n41928 = ~n10883 & n28945 ;
  assign n41929 = n4948 & ~n9939 ;
  assign n41930 = n134 & ~n5882 ;
  assign n41931 = n7882 & n41930 ;
  assign n41932 = n16717 | n41931 ;
  assign n41933 = n6442 | n41932 ;
  assign n41934 = n11777 ^ n9805 ^ 1'b0 ;
  assign n41935 = n12991 & ~n41934 ;
  assign n41936 = n35136 ^ n17323 ^ 1'b0 ;
  assign n41937 = ~n13771 & n36707 ;
  assign n41938 = ~n36707 & n41937 ;
  assign n41939 = n41938 ^ n33058 ^ 1'b0 ;
  assign n41940 = n41939 ^ n3428 ^ 1'b0 ;
  assign n41941 = ~n16829 & n18690 ;
  assign n41942 = ~n26656 & n41941 ;
  assign n41943 = n30637 ^ n23670 ^ 1'b0 ;
  assign n41944 = n27927 & n41943 ;
  assign n41945 = n41944 ^ n12178 ^ 1'b0 ;
  assign n41946 = n41942 & ~n41945 ;
  assign n41947 = n19097 & ~n37664 ;
  assign n41948 = n16089 & n41947 ;
  assign n41949 = ~n24041 & n41948 ;
  assign n41950 = n41949 ^ n26051 ^ 1'b0 ;
  assign n41951 = n11123 | n16445 ;
  assign n41952 = ( n4847 & n13879 ) | ( n4847 & ~n35301 ) | ( n13879 & ~n35301 ) ;
  assign n41953 = ~n26440 & n41952 ;
  assign n41955 = n35904 ^ n31369 ^ 1'b0 ;
  assign n41954 = n17863 | n20688 ;
  assign n41956 = n41955 ^ n41954 ^ 1'b0 ;
  assign n41957 = ( n13771 & ~n38787 ) | ( n13771 & n39943 ) | ( ~n38787 & n39943 ) ;
  assign n41958 = n31636 ^ n7729 ^ n2797 ;
  assign n41959 = n24481 ^ n6866 ^ 1'b0 ;
  assign n41960 = ~n4503 & n32573 ;
  assign n41961 = ~n8463 & n41960 ;
  assign n41962 = n39994 ^ n11213 ^ n2617 ;
  assign n41963 = n39231 ^ n5418 ^ n3404 ;
  assign n41964 = n11542 | n31491 ;
  assign n41965 = n7747 | n41964 ;
  assign n41966 = n41965 ^ n4678 ^ 1'b0 ;
  assign n41967 = n17909 ^ n13721 ^ 1'b0 ;
  assign n41968 = ~n15401 & n41967 ;
  assign n41969 = n9621 ^ n2511 ^ 1'b0 ;
  assign n41970 = n34508 & n41969 ;
  assign n41971 = n28635 & n41970 ;
  assign n41972 = n41971 ^ n33775 ^ 1'b0 ;
  assign n41973 = n22191 & ~n41972 ;
  assign n41974 = n31692 ^ n5484 ^ 1'b0 ;
  assign n41975 = ~n13862 & n28819 ;
  assign n41976 = ~n1996 & n5175 ;
  assign n41977 = ~n19334 & n28455 ;
  assign n41978 = ~n41976 & n41977 ;
  assign n41979 = n32972 ^ n10994 ^ n8397 ;
  assign n41980 = n41979 ^ n32124 ^ 1'b0 ;
  assign n41981 = n41978 | n41980 ;
  assign n41982 = n22440 ^ n4760 ^ 1'b0 ;
  assign n41983 = n27878 & n41982 ;
  assign n41984 = n36021 & n41983 ;
  assign n41985 = n41984 ^ n20734 ^ 1'b0 ;
  assign n41986 = n5639 & ~n41985 ;
  assign n41987 = n12588 | n17838 ;
  assign n41988 = ( n3554 & n5911 ) | ( n3554 & n29704 ) | ( n5911 & n29704 ) ;
  assign n41989 = ( ~n3557 & n24001 ) | ( ~n3557 & n41988 ) | ( n24001 & n41988 ) ;
  assign n41990 = n17994 ^ n13678 ^ 1'b0 ;
  assign n41991 = n25957 | n41990 ;
  assign n41992 = n14802 ^ n1721 ^ 1'b0 ;
  assign n41993 = n9463 & ~n41436 ;
  assign n41994 = n41992 & n41993 ;
  assign n41995 = n37652 ^ n37278 ^ n21918 ;
  assign n41996 = n18690 ^ n15979 ^ n1105 ;
  assign n41997 = n7956 | n41996 ;
  assign n41998 = ~n16545 & n30907 ;
  assign n41999 = n2815 & n41998 ;
  assign n42000 = n41999 ^ n10929 ^ 1'b0 ;
  assign n42001 = n10344 ^ n9941 ^ 1'b0 ;
  assign n42002 = n7406 & n42001 ;
  assign n42003 = n42002 ^ n33406 ^ 1'b0 ;
  assign n42004 = n37912 | n42003 ;
  assign n42005 = n2486 | n33644 ;
  assign n42006 = n34684 & ~n42005 ;
  assign n42007 = n42006 ^ n17508 ^ 1'b0 ;
  assign n42008 = n14632 & n42007 ;
  assign n42009 = n15781 & n25194 ;
  assign n42010 = ~n42008 & n42009 ;
  assign n42013 = n8998 & n17999 ;
  assign n42011 = n13331 ^ n437 ^ 1'b0 ;
  assign n42012 = ~n12162 & n42011 ;
  assign n42014 = n42013 ^ n42012 ^ n32891 ;
  assign n42015 = n42014 ^ n11516 ^ 1'b0 ;
  assign n42016 = n18363 ^ n8193 ^ 1'b0 ;
  assign n42017 = n11251 | n42016 ;
  assign n42018 = n15537 & ~n20382 ;
  assign n42019 = n30472 & n42018 ;
  assign n42020 = ~n29390 & n39920 ;
  assign n42021 = n8426 & n42020 ;
  assign n42022 = n8826 ^ n6375 ^ 1'b0 ;
  assign n42023 = n12861 | n42022 ;
  assign n42024 = n42023 ^ n2736 ^ 1'b0 ;
  assign n42025 = ~n28108 & n42024 ;
  assign n42026 = n1509 | n42025 ;
  assign n42027 = n8277 | n37031 ;
  assign n42028 = n21694 ^ n11107 ^ 1'b0 ;
  assign n42029 = n4569 & ~n24235 ;
  assign n42030 = n31258 ^ n11763 ^ n6582 ;
  assign n42031 = n11672 & n15396 ;
  assign n42032 = n42030 & n42031 ;
  assign n42033 = n42032 ^ n7028 ^ 1'b0 ;
  assign n42034 = n1082 & n20925 ;
  assign n42035 = n3761 & n42034 ;
  assign n42036 = n7600 & n25425 ;
  assign n42037 = n42036 ^ n37393 ^ 1'b0 ;
  assign n42038 = n29177 ^ n22304 ^ 1'b0 ;
  assign n42039 = n4105 & ~n42038 ;
  assign n42040 = ( n1238 & ~n1628 ) | ( n1238 & n5481 ) | ( ~n1628 & n5481 ) ;
  assign n42041 = n17079 ^ n3620 ^ 1'b0 ;
  assign n42042 = n42040 & n42041 ;
  assign n42043 = ~n42039 & n42042 ;
  assign n42044 = n6167 | n42043 ;
  assign n42045 = n39455 | n42044 ;
  assign n42046 = n12984 | n42045 ;
  assign n42047 = ( n3745 & n14833 ) | ( n3745 & n23075 ) | ( n14833 & n23075 ) ;
  assign n42048 = n42047 ^ n40648 ^ n8539 ;
  assign n42049 = n28235 & ~n28857 ;
  assign n42050 = n20614 & n21290 ;
  assign n42051 = n4922 & n28520 ;
  assign n42052 = n21355 & ~n22381 ;
  assign n42053 = n30558 & n42052 ;
  assign n42054 = n19771 ^ n8382 ^ n5318 ;
  assign n42055 = ( n13760 & n19580 ) | ( n13760 & n37531 ) | ( n19580 & n37531 ) ;
  assign n42056 = ~n30685 & n42055 ;
  assign n42057 = ~n3997 & n4769 ;
  assign n42058 = n42057 ^ n10263 ^ 1'b0 ;
  assign n42059 = n10341 & n15194 ;
  assign n42060 = ~n40251 & n42059 ;
  assign n42067 = n9221 ^ n7559 ^ 1'b0 ;
  assign n42064 = ( n3564 & ~n23392 ) | ( n3564 & n38296 ) | ( ~n23392 & n38296 ) ;
  assign n42061 = n29119 & n32276 ;
  assign n42062 = n11633 | n42061 ;
  assign n42063 = n16154 | n42062 ;
  assign n42065 = n42064 ^ n42063 ^ 1'b0 ;
  assign n42066 = n7055 & n42065 ;
  assign n42068 = n42067 ^ n42066 ^ 1'b0 ;
  assign n42069 = n5699 & n25372 ;
  assign n42070 = ~n3959 & n42069 ;
  assign n42077 = n17418 ^ n4115 ^ 1'b0 ;
  assign n42071 = n6808 ^ n2556 ^ 1'b0 ;
  assign n42072 = n11220 & ~n42071 ;
  assign n42073 = ~n9050 & n42072 ;
  assign n42074 = n119 & n127 ;
  assign n42075 = ~n42073 & n42074 ;
  assign n42076 = n23295 & ~n42075 ;
  assign n42078 = n42077 ^ n42076 ^ 1'b0 ;
  assign n42079 = ~n1182 & n5437 ;
  assign n42080 = ( n27149 & ~n31320 ) | ( n27149 & n42079 ) | ( ~n31320 & n42079 ) ;
  assign n42081 = n22379 ^ n7163 ^ 1'b0 ;
  assign n42082 = n15244 & n42081 ;
  assign n42083 = ~n27840 & n42082 ;
  assign n42084 = n6491 | n17818 ;
  assign n42085 = n42084 ^ n31784 ^ 1'b0 ;
  assign n42086 = n30805 & n42085 ;
  assign n42087 = n37916 & n39762 ;
  assign n42088 = ~n36343 & n42087 ;
  assign n42089 = n16666 ^ n1903 ^ 1'b0 ;
  assign n42090 = n10738 & ~n41444 ;
  assign n42095 = n36 & ~n4186 ;
  assign n42091 = ~n17602 & n20295 ;
  assign n42092 = n42091 ^ n10721 ^ 1'b0 ;
  assign n42093 = n42092 ^ n39735 ^ 1'b0 ;
  assign n42094 = n22250 | n42093 ;
  assign n42096 = n42095 ^ n42094 ^ 1'b0 ;
  assign n42097 = n4789 & n24873 ;
  assign n42098 = n16616 ^ n13858 ^ 1'b0 ;
  assign n42099 = n13859 & ~n42098 ;
  assign n42100 = n36640 & n42099 ;
  assign n42101 = n42097 & n42100 ;
  assign n42102 = n17346 & ~n26405 ;
  assign n42103 = n42102 ^ n24229 ^ 1'b0 ;
  assign n42104 = n34757 & n40823 ;
  assign n42105 = n5837 & ~n11890 ;
  assign n42106 = n42105 ^ n24644 ^ 1'b0 ;
  assign n42107 = ( x8 & n7854 ) | ( x8 & n42106 ) | ( n7854 & n42106 ) ;
  assign n42108 = n9100 & ~n34251 ;
  assign n42109 = n11413 & n42108 ;
  assign n42110 = n42109 ^ n35675 ^ n6473 ;
  assign n42111 = n15872 & n27877 ;
  assign n42112 = ~n5759 & n42111 ;
  assign n42113 = n24110 ^ n12836 ^ 1'b0 ;
  assign n42114 = n42112 | n42113 ;
  assign n42115 = n26956 | n42114 ;
  assign n42116 = n7880 & ~n42115 ;
  assign n42117 = n3087 ^ n2181 ^ 1'b0 ;
  assign n42118 = ~n2841 & n42117 ;
  assign n42119 = n21348 ^ n4993 ^ 1'b0 ;
  assign n42120 = n797 | n2677 ;
  assign n42121 = n42120 ^ n32695 ^ n5634 ;
  assign n42122 = n11072 & n37601 ;
  assign n42123 = n9504 & ~n12893 ;
  assign n42124 = n42123 ^ n29869 ^ 1'b0 ;
  assign n42125 = n3237 & n14934 ;
  assign n42126 = n22761 & n42125 ;
  assign n42127 = n28828 ^ n303 ^ 1'b0 ;
  assign n42128 = n15861 & ~n42127 ;
  assign n42129 = n36621 ^ n3658 ^ 1'b0 ;
  assign n42130 = n18956 ^ n3321 ^ 1'b0 ;
  assign n42131 = ( n22369 & ~n32823 ) | ( n22369 & n42130 ) | ( ~n32823 & n42130 ) ;
  assign n42132 = n8403 & ~n19482 ;
  assign n42133 = n42132 ^ n5653 ^ 1'b0 ;
  assign n42134 = ~n12629 & n20776 ;
  assign n42135 = n3313 & n42134 ;
  assign n42136 = ~n7856 & n30593 ;
  assign n42137 = n27675 & n42136 ;
  assign n42138 = ~n25723 & n42137 ;
  assign n42139 = n6223 ^ n5675 ^ 1'b0 ;
  assign n42140 = n1167 & ~n42139 ;
  assign n42141 = n25323 ^ n3528 ^ 1'b0 ;
  assign n42142 = n42140 & n42141 ;
  assign n42143 = ~n16514 & n42142 ;
  assign n42144 = n35752 ^ n18105 ^ 1'b0 ;
  assign n42152 = n197 & ~n4862 ;
  assign n42153 = ~n13069 & n42152 ;
  assign n42145 = n1400 & ~n23833 ;
  assign n42146 = ~n2126 & n24259 ;
  assign n42147 = n21030 & n42146 ;
  assign n42148 = n42147 ^ n27600 ^ 1'b0 ;
  assign n42149 = n42148 ^ n5290 ^ 1'b0 ;
  assign n42150 = n11355 | n42149 ;
  assign n42151 = n42145 & ~n42150 ;
  assign n42154 = n42153 ^ n42151 ^ 1'b0 ;
  assign n42155 = n30058 & ~n36848 ;
  assign n42156 = n31010 ^ n29268 ^ 1'b0 ;
  assign n42157 = n42156 ^ n19283 ^ 1'b0 ;
  assign n42158 = n36683 ^ n17256 ^ 1'b0 ;
  assign n42159 = n42157 | n42158 ;
  assign n42160 = n33059 ^ n8978 ^ 1'b0 ;
  assign n42161 = ( n16888 & n28876 ) | ( n16888 & n29303 ) | ( n28876 & n29303 ) ;
  assign n42162 = ~n3881 & n30317 ;
  assign n42163 = ( n4688 & ~n42161 ) | ( n4688 & n42162 ) | ( ~n42161 & n42162 ) ;
  assign n42164 = ( n7357 & n19780 ) | ( n7357 & n34775 ) | ( n19780 & n34775 ) ;
  assign n42165 = n28165 & ~n33749 ;
  assign n42166 = n12668 & n36539 ;
  assign n42167 = n23 & n14378 ;
  assign n42168 = n42167 ^ n11558 ^ 1'b0 ;
  assign n42169 = ~n4246 & n42168 ;
  assign n42170 = n42169 ^ n28872 ^ n23771 ;
  assign n42171 = n4773 & ~n13222 ;
  assign n42172 = n24380 ^ n1875 ^ 1'b0 ;
  assign n42173 = ~n1032 & n42172 ;
  assign n42174 = n42173 ^ n4204 ^ 1'b0 ;
  assign n42175 = n38319 ^ n17565 ^ 1'b0 ;
  assign n42176 = n18470 & n42175 ;
  assign n42177 = n1848 & n10379 ;
  assign n42178 = n42177 ^ n17313 ^ 1'b0 ;
  assign n42179 = n12470 ^ n12333 ^ n10829 ;
  assign n42180 = ~n42178 & n42179 ;
  assign n42181 = n42180 ^ n5954 ^ 1'b0 ;
  assign n42182 = n9105 ^ n8002 ^ 1'b0 ;
  assign n42183 = n4773 ^ n2341 ^ 1'b0 ;
  assign n42184 = n14392 & ~n42183 ;
  assign n42185 = n34705 ^ n3120 ^ 1'b0 ;
  assign n42186 = n1627 & ~n42185 ;
  assign n42187 = n1815 & n42186 ;
  assign n42188 = n19596 ^ n19079 ^ 1'b0 ;
  assign n42189 = n6352 & ~n12701 ;
  assign n42190 = ~n12908 & n42189 ;
  assign n42191 = n14961 & n17523 ;
  assign n42192 = ~n601 & n42191 ;
  assign n42193 = n18853 & n42192 ;
  assign n42194 = n1957 | n5706 ;
  assign n42195 = n1898 & n10533 ;
  assign n42196 = n42194 & n42195 ;
  assign n42197 = n1591 ^ n534 ^ 1'b0 ;
  assign n42198 = n42196 | n42197 ;
  assign n42199 = n42198 ^ n23252 ^ 1'b0 ;
  assign n42200 = n4338 & n24014 ;
  assign n42201 = n42200 ^ n26286 ^ 1'b0 ;
  assign n42202 = n8777 & ~n14200 ;
  assign n42203 = n9879 & ~n42202 ;
  assign n42204 = ( n5428 & ~n6396 ) | ( n5428 & n11466 ) | ( ~n6396 & n11466 ) ;
  assign n42205 = n11445 & ~n28945 ;
  assign n42206 = n42204 & n42205 ;
  assign n42207 = n5151 ^ n1340 ^ 1'b0 ;
  assign n42208 = n7657 & ~n20206 ;
  assign n42209 = n12670 & n42208 ;
  assign n42210 = n41590 ^ n2002 ^ 1'b0 ;
  assign n42211 = n318 & n42210 ;
  assign n42212 = ( n12894 & ~n16010 ) | ( n12894 & n20764 ) | ( ~n16010 & n20764 ) ;
  assign n42213 = n42212 ^ n15955 ^ 1'b0 ;
  assign n42214 = n37813 ^ n21365 ^ 1'b0 ;
  assign n42215 = n2479 & n6153 ;
  assign n42216 = n42215 ^ n22917 ^ 1'b0 ;
  assign n42217 = n42216 ^ n17630 ^ 1'b0 ;
  assign n42218 = ( n2508 & ~n5222 ) | ( n2508 & n35882 ) | ( ~n5222 & n35882 ) ;
  assign n42219 = n13338 ^ n7137 ^ 1'b0 ;
  assign n42220 = n42219 ^ n18110 ^ 1'b0 ;
  assign n42221 = ( ~n12887 & n16419 ) | ( ~n12887 & n22422 ) | ( n16419 & n22422 ) ;
  assign n42222 = ( n20430 & n30543 ) | ( n20430 & n42221 ) | ( n30543 & n42221 ) ;
  assign n42223 = ~n23517 & n24051 ;
  assign n42224 = n42223 ^ n3173 ^ 1'b0 ;
  assign n42225 = n3128 & n20396 ;
  assign n42226 = n19032 & n42225 ;
  assign n42227 = n2944 | n42226 ;
  assign n42228 = n42227 ^ n19983 ^ 1'b0 ;
  assign n42229 = n42228 ^ n17938 ^ n12603 ;
  assign n42230 = ( n11100 & ~n42224 ) | ( n11100 & n42229 ) | ( ~n42224 & n42229 ) ;
  assign n42231 = n32331 ^ n16909 ^ 1'b0 ;
  assign n42232 = n14656 & ~n42231 ;
  assign n42233 = n42232 ^ n16737 ^ n4185 ;
  assign n42234 = n12360 ^ n12008 ^ n2982 ;
  assign n42235 = n42234 ^ n17325 ^ n3306 ;
  assign n42236 = n9793 | n41664 ;
  assign n42237 = n42236 ^ n3645 ^ 1'b0 ;
  assign n42238 = n8052 ^ n5342 ^ 1'b0 ;
  assign n42239 = n30240 | n42238 ;
  assign n42240 = n42239 ^ n10814 ^ 1'b0 ;
  assign n42241 = n1529 & n12966 ;
  assign n42242 = n42241 ^ n4872 ^ 1'b0 ;
  assign n42245 = n26624 | n39526 ;
  assign n42246 = n37072 & ~n42245 ;
  assign n42243 = n38697 ^ n25673 ^ 1'b0 ;
  assign n42244 = n40264 & ~n42243 ;
  assign n42247 = n42246 ^ n42244 ^ 1'b0 ;
  assign n42248 = n139 | n36361 ;
  assign n42249 = n1613 & ~n42248 ;
  assign n42250 = n935 & ~n1170 ;
  assign n42251 = n42250 ^ n2326 ^ 1'b0 ;
  assign n42252 = ( ~n16138 & n28855 ) | ( ~n16138 & n42251 ) | ( n28855 & n42251 ) ;
  assign n42254 = n19491 ^ n12715 ^ 1'b0 ;
  assign n42253 = n21868 ^ n4431 ^ 1'b0 ;
  assign n42255 = n42254 ^ n42253 ^ 1'b0 ;
  assign n42256 = n38896 ^ n10685 ^ 1'b0 ;
  assign n42258 = n22477 & ~n28290 ;
  assign n42259 = ~n11233 & n42258 ;
  assign n42257 = n471 | n13626 ;
  assign n42260 = n42259 ^ n42257 ^ 1'b0 ;
  assign n42261 = n33788 ^ n12439 ^ 1'b0 ;
  assign n42262 = n15441 | n42261 ;
  assign n42263 = n42262 ^ n28944 ^ n23941 ;
  assign n42264 = n20426 ^ n15846 ^ n3713 ;
  assign n42265 = n6348 & ~n42264 ;
  assign n42266 = n42265 ^ n27024 ^ 1'b0 ;
  assign n42267 = ~n177 & n6143 ;
  assign n42268 = n42267 ^ n37907 ^ 1'b0 ;
  assign n42269 = n42268 ^ n10512 ^ 1'b0 ;
  assign n42270 = n42269 ^ n3817 ^ n878 ;
  assign n42271 = n42270 ^ n39544 ^ n17224 ;
  assign n42272 = n31070 ^ n22437 ^ 1'b0 ;
  assign n42273 = n12233 & n41106 ;
  assign n42274 = n1344 | n42273 ;
  assign n42275 = n350 & ~n5844 ;
  assign n42276 = n30589 ^ n6629 ^ 1'b0 ;
  assign n42277 = n3123 & n42276 ;
  assign n42278 = n42277 ^ n2735 ^ 1'b0 ;
  assign n42279 = n2055 | n42278 ;
  assign n42282 = n22945 | n32157 ;
  assign n42283 = n42282 ^ n25555 ^ 1'b0 ;
  assign n42280 = n39357 ^ n10282 ^ n572 ;
  assign n42281 = n23258 & ~n42280 ;
  assign n42284 = n42283 ^ n42281 ^ 1'b0 ;
  assign n42285 = n4704 & ~n17510 ;
  assign n42286 = n21520 ^ n13565 ^ 1'b0 ;
  assign n42287 = n1779 | n6825 ;
  assign n42288 = n2363 | n42287 ;
  assign n42289 = n42288 ^ n1040 ^ 1'b0 ;
  assign n42293 = n3156 & ~n19493 ;
  assign n42294 = ~n8486 & n42293 ;
  assign n42290 = ~n4263 & n9716 ;
  assign n42291 = ~n5346 & n42290 ;
  assign n42292 = n40691 & ~n42291 ;
  assign n42295 = n42294 ^ n42292 ^ 1'b0 ;
  assign n42296 = ( n6262 & ~n11042 ) | ( n6262 & n14624 ) | ( ~n11042 & n14624 ) ;
  assign n42297 = n36683 ^ n26778 ^ 1'b0 ;
  assign n42298 = n11723 ^ n8759 ^ 1'b0 ;
  assign n42299 = n860 & ~n42298 ;
  assign n42300 = n42299 ^ n8662 ^ 1'b0 ;
  assign n42301 = ( n3422 & ~n4091 ) | ( n3422 & n33115 ) | ( ~n4091 & n33115 ) ;
  assign n42302 = n42301 ^ n19352 ^ 1'b0 ;
  assign n42303 = n5324 & ~n29578 ;
  assign n42304 = ( n4067 & n10861 ) | ( n4067 & n11672 ) | ( n10861 & n11672 ) ;
  assign n42305 = n42304 ^ n12296 ^ n9757 ;
  assign n42306 = n42305 ^ n14177 ^ 1'b0 ;
  assign n42307 = ( n1010 & ~n2135 ) | ( n1010 & n8829 ) | ( ~n2135 & n8829 ) ;
  assign n42308 = ~n6614 & n6762 ;
  assign n42309 = n19982 & ~n42308 ;
  assign n42310 = n5242 & n28419 ;
  assign n42311 = ~n5924 & n27909 ;
  assign n42312 = n42311 ^ n20056 ^ 1'b0 ;
  assign n42313 = n32680 ^ n11440 ^ 1'b0 ;
  assign n42314 = n304 | n42313 ;
  assign n42315 = ~n5239 & n9300 ;
  assign n42316 = n19203 | n20196 ;
  assign n42317 = ~n9765 & n17740 ;
  assign n42318 = n11877 & ~n42317 ;
  assign n42319 = n26586 & n42318 ;
  assign n42320 = ( n13374 & ~n16801 ) | ( n13374 & n38852 ) | ( ~n16801 & n38852 ) ;
  assign n42321 = n6966 | n38551 ;
  assign n42322 = n20351 & ~n42321 ;
  assign n42323 = n7225 | n42322 ;
  assign n42324 = n8566 & n42323 ;
  assign n42325 = n42324 ^ n33703 ^ 1'b0 ;
  assign n42326 = n7639 & ~n12681 ;
  assign n42327 = n8751 & n42326 ;
  assign n42328 = n19354 & n42327 ;
  assign n42329 = n38204 & n42328 ;
  assign n42330 = ~n7008 & n33646 ;
  assign n42331 = ~n16812 & n17848 ;
  assign n42332 = n28904 ^ n17302 ^ 1'b0 ;
  assign n42333 = n26171 | n42332 ;
  assign n42337 = n1836 | n24984 ;
  assign n42338 = n42337 ^ n25283 ^ 1'b0 ;
  assign n42339 = n42338 ^ n6487 ^ 1'b0 ;
  assign n42334 = ~n19189 & n23065 ;
  assign n42335 = ~n11094 & n42334 ;
  assign n42336 = n42335 ^ n25707 ^ 1'b0 ;
  assign n42340 = n42339 ^ n42336 ^ n2766 ;
  assign n42341 = n13620 | n20111 ;
  assign n42342 = n42341 ^ n17042 ^ 1'b0 ;
  assign n42343 = n37379 & n41292 ;
  assign n42344 = n18319 ^ n14197 ^ 1'b0 ;
  assign n42345 = n2566 & n42344 ;
  assign n42348 = n1808 & ~n30634 ;
  assign n42346 = n20250 ^ n8446 ^ 1'b0 ;
  assign n42347 = n32573 & n42346 ;
  assign n42349 = n42348 ^ n42347 ^ 1'b0 ;
  assign n42350 = ~n1351 & n29140 ;
  assign n42353 = n22131 ^ n6343 ^ 1'b0 ;
  assign n42352 = n31070 ^ n22956 ^ n12591 ;
  assign n42351 = n7523 | n17214 ;
  assign n42354 = n42353 ^ n42352 ^ n42351 ;
  assign n42355 = n4207 & ~n38007 ;
  assign n42356 = n42355 ^ n13580 ^ 1'b0 ;
  assign n42357 = n13312 & n31862 ;
  assign n42358 = n42357 ^ n4405 ^ 1'b0 ;
  assign n42359 = n5175 ^ n2569 ^ 1'b0 ;
  assign n42360 = n3578 | n42359 ;
  assign n42361 = n42360 ^ n18534 ^ n7070 ;
  assign n42362 = n37029 ^ n19226 ^ 1'b0 ;
  assign n42363 = ~n4372 & n39334 ;
  assign n42364 = n21054 | n32530 ;
  assign n42366 = n19360 & ~n21510 ;
  assign n42367 = n42366 ^ n8046 ^ 1'b0 ;
  assign n42368 = ( n9263 & n14067 ) | ( n9263 & ~n42367 ) | ( n14067 & ~n42367 ) ;
  assign n42365 = ~n19009 & n20038 ;
  assign n42369 = n42368 ^ n42365 ^ 1'b0 ;
  assign n42370 = n17175 & n17378 ;
  assign n42371 = n7368 & n42370 ;
  assign n42372 = n1397 | n42371 ;
  assign n42373 = n42372 ^ n20819 ^ 1'b0 ;
  assign n42374 = n21328 & ~n42373 ;
  assign n42375 = n42374 ^ n40266 ^ 1'b0 ;
  assign n42376 = n5977 | n14847 ;
  assign n42377 = n9683 & ~n42376 ;
  assign n42378 = n42377 ^ n3214 ^ 1'b0 ;
  assign n42379 = n33584 ^ n25242 ^ n17792 ;
  assign n42380 = n19343 | n20057 ;
  assign n42381 = n20392 & n25135 ;
  assign n42382 = n42381 ^ n34111 ^ n11162 ;
  assign n42383 = n13539 & ~n20364 ;
  assign n42384 = n42383 ^ n20294 ^ 1'b0 ;
  assign n42385 = n4226 & ~n20237 ;
  assign n42386 = n37670 & n42385 ;
  assign n42387 = n30331 ^ n27055 ^ 1'b0 ;
  assign n42388 = n25957 ^ n24058 ^ 1'b0 ;
  assign n42389 = n9076 | n42388 ;
  assign n42390 = n20299 & ~n23035 ;
  assign n42391 = n28161 & n42390 ;
  assign n42392 = ~n9224 & n20295 ;
  assign n42393 = n42392 ^ n24797 ^ 1'b0 ;
  assign n42394 = ( n14007 & n15693 ) | ( n14007 & ~n42393 ) | ( n15693 & ~n42393 ) ;
  assign n42395 = n2313 & ~n29000 ;
  assign n42396 = n10465 ^ n2580 ^ 1'b0 ;
  assign n42397 = n11118 ^ n8379 ^ 1'b0 ;
  assign n42398 = n22315 ^ n3135 ^ 1'b0 ;
  assign n42399 = n3730 & n9586 ;
  assign n42400 = n22645 ^ n9614 ^ 1'b0 ;
  assign n42401 = ~n557 & n20638 ;
  assign n42402 = n42401 ^ n30478 ^ 1'b0 ;
  assign n42403 = n17459 ^ n15228 ^ 1'b0 ;
  assign n42404 = ~n10407 & n17875 ;
  assign n42405 = n42403 & n42404 ;
  assign n42406 = n16830 | n42405 ;
  assign n42407 = ~n3027 & n10094 ;
  assign n42408 = ~n4416 & n36831 ;
  assign n42409 = n42408 ^ n39049 ^ 1'b0 ;
  assign n42410 = n11548 & ~n31035 ;
  assign n42411 = n28641 ^ n9146 ^ 1'b0 ;
  assign n42412 = n11935 & n42411 ;
  assign n42413 = n42410 & n42412 ;
  assign n42414 = n27514 ^ n18486 ^ 1'b0 ;
  assign n42415 = n42413 & n42414 ;
  assign n42416 = n30244 ^ n18272 ^ 1'b0 ;
  assign n42417 = n17499 | n42416 ;
  assign n42418 = n14824 ^ n13329 ^ 1'b0 ;
  assign n42419 = ~n8103 & n19155 ;
  assign n42420 = n16000 ^ n12383 ^ 1'b0 ;
  assign n42421 = n4165 & ~n9678 ;
  assign n42422 = n17973 ^ n299 ^ 1'b0 ;
  assign n42423 = n3784 | n42422 ;
  assign n42424 = n32372 | n42423 ;
  assign n42425 = n4105 & n42424 ;
  assign n42426 = n36346 & n42425 ;
  assign n42427 = ~n16232 & n29769 ;
  assign n42428 = n25111 ^ n11185 ^ 1'b0 ;
  assign n42429 = n6139 & ~n24394 ;
  assign n42430 = n31418 & n42429 ;
  assign n42431 = n17939 ^ n2147 ^ 1'b0 ;
  assign n42432 = ~n8379 & n42431 ;
  assign n42433 = n42432 ^ n10543 ^ 1'b0 ;
  assign n42434 = n42430 & ~n42433 ;
  assign n42435 = ( n1021 & n18270 ) | ( n1021 & ~n42434 ) | ( n18270 & ~n42434 ) ;
  assign n42440 = n9848 ^ n5996 ^ 1'b0 ;
  assign n42441 = n16 & ~n42440 ;
  assign n42442 = ~n27700 & n42441 ;
  assign n42436 = ~n4110 & n12578 ;
  assign n42437 = n42436 ^ n2254 ^ 1'b0 ;
  assign n42438 = n9520 & n42437 ;
  assign n42439 = n42438 ^ n14831 ^ 1'b0 ;
  assign n42443 = n42442 ^ n42439 ^ 1'b0 ;
  assign n42446 = n469 ^ n134 ^ n26 ;
  assign n42444 = n2510 & n18910 ;
  assign n42445 = ~n37542 & n42444 ;
  assign n42447 = n42446 ^ n42445 ^ 1'b0 ;
  assign n42448 = n7914 ^ n3131 ^ 1'b0 ;
  assign n42449 = ( n530 & n15962 ) | ( n530 & ~n42448 ) | ( n15962 & ~n42448 ) ;
  assign n42450 = ~n20623 & n21873 ;
  assign n42451 = ~n42449 & n42450 ;
  assign n42452 = n30602 ^ n1893 ^ 1'b0 ;
  assign n42453 = n10432 & ~n27608 ;
  assign n42454 = ~n12053 & n42453 ;
  assign n42455 = n9360 & ~n15401 ;
  assign n42456 = n28688 ^ n20226 ^ 1'b0 ;
  assign n42457 = ~n22503 & n42456 ;
  assign n42459 = n10200 ^ n8398 ^ n3365 ;
  assign n42460 = n21654 ^ n819 ^ 1'b0 ;
  assign n42461 = n42459 & ~n42460 ;
  assign n42462 = ( n14807 & ~n17304 ) | ( n14807 & n42461 ) | ( ~n17304 & n42461 ) ;
  assign n42458 = n5517 & ~n15026 ;
  assign n42463 = n42462 ^ n42458 ^ n31953 ;
  assign n42464 = n7225 & ~n11763 ;
  assign n42465 = n20371 & n42464 ;
  assign n42466 = ( ~n8638 & n17499 ) | ( ~n8638 & n42465 ) | ( n17499 & n42465 ) ;
  assign n42467 = n25518 & ~n35777 ;
  assign n42468 = ~n37536 & n42467 ;
  assign n42469 = n2798 ^ n997 ^ 1'b0 ;
  assign n42470 = n11498 & n42469 ;
  assign n42471 = n42470 ^ n6692 ^ 1'b0 ;
  assign n42472 = n39488 ^ n18695 ^ 1'b0 ;
  assign n42473 = n42471 | n42472 ;
  assign n42474 = n15919 & ~n27863 ;
  assign n42475 = n10670 & n20515 ;
  assign n42476 = n42474 & n42475 ;
  assign n42477 = n914 & n4717 ;
  assign n42478 = n42477 ^ n7477 ^ 1'b0 ;
  assign n42479 = n17094 & n42478 ;
  assign n42480 = n811 | n14452 ;
  assign n42481 = n42480 ^ n3105 ^ 1'b0 ;
  assign n42482 = n9663 & n19940 ;
  assign n42483 = ( ~n10330 & n15066 ) | ( ~n10330 & n42482 ) | ( n15066 & n42482 ) ;
  assign n42484 = ~n17185 & n27808 ;
  assign n42485 = ~n10676 & n42484 ;
  assign n42486 = x11 | n42485 ;
  assign n42487 = n15708 ^ n455 ^ 1'b0 ;
  assign n42488 = n29512 | n42487 ;
  assign n42489 = n12391 & n42488 ;
  assign n42490 = n19482 ^ n16737 ^ 1'b0 ;
  assign n42491 = n17727 & ~n38309 ;
  assign n42492 = n42491 ^ n10670 ^ 1'b0 ;
  assign n42493 = n3824 & n7289 ;
  assign n42494 = n42492 & ~n42493 ;
  assign n42495 = n17781 ^ n16228 ^ 1'b0 ;
  assign n42496 = n16556 & n19653 ;
  assign n42497 = n37187 ^ n5535 ^ 1'b0 ;
  assign n42498 = ~n42496 & n42497 ;
  assign n42499 = n17037 & n26540 ;
  assign n42500 = n15189 & n17452 ;
  assign n42501 = n42500 ^ n19269 ^ 1'b0 ;
  assign n42502 = n40162 ^ n32073 ^ 1'b0 ;
  assign n42503 = n16735 ^ n14593 ^ 1'b0 ;
  assign n42504 = ( n3949 & n4275 ) | ( n3949 & ~n4673 ) | ( n4275 & ~n4673 ) ;
  assign n42505 = n23268 | n35571 ;
  assign n42506 = n42504 & ~n42505 ;
  assign n42507 = n42506 ^ n32821 ^ 1'b0 ;
  assign n42508 = ( ~n15638 & n42503 ) | ( ~n15638 & n42507 ) | ( n42503 & n42507 ) ;
  assign n42509 = n1661 | n25741 ;
  assign n42510 = n3786 & ~n9669 ;
  assign n42511 = ~n8076 & n42510 ;
  assign n42512 = n600 & n42511 ;
  assign n42513 = n1625 & n42512 ;
  assign n42514 = n42513 ^ n18522 ^ 1'b0 ;
  assign n42515 = n14460 | n42514 ;
  assign n42516 = n42515 ^ n8356 ^ 1'b0 ;
  assign n42517 = n7661 & n23492 ;
  assign n42518 = n23723 & ~n39996 ;
  assign n42519 = ~n26573 & n42518 ;
  assign n42521 = n12725 & n13019 ;
  assign n42522 = n42521 ^ n5333 ^ 1'b0 ;
  assign n42520 = n3821 & ~n10723 ;
  assign n42523 = n42522 ^ n42520 ^ 1'b0 ;
  assign n42524 = ~n36625 & n42523 ;
  assign n42525 = n15737 | n23035 ;
  assign n42526 = n21657 & ~n42525 ;
  assign n42527 = n20264 & n23479 ;
  assign n42528 = n6037 & n23982 ;
  assign n42529 = n10598 & n42528 ;
  assign n42530 = n42529 ^ n4427 ^ 1'b0 ;
  assign n42531 = ( n18920 & n42527 ) | ( n18920 & ~n42530 ) | ( n42527 & ~n42530 ) ;
  assign n42532 = n40327 ^ n12952 ^ 1'b0 ;
  assign n42536 = n17869 ^ n13028 ^ 1'b0 ;
  assign n42537 = n13327 | n42536 ;
  assign n42533 = n12533 ^ n11591 ^ 1'b0 ;
  assign n42534 = n39417 & n42533 ;
  assign n42535 = ~n7938 & n42534 ;
  assign n42538 = n42537 ^ n42535 ^ 1'b0 ;
  assign n42539 = ~n31286 & n32621 ;
  assign n42540 = n7659 & ~n34612 ;
  assign n42541 = ~n10007 & n27875 ;
  assign n42542 = n4180 & n42541 ;
  assign n42543 = n42540 | n42542 ;
  assign n42544 = n7099 & ~n11824 ;
  assign n42545 = n42544 ^ n2843 ^ 1'b0 ;
  assign n42546 = ( ~n6109 & n12337 ) | ( ~n6109 & n42545 ) | ( n12337 & n42545 ) ;
  assign n42547 = n42546 ^ n37180 ^ n28538 ;
  assign n42548 = ~n8234 & n10849 ;
  assign n42549 = ~n27978 & n38142 ;
  assign n42550 = n42548 & n42549 ;
  assign n42551 = n5421 | n27272 ;
  assign n42552 = n42551 ^ n481 ^ 1'b0 ;
  assign n42553 = n16081 | n41043 ;
  assign n42554 = n42552 & ~n42553 ;
  assign n42555 = n38827 ^ n20091 ^ n17406 ;
  assign n42558 = ( n12989 & n17513 ) | ( n12989 & n21064 ) | ( n17513 & n21064 ) ;
  assign n42556 = ~n4447 & n12965 ;
  assign n42557 = ~n22985 & n42556 ;
  assign n42559 = n42558 ^ n42557 ^ n4345 ;
  assign n42560 = ~n9033 & n17443 ;
  assign n42561 = n39432 ^ n8298 ^ 1'b0 ;
  assign n42562 = n13218 ^ n3510 ^ 1'b0 ;
  assign n42563 = n22871 & ~n29426 ;
  assign n42564 = n316 | n22312 ;
  assign n42565 = n42564 ^ n24028 ^ 1'b0 ;
  assign n42566 = n42565 ^ n16781 ^ 1'b0 ;
  assign n42567 = n14365 & ~n18723 ;
  assign n42568 = n15405 ^ n1746 ^ 1'b0 ;
  assign n42569 = n2114 & ~n34915 ;
  assign n42570 = n3299 | n40161 ;
  assign n42571 = ~n4134 & n22862 ;
  assign n42572 = ( n6754 & n9378 ) | ( n6754 & n42571 ) | ( n9378 & n42571 ) ;
  assign n42573 = ~n2784 & n42572 ;
  assign n42574 = n17576 ^ n14244 ^ 1'b0 ;
  assign n42575 = ~n11202 & n42574 ;
  assign n42579 = n14509 ^ n3135 ^ n130 ;
  assign n42576 = n5051 ^ n3071 ^ 1'b0 ;
  assign n42577 = n5333 & n9253 ;
  assign n42578 = n42576 & n42577 ;
  assign n42580 = n42579 ^ n42578 ^ n3698 ;
  assign n42581 = n42580 ^ n12002 ^ 1'b0 ;
  assign n42582 = ( n9730 & n11059 ) | ( n9730 & n20494 ) | ( n11059 & n20494 ) ;
  assign n42583 = n9388 & n16061 ;
  assign n42584 = n23171 ^ n18270 ^ 1'b0 ;
  assign n42585 = n2419 & ~n12791 ;
  assign n42586 = ~n15285 & n42585 ;
  assign n42587 = n14228 ^ n10147 ^ 1'b0 ;
  assign n42588 = n17079 & n42587 ;
  assign n42589 = n40022 ^ n21167 ^ 1'b0 ;
  assign n42590 = n42588 & ~n42589 ;
  assign n42591 = n10344 ^ n10052 ^ 1'b0 ;
  assign n42592 = ~n10001 & n42591 ;
  assign n42593 = n11688 & ~n23900 ;
  assign n42594 = ( ~n18753 & n20349 ) | ( ~n18753 & n37783 ) | ( n20349 & n37783 ) ;
  assign n42595 = n9811 ^ n9644 ^ 1'b0 ;
  assign n42596 = ~n4851 & n29705 ;
  assign n42597 = n42596 ^ n3022 ^ 1'b0 ;
  assign n42598 = n8950 & ~n11079 ;
  assign n42599 = n42597 | n42598 ;
  assign n42600 = n42599 ^ n23455 ^ 1'b0 ;
  assign n42601 = n3489 ^ n968 ^ 1'b0 ;
  assign n42602 = ~n20382 & n42601 ;
  assign n42603 = n4104 & n42602 ;
  assign n42604 = n42603 ^ n30944 ^ n26567 ;
  assign n42605 = n31712 ^ n22457 ^ 1'b0 ;
  assign n42606 = n17357 ^ n648 ^ 1'b0 ;
  assign n42607 = n11111 | n42606 ;
  assign n42608 = n29054 | n41931 ;
  assign n42609 = n5052 & ~n42608 ;
  assign n42610 = n6353 & n38445 ;
  assign n42611 = ( n35794 & n42609 ) | ( n35794 & ~n42610 ) | ( n42609 & ~n42610 ) ;
  assign n42612 = n21408 ^ n10054 ^ 1'b0 ;
  assign n42613 = ~n30800 & n36567 ;
  assign n42614 = ~n40654 & n42613 ;
  assign n42615 = n428 & ~n26151 ;
  assign n42616 = n3588 & n42615 ;
  assign n42617 = n614 & ~n17243 ;
  assign n42618 = n42617 ^ n34933 ^ 1'b0 ;
  assign n42619 = ~n3768 & n10827 ;
  assign n42620 = n35808 ^ n7144 ^ 1'b0 ;
  assign n42621 = n35761 | n42620 ;
  assign n42622 = n42619 & ~n42621 ;
  assign n42623 = n17804 ^ n10973 ^ 1'b0 ;
  assign n42624 = ~n10331 & n42623 ;
  assign n42625 = n3358 & ~n42624 ;
  assign n42626 = n42625 ^ n3817 ^ 1'b0 ;
  assign n42627 = n41793 ^ n9086 ^ 1'b0 ;
  assign n42628 = n22263 ^ n20771 ^ 1'b0 ;
  assign n42629 = ~n596 & n42628 ;
  assign n42630 = ( n7462 & ~n33367 ) | ( n7462 & n42629 ) | ( ~n33367 & n42629 ) ;
  assign n42631 = n15013 | n37877 ;
  assign n42632 = n16534 | n23573 ;
  assign n42633 = n6745 & n42632 ;
  assign n42634 = n7337 | n28551 ;
  assign n42635 = n42634 ^ n9935 ^ 1'b0 ;
  assign n42636 = n1932 | n7895 ;
  assign n42637 = n8582 & ~n22119 ;
  assign n42638 = ( n32717 & n34266 ) | ( n32717 & n42291 ) | ( n34266 & n42291 ) ;
  assign n42639 = n20965 | n35679 ;
  assign n42640 = n35521 | n42639 ;
  assign n42641 = ~n809 & n30445 ;
  assign n42642 = n13813 ^ n6022 ^ 1'b0 ;
  assign n42643 = n12303 & n42642 ;
  assign n42644 = n16650 & n42643 ;
  assign n42645 = n19996 & ~n35364 ;
  assign n42646 = n40108 ^ n25042 ^ n19793 ;
  assign n42647 = n32163 ^ n7307 ^ 1'b0 ;
  assign n42648 = ~n21913 & n42647 ;
  assign n42649 = n3918 & n10297 ;
  assign n42650 = n33803 ^ n32716 ^ n14207 ;
  assign n42651 = ~n102 & n1701 ;
  assign n42652 = n102 & n42651 ;
  assign n42653 = n115 & n42652 ;
  assign n42654 = ~n3658 & n23864 ;
  assign n42655 = n42653 & n42654 ;
  assign n42656 = n42655 ^ n8125 ^ n4041 ;
  assign n42657 = n19693 & n42656 ;
  assign n42658 = n42650 & ~n42657 ;
  assign n42659 = n42658 ^ n13307 ^ 1'b0 ;
  assign n42660 = n18625 | n42659 ;
  assign n42661 = n8334 | n42660 ;
  assign n42662 = n15394 & ~n42661 ;
  assign n42663 = n11273 & ~n26319 ;
  assign n42664 = ~n23055 & n42663 ;
  assign n42665 = n15436 ^ n14721 ^ 1'b0 ;
  assign n42666 = n42664 & n42665 ;
  assign n42667 = n24130 ^ n14880 ^ n12486 ;
  assign n42668 = n42667 ^ n37995 ^ n31727 ;
  assign n42669 = n15774 ^ n13671 ^ 1'b0 ;
  assign n42670 = ( n3600 & n7968 ) | ( n3600 & ~n42669 ) | ( n7968 & ~n42669 ) ;
  assign n42671 = n7807 | n31515 ;
  assign n42672 = n2954 ^ n1283 ^ 1'b0 ;
  assign n42673 = n24493 & ~n42672 ;
  assign n42674 = n21813 ^ n14071 ^ 1'b0 ;
  assign n42675 = n8950 & n12010 ;
  assign n42676 = n15700 ^ n14993 ^ 1'b0 ;
  assign n42677 = n1138 | n23118 ;
  assign n42678 = n42677 ^ n25766 ^ 1'b0 ;
  assign n42679 = n13205 | n42678 ;
  assign n42680 = n7976 ^ n3094 ^ 1'b0 ;
  assign n42681 = n30851 & ~n41959 ;
  assign n42682 = n9363 ^ n127 ^ 1'b0 ;
  assign n42683 = n31858 & n42682 ;
  assign n42684 = n4961 ^ n2317 ^ 1'b0 ;
  assign n42685 = ~n32928 & n42684 ;
  assign n42686 = n30798 ^ n6045 ^ 1'b0 ;
  assign n42687 = n25741 & n42686 ;
  assign n42688 = n17389 | n36742 ;
  assign n42689 = n42688 ^ n15777 ^ 1'b0 ;
  assign n42690 = n42689 ^ n10145 ^ 1'b0 ;
  assign n42691 = n42690 ^ n41653 ^ n39077 ;
  assign n42692 = ~n11628 & n35445 ;
  assign n42693 = n42692 ^ n31837 ^ 1'b0 ;
  assign n42694 = n18542 | n31682 ;
  assign n42695 = n24290 & ~n42694 ;
  assign n42696 = n15101 & ~n21174 ;
  assign n42697 = n39843 ^ n28185 ^ 1'b0 ;
  assign n42698 = n34377 ^ n11911 ^ 1'b0 ;
  assign n42699 = n25347 & n42698 ;
  assign n42701 = n12751 ^ n2104 ^ n740 ;
  assign n42702 = n11503 | n42701 ;
  assign n42703 = n42702 ^ n12449 ^ 1'b0 ;
  assign n42700 = n4829 & n5961 ;
  assign n42704 = n42703 ^ n42700 ^ 1'b0 ;
  assign n42705 = n17121 | n42704 ;
  assign n42706 = n6406 & ~n12955 ;
  assign n42707 = n42706 ^ n23491 ^ 1'b0 ;
  assign n42708 = ( n1526 & n15871 ) | ( n1526 & n42707 ) | ( n15871 & n42707 ) ;
  assign n42711 = n21868 ^ n345 ^ 1'b0 ;
  assign n42710 = ~n4231 & n32198 ;
  assign n42709 = ~n34051 & n34251 ;
  assign n42712 = n42711 ^ n42710 ^ n42709 ;
  assign n42713 = n19148 & ~n25900 ;
  assign n42714 = n30113 & n42713 ;
  assign n42715 = ~n25184 & n27247 ;
  assign n42716 = n8243 ^ n6659 ^ 1'b0 ;
  assign n42717 = n8039 | n42716 ;
  assign n42718 = n16488 ^ n9218 ^ 1'b0 ;
  assign n42719 = ~n42717 & n42718 ;
  assign n42720 = n42715 & n42719 ;
  assign n42721 = n18243 | n27806 ;
  assign n42722 = n17162 ^ n16332 ^ 1'b0 ;
  assign n42723 = n26505 | n42722 ;
  assign n42724 = n445 & n1167 ;
  assign n42725 = n5550 & n42724 ;
  assign n42726 = n2946 & n4195 ;
  assign n42727 = ~n14847 & n42726 ;
  assign n42728 = n7773 & n37528 ;
  assign n42729 = n42728 ^ n26618 ^ 1'b0 ;
  assign n42730 = n34021 & ~n42729 ;
  assign n42731 = n42730 ^ n2262 ^ 1'b0 ;
  assign n42732 = n37111 ^ n1481 ^ 1'b0 ;
  assign n42733 = n42731 & ~n42732 ;
  assign n42734 = n42099 ^ n26450 ^ n10206 ;
  assign n42735 = n24502 | n28543 ;
  assign n42736 = n6639 & n21742 ;
  assign n42737 = ~n14375 & n42736 ;
  assign n42738 = ( n12106 & n42735 ) | ( n12106 & ~n42737 ) | ( n42735 & ~n42737 ) ;
  assign n42739 = ~n12923 & n19097 ;
  assign n42740 = n42739 ^ n2945 ^ 1'b0 ;
  assign n42741 = n9768 & n38960 ;
  assign n42742 = ~n42740 & n42741 ;
  assign n42743 = n42742 ^ n15590 ^ n6544 ;
  assign n42744 = n38581 ^ n24053 ^ 1'b0 ;
  assign n42745 = n6983 & ~n42744 ;
  assign n42746 = n9750 & n22539 ;
  assign n42747 = n42746 ^ n18587 ^ 1'b0 ;
  assign n42748 = n31139 ^ n18715 ^ 1'b0 ;
  assign n42749 = n42747 | n42748 ;
  assign n42750 = n42749 ^ n1848 ^ 1'b0 ;
  assign n42751 = ~n1481 & n42750 ;
  assign n42752 = n5879 | n10020 ;
  assign n42753 = n42752 ^ n23158 ^ 1'b0 ;
  assign n42754 = ~n4427 & n42753 ;
  assign n42755 = n1531 & ~n26400 ;
  assign n42756 = ~n5824 & n17771 ;
  assign n42757 = n42756 ^ n432 ^ 1'b0 ;
  assign n42758 = n42755 & n42757 ;
  assign n42759 = n6595 | n36899 ;
  assign n42760 = n25187 ^ n6787 ^ 1'b0 ;
  assign n42761 = n42760 ^ n9149 ^ n2397 ;
  assign n42762 = n2594 & ~n9911 ;
  assign n42763 = n42762 ^ n17897 ^ 1'b0 ;
  assign n42764 = n4765 | n9571 ;
  assign n42765 = n25728 & n42764 ;
  assign n42766 = n27474 | n30944 ;
  assign n42767 = n42766 ^ n220 ^ 1'b0 ;
  assign n42768 = n17652 & ~n42767 ;
  assign n42769 = ~n42765 & n42768 ;
  assign n42770 = n3389 | n20371 ;
  assign n42771 = n9246 | n42770 ;
  assign n42772 = n25621 ^ n13745 ^ n7181 ;
  assign n42773 = n7130 & ~n12840 ;
  assign n42774 = n42773 ^ n4055 ^ n2434 ;
  assign n42775 = n22465 ^ n12049 ^ 1'b0 ;
  assign n42776 = n3564 & n31615 ;
  assign n42777 = n11285 & ~n42776 ;
  assign n42778 = ~n42701 & n42777 ;
  assign n42779 = n42778 ^ n25400 ^ 1'b0 ;
  assign n42780 = n22147 & n42779 ;
  assign n42781 = n40799 ^ n23406 ^ 1'b0 ;
  assign n42782 = n33571 ^ n22 ^ 1'b0 ;
  assign n42783 = n42781 | n42782 ;
  assign n42787 = n11344 | n14516 ;
  assign n42788 = n16129 | n42787 ;
  assign n42784 = n15914 ^ n890 ^ 1'b0 ;
  assign n42785 = n9032 & n42784 ;
  assign n42786 = n1277 & n42785 ;
  assign n42789 = n42788 ^ n42786 ^ 1'b0 ;
  assign n42790 = ( n11037 & n23464 ) | ( n11037 & ~n42789 ) | ( n23464 & ~n42789 ) ;
  assign n42791 = n42790 ^ n3898 ^ 1'b0 ;
  assign n42792 = ~n24779 & n42791 ;
  assign n42793 = n4436 | n12583 ;
  assign n42798 = n6201 | n16591 ;
  assign n42799 = n2764 | n42798 ;
  assign n42795 = n6042 & n23025 ;
  assign n42796 = ( n17913 & n37510 ) | ( n17913 & ~n42795 ) | ( n37510 & ~n42795 ) ;
  assign n42794 = n17771 & ~n26523 ;
  assign n42797 = n42796 ^ n42794 ^ 1'b0 ;
  assign n42800 = n42799 ^ n42797 ^ 1'b0 ;
  assign n42801 = n42793 & ~n42800 ;
  assign n42802 = n31854 ^ n27899 ^ 1'b0 ;
  assign n42803 = n11451 | n22867 ;
  assign n42804 = n5377 | n6915 ;
  assign n42805 = n2670 | n42804 ;
  assign n42806 = n42805 ^ n9217 ^ 1'b0 ;
  assign n42807 = ( n3700 & ~n7943 ) | ( n3700 & n42806 ) | ( ~n7943 & n42806 ) ;
  assign n42810 = n7838 | n9392 ;
  assign n42808 = n19436 ^ n6417 ^ 1'b0 ;
  assign n42809 = n42808 ^ n17830 ^ n12929 ;
  assign n42811 = n42810 ^ n42809 ^ 1'b0 ;
  assign n42812 = n25508 ^ n1909 ^ 1'b0 ;
  assign n42813 = ~n1918 & n4215 ;
  assign n42814 = n42813 ^ n3163 ^ 1'b0 ;
  assign n42815 = ~n44 & n34673 ;
  assign n42816 = n42815 ^ n5720 ^ 1'b0 ;
  assign n42817 = ~n5305 & n12730 ;
  assign n42818 = n28182 & ~n42817 ;
  assign n42819 = ~n42816 & n42818 ;
  assign n42820 = n6095 ^ n2515 ^ 1'b0 ;
  assign n42821 = n42820 ^ n9964 ^ 1'b0 ;
  assign n42822 = n21475 | n42821 ;
  assign n42823 = n42822 ^ n21326 ^ 1'b0 ;
  assign n42824 = n4551 | n26985 ;
  assign n42825 = n22540 & ~n42824 ;
  assign n42826 = ( n11243 & ~n37128 ) | ( n11243 & n42825 ) | ( ~n37128 & n42825 ) ;
  assign n42827 = n14439 ^ n11540 ^ n11366 ;
  assign n42828 = ( n18229 & n41428 ) | ( n18229 & n42827 ) | ( n41428 & n42827 ) ;
  assign n42829 = ~n1195 & n12662 ;
  assign n42830 = n12851 | n42829 ;
  assign n42831 = n41190 & ~n42830 ;
  assign n42832 = n20896 ^ n1511 ^ 1'b0 ;
  assign n42833 = n18448 & n42832 ;
  assign n42834 = n9308 ^ n7823 ^ 1'b0 ;
  assign n42835 = ~n7900 & n42834 ;
  assign n42836 = ( n33756 & n37918 ) | ( n33756 & ~n42835 ) | ( n37918 & ~n42835 ) ;
  assign n42837 = ~n1868 & n5691 ;
  assign n42838 = n5656 | n11870 ;
  assign n42839 = n42838 ^ n9072 ^ 1'b0 ;
  assign n42840 = ( n13605 & n42837 ) | ( n13605 & ~n42839 ) | ( n42837 & ~n42839 ) ;
  assign n42841 = ~n4867 & n23368 ;
  assign n42842 = n42841 ^ n9292 ^ 1'b0 ;
  assign n42843 = ~n30993 & n42842 ;
  assign n42844 = ~n10711 & n42843 ;
  assign n42845 = n601 & ~n6710 ;
  assign n42846 = n4723 | n18777 ;
  assign n42847 = n42846 ^ n36296 ^ 1'b0 ;
  assign n42848 = n1099 & n18210 ;
  assign n42849 = ~n42847 & n42848 ;
  assign n42852 = n37273 ^ n15864 ^ n172 ;
  assign n42850 = n29516 ^ n1031 ^ 1'b0 ;
  assign n42851 = n19321 & n42850 ;
  assign n42853 = n42852 ^ n42851 ^ 1'b0 ;
  assign n42854 = n8204 ^ n7915 ^ 1'b0 ;
  assign n42855 = n7342 | n12885 ;
  assign n42856 = n11666 & ~n42855 ;
  assign n42857 = n42856 ^ n14416 ^ 1'b0 ;
  assign n42858 = n11964 & ~n42857 ;
  assign n42859 = n42858 ^ n21198 ^ n9409 ;
  assign n42860 = ( n24395 & n32054 ) | ( n24395 & n34037 ) | ( n32054 & n34037 ) ;
  assign n42861 = n27168 ^ n23095 ^ 1'b0 ;
  assign n42862 = ~n3949 & n5354 ;
  assign n42863 = ~n6614 & n42862 ;
  assign n42864 = n517 & n794 ;
  assign n42865 = n42864 ^ n42850 ^ 1'b0 ;
  assign n42866 = ~n5008 & n42865 ;
  assign n42867 = n18069 & n42866 ;
  assign n42868 = n42867 ^ n20989 ^ 1'b0 ;
  assign n42869 = n13795 | n42868 ;
  assign n42870 = n2471 & n9872 ;
  assign n42871 = n24885 ^ n14697 ^ 1'b0 ;
  assign n42872 = n25900 ^ n20475 ^ n20394 ;
  assign n42873 = n42872 ^ n10502 ^ 1'b0 ;
  assign n42874 = n9339 ^ n8520 ^ n3745 ;
  assign n42875 = n5533 & n26929 ;
  assign n42876 = n7941 & n42875 ;
  assign n42877 = n6128 & n25633 ;
  assign n42878 = ~n1083 & n42877 ;
  assign n42879 = n6535 & ~n42878 ;
  assign n42880 = n42879 ^ n23571 ^ 1'b0 ;
  assign n42881 = n42880 ^ n37839 ^ 1'b0 ;
  assign n42882 = n36459 & n42881 ;
  assign n42883 = n4272 & ~n39719 ;
  assign n42884 = n23821 ^ n18432 ^ 1'b0 ;
  assign n42885 = ~n5583 & n22094 ;
  assign n42886 = n15770 | n21054 ;
  assign n42887 = n2944 & ~n42886 ;
  assign n42888 = n12330 | n42887 ;
  assign n42889 = n16721 | n42888 ;
  assign n42890 = n42889 ^ n20885 ^ 1'b0 ;
  assign n42892 = n7185 | n15564 ;
  assign n42893 = n42892 ^ n3350 ^ 1'b0 ;
  assign n42891 = ( n2206 & n7084 ) | ( n2206 & n10601 ) | ( n7084 & n10601 ) ;
  assign n42894 = n42893 ^ n42891 ^ n30483 ;
  assign n42895 = n34690 ^ n22391 ^ n7110 ;
  assign n42896 = n21269 ^ n2186 ^ 1'b0 ;
  assign n42897 = n8509 | n34046 ;
  assign n42898 = n8927 & n18448 ;
  assign n42899 = ~n42897 & n42898 ;
  assign n42900 = n35276 ^ n617 ^ 1'b0 ;
  assign n42901 = ~n3578 & n16525 ;
  assign n42902 = n42901 ^ n9643 ^ 1'b0 ;
  assign n42903 = n21410 ^ n7808 ^ 1'b0 ;
  assign n42904 = ( ~n2882 & n39841 ) | ( ~n2882 & n42485 ) | ( n39841 & n42485 ) ;
  assign n42905 = n16021 & n41169 ;
  assign n42906 = ~n5924 & n42905 ;
  assign n42907 = n42906 ^ n395 ^ 1'b0 ;
  assign n42908 = n13574 & ~n42907 ;
  assign n42909 = n8619 & n20460 ;
  assign n42910 = n42909 ^ n11744 ^ 1'b0 ;
  assign n42911 = n42908 & ~n42910 ;
  assign n42912 = n10424 & ~n42911 ;
  assign n42913 = n1364 & n16271 ;
  assign n42914 = n42913 ^ n5363 ^ 1'b0 ;
  assign n42915 = n7842 & ~n13282 ;
  assign n42916 = ( n6094 & n16204 ) | ( n6094 & n19409 ) | ( n16204 & n19409 ) ;
  assign n42917 = n12875 ^ n1000 ^ 1'b0 ;
  assign n42918 = ( n17772 & n39292 ) | ( n17772 & ~n42917 ) | ( n39292 & ~n42917 ) ;
  assign n42919 = n4010 & ~n12428 ;
  assign n42920 = n42919 ^ n12877 ^ 1'b0 ;
  assign n42921 = n14666 & n42920 ;
  assign n42922 = ~n5284 & n42449 ;
  assign n42923 = n11040 & ~n42401 ;
  assign n42924 = n16484 | n42923 ;
  assign n42925 = n1456 | n42924 ;
  assign n42926 = ~n4786 & n16422 ;
  assign n42927 = n42926 ^ n2846 ^ 1'b0 ;
  assign n42928 = ~n13379 & n42927 ;
  assign n42929 = n42928 ^ n3439 ^ 1'b0 ;
  assign n42930 = n39405 ^ n11841 ^ 1'b0 ;
  assign n42931 = n42929 & ~n42930 ;
  assign n42932 = ~n10548 & n13307 ;
  assign n42933 = n42932 ^ n8801 ^ 1'b0 ;
  assign n42934 = n25549 & n28020 ;
  assign n42935 = n21165 ^ n8164 ^ 1'b0 ;
  assign n42936 = n28229 | n35429 ;
  assign n42937 = n17844 | n38023 ;
  assign n42938 = n10578 & n15716 ;
  assign n42939 = n28983 | n31418 ;
  assign n42940 = n788 | n42939 ;
  assign n42941 = ( n1393 & ~n23630 ) | ( n1393 & n42940 ) | ( ~n23630 & n42940 ) ;
  assign n42946 = n1225 | n5704 ;
  assign n42947 = n398 & ~n42946 ;
  assign n42944 = n14710 & n40748 ;
  assign n42945 = n42944 ^ n29713 ^ 1'b0 ;
  assign n42942 = n9171 & n29543 ;
  assign n42943 = ~n6589 & n42942 ;
  assign n42948 = n42947 ^ n42945 ^ n42943 ;
  assign n42949 = n4270 ^ n1200 ^ 1'b0 ;
  assign n42950 = n8041 | n42949 ;
  assign n42951 = ~n9826 & n23257 ;
  assign n42952 = n24108 & n42951 ;
  assign n42953 = ~n529 & n15654 ;
  assign n42954 = n42953 ^ n14319 ^ 1'b0 ;
  assign n42955 = n7141 & ~n40242 ;
  assign n42956 = n42955 ^ n17498 ^ 1'b0 ;
  assign n42957 = n5672 | n36606 ;
  assign n42958 = n42957 ^ n15448 ^ 1'b0 ;
  assign n42959 = n36775 ^ n1182 ^ 1'b0 ;
  assign n42960 = n3995 ^ n704 ^ 1'b0 ;
  assign n42961 = ( ~n21837 & n24900 ) | ( ~n21837 & n34700 ) | ( n24900 & n34700 ) ;
  assign n42962 = n4863 | n42961 ;
  assign n42963 = n42960 & ~n42962 ;
  assign n42964 = n15189 | n42963 ;
  assign n42965 = n17556 & n42964 ;
  assign n42966 = n30685 & ~n34956 ;
  assign n42967 = n6456 & n42966 ;
  assign n42968 = n42967 ^ n24164 ^ n12449 ;
  assign n42969 = n3858 & ~n42968 ;
  assign n42971 = n2114 & ~n7479 ;
  assign n42972 = n126 & n42971 ;
  assign n42973 = n42972 ^ n18119 ^ 1'b0 ;
  assign n42974 = n10786 & ~n42973 ;
  assign n42975 = n1088 & n42974 ;
  assign n42976 = n2111 & n42975 ;
  assign n42970 = n8866 & n18530 ;
  assign n42977 = n42976 ^ n42970 ^ 1'b0 ;
  assign n42978 = n6511 & n42977 ;
  assign n42979 = n42978 ^ n36592 ^ 1'b0 ;
  assign n42980 = n42979 ^ n2517 ^ 1'b0 ;
  assign n42984 = n2157 | n19028 ;
  assign n42985 = n42984 ^ n257 ^ 1'b0 ;
  assign n42981 = n9833 & n38621 ;
  assign n42982 = n30260 & n42981 ;
  assign n42983 = n32637 & ~n42982 ;
  assign n42986 = n42985 ^ n42983 ^ 1'b0 ;
  assign n42987 = n16605 ^ n3626 ^ 1'b0 ;
  assign n42988 = ~n27885 & n42987 ;
  assign n42989 = n42988 ^ n18044 ^ 1'b0 ;
  assign n42990 = ( n15276 & n27159 ) | ( n15276 & n42989 ) | ( n27159 & n42989 ) ;
  assign n42991 = n21555 & n41169 ;
  assign n42992 = n42991 ^ n41444 ^ 1'b0 ;
  assign n42994 = n25171 & n26820 ;
  assign n42995 = n42994 ^ n24622 ^ 1'b0 ;
  assign n42993 = n3332 & ~n32905 ;
  assign n42996 = n42995 ^ n42993 ^ 1'b0 ;
  assign n42997 = n42996 ^ n11813 ^ 1'b0 ;
  assign n42998 = ~n13825 & n19782 ;
  assign n42999 = n10134 & n42998 ;
  assign n43000 = n15384 ^ n3312 ^ 1'b0 ;
  assign n43001 = n39621 ^ n32180 ^ n3043 ;
  assign n43002 = ( n2592 & n5236 ) | ( n2592 & n14174 ) | ( n5236 & n14174 ) ;
  assign n43003 = n22923 & ~n23091 ;
  assign n43004 = n10313 & n43003 ;
  assign n43005 = n18866 & ~n43004 ;
  assign n43006 = ( n15353 & ~n43002 ) | ( n15353 & n43005 ) | ( ~n43002 & n43005 ) ;
  assign n43007 = n33312 ^ n2322 ^ 1'b0 ;
  assign n43008 = ~n10305 & n43007 ;
  assign n43009 = ~n1505 & n43008 ;
  assign n43010 = n43009 ^ n37951 ^ 1'b0 ;
  assign n43011 = n18242 & n42595 ;
  assign n43012 = n19658 | n23036 ;
  assign n43013 = n43012 ^ n33776 ^ 1'b0 ;
  assign n43014 = n30521 & ~n38206 ;
  assign n43015 = n18211 ^ n8681 ^ 1'b0 ;
  assign n43016 = n43015 ^ n40674 ^ 1'b0 ;
  assign n43017 = ( n11709 & n15511 ) | ( n11709 & n21935 ) | ( n15511 & n21935 ) ;
  assign n43018 = n773 | n5963 ;
  assign n43019 = n43018 ^ n38976 ^ 1'b0 ;
  assign n43020 = n22886 ^ n6010 ^ 1'b0 ;
  assign n43021 = n43020 ^ n23970 ^ 1'b0 ;
  assign n43022 = n23963 & ~n43021 ;
  assign n43023 = n6985 | n13215 ;
  assign n43024 = n43023 ^ n14152 ^ 1'b0 ;
  assign n43025 = ~n6493 & n43024 ;
  assign n43026 = n11563 & ~n24996 ;
  assign n43027 = n43026 ^ n24699 ^ 1'b0 ;
  assign n43028 = n30712 & n43027 ;
  assign n43029 = n43028 ^ n42186 ^ n10861 ;
  assign n43030 = n15193 & ~n25164 ;
  assign n43031 = n43030 ^ n7944 ^ n1636 ;
  assign n43033 = n7678 | n10111 ;
  assign n43034 = n10211 | n43033 ;
  assign n43032 = n3061 & n31757 ;
  assign n43035 = n43034 ^ n43032 ^ n35186 ;
  assign n43036 = n13449 ^ n7847 ^ 1'b0 ;
  assign n43037 = n42237 ^ n2502 ^ 1'b0 ;
  assign n43038 = ~n41775 & n43037 ;
  assign n43039 = n8347 & n15424 ;
  assign n43040 = n14735 & ~n18277 ;
  assign n43041 = n6360 & ~n13850 ;
  assign n43042 = n25341 ^ n10122 ^ 1'b0 ;
  assign n43043 = ~n43041 & n43042 ;
  assign n43044 = ~n4985 & n43043 ;
  assign n43045 = n18806 & n43044 ;
  assign n43046 = ~n2347 & n2596 ;
  assign n43047 = ~n20453 & n29006 ;
  assign n43048 = n37219 & n39168 ;
  assign n43049 = n861 & ~n34624 ;
  assign n43050 = n30583 & n43049 ;
  assign n43051 = n36 & n43050 ;
  assign n43052 = n20272 & ~n43051 ;
  assign n43053 = n6558 ^ n1886 ^ 1'b0 ;
  assign n43054 = ( n22917 & ~n27596 ) | ( n22917 & n43053 ) | ( ~n27596 & n43053 ) ;
  assign n43055 = n43054 ^ n1729 ^ n514 ;
  assign n43056 = ~n2425 & n25600 ;
  assign n43057 = ~n43055 & n43056 ;
  assign n43058 = n5449 ^ n4631 ^ 1'b0 ;
  assign n43059 = ~n2047 & n43058 ;
  assign n43060 = ( n22850 & n26034 ) | ( n22850 & ~n43059 ) | ( n26034 & ~n43059 ) ;
  assign n43061 = n26064 & ~n33042 ;
  assign n43062 = ~n2130 & n43061 ;
  assign n43066 = n17310 ^ n12393 ^ 1'b0 ;
  assign n43067 = n28245 ^ n24220 ^ 1'b0 ;
  assign n43068 = ~n43066 & n43067 ;
  assign n43069 = n43068 ^ n20484 ^ 1'b0 ;
  assign n43063 = n13165 ^ n12237 ^ 1'b0 ;
  assign n43064 = n6452 & ~n43063 ;
  assign n43065 = n10274 & n43064 ;
  assign n43070 = n43069 ^ n43065 ^ 1'b0 ;
  assign n43071 = n34761 ^ n2945 ^ 1'b0 ;
  assign n43072 = n12454 & n43071 ;
  assign n43073 = ~n8891 & n23565 ;
  assign n43074 = n3488 & n43073 ;
  assign n43075 = ~n8807 & n43074 ;
  assign n43076 = n43072 & ~n43075 ;
  assign n43077 = n12954 ^ n2816 ^ 1'b0 ;
  assign n43078 = n11288 | n43077 ;
  assign n43079 = ~n4097 & n6336 ;
  assign n43080 = n23333 & n43079 ;
  assign n43081 = n20015 ^ n580 ^ 1'b0 ;
  assign n43082 = n43081 ^ n42471 ^ 1'b0 ;
  assign n43083 = n22687 ^ n20836 ^ 1'b0 ;
  assign n43084 = n18875 & n43083 ;
  assign n43085 = ( n8721 & n25750 ) | ( n8721 & n43084 ) | ( n25750 & n43084 ) ;
  assign n43086 = n18987 & ~n33144 ;
  assign n43087 = n3519 & ~n20149 ;
  assign n43089 = n11569 & n29105 ;
  assign n43090 = n6784 & ~n43089 ;
  assign n43091 = n43090 ^ n23308 ^ 1'b0 ;
  assign n43092 = n2953 & n43091 ;
  assign n43093 = n2044 & n43092 ;
  assign n43088 = n10442 & n30275 ;
  assign n43094 = n43093 ^ n43088 ^ n1300 ;
  assign n43095 = n21646 & ~n28928 ;
  assign n43096 = n787 | n27156 ;
  assign n43097 = ( n6922 & ~n9487 ) | ( n6922 & n29877 ) | ( ~n9487 & n29877 ) ;
  assign n43098 = ~n42194 & n43097 ;
  assign n43099 = ~n19616 & n38446 ;
  assign n43100 = ~n39029 & n43099 ;
  assign n43101 = n43100 ^ n13388 ^ 1'b0 ;
  assign n43102 = n43101 ^ n28773 ^ 1'b0 ;
  assign n43103 = n4129 ^ n38 ^ 1'b0 ;
  assign n43104 = n26233 ^ n9221 ^ 1'b0 ;
  assign n43105 = n43103 | n43104 ;
  assign n43106 = ( n5069 & n38244 ) | ( n5069 & ~n43105 ) | ( n38244 & ~n43105 ) ;
  assign n43107 = n29660 ^ n29341 ^ n1334 ;
  assign n43108 = n43107 ^ n37616 ^ 1'b0 ;
  assign n43109 = n7154 | n42550 ;
  assign n43110 = n7255 | n43109 ;
  assign n43111 = ( n22876 & ~n35242 ) | ( n22876 & n38631 ) | ( ~n35242 & n38631 ) ;
  assign n43112 = ~n2603 & n10161 ;
  assign n43113 = n43111 & n43112 ;
  assign n43114 = n11854 ^ n1022 ^ 1'b0 ;
  assign n43115 = n27043 & ~n43114 ;
  assign n43116 = n16750 ^ n11383 ^ 1'b0 ;
  assign n43117 = n41849 | n43116 ;
  assign n43118 = ( n20285 & n31688 ) | ( n20285 & ~n43117 ) | ( n31688 & ~n43117 ) ;
  assign n43119 = n34034 ^ n10531 ^ 1'b0 ;
  assign n43120 = n2148 & n21851 ;
  assign n43121 = n43119 & n43120 ;
  assign n43122 = n24619 & ~n43121 ;
  assign n43123 = ~n3867 & n43122 ;
  assign n43124 = ~n80 & n10218 ;
  assign n43125 = n9127 | n20364 ;
  assign n43126 = n4025 & n30398 ;
  assign n43127 = n4751 & n41460 ;
  assign n43128 = n4202 | n11668 ;
  assign n43129 = ~n5312 & n22684 ;
  assign n43130 = n25796 ^ n11042 ^ 1'b0 ;
  assign n43131 = ~n24537 & n43130 ;
  assign n43134 = n18093 ^ n1906 ^ 1'b0 ;
  assign n43135 = n27516 & ~n43134 ;
  assign n43132 = n22421 | n24705 ;
  assign n43133 = n43132 ^ n19372 ^ 1'b0 ;
  assign n43136 = n43135 ^ n43133 ^ 1'b0 ;
  assign n43137 = ~n20476 & n33235 ;
  assign n43138 = n43137 ^ n41848 ^ 1'b0 ;
  assign n43139 = n28295 & ~n29251 ;
  assign n43140 = n43139 ^ n36508 ^ 1'b0 ;
  assign n43141 = ~n5846 & n8476 ;
  assign n43143 = n11690 ^ n5176 ^ 1'b0 ;
  assign n43144 = ~n25738 & n43143 ;
  assign n43145 = n20605 & ~n38170 ;
  assign n43146 = ~n43144 & n43145 ;
  assign n43142 = n17712 | n22079 ;
  assign n43147 = n43146 ^ n43142 ^ n8323 ;
  assign n43148 = n25161 ^ n17199 ^ n16207 ;
  assign n43149 = n1272 & n43148 ;
  assign n43150 = n43149 ^ n28120 ^ 1'b0 ;
  assign n43152 = ~n5203 & n17842 ;
  assign n43153 = n43152 ^ n14135 ^ 1'b0 ;
  assign n43154 = n43153 ^ n29575 ^ n13509 ;
  assign n43151 = n22734 ^ n3691 ^ 1'b0 ;
  assign n43155 = n43154 ^ n43151 ^ 1'b0 ;
  assign n43156 = n9125 & ~n23866 ;
  assign n43157 = n43156 ^ n5024 ^ 1'b0 ;
  assign n43158 = n19352 & n32954 ;
  assign n43159 = n43158 ^ n31607 ^ 1'b0 ;
  assign n43160 = ( n9224 & ~n13772 ) | ( n9224 & n16743 ) | ( ~n13772 & n16743 ) ;
  assign n43161 = ( n2071 & n27295 ) | ( n2071 & n28769 ) | ( n27295 & n28769 ) ;
  assign n43162 = n30679 & ~n43161 ;
  assign n43163 = n3793 & ~n8706 ;
  assign n43164 = n43163 ^ n13252 ^ n10453 ;
  assign n43165 = n8934 ^ n5942 ^ 1'b0 ;
  assign n43166 = ~n8054 & n12319 ;
  assign n43167 = ~n70 & n43166 ;
  assign n43168 = n4857 & ~n43167 ;
  assign n43169 = n43168 ^ n10422 ^ 1'b0 ;
  assign n43170 = n1746 & ~n43169 ;
  assign n43171 = ~n7186 & n13875 ;
  assign n43172 = ~n4545 & n43171 ;
  assign n43173 = n10682 & n43172 ;
  assign n43174 = ~n8070 & n43173 ;
  assign n43175 = n1832 & ~n43174 ;
  assign n43176 = n43174 & n43175 ;
  assign n43177 = ~n18239 & n18465 ;
  assign n43178 = ~n18465 & n43177 ;
  assign n43179 = n43176 | n43178 ;
  assign n43180 = n22200 & ~n43179 ;
  assign n43181 = n36043 ^ n16325 ^ 1'b0 ;
  assign n43182 = n9191 & n19172 ;
  assign n43183 = n31556 & n43182 ;
  assign n43184 = ~n6667 & n30321 ;
  assign n43185 = n43184 ^ n18683 ^ 1'b0 ;
  assign n43186 = n12018 ^ n230 ^ 1'b0 ;
  assign n43187 = n23 & n2992 ;
  assign n43188 = n43187 ^ n14106 ^ 1'b0 ;
  assign n43189 = ~n2434 & n36699 ;
  assign n43190 = ~n1348 & n6562 ;
  assign n43191 = n43190 ^ n7779 ^ 1'b0 ;
  assign n43192 = ~n1022 & n17737 ;
  assign n43193 = n4911 ^ n3546 ^ 1'b0 ;
  assign n43194 = n15122 & ~n43193 ;
  assign n43195 = n43194 ^ n5249 ^ 1'b0 ;
  assign n43196 = n43195 ^ n26317 ^ 1'b0 ;
  assign n43197 = ~n22512 & n43196 ;
  assign n43198 = ~n15112 & n15690 ;
  assign n43199 = ~n38710 & n43198 ;
  assign n43200 = n43199 ^ n9776 ^ 1'b0 ;
  assign n43201 = ( n1991 & n8891 ) | ( n1991 & n20720 ) | ( n8891 & n20720 ) ;
  assign n43202 = n17477 ^ n6531 ^ 1'b0 ;
  assign n43203 = n22734 & ~n43202 ;
  assign n43205 = n7627 | n8656 ;
  assign n43206 = n23089 | n43205 ;
  assign n43207 = n26584 ^ n12198 ^ 1'b0 ;
  assign n43208 = n15653 & ~n43207 ;
  assign n43209 = ~n43206 & n43208 ;
  assign n43210 = n43209 ^ n28868 ^ n12000 ;
  assign n43204 = n12531 | n16675 ;
  assign n43211 = n43210 ^ n43204 ^ 1'b0 ;
  assign n43212 = n17886 & n31078 ;
  assign n43213 = n19435 ^ n18950 ^ n7776 ;
  assign n43214 = n43213 ^ n39250 ^ 1'b0 ;
  assign n43215 = n7654 & n26094 ;
  assign n43216 = ( n2946 & n11267 ) | ( n2946 & n43215 ) | ( n11267 & n43215 ) ;
  assign n43217 = n6498 | n6503 ;
  assign n43218 = ( n19738 & ~n43216 ) | ( n19738 & n43217 ) | ( ~n43216 & n43217 ) ;
  assign n43219 = n5318 | n35820 ;
  assign n43220 = n43219 ^ n12630 ^ n2758 ;
  assign n43221 = ~n29242 & n34372 ;
  assign n43222 = n24418 ^ n11690 ^ 1'b0 ;
  assign n43223 = n25603 ^ n14019 ^ 1'b0 ;
  assign n43224 = n35242 | n43223 ;
  assign n43226 = n27932 & n35593 ;
  assign n43225 = n8355 & ~n41188 ;
  assign n43227 = n43226 ^ n43225 ^ 1'b0 ;
  assign n43228 = n39449 ^ n2953 ^ 1'b0 ;
  assign n43230 = n20969 ^ n4422 ^ n3988 ;
  assign n43229 = n6852 | n36834 ;
  assign n43231 = n43230 ^ n43229 ^ 1'b0 ;
  assign n43232 = n6710 | n23861 ;
  assign n43233 = n23902 & ~n43232 ;
  assign n43234 = n43233 ^ n28637 ^ n3647 ;
  assign n43235 = n43234 ^ n36349 ^ n2994 ;
  assign n43241 = n9624 ^ n8249 ^ 1'b0 ;
  assign n43236 = n16252 ^ n15103 ^ 1'b0 ;
  assign n43237 = ~n3473 & n43236 ;
  assign n43238 = n29548 ^ n12596 ^ 1'b0 ;
  assign n43239 = n43237 & ~n43238 ;
  assign n43240 = ~n6729 & n43239 ;
  assign n43242 = n43241 ^ n43240 ^ 1'b0 ;
  assign n43243 = n8291 & ~n28886 ;
  assign n43244 = n18238 & ~n24210 ;
  assign n43245 = n4614 & n15381 ;
  assign n43246 = ~n34266 & n43245 ;
  assign n43247 = n21544 ^ n8832 ^ 1'b0 ;
  assign n43248 = n3581 & n43247 ;
  assign n43249 = n35197 ^ n21577 ^ 1'b0 ;
  assign n43250 = n23042 | n43249 ;
  assign n43251 = n5323 & n26630 ;
  assign n43252 = n43251 ^ n9563 ^ 1'b0 ;
  assign n43253 = n18966 ^ n8756 ^ 1'b0 ;
  assign n43254 = n9178 & n43253 ;
  assign n43255 = n43254 ^ n29230 ^ 1'b0 ;
  assign n43256 = n14075 & n39568 ;
  assign n43257 = ( n23546 & n23839 ) | ( n23546 & n29040 ) | ( n23839 & n29040 ) ;
  assign n43258 = n28454 ^ n27951 ^ n9552 ;
  assign n43259 = n40932 ^ n33059 ^ 1'b0 ;
  assign n43260 = n13812 ^ n4208 ^ n1531 ;
  assign n43261 = n43260 ^ n27475 ^ n3618 ;
  assign n43262 = n14851 | n43261 ;
  assign n43263 = n8371 | n43262 ;
  assign n43264 = n9818 ^ n685 ^ 1'b0 ;
  assign n43265 = n12139 & ~n39430 ;
  assign n43266 = n4396 & n43265 ;
  assign n43267 = n6650 & ~n43266 ;
  assign n43268 = n43264 & n43267 ;
  assign n43269 = n19664 & n25278 ;
  assign n43270 = n1324 & n43269 ;
  assign n43271 = n4308 | n9141 ;
  assign n43272 = n9760 | n43271 ;
  assign n43273 = n772 & ~n36011 ;
  assign n43274 = ~n43272 & n43273 ;
  assign n43275 = ~n9669 & n31858 ;
  assign n43276 = n43275 ^ n31599 ^ 1'b0 ;
  assign n43277 = ( ~n11549 & n12460 ) | ( ~n11549 & n43276 ) | ( n12460 & n43276 ) ;
  assign n43278 = ~n22173 & n43277 ;
  assign n43279 = n43278 ^ n4728 ^ 1'b0 ;
  assign n43280 = n1363 | n4549 ;
  assign n43281 = n43280 ^ n661 ^ 1'b0 ;
  assign n43282 = ~n32611 & n43281 ;
  assign n43283 = ~n17351 & n43282 ;
  assign n43284 = n78 | n29847 ;
  assign n43286 = n20294 ^ n11954 ^ 1'b0 ;
  assign n43287 = ~n10660 & n43286 ;
  assign n43285 = ~n20970 & n35752 ;
  assign n43288 = n43287 ^ n43285 ^ n1197 ;
  assign n43289 = ~n43284 & n43288 ;
  assign n43290 = n2037 & n7657 ;
  assign n43291 = n12402 & n43290 ;
  assign n43292 = n43291 ^ n2979 ^ 1'b0 ;
  assign n43293 = n31144 & n43292 ;
  assign n43294 = ~n3084 & n43293 ;
  assign n43297 = ( n2595 & n3024 ) | ( n2595 & ~n33153 ) | ( n3024 & ~n33153 ) ;
  assign n43295 = n19409 ^ n11374 ^ n162 ;
  assign n43296 = n43295 ^ n21607 ^ 1'b0 ;
  assign n43298 = n43297 ^ n43296 ^ 1'b0 ;
  assign n43299 = n3192 & n16047 ;
  assign n43300 = n25914 ^ n24628 ^ n3056 ;
  assign n43301 = n43300 ^ n17475 ^ 1'b0 ;
  assign n43302 = n169 & n43301 ;
  assign n43307 = n16373 | n29725 ;
  assign n43303 = n4110 | n9490 ;
  assign n43304 = n43303 ^ n7525 ^ 1'b0 ;
  assign n43305 = n17898 ^ n10459 ^ 1'b0 ;
  assign n43306 = n43304 & n43305 ;
  assign n43308 = n43307 ^ n43306 ^ 1'b0 ;
  assign n43309 = ~n2002 & n13260 ;
  assign n43310 = n10626 & n43309 ;
  assign n43313 = n24131 ^ n15687 ^ n6353 ;
  assign n43311 = ~n11678 & n12187 ;
  assign n43312 = n17493 & ~n43311 ;
  assign n43314 = n43313 ^ n43312 ^ 1'b0 ;
  assign n43315 = n12617 & ~n29872 ;
  assign n43316 = n19564 ^ n1036 ^ 1'b0 ;
  assign n43317 = n13265 & n43316 ;
  assign n43321 = n41564 | n42610 ;
  assign n43318 = n15184 & n22694 ;
  assign n43319 = ~n16207 & n43318 ;
  assign n43320 = n7471 & ~n43319 ;
  assign n43322 = n43321 ^ n43320 ^ 1'b0 ;
  assign n43323 = ~n5634 & n13377 ;
  assign n43324 = n43323 ^ n8240 ^ 1'b0 ;
  assign n43325 = n19356 ^ n9435 ^ n176 ;
  assign n43326 = n15210 | n43325 ;
  assign n43327 = n43324 & ~n43326 ;
  assign n43328 = n20216 & ~n34220 ;
  assign n43329 = n2135 & n19364 ;
  assign n43330 = n41765 ^ n40593 ^ n19212 ;
  assign n43331 = n17518 & n27802 ;
  assign n43332 = ( n11465 & n14657 ) | ( n11465 & ~n17467 ) | ( n14657 & ~n17467 ) ;
  assign n43333 = n10910 & ~n43332 ;
  assign n43334 = n11243 & n29192 ;
  assign n43335 = n5522 & ~n33372 ;
  assign n43336 = n43335 ^ n13870 ^ 1'b0 ;
  assign n43337 = n43334 | n43336 ;
  assign n43338 = n8840 | n19695 ;
  assign n43339 = n43338 ^ n5914 ^ 1'b0 ;
  assign n43340 = n26912 ^ n16950 ^ 1'b0 ;
  assign n43341 = n43339 | n43340 ;
  assign n43342 = n43341 ^ n18828 ^ 1'b0 ;
  assign n43343 = n16611 & n18443 ;
  assign n43344 = ~n26371 & n43343 ;
  assign n43345 = n43344 ^ n39134 ^ 1'b0 ;
  assign n43346 = n4294 & ~n29724 ;
  assign n43347 = n43345 & n43346 ;
  assign n43348 = ~n13063 & n22110 ;
  assign n43349 = n16023 & n25971 ;
  assign n43350 = ~n5747 & n43349 ;
  assign n43351 = n21941 ^ n16523 ^ n511 ;
  assign n43352 = n43351 ^ n36346 ^ n34901 ;
  assign n43353 = n12186 ^ n8656 ^ 1'b0 ;
  assign n43354 = n20423 & ~n43353 ;
  assign n43357 = ~n5672 & n15126 ;
  assign n43358 = ~n18785 & n43357 ;
  assign n43355 = n7977 & ~n16882 ;
  assign n43356 = n43355 ^ n32939 ^ 1'b0 ;
  assign n43359 = n43358 ^ n43356 ^ n676 ;
  assign n43361 = n1265 & ~n6790 ;
  assign n43360 = n5012 | n40565 ;
  assign n43362 = n43361 ^ n43360 ^ 1'b0 ;
  assign n43363 = n9939 & n27605 ;
  assign n43364 = ~n28224 & n42838 ;
  assign n43365 = ( ~n21867 & n32308 ) | ( ~n21867 & n33105 ) | ( n32308 & n33105 ) ;
  assign n43366 = n24793 & ~n38357 ;
  assign n43367 = n43365 & n43366 ;
  assign n43368 = n15394 ^ n14129 ^ 1'b0 ;
  assign n43369 = n12575 ^ n8424 ^ 1'b0 ;
  assign n43370 = n14706 & ~n43369 ;
  assign n43372 = ( n2993 & ~n22479 ) | ( n2993 & n28273 ) | ( ~n22479 & n28273 ) ;
  assign n43371 = n20824 & ~n42809 ;
  assign n43373 = n43372 ^ n43371 ^ 1'b0 ;
  assign n43374 = n38346 ^ n20083 ^ n3626 ;
  assign n43375 = ( n8347 & n35503 ) | ( n8347 & ~n42392 ) | ( n35503 & ~n42392 ) ;
  assign n43376 = n42915 ^ n17360 ^ 1'b0 ;
  assign n43377 = ~n2722 & n43376 ;
  assign n43378 = n2861 ^ n1715 ^ 1'b0 ;
  assign n43379 = n31500 & ~n41487 ;
  assign n43380 = n43379 ^ n30407 ^ 1'b0 ;
  assign n43383 = n7069 & ~n20356 ;
  assign n43381 = n2108 | n2722 ;
  assign n43382 = n14736 & ~n43381 ;
  assign n43384 = n43383 ^ n43382 ^ n6042 ;
  assign n43385 = n43384 ^ n177 ^ 1'b0 ;
  assign n43386 = n24531 ^ n21665 ^ 1'b0 ;
  assign n43387 = ~n43385 & n43386 ;
  assign n43388 = n27799 ^ n16356 ^ 1'b0 ;
  assign n43389 = ~n4917 & n32782 ;
  assign n43390 = ~n17994 & n18061 ;
  assign n43391 = n43390 ^ n22469 ^ n2169 ;
  assign n43392 = ( ~n9184 & n13667 ) | ( ~n9184 & n15134 ) | ( n13667 & n15134 ) ;
  assign n43393 = n43392 ^ n4280 ^ 1'b0 ;
  assign n43394 = n43391 & ~n43393 ;
  assign n43395 = n8789 ^ n561 ^ 1'b0 ;
  assign n43396 = ~n21838 & n43395 ;
  assign n43397 = n39145 ^ n32937 ^ 1'b0 ;
  assign n43398 = ~n3455 & n31635 ;
  assign n43399 = n30107 ^ n28327 ^ n5135 ;
  assign n43400 = ( n13473 & ~n27946 ) | ( n13473 & n43399 ) | ( ~n27946 & n43399 ) ;
  assign n43402 = n12286 ^ n2827 ^ 1'b0 ;
  assign n43401 = n29882 ^ n7268 ^ 1'b0 ;
  assign n43403 = n43402 ^ n43401 ^ n27548 ;
  assign n43404 = n29863 ^ n7001 ^ n6358 ;
  assign n43405 = n42 | n5718 ;
  assign n43406 = n43405 ^ n9168 ^ 1'b0 ;
  assign n43407 = n29382 | n43406 ;
  assign n43408 = n14016 ^ n13730 ^ 1'b0 ;
  assign n43409 = n26216 & ~n43408 ;
  assign n43410 = ~n2287 & n7332 ;
  assign n43411 = n8356 & n43410 ;
  assign n43412 = ~n36824 & n43411 ;
  assign n43413 = n43412 ^ n3130 ^ 1'b0 ;
  assign n43414 = n19080 | n43413 ;
  assign n43415 = n28375 & ~n43414 ;
  assign n43416 = ( n25042 & ~n29788 ) | ( n25042 & n40904 ) | ( ~n29788 & n40904 ) ;
  assign n43419 = n38683 ^ n12883 ^ n3165 ;
  assign n43420 = n43261 & n43419 ;
  assign n43417 = ~n517 & n22429 ;
  assign n43418 = n43417 ^ n14829 ^ 1'b0 ;
  assign n43421 = n43420 ^ n43418 ^ n19294 ;
  assign n43422 = n40615 ^ n21842 ^ n8891 ;
  assign n43423 = n11233 | n23108 ;
  assign n43424 = n23528 & ~n29391 ;
  assign n43425 = ~n5101 & n14216 ;
  assign n43426 = ~n5139 & n43425 ;
  assign n43427 = n27882 ^ n9860 ^ 1'b0 ;
  assign n43428 = n17160 | n43427 ;
  assign n43429 = n25878 ^ n20496 ^ 1'b0 ;
  assign n43430 = n521 | n3273 ;
  assign n43431 = n7853 & ~n43430 ;
  assign n43432 = n43431 ^ n875 ^ 1'b0 ;
  assign n43433 = n28071 ^ n2214 ^ 1'b0 ;
  assign n43434 = n9012 | n23787 ;
  assign n43435 = n11010 & ~n25958 ;
  assign n43436 = n20727 ^ n11454 ^ 1'b0 ;
  assign n43437 = n32077 ^ n6389 ^ 1'b0 ;
  assign n43438 = n43436 | n43437 ;
  assign n43439 = n28323 ^ n11544 ^ 1'b0 ;
  assign n43440 = n43438 | n43439 ;
  assign n43441 = n31622 & ~n42614 ;
  assign n43442 = ~n8142 & n43441 ;
  assign n43443 = n19191 ^ n8952 ^ 1'b0 ;
  assign n43444 = n15981 ^ n15145 ^ 1'b0 ;
  assign n43445 = n43443 & ~n43444 ;
  assign n43446 = n26105 ^ n1177 ^ 1'b0 ;
  assign n43447 = n41918 | n43446 ;
  assign n43448 = n43445 & n43447 ;
  assign n43449 = n8150 ^ n2693 ^ 1'b0 ;
  assign n43450 = n3566 & ~n19638 ;
  assign n43451 = n16453 & n43450 ;
  assign n43452 = n43449 & ~n43451 ;
  assign n43453 = ~n1330 & n8925 ;
  assign n43454 = n43453 ^ n3660 ^ 1'b0 ;
  assign n43455 = n32174 ^ n6916 ^ 1'b0 ;
  assign n43456 = ~n1682 & n43455 ;
  assign n43457 = ( n41496 & n43454 ) | ( n41496 & ~n43456 ) | ( n43454 & ~n43456 ) ;
  assign n43458 = ( n2135 & n4110 ) | ( n2135 & n23963 ) | ( n4110 & n23963 ) ;
  assign n43459 = n6703 & n8278 ;
  assign n43460 = n5113 & n43459 ;
  assign n43461 = n18001 & ~n43460 ;
  assign n43462 = ~n16258 & n43461 ;
  assign n43463 = n1812 & ~n15932 ;
  assign n43464 = n5092 & n43463 ;
  assign n43465 = n9939 | n43464 ;
  assign n43466 = n22721 & n26317 ;
  assign n43467 = n18242 | n35951 ;
  assign n43468 = ~n35663 & n43467 ;
  assign n43469 = n35461 ^ n19062 ^ 1'b0 ;
  assign n43470 = n3327 | n19974 ;
  assign n43471 = n4328 & ~n43470 ;
  assign n43472 = n4693 ^ n45 ^ 1'b0 ;
  assign n43473 = n2370 & ~n15803 ;
  assign n43474 = n43473 ^ n16298 ^ 1'b0 ;
  assign n43476 = n11794 & n36661 ;
  assign n43477 = ~n15933 & n43476 ;
  assign n43478 = n43477 ^ n2214 ^ 1'b0 ;
  assign n43475 = ( n3009 & ~n6361 ) | ( n3009 & n10239 ) | ( ~n6361 & n10239 ) ;
  assign n43479 = n43478 ^ n43475 ^ n8183 ;
  assign n43480 = n34351 ^ n350 ^ 1'b0 ;
  assign n43481 = n43479 | n43480 ;
  assign n43482 = n28524 | n43481 ;
  assign n43483 = n6316 ^ x10 ^ 1'b0 ;
  assign n43484 = n33415 & ~n43483 ;
  assign n43485 = n24040 ^ n691 ^ 1'b0 ;
  assign n43486 = n38901 ^ n10059 ^ 1'b0 ;
  assign n43487 = n5099 & ~n43486 ;
  assign n43488 = ~n43485 & n43487 ;
  assign n43489 = n43488 ^ n37831 ^ 1'b0 ;
  assign n43490 = n43489 ^ n12570 ^ 1'b0 ;
  assign n43491 = n1336 & n25615 ;
  assign n43492 = n43491 ^ n27347 ^ 1'b0 ;
  assign n43493 = n10977 & ~n37629 ;
  assign n43494 = n43493 ^ n17455 ^ 1'b0 ;
  assign n43495 = n29276 & ~n43427 ;
  assign n43499 = n3652 & n14776 ;
  assign n43500 = n43499 ^ n12742 ^ 1'b0 ;
  assign n43496 = n40738 ^ n9729 ^ 1'b0 ;
  assign n43497 = ~n8838 & n43496 ;
  assign n43498 = ~n9095 & n43497 ;
  assign n43501 = n43500 ^ n43498 ^ 1'b0 ;
  assign n43502 = n14433 & ~n37607 ;
  assign n43503 = n43502 ^ n3367 ^ 1'b0 ;
  assign n43504 = n7534 | n18008 ;
  assign n43505 = n43503 | n43504 ;
  assign n43507 = ~n11690 & n25624 ;
  assign n43508 = n43507 ^ n7428 ^ 1'b0 ;
  assign n43509 = n20578 & ~n43508 ;
  assign n43506 = n8663 & ~n25955 ;
  assign n43510 = n43509 ^ n43506 ^ 1'b0 ;
  assign n43511 = ~n17164 & n31657 ;
  assign n43512 = n4097 & n43511 ;
  assign n43513 = ~n3899 & n43512 ;
  assign n43514 = n20246 ^ n7001 ^ 1'b0 ;
  assign n43518 = n3641 | n22003 ;
  assign n43515 = ~n1668 & n5909 ;
  assign n43516 = n6833 & n43515 ;
  assign n43517 = n7165 & n43516 ;
  assign n43519 = n43518 ^ n43517 ^ 1'b0 ;
  assign n43520 = n43519 ^ n29842 ^ 1'b0 ;
  assign n43521 = n43520 ^ n43487 ^ n1262 ;
  assign n43522 = n40492 ^ n35201 ^ n22424 ;
  assign n43523 = n5442 & n14996 ;
  assign n43524 = n7344 & n43523 ;
  assign n43525 = n21931 | n43524 ;
  assign n43526 = n43525 ^ n28819 ^ 1'b0 ;
  assign n43527 = n16630 ^ n8140 ^ 1'b0 ;
  assign n43528 = n25445 ^ n15821 ^ n13479 ;
  assign n43529 = n43528 ^ n16637 ^ 1'b0 ;
  assign n43530 = n43529 ^ n30576 ^ 1'b0 ;
  assign n43531 = ~n43527 & n43530 ;
  assign n43532 = n1961 ^ n1709 ^ 1'b0 ;
  assign n43533 = n9503 | n12088 ;
  assign n43534 = n43533 ^ n13841 ^ 1'b0 ;
  assign n43535 = n17366 & ~n43534 ;
  assign n43536 = n43535 ^ n11466 ^ n7864 ;
  assign n43538 = n18339 ^ n13477 ^ 1'b0 ;
  assign n43539 = ~n5909 & n43538 ;
  assign n43540 = ~n4505 & n43539 ;
  assign n43541 = n10197 ^ n8073 ^ 1'b0 ;
  assign n43542 = n43540 & n43541 ;
  assign n43537 = n21991 ^ n15857 ^ 1'b0 ;
  assign n43543 = n43542 ^ n43537 ^ 1'b0 ;
  assign n43544 = n4001 & ~n16155 ;
  assign n43545 = ~n21045 & n43544 ;
  assign n43546 = n38655 ^ n7534 ^ 1'b0 ;
  assign n43547 = n43545 | n43546 ;
  assign n43549 = ~n313 & n16323 ;
  assign n43548 = n16678 & n32501 ;
  assign n43550 = n43549 ^ n43548 ^ 1'b0 ;
  assign n43551 = ~n5873 & n43550 ;
  assign n43552 = n11652 & ~n39081 ;
  assign n43553 = n43552 ^ n10780 ^ 1'b0 ;
  assign n43554 = n7722 | n9666 ;
  assign n43555 = n43554 ^ n2095 ^ 1'b0 ;
  assign n43556 = ( ~n20543 & n35569 ) | ( ~n20543 & n43555 ) | ( n35569 & n43555 ) ;
  assign n43557 = n9184 ^ n4290 ^ 1'b0 ;
  assign n43558 = n14706 & ~n43557 ;
  assign n43559 = n2020 & ~n5652 ;
  assign n43560 = n5652 & n43559 ;
  assign n43561 = ~n1032 & n43560 ;
  assign n43562 = n41365 ^ n9560 ^ n3747 ;
  assign n43563 = ( n18210 & ~n43561 ) | ( n18210 & n43562 ) | ( ~n43561 & n43562 ) ;
  assign n43564 = n5641 & n8265 ;
  assign n43565 = n43564 ^ n5001 ^ 1'b0 ;
  assign n43566 = n2698 & n43565 ;
  assign n43567 = n28080 & ~n32545 ;
  assign n43568 = n36963 ^ n21646 ^ 1'b0 ;
  assign n43569 = n15702 ^ n384 ^ 1'b0 ;
  assign n43570 = n20157 & n43569 ;
  assign n43571 = ~n14129 & n15420 ;
  assign n43572 = n7160 & ~n43571 ;
  assign n43573 = n43572 ^ n32827 ^ n927 ;
  assign n43574 = n43570 & ~n43573 ;
  assign n43575 = n20470 ^ n15849 ^ 1'b0 ;
  assign n43576 = n10190 ^ n2259 ^ 1'b0 ;
  assign n43577 = n22171 & n43576 ;
  assign n43578 = n43577 ^ n17811 ^ 1'b0 ;
  assign n43579 = ~n29685 & n43578 ;
  assign n43580 = n23411 ^ n16661 ^ 1'b0 ;
  assign n43581 = n36035 ^ n16381 ^ n13218 ;
  assign n43582 = ~n5370 & n43581 ;
  assign n43583 = n43582 ^ n12952 ^ 1'b0 ;
  assign n43584 = n13298 & n34728 ;
  assign n43585 = n15401 | n16480 ;
  assign n43586 = n30094 ^ n24695 ^ 1'b0 ;
  assign n43587 = n15498 ^ n6107 ^ 1'b0 ;
  assign n43588 = n4247 | n43587 ;
  assign n43589 = n17859 ^ n1697 ^ 1'b0 ;
  assign n43590 = ( ~n19973 & n37672 ) | ( ~n19973 & n43589 ) | ( n37672 & n43589 ) ;
  assign n43591 = n15259 | n43590 ;
  assign n43592 = n43591 ^ n16476 ^ 1'b0 ;
  assign n43593 = ~n22664 & n43592 ;
  assign n43594 = n43588 & n43593 ;
  assign n43595 = ~n17854 & n25283 ;
  assign n43596 = ( n4862 & n5578 ) | ( n4862 & n43595 ) | ( n5578 & n43595 ) ;
  assign n43597 = n43596 ^ n24447 ^ 1'b0 ;
  assign n43598 = n14488 ^ n3386 ^ 1'b0 ;
  assign n43599 = ~n919 & n43598 ;
  assign n43600 = ( ~n35600 & n38133 ) | ( ~n35600 & n43599 ) | ( n38133 & n43599 ) ;
  assign n43601 = n37820 ^ n22562 ^ n13023 ;
  assign n43602 = n4906 & n24400 ;
  assign n43603 = n43602 ^ n28972 ^ 1'b0 ;
  assign n43604 = n27382 ^ n3238 ^ 1'b0 ;
  assign n43605 = n2991 & n25090 ;
  assign n43606 = n43605 ^ n12466 ^ 1'b0 ;
  assign n43608 = n7586 | n20819 ;
  assign n43609 = n26518 | n43608 ;
  assign n43607 = ~n1177 & n22202 ;
  assign n43610 = n43609 ^ n43607 ^ n11534 ;
  assign n43620 = ~n10212 & n12459 ;
  assign n43611 = n11046 & n16966 ;
  assign n43612 = n43611 ^ n9363 ^ 1'b0 ;
  assign n43614 = n3398 & ~n8288 ;
  assign n43615 = ~n3398 & n43614 ;
  assign n43616 = n12481 & n43615 ;
  assign n43613 = n7650 & n40822 ;
  assign n43617 = n43616 ^ n43613 ^ 1'b0 ;
  assign n43618 = n43617 ^ n774 ^ 1'b0 ;
  assign n43619 = ~n43612 & n43618 ;
  assign n43621 = n43620 ^ n43619 ^ 1'b0 ;
  assign n43622 = n37403 ^ n35982 ^ n33885 ;
  assign n43623 = n29653 ^ n14545 ^ 1'b0 ;
  assign n43624 = n37009 & n43623 ;
  assign n43625 = n43624 ^ n8024 ^ n2492 ;
  assign n43626 = n15092 & ~n17015 ;
  assign n43627 = ~n43625 & n43626 ;
  assign n43629 = n42805 ^ n1639 ^ 1'b0 ;
  assign n43630 = ~n26139 & n43629 ;
  assign n43628 = ~n14460 & n36056 ;
  assign n43631 = n43630 ^ n43628 ^ 1'b0 ;
  assign n43632 = n33836 ^ n22220 ^ 1'b0 ;
  assign n43633 = n5538 | n13154 ;
  assign n43634 = n43633 ^ n3814 ^ 1'b0 ;
  assign n43635 = ( ~n14775 & n34793 ) | ( ~n14775 & n43634 ) | ( n34793 & n43634 ) ;
  assign n43636 = ( n17377 & n25312 ) | ( n17377 & ~n27619 ) | ( n25312 & ~n27619 ) ;
  assign n43637 = n17991 & ~n32623 ;
  assign n43638 = ~n43636 & n43637 ;
  assign n43639 = ( ~n10718 & n24252 ) | ( ~n10718 & n43638 ) | ( n24252 & n43638 ) ;
  assign n43640 = n15442 ^ n1202 ^ 1'b0 ;
  assign n43641 = n42268 & ~n43640 ;
  assign n43642 = n43641 ^ n26556 ^ 1'b0 ;
  assign n43643 = n7831 & n43642 ;
  assign n43644 = n8195 ^ n5602 ^ 1'b0 ;
  assign n43645 = n42140 & n43644 ;
  assign n43646 = n43645 ^ n5294 ^ 1'b0 ;
  assign n43647 = n426 | n43646 ;
  assign n43648 = n7932 & n20356 ;
  assign n43649 = n13632 & n43648 ;
  assign n43650 = n8624 & ~n43649 ;
  assign n43652 = n21296 ^ n10141 ^ 1'b0 ;
  assign n43651 = n3679 & n36194 ;
  assign n43653 = n43652 ^ n43651 ^ 1'b0 ;
  assign n43654 = ~n2372 & n24332 ;
  assign n43655 = n43654 ^ n16451 ^ 1'b0 ;
  assign n43656 = n38827 ^ n29490 ^ n19957 ;
  assign n43657 = ( n14571 & n38481 ) | ( n14571 & ~n43656 ) | ( n38481 & ~n43656 ) ;
  assign n43658 = n16177 & n16758 ;
  assign n43659 = n12353 | n14443 ;
  assign n43660 = n4590 | n43659 ;
  assign n43661 = n2174 & ~n43660 ;
  assign n43662 = n43661 ^ n10348 ^ 1'b0 ;
  assign n43663 = n11648 & n32073 ;
  assign n43664 = ~n14895 & n43663 ;
  assign n43665 = n31084 ^ n6163 ^ 1'b0 ;
  assign n43666 = n14712 & n43665 ;
  assign n43667 = n5808 | n43666 ;
  assign n43668 = n11956 ^ n366 ^ 1'b0 ;
  assign n43669 = n43667 & ~n43668 ;
  assign n43670 = n23611 ^ n9548 ^ 1'b0 ;
  assign n43671 = n2108 & n43670 ;
  assign n43672 = n2789 | n10090 ;
  assign n43673 = n21985 & n39993 ;
  assign n43674 = n43673 ^ n19530 ^ 1'b0 ;
  assign n43675 = ( n3961 & ~n23379 ) | ( n3961 & n43674 ) | ( ~n23379 & n43674 ) ;
  assign n43676 = n3142 & n10385 ;
  assign n43677 = n2294 & n2409 ;
  assign n43678 = ( n14873 & n23885 ) | ( n14873 & n43677 ) | ( n23885 & n43677 ) ;
  assign n43679 = n43678 ^ n6804 ^ 1'b0 ;
  assign n43680 = n43676 | n43679 ;
  assign n43681 = n28078 ^ n12357 ^ n8683 ;
  assign n43682 = n18301 ^ n12994 ^ 1'b0 ;
  assign n43683 = n23124 | n30206 ;
  assign n43684 = n36000 | n43683 ;
  assign n43685 = n3496 & ~n36966 ;
  assign n43686 = n5353 ^ n1784 ^ 1'b0 ;
  assign n43687 = n5414 ^ n1736 ^ 1'b0 ;
  assign n43688 = n7457 & ~n43687 ;
  assign n43689 = n15341 | n43688 ;
  assign n43690 = ~n13172 & n34398 ;
  assign n43691 = n43690 ^ n22626 ^ 1'b0 ;
  assign n43692 = n43691 ^ n36973 ^ n11891 ;
  assign n43693 = n14665 ^ n10055 ^ 1'b0 ;
  assign n43694 = n15774 & ~n37510 ;
  assign n43695 = n42530 ^ n5331 ^ 1'b0 ;
  assign n43696 = ~n43694 & n43695 ;
  assign n43698 = n16343 | n19083 ;
  assign n43699 = n43698 ^ n34227 ^ 1'b0 ;
  assign n43697 = n5919 & ~n34752 ;
  assign n43700 = n43699 ^ n43697 ^ 1'b0 ;
  assign n43704 = n4543 & ~n12102 ;
  assign n43705 = ( n2504 & ~n15473 ) | ( n2504 & n43704 ) | ( ~n15473 & n43704 ) ;
  assign n43701 = ~n5952 & n36376 ;
  assign n43702 = ~n842 & n3390 ;
  assign n43703 = n43701 & ~n43702 ;
  assign n43706 = n43705 ^ n43703 ^ 1'b0 ;
  assign n43707 = n570 ^ n101 ^ 1'b0 ;
  assign n43708 = n694 | n43707 ;
  assign n43709 = n14195 & ~n43708 ;
  assign n43710 = n7920 & ~n43709 ;
  assign n43711 = ~n28801 & n43710 ;
  assign n43712 = n10822 ^ n4097 ^ n2466 ;
  assign n43713 = n43712 ^ n9824 ^ 1'b0 ;
  assign n43714 = n43711 | n43713 ;
  assign n43715 = ~n12672 & n35855 ;
  assign n43716 = n43715 ^ n29942 ^ 1'b0 ;
  assign n43717 = ~n16117 & n43716 ;
  assign n43718 = n27989 ^ n20759 ^ 1'b0 ;
  assign n43719 = n9947 | n43718 ;
  assign n43720 = n43719 ^ n7650 ^ n4264 ;
  assign n43721 = n11725 & n43720 ;
  assign n43722 = n32002 ^ n22556 ^ 1'b0 ;
  assign n43723 = n2813 ^ n2657 ^ 1'b0 ;
  assign n43724 = ( n9404 & ~n15866 ) | ( n9404 & n43723 ) | ( ~n15866 & n43723 ) ;
  assign n43725 = n2693 & ~n43724 ;
  assign n43726 = ~n11264 & n43667 ;
  assign n43727 = n23012 ^ n15060 ^ 1'b0 ;
  assign n43728 = n26190 & ~n43727 ;
  assign n43729 = n32413 ^ n17964 ^ 1'b0 ;
  assign n43730 = n14175 & ~n43729 ;
  assign n43731 = ( n11420 & n38348 ) | ( n11420 & n43730 ) | ( n38348 & n43730 ) ;
  assign n43732 = n43731 ^ n4048 ^ 1'b0 ;
  assign n43733 = ( n5794 & n20340 ) | ( n5794 & ~n22878 ) | ( n20340 & ~n22878 ) ;
  assign n43734 = n3035 & ~n9933 ;
  assign n43735 = n43734 ^ n36035 ^ n19800 ;
  assign n43736 = ~n28108 & n43735 ;
  assign n43737 = n13943 ^ n6979 ^ 1'b0 ;
  assign n43738 = n43737 ^ n1341 ^ 1'b0 ;
  assign n43739 = n41261 ^ n26965 ^ 1'b0 ;
  assign n43740 = n13488 & ~n13633 ;
  assign n43741 = ( ~n25508 & n43739 ) | ( ~n25508 & n43740 ) | ( n43739 & n43740 ) ;
  assign n43742 = n19044 & n41793 ;
  assign n43743 = n43742 ^ n2595 ^ 1'b0 ;
  assign n43744 = ~n20061 & n39961 ;
  assign n43745 = n3123 & n43744 ;
  assign n43746 = n9739 ^ n1716 ^ 1'b0 ;
  assign n43747 = ~n16047 & n43746 ;
  assign n43748 = n31315 ^ n6609 ^ 1'b0 ;
  assign n43749 = n43748 ^ n7208 ^ 1'b0 ;
  assign n43750 = n7873 | n43749 ;
  assign n43751 = n4288 & n33989 ;
  assign n43752 = n43751 ^ n30160 ^ 1'b0 ;
  assign n43753 = n42040 ^ n26857 ^ n16179 ;
  assign n43754 = n43753 ^ n12539 ^ n11910 ;
  assign n43755 = ( n4463 & n19108 ) | ( n4463 & n43754 ) | ( n19108 & n43754 ) ;
  assign n43757 = ( n3537 & n20793 ) | ( n3537 & ~n28548 ) | ( n20793 & ~n28548 ) ;
  assign n43756 = n27991 ^ n14914 ^ n13198 ;
  assign n43758 = n43757 ^ n43756 ^ n22071 ;
  assign n43759 = n35847 ^ n29467 ^ n13616 ;
  assign n43760 = n43759 ^ n14298 ^ 1'b0 ;
  assign n43761 = n1411 & ~n43760 ;
  assign n43762 = n21804 ^ n2784 ^ 1'b0 ;
  assign n43763 = ( ~n6079 & n13881 ) | ( ~n6079 & n31457 ) | ( n13881 & n31457 ) ;
  assign n43764 = n43763 ^ n22292 ^ n7962 ;
  assign n43765 = n7047 & ~n19712 ;
  assign n43766 = n43765 ^ n18559 ^ 1'b0 ;
  assign n43767 = n5139 | n14457 ;
  assign n43768 = ~n42507 & n43767 ;
  assign n43769 = n43768 ^ n16648 ^ 1'b0 ;
  assign n43770 = ~n34081 & n40251 ;
  assign n43771 = n14555 & n43770 ;
  assign n43772 = n12082 ^ n8993 ^ 1'b0 ;
  assign n43773 = n38637 ^ n5955 ^ 1'b0 ;
  assign n43774 = n43772 & n43773 ;
  assign n43775 = n36746 ^ n2165 ^ 1'b0 ;
  assign n43778 = n461 & ~n6660 ;
  assign n43777 = ~n1421 & n16728 ;
  assign n43779 = n43778 ^ n43777 ^ 1'b0 ;
  assign n43776 = n8907 & ~n10652 ;
  assign n43780 = n43779 ^ n43776 ^ 1'b0 ;
  assign n43781 = n23737 | n43780 ;
  assign n43782 = ~n14758 & n22613 ;
  assign n43783 = n43782 ^ n14967 ^ 1'b0 ;
  assign n43784 = n19300 ^ n4869 ^ 1'b0 ;
  assign n43785 = n20532 ^ n2841 ^ 1'b0 ;
  assign n43786 = ~n39061 & n43785 ;
  assign n43787 = n43786 ^ n3971 ^ 1'b0 ;
  assign n43788 = ~n6312 & n14132 ;
  assign n43789 = ~n32157 & n43788 ;
  assign n43790 = n43789 ^ n16453 ^ 1'b0 ;
  assign n43791 = n15382 & ~n43199 ;
  assign n43793 = n1108 & ~n9919 ;
  assign n43792 = ~n15525 & n32796 ;
  assign n43794 = n43793 ^ n43792 ^ 1'b0 ;
  assign n43795 = n33170 | n43794 ;
  assign n43796 = ~n3375 & n5696 ;
  assign n43797 = n43796 ^ n30050 ^ 1'b0 ;
  assign n43798 = ~n1842 & n15468 ;
  assign n43799 = n19191 ^ n17883 ^ 1'b0 ;
  assign n43800 = n17287 & ~n43799 ;
  assign n43801 = n43800 ^ n15590 ^ 1'b0 ;
  assign n43802 = n39365 & n43801 ;
  assign n43803 = n7641 & n22521 ;
  assign n43804 = ~n18613 & n40423 ;
  assign n43805 = ~n3866 & n15046 ;
  assign n43806 = n43805 ^ n5537 ^ 1'b0 ;
  assign n43810 = n8265 | n18454 ;
  assign n43807 = n1699 | n15657 ;
  assign n43808 = n32676 | n43807 ;
  assign n43809 = n43808 ^ n32696 ^ 1'b0 ;
  assign n43811 = n43810 ^ n43809 ^ n8160 ;
  assign n43812 = n15679 & ~n43811 ;
  assign n43813 = n43812 ^ n8790 ^ 1'b0 ;
  assign n43814 = n25978 & n43277 ;
  assign n43816 = n37534 ^ n4129 ^ 1'b0 ;
  assign n43815 = ~n19891 & n25420 ;
  assign n43817 = n43816 ^ n43815 ^ 1'b0 ;
  assign n43818 = n8128 | n43817 ;
  assign n43819 = n43818 ^ n17702 ^ 1'b0 ;
  assign n43820 = n491 & n25045 ;
  assign n43821 = n10827 & n43820 ;
  assign n43822 = n16805 ^ n16075 ^ 1'b0 ;
  assign n43823 = n1056 & n43822 ;
  assign n43824 = n8575 ^ n2655 ^ 1'b0 ;
  assign n43825 = ~n1589 & n43824 ;
  assign n43826 = ~n43823 & n43825 ;
  assign n43827 = n15391 | n17472 ;
  assign n43828 = n7968 | n43827 ;
  assign n43829 = n21954 ^ n10568 ^ 1'b0 ;
  assign n43830 = n37589 & n43829 ;
  assign n43831 = ( ~n13610 & n14664 ) | ( ~n13610 & n43830 ) | ( n14664 & n43830 ) ;
  assign n43832 = n77 & ~n32446 ;
  assign n43833 = n19903 & ~n19986 ;
  assign n43834 = n40723 & n43833 ;
  assign n43835 = n43834 ^ n5595 ^ 1'b0 ;
  assign n43836 = n16548 & n26239 ;
  assign n43837 = n43836 ^ n41941 ^ 1'b0 ;
  assign n43838 = n18273 & ~n43837 ;
  assign n43839 = n43838 ^ n45 ^ 1'b0 ;
  assign n43840 = ( n4560 & n18453 ) | ( n4560 & ~n22918 ) | ( n18453 & ~n22918 ) ;
  assign n43841 = n36113 ^ n30704 ^ 1'b0 ;
  assign n43842 = n43840 | n43841 ;
  assign n43843 = ~n6765 & n42630 ;
  assign n43844 = ~n21482 & n43843 ;
  assign n43845 = ~n1247 & n41100 ;
  assign n43846 = n43844 & n43845 ;
  assign n43847 = n7975 & ~n41772 ;
  assign n43848 = n43847 ^ n33091 ^ 1'b0 ;
  assign n43849 = n10764 | n18598 ;
  assign n43851 = n1856 & n27612 ;
  assign n43850 = n8299 & ~n29931 ;
  assign n43852 = n43851 ^ n43850 ^ 1'b0 ;
  assign n43853 = n43852 ^ n29163 ^ n9135 ;
  assign n43854 = n16309 ^ n1421 ^ 1'b0 ;
  assign n43855 = n886 | n43854 ;
  assign n43856 = n43855 ^ n23845 ^ 1'b0 ;
  assign n43857 = n16129 & n17402 ;
  assign n43858 = n43857 ^ n12090 ^ 1'b0 ;
  assign n43859 = ~n26620 & n43858 ;
  assign n43860 = n361 & ~n43859 ;
  assign n43861 = ~n863 & n12926 ;
  assign n43862 = n30398 & ~n36536 ;
  assign n43863 = n33405 | n37559 ;
  assign n43864 = n4281 | n43863 ;
  assign n43865 = n1118 & ~n14491 ;
  assign n43866 = n42707 ^ n37854 ^ 1'b0 ;
  assign n43867 = n7992 | n43866 ;
  assign n43868 = ( n9369 & n42602 ) | ( n9369 & n43867 ) | ( n42602 & n43867 ) ;
  assign n43869 = n40427 ^ n2256 ^ 1'b0 ;
  assign n43870 = ~n5298 & n36301 ;
  assign n43871 = n15531 ^ n14425 ^ 1'b0 ;
  assign n43872 = n10816 & n43871 ;
  assign n43873 = n9195 ^ n2070 ^ 1'b0 ;
  assign n43874 = n43872 & ~n43873 ;
  assign n43875 = n39068 ^ n29892 ^ 1'b0 ;
  assign n43876 = n29238 & n43875 ;
  assign n43877 = n18877 ^ n15958 ^ n2327 ;
  assign n43878 = ( ~n18069 & n21932 ) | ( ~n18069 & n43877 ) | ( n21932 & n43877 ) ;
  assign n43879 = ~n9577 & n21892 ;
  assign n43880 = n43878 & n43879 ;
  assign n43881 = n38845 & ~n43880 ;
  assign n43882 = n20086 | n21172 ;
  assign n43883 = n43882 ^ n13693 ^ 1'b0 ;
  assign n43884 = n2650 | n41061 ;
  assign n43885 = n5137 & ~n43884 ;
  assign n43886 = ( n3191 & n7726 ) | ( n3191 & ~n34958 ) | ( n7726 & ~n34958 ) ;
  assign n43887 = n43886 ^ n20282 ^ 1'b0 ;
  assign n43888 = n22453 ^ n303 ^ 1'b0 ;
  assign n43889 = n8965 & ~n43888 ;
  assign n43890 = n24290 & ~n43889 ;
  assign n43891 = n1448 | n7008 ;
  assign n43892 = ~n29697 & n32995 ;
  assign n43893 = n43892 ^ n3290 ^ 1'b0 ;
  assign n43894 = n43893 ^ n15744 ^ n6333 ;
  assign n43899 = n2563 & n21820 ;
  assign n43900 = n43899 ^ n757 ^ 1'b0 ;
  assign n43897 = n5444 & n11647 ;
  assign n43895 = n16269 ^ n8945 ^ 1'b0 ;
  assign n43896 = n30964 | n43895 ;
  assign n43898 = n43897 ^ n43896 ^ 1'b0 ;
  assign n43901 = n43900 ^ n43898 ^ n14414 ;
  assign n43902 = n16481 ^ n2201 ^ 1'b0 ;
  assign n43903 = n21742 & n43902 ;
  assign n43906 = n14640 | n42294 ;
  assign n43907 = n14572 | n43906 ;
  assign n43904 = n14979 ^ n6451 ^ n1213 ;
  assign n43905 = n40405 | n43904 ;
  assign n43908 = n43907 ^ n43905 ^ 1'b0 ;
  assign n43909 = ~n10572 & n13161 ;
  assign n43910 = ~n6679 & n43909 ;
  assign n43911 = n40659 | n43910 ;
  assign n43912 = n43911 ^ n1386 ^ 1'b0 ;
  assign n43913 = n7130 ^ n6605 ^ 1'b0 ;
  assign n43914 = n39546 & ~n43913 ;
  assign n43915 = n30514 ^ n14504 ^ 1'b0 ;
  assign n43916 = n29664 | n43915 ;
  assign n43917 = n43449 ^ n12422 ^ n11272 ;
  assign n43918 = n43917 ^ n12941 ^ 1'b0 ;
  assign n43919 = n37626 ^ n20470 ^ n3040 ;
  assign n43920 = n43919 ^ n24939 ^ n4283 ;
  assign n43921 = n19135 & n31063 ;
  assign n43922 = n15243 & n24888 ;
  assign n43923 = n43921 & n43922 ;
  assign n43924 = n4297 & n12449 ;
  assign n43925 = n4308 & ~n43924 ;
  assign n43926 = n8348 ^ n4557 ^ 1'b0 ;
  assign n43927 = n27789 & n43926 ;
  assign n43928 = n27041 & ~n28629 ;
  assign n43929 = ~n22012 & n43928 ;
  assign n43930 = n16802 | n32500 ;
  assign n43931 = n7858 | n14207 ;
  assign n43932 = n43931 ^ n20 ^ 1'b0 ;
  assign n43933 = ~n17694 & n18060 ;
  assign n43934 = n43933 ^ n17112 ^ 1'b0 ;
  assign n43935 = n25504 & n33154 ;
  assign n43936 = n1869 | n38468 ;
  assign n43937 = n20142 ^ n8184 ^ 1'b0 ;
  assign n43938 = n34369 & ~n43937 ;
  assign n43939 = ~n4576 & n43938 ;
  assign n43940 = n30850 | n43939 ;
  assign n43941 = n17732 & ~n43940 ;
  assign n43944 = n3510 & n24251 ;
  assign n43942 = n3408 & ~n30432 ;
  assign n43943 = n1483 & ~n43942 ;
  assign n43945 = n43944 ^ n43943 ^ 1'b0 ;
  assign n43948 = n5014 & ~n27543 ;
  assign n43946 = n28847 ^ n27920 ^ 1'b0 ;
  assign n43947 = n16256 | n43946 ;
  assign n43949 = n43948 ^ n43947 ^ n26189 ;
  assign n43950 = n6261 & n37285 ;
  assign n43951 = n7104 ^ n1972 ^ 1'b0 ;
  assign n43952 = n30260 ^ n9526 ^ 1'b0 ;
  assign n43953 = n38018 & ~n43952 ;
  assign n43954 = n20698 & n33895 ;
  assign n43955 = n43954 ^ n2861 ^ 1'b0 ;
  assign n43956 = n5344 & ~n12111 ;
  assign n43957 = n9936 | n38041 ;
  assign n43958 = n32931 ^ n15533 ^ 1'b0 ;
  assign n43959 = n11558 | n43958 ;
  assign n43960 = ~n15544 & n36279 ;
  assign n43961 = n33690 & n43960 ;
  assign n43962 = ~n43959 & n43961 ;
  assign n43963 = n43962 ^ n20646 ^ 1'b0 ;
  assign n43964 = n24942 | n37396 ;
  assign n43965 = n43964 ^ n15841 ^ 1'b0 ;
  assign n43966 = n3918 | n17988 ;
  assign n43967 = n3603 & ~n5233 ;
  assign n43968 = n26611 & ~n43967 ;
  assign n43969 = n5001 & n29453 ;
  assign n43970 = ~n31005 & n43969 ;
  assign n43971 = ( n25292 & n28652 ) | ( n25292 & ~n40822 ) | ( n28652 & ~n40822 ) ;
  assign n43972 = n22147 | n43971 ;
  assign n43975 = ( n7006 & n12013 ) | ( n7006 & ~n27959 ) | ( n12013 & ~n27959 ) ;
  assign n43973 = ( n39 & n358 ) | ( n39 & n31245 ) | ( n358 & n31245 ) ;
  assign n43974 = n10665 | n43973 ;
  assign n43976 = n43975 ^ n43974 ^ 1'b0 ;
  assign n43977 = n22606 ^ n15244 ^ 1'b0 ;
  assign n43978 = ~n18288 & n43977 ;
  assign n43979 = ( n8830 & ~n16628 ) | ( n8830 & n43978 ) | ( ~n16628 & n43978 ) ;
  assign n43980 = n30634 ^ n6246 ^ 1'b0 ;
  assign n43981 = n31495 ^ n9101 ^ 1'b0 ;
  assign n43982 = n2340 | n5847 ;
  assign n43983 = n43981 & ~n43982 ;
  assign n43984 = n7645 & n9557 ;
  assign n43985 = ~n11818 & n43984 ;
  assign n43986 = n10744 ^ n4498 ^ 1'b0 ;
  assign n43987 = n24812 & n43986 ;
  assign n43988 = n19356 ^ n5376 ^ 1'b0 ;
  assign n43989 = ~n23963 & n43988 ;
  assign n43990 = ( n41083 & n41618 ) | ( n41083 & n43989 ) | ( n41618 & n43989 ) ;
  assign n43991 = ~n24883 & n30898 ;
  assign n43992 = n43991 ^ n39277 ^ 1'b0 ;
  assign n43993 = n22961 ^ n9670 ^ 1'b0 ;
  assign n43994 = n2225 | n11760 ;
  assign n43995 = n43994 ^ n15013 ^ 1'b0 ;
  assign n43996 = n12933 | n22026 ;
  assign n43997 = n43996 ^ n40150 ^ 1'b0 ;
  assign n43998 = ~n23443 & n43997 ;
  assign n44000 = ( n5241 & n14415 ) | ( n5241 & ~n19256 ) | ( n14415 & ~n19256 ) ;
  assign n43999 = n1078 & n34087 ;
  assign n44001 = n44000 ^ n43999 ^ 1'b0 ;
  assign n44002 = n33213 & n39592 ;
  assign n44003 = n44001 & n44002 ;
  assign n44004 = n32158 ^ n21918 ^ n8882 ;
  assign n44005 = n35734 ^ n17304 ^ 1'b0 ;
  assign n44006 = n41515 ^ n13804 ^ 1'b0 ;
  assign n44007 = n30389 ^ n17190 ^ 1'b0 ;
  assign n44008 = n2460 & ~n21770 ;
  assign n44009 = n13706 ^ n11671 ^ 1'b0 ;
  assign n44010 = ~n8700 & n44009 ;
  assign n44011 = n43435 ^ n39351 ^ 1'b0 ;
  assign n44012 = n4710 | n44011 ;
  assign n44013 = n31459 ^ n14674 ^ 1'b0 ;
  assign n44014 = n24665 ^ n21637 ^ n1276 ;
  assign n44015 = ~n44013 & n44014 ;
  assign n44016 = n44015 ^ n850 ^ 1'b0 ;
  assign n44017 = n5418 & n6909 ;
  assign n44018 = n16816 & n44017 ;
  assign n44019 = n13489 & n34617 ;
  assign n44020 = ~n700 & n29210 ;
  assign n44021 = n44019 | n44020 ;
  assign n44022 = n18694 & n19344 ;
  assign n44023 = n15956 ^ n6051 ^ 1'b0 ;
  assign n44024 = ~n19065 & n44023 ;
  assign n44025 = ~n10919 & n31229 ;
  assign n44026 = n26451 ^ n8753 ^ 1'b0 ;
  assign n44027 = ~n44025 & n44026 ;
  assign n44028 = n26400 ^ n12869 ^ 1'b0 ;
  assign n44029 = ~n31515 & n44028 ;
  assign n44030 = n44029 ^ n16835 ^ 1'b0 ;
  assign n44031 = n4675 & ~n6189 ;
  assign n44033 = n39259 ^ n24825 ^ 1'b0 ;
  assign n44032 = n15991 | n39259 ;
  assign n44034 = n44033 ^ n44032 ^ 1'b0 ;
  assign n44035 = n44034 ^ n13031 ^ 1'b0 ;
  assign n44036 = n1926 | n10391 ;
  assign n44037 = n33585 | n44036 ;
  assign n44038 = n22282 | n29558 ;
  assign n44039 = n12058 ^ n4173 ^ 1'b0 ;
  assign n44040 = n37897 | n44039 ;
  assign n44041 = ~n8888 & n9086 ;
  assign n44043 = n1149 & n4064 ;
  assign n44044 = n44043 ^ n12712 ^ 1'b0 ;
  assign n44045 = ( n5073 & n19898 ) | ( n5073 & ~n44044 ) | ( n19898 & ~n44044 ) ;
  assign n44046 = n44045 ^ n5744 ^ 1'b0 ;
  assign n44047 = ~n624 & n3864 ;
  assign n44048 = n496 | n44047 ;
  assign n44049 = ~n11610 & n44048 ;
  assign n44050 = ~n44046 & n44049 ;
  assign n44042 = ~n29429 & n42237 ;
  assign n44051 = n44050 ^ n44042 ^ 1'b0 ;
  assign n44052 = n10196 & ~n25543 ;
  assign n44053 = n6196 & ~n16787 ;
  assign n44054 = n34291 ^ n27888 ^ n3663 ;
  assign n44055 = n41818 ^ n20508 ^ 1'b0 ;
  assign n44056 = n3464 | n13325 ;
  assign n44057 = n8398 | n10321 ;
  assign n44058 = n1153 & ~n44057 ;
  assign n44059 = n5092 & n44058 ;
  assign n44060 = n1602 | n2769 ;
  assign n44061 = n38660 & ~n44060 ;
  assign n44062 = n21393 ^ n18560 ^ 1'b0 ;
  assign n44063 = n44062 ^ n10543 ^ 1'b0 ;
  assign n44064 = ~n44061 & n44063 ;
  assign n44065 = n11546 | n23861 ;
  assign n44066 = n44065 ^ n21381 ^ 1'b0 ;
  assign n44067 = n5785 ^ n978 ^ 1'b0 ;
  assign n44068 = n8489 & n34399 ;
  assign n44069 = n44068 ^ n15870 ^ 1'b0 ;
  assign n44070 = n44067 | n44069 ;
  assign n44071 = n44070 ^ n15535 ^ 1'b0 ;
  assign n44072 = n16316 ^ n2169 ^ 1'b0 ;
  assign n44073 = n37130 & n44072 ;
  assign n44075 = n10851 & n22458 ;
  assign n44076 = n44075 ^ n26360 ^ n10436 ;
  assign n44074 = n15183 & ~n31157 ;
  assign n44077 = n44076 ^ n44074 ^ 1'b0 ;
  assign n44078 = n44077 ^ n23731 ^ n3256 ;
  assign n44079 = n26576 ^ n9131 ^ 1'b0 ;
  assign n44080 = n12235 ^ n8143 ^ n1269 ;
  assign n44081 = n626 & ~n16170 ;
  assign n44082 = n8205 & n44081 ;
  assign n44083 = n26404 & n32573 ;
  assign n44084 = n44082 & n44083 ;
  assign n44085 = n44084 ^ n7782 ^ 1'b0 ;
  assign n44086 = ( n35097 & ~n44080 ) | ( n35097 & n44085 ) | ( ~n44080 & n44085 ) ;
  assign n44087 = n17162 ^ n15855 ^ 1'b0 ;
  assign n44088 = n44045 & n44087 ;
  assign n44089 = n35515 ^ n12955 ^ 1'b0 ;
  assign n44090 = n44088 & ~n44089 ;
  assign n44091 = n7727 & ~n14854 ;
  assign n44092 = n44091 ^ n12420 ^ 1'b0 ;
  assign n44093 = n2726 | n21965 ;
  assign n44094 = n34847 ^ n14471 ^ 1'b0 ;
  assign n44095 = n44093 & ~n44094 ;
  assign n44096 = ~n44092 & n44095 ;
  assign n44097 = ~n1793 & n10632 ;
  assign n44098 = n21060 ^ n6167 ^ 1'b0 ;
  assign n44099 = n44098 ^ n39309 ^ n27846 ;
  assign n44100 = n254 | n4567 ;
  assign n44101 = ~n9713 & n44100 ;
  assign n44102 = n13391 & ~n17174 ;
  assign n44103 = ( n13421 & n33115 ) | ( n13421 & ~n44102 ) | ( n33115 & ~n44102 ) ;
  assign n44104 = n17438 | n44103 ;
  assign n44105 = n44104 ^ n15420 ^ 1'b0 ;
  assign n44106 = n7397 & n29217 ;
  assign n44107 = n20711 & n37311 ;
  assign n44108 = n25775 & n44107 ;
  assign n44109 = ~n9789 & n10648 ;
  assign n44110 = n44109 ^ n19005 ^ 1'b0 ;
  assign n44113 = ( n126 & n20600 ) | ( n126 & ~n34881 ) | ( n20600 & ~n34881 ) ;
  assign n44111 = n12163 & n24835 ;
  assign n44112 = n44111 ^ n34351 ^ n23376 ;
  assign n44114 = n44113 ^ n44112 ^ 1'b0 ;
  assign n44116 = n31769 ^ n8751 ^ 1'b0 ;
  assign n44117 = ~n14881 & n44116 ;
  assign n44115 = n10498 & n19145 ;
  assign n44118 = n44117 ^ n44115 ^ 1'b0 ;
  assign n44119 = n10824 & ~n44118 ;
  assign n44120 = ~n2581 & n44119 ;
  assign n44121 = n44120 ^ n31460 ^ n20974 ;
  assign n44122 = n27816 ^ n8551 ^ 1'b0 ;
  assign n44123 = n5090 & ~n44122 ;
  assign n44124 = ~n7739 & n9043 ;
  assign n44125 = n44124 ^ n34690 ^ 1'b0 ;
  assign n44126 = n25131 ^ n7003 ^ 1'b0 ;
  assign n44127 = n3656 & n9481 ;
  assign n44128 = n44127 ^ n5464 ^ n3439 ;
  assign n44129 = n1926 & n44128 ;
  assign n44130 = n33112 ^ n13673 ^ 1'b0 ;
  assign n44131 = ~n22834 & n44130 ;
  assign n44132 = ~n11190 & n20453 ;
  assign n44133 = n20856 ^ n9186 ^ n7652 ;
  assign n44134 = n2835 | n44133 ;
  assign n44135 = n9514 & ~n44134 ;
  assign n44136 = n44135 ^ n38875 ^ n22472 ;
  assign n44137 = n25992 ^ n5626 ^ 1'b0 ;
  assign n44138 = n31524 & ~n44137 ;
  assign n44139 = n44138 ^ n21832 ^ 1'b0 ;
  assign n44140 = n18382 ^ n6330 ^ 1'b0 ;
  assign n44141 = ~n6462 & n32353 ;
  assign n44142 = n24978 ^ n1186 ^ 1'b0 ;
  assign n44143 = ( n7614 & ~n13678 ) | ( n7614 & n37393 ) | ( ~n13678 & n37393 ) ;
  assign n44144 = n43478 ^ n7672 ^ 1'b0 ;
  assign n44145 = ~n6227 & n44144 ;
  assign n44146 = n44145 ^ n28620 ^ 1'b0 ;
  assign n44147 = n44143 & n44146 ;
  assign n44148 = n29358 ^ n14423 ^ n45 ;
  assign n44149 = n44148 ^ n38151 ^ n37110 ;
  assign n44150 = n44149 ^ n30765 ^ 1'b0 ;
  assign n44151 = n5874 | n30188 ;
  assign n44152 = n44151 ^ n28204 ^ 1'b0 ;
  assign n44153 = n1091 & n3685 ;
  assign n44154 = n44153 ^ n9765 ^ 1'b0 ;
  assign n44155 = ( n4034 & ~n4343 ) | ( n4034 & n44154 ) | ( ~n4343 & n44154 ) ;
  assign n44156 = n20356 & ~n44155 ;
  assign n44157 = n44156 ^ n16776 ^ 1'b0 ;
  assign n44158 = n14213 ^ n1109 ^ 1'b0 ;
  assign n44159 = ~n14711 & n44158 ;
  assign n44160 = ~n4403 & n25050 ;
  assign n44161 = n44160 ^ n14678 ^ 1'b0 ;
  assign n44162 = n13402 ^ n8517 ^ 1'b0 ;
  assign n44163 = ~n9110 & n44162 ;
  assign n44164 = n11700 & n44163 ;
  assign n44165 = ~n14135 & n44164 ;
  assign n44166 = n44165 ^ n1143 ^ 1'b0 ;
  assign n44167 = n1151 & n13263 ;
  assign n44168 = n12867 | n41655 ;
  assign n44169 = ~n5273 & n7096 ;
  assign n44170 = ~n15972 & n44169 ;
  assign n44171 = n44170 ^ n7383 ^ 1'b0 ;
  assign n44172 = n11088 | n14567 ;
  assign n44173 = n14168 & ~n44172 ;
  assign n44174 = n6945 ^ n5757 ^ 1'b0 ;
  assign n44175 = n9753 & n44174 ;
  assign n44176 = ~n20285 & n44175 ;
  assign n44177 = n44176 ^ n5908 ^ 1'b0 ;
  assign n44178 = n32565 ^ n30405 ^ n19875 ;
  assign n44179 = n44178 ^ n30564 ^ 1'b0 ;
  assign n44180 = n44177 | n44179 ;
  assign n44181 = n542 | n44180 ;
  assign n44182 = n24926 ^ n2759 ^ 1'b0 ;
  assign n44183 = n33057 ^ n9164 ^ 1'b0 ;
  assign n44184 = n5458 | n44183 ;
  assign n44185 = ~n5822 & n10814 ;
  assign n44186 = n44185 ^ n41327 ^ 1'b0 ;
  assign n44187 = n11326 | n26514 ;
  assign n44188 = n1302 & ~n1771 ;
  assign n44189 = n44188 ^ n20314 ^ n6076 ;
  assign n44190 = n8195 & n44189 ;
  assign n44191 = ~n23837 & n44190 ;
  assign n44193 = n11247 | n14110 ;
  assign n44194 = n44193 ^ n3027 ^ 1'b0 ;
  assign n44192 = n2138 | n23856 ;
  assign n44195 = n44194 ^ n44192 ^ 1'b0 ;
  assign n44196 = n5329 | n38373 ;
  assign n44197 = n9811 ^ n9750 ^ 1'b0 ;
  assign n44198 = n17459 | n44197 ;
  assign n44199 = n9658 | n10223 ;
  assign n44200 = n5009 | n44199 ;
  assign n44201 = n44198 & ~n44200 ;
  assign n44202 = n14978 ^ n281 ^ 1'b0 ;
  assign n44203 = n39307 ^ n7039 ^ 1'b0 ;
  assign n44204 = n5236 | n44203 ;
  assign n44205 = ( n11071 & n16481 ) | ( n11071 & n44204 ) | ( n16481 & n44204 ) ;
  assign n44206 = n44205 ^ n4977 ^ n4383 ;
  assign n44207 = ( n1188 & n8048 ) | ( n1188 & ~n13923 ) | ( n8048 & ~n13923 ) ;
  assign n44208 = n3387 & ~n7610 ;
  assign n44209 = n44208 ^ n4147 ^ 1'b0 ;
  assign n44210 = n30575 | n32545 ;
  assign n44211 = ~n28024 & n28499 ;
  assign n44212 = n30531 | n31976 ;
  assign n44213 = n41344 & ~n44212 ;
  assign n44214 = n30989 ^ n10313 ^ 1'b0 ;
  assign n44215 = n24743 & n44214 ;
  assign n44216 = n44215 ^ n2561 ^ 1'b0 ;
  assign n44217 = n6135 & n35585 ;
  assign n44218 = n44217 ^ n43931 ^ n22087 ;
  assign n44219 = n7260 ^ n5447 ^ 1'b0 ;
  assign n44220 = ~n5044 & n44219 ;
  assign n44221 = n10739 ^ n9483 ^ 1'b0 ;
  assign n44222 = n29527 ^ n13201 ^ 1'b0 ;
  assign n44223 = n36412 ^ n31334 ^ n16625 ;
  assign n44224 = ( n21054 & ~n32495 ) | ( n21054 & n41255 ) | ( ~n32495 & n41255 ) ;
  assign n44225 = n10503 ^ n6666 ^ 1'b0 ;
  assign n44228 = n9912 | n36935 ;
  assign n44229 = n44228 ^ n30847 ^ 1'b0 ;
  assign n44226 = n25048 ^ n13331 ^ 1'b0 ;
  assign n44227 = ~n8446 & n44226 ;
  assign n44230 = n44229 ^ n44227 ^ 1'b0 ;
  assign n44231 = n3823 & n32378 ;
  assign n44232 = n15274 & n44231 ;
  assign n44233 = n18741 ^ n9222 ^ 1'b0 ;
  assign n44234 = n13068 ^ n9863 ^ n6568 ;
  assign n44235 = n44233 | n44234 ;
  assign n44236 = ( n8456 & n29022 ) | ( n8456 & ~n42972 ) | ( n29022 & ~n42972 ) ;
  assign n44237 = n17064 & ~n34765 ;
  assign n44238 = n44237 ^ n26091 ^ 1'b0 ;
  assign n44239 = ~n7054 & n44238 ;
  assign n44240 = n836 & ~n27755 ;
  assign n44241 = n9476 & n44240 ;
  assign n44242 = n38390 ^ n24396 ^ 1'b0 ;
  assign n44243 = n25429 & ~n44242 ;
  assign n44244 = ~n1818 & n2234 ;
  assign n44245 = ~n7572 & n44244 ;
  assign n44246 = n9315 ^ n478 ^ 1'b0 ;
  assign n44247 = ( ~n7481 & n9462 ) | ( ~n7481 & n21031 ) | ( n9462 & n21031 ) ;
  assign n44248 = n9103 & ~n44247 ;
  assign n44249 = n44248 ^ n36337 ^ 1'b0 ;
  assign n44250 = n28078 & n40001 ;
  assign n44251 = ~n5050 & n36876 ;
  assign n44252 = n44251 ^ n14597 ^ 1'b0 ;
  assign n44253 = n2841 & ~n44252 ;
  assign n44254 = ~n23554 & n24952 ;
  assign n44255 = ~n23312 & n44254 ;
  assign n44256 = n22367 | n26533 ;
  assign n44257 = n32995 & n44133 ;
  assign n44258 = n44257 ^ n17003 ^ 1'b0 ;
  assign n44260 = n2750 | n3989 ;
  assign n44259 = n31501 ^ n4708 ^ 1'b0 ;
  assign n44261 = n44260 ^ n44259 ^ n40009 ;
  assign n44262 = n1182 & ~n1527 ;
  assign n44263 = n44262 ^ n39067 ^ 1'b0 ;
  assign n44264 = n29685 ^ n18508 ^ 1'b0 ;
  assign n44265 = n11744 ^ n4417 ^ n3128 ;
  assign n44266 = n13116 & n44265 ;
  assign n44267 = ~n181 & n23531 ;
  assign n44269 = n35198 & ~n35983 ;
  assign n44268 = n25877 | n30765 ;
  assign n44270 = n44269 ^ n44268 ^ 1'b0 ;
  assign n44271 = n28796 ^ n6634 ^ 1'b0 ;
  assign n44272 = n3508 & n44271 ;
  assign n44273 = n3191 & n28524 ;
  assign n44274 = n9667 & n44273 ;
  assign n44275 = n10772 & ~n44274 ;
  assign n44276 = n24118 | n44275 ;
  assign n44277 = n25652 & n36413 ;
  assign n44278 = n44277 ^ n6152 ^ 1'b0 ;
  assign n44279 = n44276 & ~n44278 ;
  assign n44280 = n4545 & ~n34143 ;
  assign n44281 = n44280 ^ n2114 ^ 1'b0 ;
  assign n44282 = n15029 ^ n8899 ^ n7939 ;
  assign n44283 = n44281 & ~n44282 ;
  assign n44284 = n32170 & n44283 ;
  assign n44285 = ( n23723 & ~n44279 ) | ( n23723 & n44284 ) | ( ~n44279 & n44284 ) ;
  assign n44286 = n10472 | n19564 ;
  assign n44287 = ~n11115 & n44286 ;
  assign n44288 = n44287 ^ n12091 ^ 1'b0 ;
  assign n44289 = ( n17401 & n27483 ) | ( n17401 & n44288 ) | ( n27483 & n44288 ) ;
  assign n44290 = ~n5513 & n17010 ;
  assign n44291 = n31106 ^ n15382 ^ n164 ;
  assign n44293 = n26152 ^ n2403 ^ 1'b0 ;
  assign n44294 = n37492 & n44293 ;
  assign n44292 = n6319 | n12987 ;
  assign n44295 = n44294 ^ n44292 ^ 1'b0 ;
  assign n44296 = n19164 ^ n11472 ^ n4331 ;
  assign n44297 = ~n25898 & n44296 ;
  assign n44298 = n42319 ^ n16948 ^ 1'b0 ;
  assign n44299 = n44297 & n44298 ;
  assign n44300 = n10187 & ~n12578 ;
  assign n44301 = n28609 ^ n24891 ^ 1'b0 ;
  assign n44302 = n21425 ^ n7935 ^ 1'b0 ;
  assign n44303 = n816 & ~n44302 ;
  assign n44304 = n22436 & ~n42726 ;
  assign n44305 = ~n22702 & n44304 ;
  assign n44306 = n36017 ^ n12050 ^ n9054 ;
  assign n44307 = ( n5001 & ~n9910 ) | ( n5001 & n44306 ) | ( ~n9910 & n44306 ) ;
  assign n44308 = ~n10391 & n40237 ;
  assign n44309 = ~n24319 & n44308 ;
  assign n44310 = n40586 | n44309 ;
  assign n44311 = n14495 ^ n691 ^ n42 ;
  assign n44312 = n44311 ^ n19175 ^ 1'b0 ;
  assign n44313 = n554 & n44312 ;
  assign n44314 = ~n18998 & n44313 ;
  assign n44315 = n26404 ^ n1026 ^ 1'b0 ;
  assign n44316 = n32195 & n44315 ;
  assign n44317 = ~n2695 & n35069 ;
  assign n44318 = ~n12174 & n25251 ;
  assign n44319 = ~n41311 & n44318 ;
  assign n44320 = n44319 ^ n13094 ^ 1'b0 ;
  assign n44321 = n44317 & n44320 ;
  assign n44322 = n29914 ^ n16887 ^ 1'b0 ;
  assign n44323 = n43233 ^ n411 ^ 1'b0 ;
  assign n44324 = n197 & n23804 ;
  assign n44325 = n615 & ~n7087 ;
  assign n44326 = n44325 ^ n14415 ^ 1'b0 ;
  assign n44327 = ~n17296 & n17440 ;
  assign n44328 = n44326 & n44327 ;
  assign n44329 = n44328 ^ n2784 ^ 1'b0 ;
  assign n44330 = n44324 | n44329 ;
  assign n44331 = n4784 | n31058 ;
  assign n44332 = n11152 ^ n10420 ^ 1'b0 ;
  assign n44333 = n25095 ^ n5616 ^ 1'b0 ;
  assign n44334 = n6185 & n11409 ;
  assign n44335 = n44333 & ~n44334 ;
  assign n44336 = n25596 ^ n17351 ^ 1'b0 ;
  assign n44337 = n31401 & n44336 ;
  assign n44338 = ~n10492 & n44337 ;
  assign n44339 = n44338 ^ n3134 ^ 1'b0 ;
  assign n44340 = n1368 & ~n3225 ;
  assign n44341 = n10551 & n44340 ;
  assign n44342 = n24715 & n44341 ;
  assign n44343 = ~n12626 & n44342 ;
  assign n44344 = ~n10950 & n18652 ;
  assign n44345 = n44344 ^ n5459 ^ 1'b0 ;
  assign n44346 = n1616 & n9772 ;
  assign n44347 = n25413 ^ n22996 ^ 1'b0 ;
  assign n44348 = n44346 & n44347 ;
  assign n44349 = ( n30858 & n44133 ) | ( n30858 & ~n44348 ) | ( n44133 & ~n44348 ) ;
  assign n44350 = ~n401 & n12445 ;
  assign n44351 = n15461 & n44350 ;
  assign n44352 = n6756 ^ n2216 ^ 1'b0 ;
  assign n44353 = n37256 & n44352 ;
  assign n44354 = n27998 ^ n5914 ^ 1'b0 ;
  assign n44355 = n11846 & n44354 ;
  assign n44356 = ~n44353 & n44355 ;
  assign n44357 = ~n11231 & n13455 ;
  assign n44358 = n4024 & n20962 ;
  assign n44359 = n44358 ^ n39322 ^ 1'b0 ;
  assign n44360 = n44357 & n44359 ;
  assign n44362 = n5780 & n11120 ;
  assign n44363 = n44362 ^ n12126 ^ n7409 ;
  assign n44361 = n28761 ^ n1609 ^ 1'b0 ;
  assign n44364 = n44363 ^ n44361 ^ 1'b0 ;
  assign n44365 = n44364 ^ n43347 ^ 1'b0 ;
  assign n44366 = n9111 ^ n5372 ^ n4159 ;
  assign n44367 = n23656 | n39313 ;
  assign n44368 = n9527 | n44367 ;
  assign n44369 = n44368 ^ n35325 ^ 1'b0 ;
  assign n44370 = n44369 ^ n20158 ^ 1'b0 ;
  assign n44371 = n2206 & ~n44370 ;
  assign n44372 = ~n44366 & n44371 ;
  assign n44373 = ~n17552 & n42140 ;
  assign n44374 = n44373 ^ n43519 ^ 1'b0 ;
  assign n44375 = n15367 ^ n11408 ^ n6284 ;
  assign n44376 = n11355 ^ n8016 ^ 1'b0 ;
  assign n44377 = ~n44375 & n44376 ;
  assign n44378 = n2733 ^ n1093 ^ 1'b0 ;
  assign n44379 = n10631 & n44378 ;
  assign n44380 = ~n44377 & n44379 ;
  assign n44381 = n42201 & n44380 ;
  assign n44382 = n14211 ^ n6275 ^ 1'b0 ;
  assign n44383 = n16488 | n44382 ;
  assign n44384 = n16601 & n21862 ;
  assign n44385 = n36258 | n44384 ;
  assign n44386 = n44385 ^ n7344 ^ 1'b0 ;
  assign n44390 = n14129 ^ n12483 ^ 1'b0 ;
  assign n44388 = n4578 | n5891 ;
  assign n44389 = n12330 | n44388 ;
  assign n44391 = n44390 ^ n44389 ^ 1'b0 ;
  assign n44387 = n1943 & n29450 ;
  assign n44392 = n44391 ^ n44387 ^ 1'b0 ;
  assign n44393 = n4400 & n31384 ;
  assign n44394 = n44392 & n44393 ;
  assign n44395 = n44394 ^ n13821 ^ 1'b0 ;
  assign n44396 = n8056 & ~n44395 ;
  assign n44397 = n6091 & n10534 ;
  assign n44398 = ~n13609 & n44397 ;
  assign n44399 = ~n9832 & n14786 ;
  assign n44400 = ~n1807 & n44399 ;
  assign n44401 = n44400 ^ n28763 ^ 1'b0 ;
  assign n44402 = n36966 & ~n44401 ;
  assign n44403 = ~n16865 & n23483 ;
  assign n44404 = n44403 ^ n39526 ^ 1'b0 ;
  assign n44405 = ( ~n7054 & n7911 ) | ( ~n7054 & n16828 ) | ( n7911 & n16828 ) ;
  assign n44406 = ( n30818 & ~n39826 ) | ( n30818 & n44405 ) | ( ~n39826 & n44405 ) ;
  assign n44407 = n35109 ^ n7494 ^ 1'b0 ;
  assign n44408 = n11911 & ~n44407 ;
  assign n44409 = ( n8402 & n35927 ) | ( n8402 & n44408 ) | ( n35927 & n44408 ) ;
  assign n44411 = n13764 ^ n5415 ^ 1'b0 ;
  assign n44412 = n13463 & ~n44411 ;
  assign n44410 = ~n645 & n11924 ;
  assign n44413 = n44412 ^ n44410 ^ 1'b0 ;
  assign n44414 = n34066 | n44413 ;
  assign n44419 = ~n1015 & n7543 ;
  assign n44415 = n22532 ^ n18547 ^ n5751 ;
  assign n44416 = n27283 & n35390 ;
  assign n44417 = ~n44415 & n44416 ;
  assign n44418 = ( ~n570 & n34599 ) | ( ~n570 & n44417 ) | ( n34599 & n44417 ) ;
  assign n44420 = n44419 ^ n44418 ^ 1'b0 ;
  assign n44421 = n21564 & ~n22189 ;
  assign n44422 = ~n5825 & n44421 ;
  assign n44423 = n3691 | n6289 ;
  assign n44424 = n44423 ^ n498 ^ 1'b0 ;
  assign n44425 = ~n44422 & n44424 ;
  assign n44426 = n5315 ^ n704 ^ 1'b0 ;
  assign n44427 = n1874 & ~n44426 ;
  assign n44428 = n14211 | n44427 ;
  assign n44429 = ~n28206 & n28500 ;
  assign n44430 = n1690 & n44429 ;
  assign n44431 = ~n28481 & n44430 ;
  assign n44432 = n33632 ^ n9446 ^ 1'b0 ;
  assign n44433 = n38890 ^ n7040 ^ 1'b0 ;
  assign n44434 = n28926 & n44433 ;
  assign n44435 = n44434 ^ n6322 ^ 1'b0 ;
  assign n44436 = n16414 ^ n9666 ^ 1'b0 ;
  assign n44437 = n18145 & n44436 ;
  assign n44438 = n601 & ~n40581 ;
  assign n44439 = n21181 ^ n12785 ^ 1'b0 ;
  assign n44440 = ~n44438 & n44439 ;
  assign n44441 = n28046 ^ n21260 ^ 1'b0 ;
  assign n44442 = n22786 | n44441 ;
  assign n44443 = ( n9043 & ~n30208 ) | ( n9043 & n41261 ) | ( ~n30208 & n41261 ) ;
  assign n44444 = n44443 ^ n237 ^ 1'b0 ;
  assign n44445 = n8857 | n29991 ;
  assign n44446 = n16500 & ~n44445 ;
  assign n44447 = n761 | n13488 ;
  assign n44448 = n44447 ^ n27673 ^ 1'b0 ;
  assign n44449 = n44448 ^ n38703 ^ 1'b0 ;
  assign n44450 = ( n26569 & n44446 ) | ( n26569 & n44449 ) | ( n44446 & n44449 ) ;
  assign n44451 = n13800 & ~n36926 ;
  assign n44452 = n26642 & n44451 ;
  assign n44453 = ~n12275 & n35892 ;
  assign n44454 = n44453 ^ n44046 ^ 1'b0 ;
  assign n44455 = ~n20034 & n44454 ;
  assign n44456 = n37929 ^ n32117 ^ 1'b0 ;
  assign n44457 = n10839 | n44456 ;
  assign n44458 = n44457 ^ n76 ^ 1'b0 ;
  assign n44459 = n28118 ^ n18766 ^ 1'b0 ;
  assign n44460 = n24372 | n44459 ;
  assign n44461 = n32202 & ~n44460 ;
  assign n44462 = n44461 ^ n31351 ^ n9517 ;
  assign n44463 = ~n4713 & n12111 ;
  assign n44464 = n27979 | n39548 ;
  assign n44465 = n44041 ^ n40742 ^ 1'b0 ;
  assign n44466 = n18432 & ~n44465 ;
  assign n44467 = ( n65 & n4018 ) | ( n65 & n12440 ) | ( n4018 & n12440 ) ;
  assign n44468 = n25504 ^ n18024 ^ n12347 ;
  assign n44470 = n4092 & n5804 ;
  assign n44471 = n28876 & n44470 ;
  assign n44469 = ~n19324 & n33652 ;
  assign n44472 = n44471 ^ n44469 ^ 1'b0 ;
  assign n44473 = n41055 ^ n2082 ^ 1'b0 ;
  assign n44474 = n24748 ^ n24314 ^ n7927 ;
  assign n44475 = n16193 | n44474 ;
  assign n44476 = n6849 | n15987 ;
  assign n44477 = n5284 | n44476 ;
  assign n44478 = n2982 | n15512 ;
  assign n44479 = n34764 | n44478 ;
  assign n44480 = n34166 ^ n16965 ^ 1'b0 ;
  assign n44481 = n44479 & n44480 ;
  assign n44482 = ~n684 & n10867 ;
  assign n44483 = n26247 ^ n15379 ^ 1'b0 ;
  assign n44484 = n25559 | n44483 ;
  assign n44485 = n44482 & n44484 ;
  assign n44486 = n91 & ~n111 ;
  assign n44487 = ~n91 & n44486 ;
  assign n44488 = n44487 ^ n887 ^ 1'b0 ;
  assign n44489 = ~n2704 & n7489 ;
  assign n44490 = n2704 & n44489 ;
  assign n44492 = ~n22525 & n23766 ;
  assign n44493 = n22525 & n44492 ;
  assign n44491 = n16743 | n21723 ;
  assign n44494 = n44493 ^ n44491 ^ 1'b0 ;
  assign n44495 = ( n10103 & n44490 ) | ( n10103 & n44494 ) | ( n44490 & n44494 ) ;
  assign n44496 = ( ~n21996 & n44488 ) | ( ~n21996 & n44495 ) | ( n44488 & n44495 ) ;
  assign n44498 = ~n2192 & n26723 ;
  assign n44499 = n16694 & n44498 ;
  assign n44497 = ~n8306 & n18570 ;
  assign n44500 = n44499 ^ n44497 ^ n24703 ;
  assign n44501 = n11491 & n31180 ;
  assign n44502 = n27076 ^ n20827 ^ n10876 ;
  assign n44503 = n44502 ^ n27791 ^ 1'b0 ;
  assign n44504 = n4901 & ~n44503 ;
  assign n44505 = n9371 | n22507 ;
  assign n44506 = n35032 | n44505 ;
  assign n44507 = n17602 | n35796 ;
  assign n44508 = n44507 ^ n4004 ^ 1'b0 ;
  assign n44509 = n122 & n33337 ;
  assign n44510 = n44509 ^ n32914 ^ n16799 ;
  assign n44511 = ~n8243 & n17222 ;
  assign n44512 = ~n16650 & n19199 ;
  assign n44513 = ~n649 & n44512 ;
  assign n44514 = ~n29492 & n43356 ;
  assign n44515 = n44514 ^ n7738 ^ 1'b0 ;
  assign n44516 = ~n10541 & n11893 ;
  assign n44517 = n25698 & ~n30887 ;
  assign n44518 = n44517 ^ n8297 ^ n2581 ;
  assign n44519 = ( ~n3898 & n5324 ) | ( ~n3898 & n18709 ) | ( n5324 & n18709 ) ;
  assign n44523 = n15356 ^ n14772 ^ n11443 ;
  assign n44524 = n2129 & ~n38402 ;
  assign n44525 = n44523 & n44524 ;
  assign n44520 = n13377 & ~n25612 ;
  assign n44521 = n10079 & n44520 ;
  assign n44522 = ~n3575 & n44521 ;
  assign n44526 = n44525 ^ n44522 ^ 1'b0 ;
  assign n44527 = n14083 & ~n41190 ;
  assign n44528 = n44527 ^ n22760 ^ 1'b0 ;
  assign n44529 = n6976 & ~n21842 ;
  assign n44530 = n44529 ^ n8919 ^ 1'b0 ;
  assign n44531 = n26088 ^ n11638 ^ n3557 ;
  assign n44532 = n44531 ^ n31822 ^ 1'b0 ;
  assign n44533 = n26231 & ~n44148 ;
  assign n44534 = n44533 ^ n5408 ^ 1'b0 ;
  assign n44535 = ~n14799 & n44534 ;
  assign n44536 = n22134 & ~n42364 ;
  assign n44537 = n10548 | n21686 ;
  assign n44538 = n23027 ^ n11547 ^ n6524 ;
  assign n44539 = n19805 ^ n17844 ^ 1'b0 ;
  assign n44540 = ( n37239 & n43084 ) | ( n37239 & ~n44400 ) | ( n43084 & ~n44400 ) ;
  assign n44541 = n6365 & n41919 ;
  assign n44542 = n39695 ^ n31471 ^ 1'b0 ;
  assign n44543 = ~n44324 & n44542 ;
  assign n44544 = n29840 & n37521 ;
  assign n44545 = n20856 & n26984 ;
  assign n44546 = ( n30538 & n36005 ) | ( n30538 & ~n44545 ) | ( n36005 & ~n44545 ) ;
  assign n44547 = n12619 ^ n7771 ^ 1'b0 ;
  assign n44548 = n8176 & ~n29068 ;
  assign n44549 = n11946 & n44548 ;
  assign n44550 = ~n15802 & n25924 ;
  assign n44551 = n18818 | n25290 ;
  assign n44552 = n44551 ^ n30834 ^ 1'b0 ;
  assign n44553 = ~n5946 & n34983 ;
  assign n44554 = n12541 & ~n15953 ;
  assign n44555 = n41 | n6771 ;
  assign n44556 = n4502 | n44555 ;
  assign n44557 = n37399 ^ n7054 ^ 1'b0 ;
  assign n44558 = n1474 | n31623 ;
  assign n44559 = n14342 | n34363 ;
  assign n44560 = n30727 | n44559 ;
  assign n44561 = n35789 ^ n4463 ^ n3698 ;
  assign n44562 = n2416 ^ n73 ^ 1'b0 ;
  assign n44563 = n42690 & ~n44562 ;
  assign n44564 = ( ~n4607 & n6668 ) | ( ~n4607 & n44563 ) | ( n6668 & n44563 ) ;
  assign n44565 = n2211 & ~n20652 ;
  assign n44566 = n24036 & n44565 ;
  assign n44567 = n21225 ^ n12219 ^ 1'b0 ;
  assign n44568 = n12307 & ~n44567 ;
  assign n44569 = n14906 ^ n4434 ^ 1'b0 ;
  assign n44570 = n44568 & n44569 ;
  assign n44571 = n7659 & ~n12225 ;
  assign n44572 = ~n4153 & n6027 ;
  assign n44573 = n44572 ^ n44078 ^ 1'b0 ;
  assign n44574 = n15685 & ~n44573 ;
  assign n44575 = ~n9934 & n17237 ;
  assign n44576 = n44575 ^ n7400 ^ 1'b0 ;
  assign n44577 = n9345 ^ n7357 ^ 1'b0 ;
  assign n44578 = ~n2793 & n44577 ;
  assign n44579 = ( n654 & ~n4954 ) | ( n654 & n36446 ) | ( ~n4954 & n36446 ) ;
  assign n44580 = ( n9713 & ~n13314 ) | ( n9713 & n28534 ) | ( ~n13314 & n28534 ) ;
  assign n44581 = ~n18851 & n44580 ;
  assign n44582 = ~n44579 & n44581 ;
  assign n44583 = n10432 ^ n3131 ^ 1'b0 ;
  assign n44584 = n34420 | n44583 ;
  assign n44585 = n19913 | n44584 ;
  assign n44586 = n44585 ^ n25506 ^ 1'b0 ;
  assign n44587 = ~n8084 & n11365 ;
  assign n44588 = ~n4892 & n44587 ;
  assign n44589 = n44588 ^ n30995 ^ n10829 ;
  assign n44590 = n37212 ^ n31933 ^ n18447 ;
  assign n44591 = n3961 ^ n2550 ^ 1'b0 ;
  assign n44592 = n23554 | n30779 ;
  assign n44593 = n44592 ^ n1109 ^ 1'b0 ;
  assign n44594 = n37946 | n44593 ;
  assign n44595 = n44594 ^ n40171 ^ 1'b0 ;
  assign n44596 = n42360 | n44595 ;
  assign n44597 = n57 & n39518 ;
  assign n44598 = n18472 ^ n5537 ^ 1'b0 ;
  assign n44599 = n14887 & ~n21883 ;
  assign n44600 = n44598 & n44599 ;
  assign n44601 = ( ~n902 & n9335 ) | ( ~n902 & n10816 ) | ( n9335 & n10816 ) ;
  assign n44602 = n10892 | n44601 ;
  assign n44603 = n3711 & ~n14174 ;
  assign n44604 = n8413 ^ n30 ^ 1'b0 ;
  assign n44605 = n36093 & ~n44604 ;
  assign n44606 = n2810 ^ n1766 ^ 1'b0 ;
  assign n44607 = n30718 & ~n44606 ;
  assign n44608 = n19482 | n34235 ;
  assign n44609 = n21313 & ~n44608 ;
  assign n44610 = ~n18910 & n44609 ;
  assign n44611 = n44610 ^ n19441 ^ 1'b0 ;
  assign n44612 = n7425 ^ n5612 ^ 1'b0 ;
  assign n44613 = n44612 ^ n25590 ^ 1'b0 ;
  assign n44614 = n13834 & n44613 ;
  assign n44615 = n19097 ^ n7544 ^ 1'b0 ;
  assign n44616 = n17125 ^ n13836 ^ n8959 ;
  assign n44617 = ~n12488 & n40068 ;
  assign n44618 = n28206 & n44617 ;
  assign n44619 = ( n20903 & n44616 ) | ( n20903 & n44618 ) | ( n44616 & n44618 ) ;
  assign n44620 = n19482 ^ n4223 ^ 1'b0 ;
  assign n44621 = n10349 & n44620 ;
  assign n44622 = n44621 ^ n27050 ^ n12539 ;
  assign n44623 = n5029 | n15666 ;
  assign n44624 = n44623 ^ n3445 ^ 1'b0 ;
  assign n44625 = n19269 | n44624 ;
  assign n44626 = n21518 & ~n44625 ;
  assign n44627 = n2546 & ~n14200 ;
  assign n44628 = n22419 ^ n3732 ^ 1'b0 ;
  assign n44629 = ( n5565 & n6257 ) | ( n5565 & ~n11082 ) | ( n6257 & ~n11082 ) ;
  assign n44630 = n33957 & n44629 ;
  assign n44631 = n44628 & n44630 ;
  assign n44632 = n26949 ^ n7279 ^ 1'b0 ;
  assign n44633 = ~n1677 & n4698 ;
  assign n44634 = n13268 & n44633 ;
  assign n44635 = n44634 ^ n2823 ^ 1'b0 ;
  assign n44636 = n24883 | n40925 ;
  assign n44637 = n5312 | n44636 ;
  assign n44638 = n41327 | n44637 ;
  assign n44639 = n34081 ^ n33078 ^ 1'b0 ;
  assign n44640 = n15537 ^ n1249 ^ 1'b0 ;
  assign n44641 = n21543 & n27117 ;
  assign n44642 = n34008 ^ n23240 ^ n11391 ;
  assign n44643 = ~n5175 & n44642 ;
  assign n44644 = n9619 ^ n4674 ^ n235 ;
  assign n44645 = n6403 ^ n3734 ^ 1'b0 ;
  assign n44646 = n44645 ^ n19613 ^ n9902 ;
  assign n44647 = ~n17974 & n44646 ;
  assign n44648 = n44028 ^ n7384 ^ 1'b0 ;
  assign n44649 = ( n12423 & n24537 ) | ( n12423 & n33003 ) | ( n24537 & n33003 ) ;
  assign n44650 = n34491 | n44649 ;
  assign n44651 = ~n5342 & n8002 ;
  assign n44652 = n44651 ^ n648 ^ 1'b0 ;
  assign n44653 = ~n6089 & n17323 ;
  assign n44654 = n44652 & n44653 ;
  assign n44655 = n1088 & ~n13017 ;
  assign n44656 = ~n6705 & n44655 ;
  assign n44657 = n44656 ^ n13081 ^ 1'b0 ;
  assign n44661 = ~n10762 & n22411 ;
  assign n44658 = ~n139 & n18307 ;
  assign n44659 = n21982 & n44658 ;
  assign n44660 = n44659 ^ n29324 ^ n709 ;
  assign n44662 = n44661 ^ n44660 ^ 1'b0 ;
  assign n44663 = n10117 & ~n44662 ;
  assign n44664 = n33480 ^ n3523 ^ 1'b0 ;
  assign n44665 = n44128 & n44664 ;
  assign n44666 = n30942 ^ n15488 ^ 1'b0 ;
  assign n44667 = n28847 & n44666 ;
  assign n44668 = n44667 ^ n14495 ^ 1'b0 ;
  assign n44669 = n34664 & ~n44668 ;
  assign n44670 = n9224 | n23531 ;
  assign n44671 = n15568 & n18648 ;
  assign n44672 = n26400 ^ n22046 ^ n13543 ;
  assign n44673 = n44672 ^ n338 ^ 1'b0 ;
  assign n44674 = n44671 & n44673 ;
  assign n44675 = n4785 & ~n28542 ;
  assign n44676 = n30726 & n33372 ;
  assign n44677 = n23133 & n44676 ;
  assign n44678 = n14570 ^ n7951 ^ n4382 ;
  assign n44679 = n44678 ^ n33265 ^ 1'b0 ;
  assign n44680 = n35961 | n44679 ;
  assign n44681 = n13312 & n43503 ;
  assign n44682 = ~n7868 & n44681 ;
  assign n44683 = n408 | n7890 ;
  assign n44684 = n34720 | n44683 ;
  assign n44685 = n1779 ^ n1515 ^ 1'b0 ;
  assign n44686 = n44685 ^ n32792 ^ 1'b0 ;
  assign n44687 = n44053 ^ n3158 ^ 1'b0 ;
  assign n44689 = n29097 | n32034 ;
  assign n44690 = n2271 | n44689 ;
  assign n44688 = n5108 & ~n5380 ;
  assign n44691 = n44690 ^ n44688 ^ 1'b0 ;
  assign n44692 = ~n2879 & n16755 ;
  assign n44693 = n3202 | n35431 ;
  assign n44694 = n11596 & n44693 ;
  assign n44696 = n16250 ^ n10633 ^ 1'b0 ;
  assign n44697 = n542 & n44696 ;
  assign n44698 = n13987 ^ n12866 ^ 1'b0 ;
  assign n44699 = ~n6003 & n44698 ;
  assign n44700 = n44699 ^ n12556 ^ 1'b0 ;
  assign n44701 = ~n44697 & n44700 ;
  assign n44695 = n13974 | n22151 ;
  assign n44702 = n44701 ^ n44695 ^ 1'b0 ;
  assign n44703 = n25785 ^ n22417 ^ n17669 ;
  assign n44704 = ( n4733 & n8287 ) | ( n4733 & ~n20512 ) | ( n8287 & ~n20512 ) ;
  assign n44705 = n36651 ^ n26082 ^ n2201 ;
  assign n44706 = n44705 ^ n40135 ^ n27449 ;
  assign n44707 = n2760 & n15025 ;
  assign n44708 = n21492 & n44707 ;
  assign n44709 = n2901 & ~n44708 ;
  assign n44710 = ~n6994 & n44709 ;
  assign n44711 = ~n4557 & n38957 ;
  assign n44712 = n44711 ^ n16750 ^ 1'b0 ;
  assign n44713 = n8282 | n8603 ;
  assign n44714 = n30553 & ~n34348 ;
  assign n44715 = n30908 ^ n252 ^ 1'b0 ;
  assign n44716 = n43248 & ~n44715 ;
  assign n44717 = ~n10647 & n44716 ;
  assign n44718 = ~n3902 & n29735 ;
  assign n44719 = ~n11508 & n44718 ;
  assign n44720 = n6725 | n17740 ;
  assign n44721 = ~n7118 & n30516 ;
  assign n44722 = ~n15424 & n27117 ;
  assign n44723 = ( n21543 & ~n27890 ) | ( n21543 & n43989 ) | ( ~n27890 & n43989 ) ;
  assign n44724 = n5118 & n7633 ;
  assign n44725 = n36090 & n44724 ;
  assign n44726 = n16357 & ~n44725 ;
  assign n44727 = ( n8793 & n31240 ) | ( n8793 & n44726 ) | ( n31240 & n44726 ) ;
  assign n44728 = n6384 | n40897 ;
  assign n44729 = n44728 ^ n2209 ^ 1'b0 ;
  assign n44730 = n19022 ^ n650 ^ 1'b0 ;
  assign n44731 = n44730 ^ n29047 ^ n13300 ;
  assign n44732 = n8659 ^ n2261 ^ 1'b0 ;
  assign n44733 = n12133 ^ n2274 ^ 1'b0 ;
  assign n44734 = n9263 & n44733 ;
  assign n44735 = ~n16487 & n44734 ;
  assign n44736 = n44735 ^ n6309 ^ 1'b0 ;
  assign n44737 = ~n9994 & n32198 ;
  assign n44738 = n11349 & n44737 ;
  assign n44739 = ( n6948 & ~n26548 ) | ( n6948 & n27210 ) | ( ~n26548 & n27210 ) ;
  assign n44740 = n713 & ~n4498 ;
  assign n44741 = n11540 ^ n1523 ^ 1'b0 ;
  assign n44742 = n6027 & n44741 ;
  assign n44743 = ( n1425 & ~n32896 ) | ( n1425 & n44742 ) | ( ~n32896 & n44742 ) ;
  assign n44744 = n7464 | n44743 ;
  assign n44745 = n34311 ^ n15173 ^ 1'b0 ;
  assign n44746 = ~n8228 & n44745 ;
  assign n44747 = n6285 & n44746 ;
  assign n44748 = n44747 ^ n17214 ^ 1'b0 ;
  assign n44749 = n44748 ^ n1866 ^ 1'b0 ;
  assign n44750 = n1481 | n5571 ;
  assign n44751 = n44750 ^ n10301 ^ 1'b0 ;
  assign n44752 = n44751 ^ n423 ^ 1'b0 ;
  assign n44753 = n43144 ^ n23373 ^ 1'b0 ;
  assign n44754 = n25509 ^ n5053 ^ 1'b0 ;
  assign n44755 = ~n10861 & n44754 ;
  assign n44756 = n44753 & n44755 ;
  assign n44757 = ~n368 & n2733 ;
  assign n44758 = n44757 ^ n10569 ^ 1'b0 ;
  assign n44759 = ( n11836 & ~n13178 ) | ( n11836 & n44758 ) | ( ~n13178 & n44758 ) ;
  assign n44760 = n16169 & ~n44759 ;
  assign n44761 = n39705 ^ n38527 ^ 1'b0 ;
  assign n44762 = n43398 ^ n11478 ^ 1'b0 ;
  assign n44763 = n5064 & ~n9050 ;
  assign n44764 = n10220 | n17408 ;
  assign n44765 = n32848 & n41487 ;
  assign n44766 = n7532 & n40322 ;
  assign n44767 = n29875 ^ n14489 ^ 1'b0 ;
  assign n44768 = n44767 ^ n34329 ^ n12764 ;
  assign n44769 = n9086 & ~n17724 ;
  assign n44770 = n8043 & n11010 ;
  assign n44771 = n4988 & ~n28763 ;
  assign n44772 = ~n44770 & n44771 ;
  assign n44773 = n44281 ^ n539 ^ 1'b0 ;
  assign n44774 = n31121 ^ n5854 ^ 1'b0 ;
  assign n44775 = n1007 ^ n448 ^ 1'b0 ;
  assign n44776 = n10134 | n44775 ;
  assign n44777 = n7002 & ~n26916 ;
  assign n44778 = n44777 ^ n21794 ^ 1'b0 ;
  assign n44779 = n44778 ^ n38221 ^ n13065 ;
  assign n44780 = n41471 ^ n35252 ^ n7228 ;
  assign n44781 = n44780 ^ n15756 ^ 1'b0 ;
  assign n44782 = n5958 & n38271 ;
  assign n44783 = n44782 ^ n16390 ^ 1'b0 ;
  assign n44784 = ~n30478 & n36688 ;
  assign n44785 = n44784 ^ n35356 ^ 1'b0 ;
  assign n44786 = n36128 ^ n19503 ^ 1'b0 ;
  assign n44790 = ( n6129 & n6886 ) | ( n6129 & ~n13903 ) | ( n6886 & ~n13903 ) ;
  assign n44791 = n33032 | n44790 ;
  assign n44787 = n41072 ^ n3971 ^ 1'b0 ;
  assign n44788 = n36859 | n44787 ;
  assign n44789 = n14098 | n44788 ;
  assign n44792 = n44791 ^ n44789 ^ 1'b0 ;
  assign n44793 = n44309 ^ n13006 ^ 1'b0 ;
  assign n44794 = n5978 & ~n44793 ;
  assign n44795 = ~n4110 & n9132 ;
  assign n44796 = n44795 ^ n8567 ^ 1'b0 ;
  assign n44797 = n44796 ^ n40436 ^ n12773 ;
  assign n44798 = n14953 ^ n7652 ^ 1'b0 ;
  assign n44799 = n8591 & ~n8820 ;
  assign n44800 = n25623 & n44799 ;
  assign n44801 = n14821 & ~n19667 ;
  assign n44802 = n44801 ^ n5713 ^ 1'b0 ;
  assign n44804 = n3192 ^ n826 ^ 1'b0 ;
  assign n44803 = ~n11646 & n26416 ;
  assign n44805 = n44804 ^ n44803 ^ 1'b0 ;
  assign n44806 = ~n20885 & n21489 ;
  assign n44808 = ~n30638 & n36626 ;
  assign n44807 = n3805 & n7358 ;
  assign n44809 = n44808 ^ n44807 ^ 1'b0 ;
  assign n44810 = n14417 & ~n30441 ;
  assign n44811 = ~n3037 & n20601 ;
  assign n44812 = ~n866 & n44811 ;
  assign n44813 = n24702 & ~n44812 ;
  assign n44814 = n44813 ^ n3223 ^ 1'b0 ;
  assign n44815 = n32587 | n44814 ;
  assign n44816 = n43296 ^ n659 ^ 1'b0 ;
  assign n44817 = n35920 ^ n15978 ^ 1'b0 ;
  assign n44818 = ( n14571 & n44701 ) | ( n14571 & ~n44817 ) | ( n44701 & ~n44817 ) ;
  assign n44819 = ~n875 & n1876 ;
  assign n44820 = n44819 ^ n101 ^ 1'b0 ;
  assign n44821 = n44820 ^ n32700 ^ n28373 ;
  assign n44822 = n3073 | n15837 ;
  assign n44823 = n44822 ^ n38170 ^ 1'b0 ;
  assign n44824 = n34091 & n44823 ;
  assign n44825 = n13719 & n36986 ;
  assign n44826 = n10883 & n14323 ;
  assign n44827 = n44826 ^ n7787 ^ 1'b0 ;
  assign n44828 = n41722 & ~n44827 ;
  assign n44829 = ( n28323 & n28637 ) | ( n28323 & n35646 ) | ( n28637 & n35646 ) ;
  assign n44830 = n41856 ^ n5324 ^ 1'b0 ;
  assign n44831 = n2787 | n44830 ;
  assign n44832 = n19070 | n44831 ;
  assign n44834 = n12952 & n20600 ;
  assign n44835 = n6091 & n44834 ;
  assign n44836 = n526 & ~n44835 ;
  assign n44833 = n18979 & n36322 ;
  assign n44837 = n44836 ^ n44833 ^ 1'b0 ;
  assign n44838 = n11652 ^ n10848 ^ 1'b0 ;
  assign n44839 = n21024 ^ n10523 ^ 1'b0 ;
  assign n44840 = n44838 & n44839 ;
  assign n44841 = n42014 ^ n24987 ^ n3906 ;
  assign n44842 = n26712 ^ n17731 ^ 1'b0 ;
  assign n44843 = n21241 ^ n3416 ^ 1'b0 ;
  assign n44844 = n27963 & n44843 ;
  assign n44845 = n15310 ^ n6747 ^ 1'b0 ;
  assign n44846 = n29932 & n44845 ;
  assign n44847 = n4665 & n44846 ;
  assign n44848 = n15772 | n44582 ;
  assign n44849 = n1134 | n44848 ;
  assign n44850 = n12963 | n13943 ;
  assign n44851 = n12943 ^ n10859 ^ 1'b0 ;
  assign n44852 = n16189 | n44851 ;
  assign n44853 = ~n6771 & n38400 ;
  assign n44854 = ~n26316 & n44853 ;
  assign n44855 = n816 | n35554 ;
  assign n44856 = n24607 | n44855 ;
  assign n44858 = ~n4239 & n18361 ;
  assign n44857 = n32265 & n35097 ;
  assign n44859 = n44858 ^ n44857 ^ n15249 ;
  assign n44860 = n7786 & n32861 ;
  assign n44861 = ~n9377 & n14365 ;
  assign n44862 = ~n20781 & n44861 ;
  assign n44863 = n17070 & n44862 ;
  assign n44864 = n28842 & ~n39009 ;
  assign n44865 = ~n31327 & n44864 ;
  assign n44866 = n5718 ^ n4633 ^ 1'b0 ;
  assign n44867 = n10140 | n37672 ;
  assign n44868 = n5725 & n8041 ;
  assign n44869 = n9500 & ~n13859 ;
  assign n44870 = n6182 & ~n19991 ;
  assign n44871 = n44870 ^ n3305 ^ 1'b0 ;
  assign n44872 = ~n5634 & n10284 ;
  assign n44873 = n44872 ^ n15195 ^ 1'b0 ;
  assign n44874 = n35247 ^ n8820 ^ 1'b0 ;
  assign n44875 = ~n1387 & n39212 ;
  assign n44876 = n838 & n44875 ;
  assign n44877 = n11105 ^ n3372 ^ 1'b0 ;
  assign n44878 = n23112 & ~n44877 ;
  assign n44879 = n24050 & n39246 ;
  assign n44880 = n5164 | n29699 ;
  assign n44881 = n44880 ^ n28063 ^ 1'b0 ;
  assign n44882 = n26109 ^ n777 ^ 1'b0 ;
  assign n44883 = n23294 & n44882 ;
  assign n44884 = ~n10390 & n44883 ;
  assign n44885 = n44881 & ~n44884 ;
  assign n44886 = ( n29534 & n44020 ) | ( n29534 & ~n44885 ) | ( n44020 & ~n44885 ) ;
  assign n44887 = ~n33209 & n39646 ;
  assign n44888 = n24793 ^ n16853 ^ 1'b0 ;
  assign n44889 = ~n27072 & n44888 ;
  assign n44890 = n6080 & ~n16934 ;
  assign n44891 = ~n7380 & n44890 ;
  assign n44892 = n33274 ^ n14855 ^ 1'b0 ;
  assign n44893 = ~n44891 & n44892 ;
  assign n44894 = ~n8747 & n9317 ;
  assign n44895 = n44894 ^ n12349 ^ 1'b0 ;
  assign n44896 = n35831 | n44895 ;
  assign n44897 = n7470 ^ n1540 ^ 1'b0 ;
  assign n44898 = n19596 | n30586 ;
  assign n44899 = n44898 ^ n17020 ^ 1'b0 ;
  assign n44900 = n35998 | n44899 ;
  assign n44901 = n5521 ^ n2716 ^ 1'b0 ;
  assign n44902 = n6131 & n44901 ;
  assign n44903 = ( ~n22104 & n22225 ) | ( ~n22104 & n24795 ) | ( n22225 & n24795 ) ;
  assign n44904 = ( n25884 & n44902 ) | ( n25884 & ~n44903 ) | ( n44902 & ~n44903 ) ;
  assign n44905 = ( n34229 & n44900 ) | ( n34229 & ~n44904 ) | ( n44900 & ~n44904 ) ;
  assign n44906 = ( n1979 & n13104 ) | ( n1979 & n16372 ) | ( n13104 & n16372 ) ;
  assign n44907 = ~n7090 & n20899 ;
  assign n44908 = n44907 ^ n7571 ^ 1'b0 ;
  assign n44909 = n9260 & n19857 ;
  assign n44910 = n44909 ^ n17395 ^ 1'b0 ;
  assign n44911 = n26775 & ~n44910 ;
  assign n44912 = n25921 ^ n13810 ^ 1'b0 ;
  assign n44913 = n30055 | n44912 ;
  assign n44914 = n3626 | n5494 ;
  assign n44915 = n38392 & ~n44914 ;
  assign n44916 = n44915 ^ n25685 ^ 1'b0 ;
  assign n44917 = n25666 ^ n4060 ^ 1'b0 ;
  assign n44918 = n3314 & n44378 ;
  assign n44919 = n3268 & ~n15426 ;
  assign n44920 = n44919 ^ n22620 ^ 1'b0 ;
  assign n44921 = n10247 & n44920 ;
  assign n44922 = ~n5834 & n5925 ;
  assign n44923 = ~n20625 & n44922 ;
  assign n44924 = n1793 ^ n889 ^ 1'b0 ;
  assign n44925 = ~n44923 & n44924 ;
  assign n44926 = n44925 ^ n23392 ^ n18495 ;
  assign n44927 = n23986 ^ n1937 ^ 1'b0 ;
  assign n44928 = n44927 ^ n3000 ^ 1'b0 ;
  assign n44929 = n32770 ^ n9439 ^ 1'b0 ;
  assign n44930 = n4854 & ~n44929 ;
  assign n44931 = ~n31288 & n42441 ;
  assign n44932 = ~n44930 & n44931 ;
  assign n44933 = n11569 & ~n44932 ;
  assign n44934 = n37094 ^ n31143 ^ 1'b0 ;
  assign n44935 = n36119 ^ n23443 ^ 1'b0 ;
  assign n44936 = n44934 | n44935 ;
  assign n44937 = n30489 ^ n21005 ^ n19545 ;
  assign n44939 = n2619 | n14781 ;
  assign n44940 = n44939 ^ n13520 ^ n906 ;
  assign n44941 = ~n33745 & n44940 ;
  assign n44938 = n2354 & ~n28424 ;
  assign n44942 = n44941 ^ n44938 ^ 1'b0 ;
  assign n44943 = n645 ^ n499 ^ 1'b0 ;
  assign n44944 = n6422 & n44943 ;
  assign n44945 = n44944 ^ n12366 ^ 1'b0 ;
  assign n44946 = n32475 ^ n24153 ^ 1'b0 ;
  assign n44947 = n32078 | n44946 ;
  assign n44948 = ( n12271 & n14616 ) | ( n12271 & n39264 ) | ( n14616 & n39264 ) ;
  assign n44949 = n44948 ^ n30791 ^ 1'b0 ;
  assign n44950 = n9481 & ~n35663 ;
  assign n44951 = ~n25502 & n27472 ;
  assign n44952 = n38645 | n40901 ;
  assign n44953 = n30830 ^ n6568 ^ 1'b0 ;
  assign n44954 = n6455 ^ n6443 ^ 1'b0 ;
  assign n44955 = n15558 | n44954 ;
  assign n44957 = x6 & ~n28 ;
  assign n44958 = n28 & n44957 ;
  assign n44959 = n97 | n44958 ;
  assign n44960 = n44958 & ~n44959 ;
  assign n44961 = n517 | n3037 ;
  assign n44962 = n517 & ~n44961 ;
  assign n44963 = n1109 & n44962 ;
  assign n44964 = n249 & ~n44963 ;
  assign n44965 = n44960 & n44964 ;
  assign n44966 = n1036 & n1149 ;
  assign n44967 = ~n1149 & n44966 ;
  assign n44968 = n44965 & ~n44967 ;
  assign n44969 = n16236 | n44968 ;
  assign n44970 = n44969 ^ n11483 ^ 1'b0 ;
  assign n44971 = ~n21803 & n44970 ;
  assign n44972 = n2712 | n11142 ;
  assign n44973 = n44971 | n44972 ;
  assign n44956 = n2374 & ~n7008 ;
  assign n44974 = n44973 ^ n44956 ^ 1'b0 ;
  assign n44976 = n5874 | n9453 ;
  assign n44975 = n1046 & n9276 ;
  assign n44977 = n44976 ^ n44975 ^ 1'b0 ;
  assign n44978 = n21506 & ~n35334 ;
  assign n44979 = n34222 & ~n44978 ;
  assign n44980 = ~n44977 & n44979 ;
  assign n44981 = n35847 ^ n7033 ^ 1'b0 ;
  assign n44982 = n29766 | n44981 ;
  assign n44983 = n42728 ^ n13091 ^ 1'b0 ;
  assign n44984 = n13213 & n41906 ;
  assign n44985 = n21607 ^ n3087 ^ 1'b0 ;
  assign n44986 = n29614 ^ n27233 ^ n585 ;
  assign n44989 = ~n13011 & n31200 ;
  assign n44987 = n12777 ^ n9908 ^ 1'b0 ;
  assign n44988 = n44373 | n44987 ;
  assign n44990 = n44989 ^ n44988 ^ 1'b0 ;
  assign n44991 = ~n15649 & n39168 ;
  assign n44992 = ~n3409 & n17782 ;
  assign n44993 = n3807 & n44992 ;
  assign n44994 = n29119 & ~n44993 ;
  assign n44995 = n2918 & ~n28805 ;
  assign n44996 = ( n3912 & n9448 ) | ( n3912 & ~n44405 ) | ( n9448 & ~n44405 ) ;
  assign n44997 = n4857 & ~n21683 ;
  assign n44998 = ~n4857 & n44997 ;
  assign n44999 = ( n27534 & n37318 ) | ( n27534 & ~n44998 ) | ( n37318 & ~n44998 ) ;
  assign n45000 = n2621 & n14371 ;
  assign n45001 = ( n13732 & ~n44999 ) | ( n13732 & n45000 ) | ( ~n44999 & n45000 ) ;
  assign n45002 = n28465 ^ n17748 ^ 1'b0 ;
  assign n45003 = n7512 | n44919 ;
  assign n45004 = n45003 ^ n31968 ^ 1'b0 ;
  assign n45005 = ( ~n6481 & n8172 ) | ( ~n6481 & n15533 ) | ( n8172 & n15533 ) ;
  assign n45006 = n8901 & n45005 ;
  assign n45007 = n45006 ^ n19030 ^ 1'b0 ;
  assign n45008 = n45007 ^ n38458 ^ n41 ;
  assign n45009 = ~n12065 & n26822 ;
  assign n45010 = n3234 | n19965 ;
  assign n45011 = n45010 ^ n22411 ^ 1'b0 ;
  assign n45012 = n30026 & n45011 ;
  assign n45016 = n19220 ^ n2447 ^ 1'b0 ;
  assign n45017 = n134 & n45016 ;
  assign n45018 = n14285 | n45017 ;
  assign n45013 = n10578 ^ n7761 ^ 1'b0 ;
  assign n45014 = n45013 ^ n35826 ^ 1'b0 ;
  assign n45015 = n18497 & n45014 ;
  assign n45019 = n45018 ^ n45015 ^ n16856 ;
  assign n45020 = n10520 | n21643 ;
  assign n45021 = n9068 | n13969 ;
  assign n45023 = ~n22310 & n29081 ;
  assign n45022 = n7866 & ~n43881 ;
  assign n45024 = n45023 ^ n45022 ^ 1'b0 ;
  assign n45025 = n30116 ^ n20773 ^ n11717 ;
  assign n45026 = n34621 ^ n25766 ^ 1'b0 ;
  assign n45027 = n29358 ^ n21803 ^ 1'b0 ;
  assign n45028 = n34844 ^ n14052 ^ 1'b0 ;
  assign n45029 = n21655 ^ n12747 ^ 1'b0 ;
  assign n45030 = n45028 | n45029 ;
  assign n45031 = n24327 & ~n39221 ;
  assign n45032 = ~n23873 & n28319 ;
  assign n45033 = n45031 & n45032 ;
  assign n45034 = n34463 ^ n16492 ^ 1'b0 ;
  assign n45035 = ~n18486 & n45034 ;
  assign n45036 = n42308 ^ n24860 ^ 1'b0 ;
  assign n45037 = n22457 & ~n45036 ;
  assign n45038 = n5350 & n45037 ;
  assign n45039 = n21546 & n45038 ;
  assign n45040 = n45039 ^ n32819 ^ 1'b0 ;
  assign n45041 = n45035 & n45040 ;
  assign n45042 = ~n19171 & n31486 ;
  assign n45043 = n16829 | n28088 ;
  assign n45044 = n22867 & ~n45043 ;
  assign n45045 = n45044 ^ n16712 ^ n5806 ;
  assign n45051 = n20619 & n22369 ;
  assign n45046 = n6227 & n9479 ;
  assign n45047 = ~n73 & n10087 ;
  assign n45048 = ~n13920 & n45047 ;
  assign n45049 = n37972 | n45048 ;
  assign n45050 = n45046 | n45049 ;
  assign n45052 = n45051 ^ n45050 ^ 1'b0 ;
  assign n45053 = ( ~n10164 & n23971 ) | ( ~n10164 & n45052 ) | ( n23971 & n45052 ) ;
  assign n45054 = n45053 ^ n18748 ^ 1'b0 ;
  assign n45055 = n22588 & ~n34987 ;
  assign n45056 = n45055 ^ n32351 ^ 1'b0 ;
  assign n45057 = n21840 | n38511 ;
  assign n45058 = n25357 | n45057 ;
  assign n45059 = n36976 ^ n14029 ^ 1'b0 ;
  assign n45060 = n6766 & ~n40680 ;
  assign n45061 = ~n8340 & n45060 ;
  assign n45062 = n4870 | n45061 ;
  assign n45063 = n45059 & ~n45062 ;
  assign n45065 = ~n14816 & n27402 ;
  assign n45066 = n37429 & n45065 ;
  assign n45064 = n17487 | n26674 ;
  assign n45067 = n45066 ^ n45064 ^ 1'b0 ;
  assign n45068 = n7002 & ~n34018 ;
  assign n45069 = n14222 & n45068 ;
  assign n45070 = n45069 ^ n17961 ^ 1'b0 ;
  assign n45071 = n24844 & ~n45070 ;
  assign n45072 = ~n151 & n9904 ;
  assign n45073 = n45072 ^ n20421 ^ 1'b0 ;
  assign n45074 = n545 & ~n9162 ;
  assign n45075 = n45074 ^ n7354 ^ 1'b0 ;
  assign n45076 = ( ~n28886 & n45073 ) | ( ~n28886 & n45075 ) | ( n45073 & n45075 ) ;
  assign n45077 = n27673 ^ n7740 ^ 1'b0 ;
  assign n45078 = n1064 | n45077 ;
  assign n45079 = n4673 ^ n4588 ^ 1'b0 ;
  assign n45080 = ( n1768 & n45078 ) | ( n1768 & ~n45079 ) | ( n45078 & ~n45079 ) ;
  assign n45081 = n4545 & n27064 ;
  assign n45082 = n45081 ^ x10 ^ 1'b0 ;
  assign n45083 = n26071 & n45082 ;
  assign n45084 = n33715 ^ n32324 ^ 1'b0 ;
  assign n45085 = n5479 & ~n8532 ;
  assign n45086 = n45085 ^ n24828 ^ 1'b0 ;
  assign n45087 = n6452 ^ n159 ^ 1'b0 ;
  assign n45088 = ~n18161 & n20269 ;
  assign n45089 = n11514 & ~n20691 ;
  assign n45090 = n25879 ^ n2846 ^ 1'b0 ;
  assign n45091 = n45089 | n45090 ;
  assign n45092 = n45091 ^ n34946 ^ n20924 ;
  assign n45093 = n37404 ^ n6877 ^ 1'b0 ;
  assign n45094 = n40165 ^ n27645 ^ n26446 ;
  assign n45095 = ~n633 & n45094 ;
  assign n45096 = ( n126 & ~n23774 ) | ( n126 & n37772 ) | ( ~n23774 & n37772 ) ;
  assign n45097 = n45095 & ~n45096 ;
  assign n45099 = n16462 & ~n33872 ;
  assign n45098 = ~n33955 & n39672 ;
  assign n45100 = n45099 ^ n45098 ^ 1'b0 ;
  assign n45101 = n40988 ^ n36100 ^ 1'b0 ;
  assign n45102 = n780 & n45101 ;
  assign n45103 = n25747 & n45102 ;
  assign n45104 = n12131 & ~n26332 ;
  assign n45105 = n34565 ^ n4848 ^ 1'b0 ;
  assign n45106 = n8920 & ~n45105 ;
  assign n45107 = n45106 ^ n8197 ^ 1'b0 ;
  assign n45108 = ( n5903 & n6904 ) | ( n5903 & ~n9755 ) | ( n6904 & ~n9755 ) ;
  assign n45109 = n10274 & ~n27876 ;
  assign n45110 = n45108 | n45109 ;
  assign n45111 = n28723 & ~n32369 ;
  assign n45112 = ~n26156 & n45111 ;
  assign n45113 = n42261 | n45112 ;
  assign n45114 = n45113 ^ n7243 ^ n1854 ;
  assign n45115 = ( n11636 & ~n17200 ) | ( n11636 & n26567 ) | ( ~n17200 & n26567 ) ;
  assign n45116 = n45115 ^ n5533 ^ 1'b0 ;
  assign n45117 = ( n12522 & n16644 ) | ( n12522 & n45116 ) | ( n16644 & n45116 ) ;
  assign n45121 = n6949 ^ n4571 ^ 1'b0 ;
  assign n45122 = n3878 | n45121 ;
  assign n45118 = n21304 ^ n7319 ^ 1'b0 ;
  assign n45119 = n37335 & ~n45118 ;
  assign n45120 = n28687 & n45119 ;
  assign n45123 = n45122 ^ n45120 ^ 1'b0 ;
  assign n45124 = n8615 ^ n7626 ^ n1260 ;
  assign n45125 = ~n396 & n10239 ;
  assign n45126 = n45125 ^ n29244 ^ 1'b0 ;
  assign n45127 = n10297 & n45126 ;
  assign n45128 = ~n31996 & n45127 ;
  assign n45129 = n45128 ^ n23758 ^ 1'b0 ;
  assign n45130 = ~n45124 & n45129 ;
  assign n45131 = n29027 ^ n18027 ^ n1423 ;
  assign n45132 = ~n26430 & n45131 ;
  assign n45133 = ~n16810 & n29423 ;
  assign n45134 = n45133 ^ n16870 ^ 1'b0 ;
  assign n45135 = ~n10941 & n26582 ;
  assign n45136 = n517 & n45135 ;
  assign n45137 = n42963 & ~n45136 ;
  assign n45138 = n42698 ^ n34166 ^ 1'b0 ;
  assign n45139 = ~n3703 & n26420 ;
  assign n45140 = n9089 | n14862 ;
  assign n45141 = n45140 ^ n37251 ^ 1'b0 ;
  assign n45142 = ~n24834 & n39246 ;
  assign n45143 = n20003 | n25247 ;
  assign n45144 = n45142 | n45143 ;
  assign n45145 = n13057 & n45144 ;
  assign n45146 = n10861 | n27334 ;
  assign n45147 = n45146 ^ n27721 ^ n18408 ;
  assign n45148 = ( n19436 & ~n23441 ) | ( n19436 & n41690 ) | ( ~n23441 & n41690 ) ;
  assign n45149 = n7296 | n41681 ;
  assign n45150 = n45149 ^ n37442 ^ 1'b0 ;
  assign n45151 = ~n45148 & n45150 ;
  assign n45152 = n27735 ^ n6186 ^ 1'b0 ;
  assign n45153 = n856 & ~n1861 ;
  assign n45154 = n21941 ^ n1235 ^ 1'b0 ;
  assign n45155 = n45153 & n45154 ;
  assign n45156 = n23018 ^ n9851 ^ 1'b0 ;
  assign n45157 = n15920 & ~n45156 ;
  assign n45158 = ( n10946 & n20547 ) | ( n10946 & n25913 ) | ( n20547 & n25913 ) ;
  assign n45159 = ~n17436 & n23996 ;
  assign n45160 = ( ~n41300 & n45158 ) | ( ~n41300 & n45159 ) | ( n45158 & n45159 ) ;
  assign n45161 = n26800 ^ n12010 ^ n3640 ;
  assign n45162 = n45161 ^ n29898 ^ n11788 ;
  assign n45163 = n9408 ^ n1944 ^ 1'b0 ;
  assign n45164 = n3640 ^ n2902 ^ 1'b0 ;
  assign n45165 = ~n45163 & n45164 ;
  assign n45166 = n17646 & n45165 ;
  assign n45167 = n45166 ^ n722 ^ 1'b0 ;
  assign n45168 = ~n753 & n9855 ;
  assign n45169 = n945 | n31224 ;
  assign n45170 = n45168 | n45169 ;
  assign n45171 = n28967 ^ n21238 ^ 1'b0 ;
  assign n45172 = ~n43503 & n45171 ;
  assign n45173 = n24036 ^ n18211 ^ 1'b0 ;
  assign n45174 = n242 | n45173 ;
  assign n45175 = n45174 ^ n10994 ^ 1'b0 ;
  assign n45176 = ( n4889 & ~n17641 ) | ( n4889 & n45175 ) | ( ~n17641 & n45175 ) ;
  assign n45177 = n14033 ^ n9009 ^ 1'b0 ;
  assign n45178 = n22340 ^ n12925 ^ 1'b0 ;
  assign n45179 = n26161 ^ n20070 ^ n18723 ;
  assign n45180 = ~n5254 & n45179 ;
  assign n45181 = n33225 ^ n19615 ^ 1'b0 ;
  assign n45182 = n14083 & ~n45181 ;
  assign n45183 = n14698 & ~n30422 ;
  assign n45184 = n40633 ^ n7328 ^ 1'b0 ;
  assign n45185 = n43737 & ~n45184 ;
  assign n45186 = n21185 ^ n465 ^ 1'b0 ;
  assign n45187 = ( ~n1470 & n27033 ) | ( ~n1470 & n45186 ) | ( n27033 & n45186 ) ;
  assign n45188 = n1261 & n26783 ;
  assign n45189 = ~n23534 & n45188 ;
  assign n45192 = n20929 ^ n9020 ^ 1'b0 ;
  assign n45190 = ~n25494 & n27690 ;
  assign n45191 = ~n2582 & n45190 ;
  assign n45193 = n45192 ^ n45191 ^ 1'b0 ;
  assign n45194 = n45189 | n45193 ;
  assign n45195 = n12404 ^ n9912 ^ n7812 ;
  assign n45196 = n12304 & ~n45195 ;
  assign n45197 = n45196 ^ n2012 ^ 1'b0 ;
  assign n45198 = n45197 ^ n8441 ^ 1'b0 ;
  assign n45199 = n3754 & ~n42712 ;
  assign n45200 = n45198 & n45199 ;
  assign n45201 = n29653 ^ n15414 ^ 1'b0 ;
  assign n45202 = n45201 ^ n28857 ^ n15630 ;
  assign n45203 = n38759 | n45202 ;
  assign n45204 = n45203 ^ n23094 ^ 1'b0 ;
  assign n45205 = n43934 ^ n40895 ^ n6041 ;
  assign n45207 = n1789 | n3991 ;
  assign n45206 = n19135 | n22001 ;
  assign n45208 = n45207 ^ n45206 ^ 1'b0 ;
  assign n45209 = n6888 & ~n45208 ;
  assign n45210 = n45209 ^ n9981 ^ 1'b0 ;
  assign n45211 = n12465 ^ n866 ^ 1'b0 ;
  assign n45212 = n45211 ^ n36019 ^ 1'b0 ;
  assign n45213 = n13508 ^ n7194 ^ 1'b0 ;
  assign n45214 = n40834 & n45213 ;
  assign n45215 = n16786 ^ n10931 ^ 1'b0 ;
  assign n45216 = n5370 | n45215 ;
  assign n45217 = n26238 ^ n16056 ^ 1'b0 ;
  assign n45218 = n2696 & ~n11722 ;
  assign n45219 = n39058 ^ n1506 ^ 1'b0 ;
  assign n45220 = ~n6942 & n10220 ;
  assign n45221 = n45220 ^ n9830 ^ 1'b0 ;
  assign n45222 = ( n18093 & n20264 ) | ( n18093 & n45221 ) | ( n20264 & n45221 ) ;
  assign n45223 = n11982 | n45222 ;
  assign n45224 = n997 & ~n12438 ;
  assign n45225 = n45223 & n45224 ;
  assign n45226 = ~n45219 & n45225 ;
  assign n45227 = ~n99 & n12431 ;
  assign n45228 = n45227 ^ n749 ^ 1'b0 ;
  assign n45229 = n27789 & n45228 ;
  assign n45230 = n6277 & n11701 ;
  assign n45231 = ~n19450 & n45230 ;
  assign n45232 = n8696 & ~n45231 ;
  assign n45233 = ~n918 & n45232 ;
  assign n45234 = n32946 ^ n10777 ^ 1'b0 ;
  assign n45235 = n5683 & n45234 ;
  assign n45236 = ~n22470 & n45235 ;
  assign n45237 = n14173 & ~n45236 ;
  assign n45238 = n25404 ^ n1481 ^ 1'b0 ;
  assign n45239 = ~n10105 & n45238 ;
  assign n45240 = ~n11136 & n25768 ;
  assign n45241 = n40042 ^ n35667 ^ n20469 ;
  assign n45242 = n5160 & ~n7158 ;
  assign n45243 = n6817 & ~n9158 ;
  assign n45244 = n11150 & n45243 ;
  assign n45245 = n45244 ^ n15928 ^ 1'b0 ;
  assign n45246 = n45245 ^ n40 ^ 1'b0 ;
  assign n45247 = n13274 ^ n11298 ^ 1'b0 ;
  assign n45248 = n33791 ^ n5069 ^ n2178 ;
  assign n45249 = n45248 ^ n17183 ^ 1'b0 ;
  assign n45250 = n5418 & n5617 ;
  assign n45251 = ~n20689 & n45250 ;
  assign n45252 = n45251 ^ n25566 ^ 1'b0 ;
  assign n45253 = n604 | n45252 ;
  assign n45254 = n13021 | n45253 ;
  assign n45255 = n8244 ^ n6332 ^ 1'b0 ;
  assign n45256 = ~n19883 & n45255 ;
  assign n45257 = ~n44743 & n45256 ;
  assign n45258 = n19994 & n40688 ;
  assign n45259 = n16035 & ~n25940 ;
  assign n45260 = n23351 & n45259 ;
  assign n45261 = n26293 & ~n45260 ;
  assign n45262 = ~n21829 & n35210 ;
  assign n45263 = n45262 ^ n23238 ^ n5312 ;
  assign n45264 = n25396 & n45263 ;
  assign n45265 = n1079 | n4160 ;
  assign n45266 = n45265 ^ n6355 ^ 1'b0 ;
  assign n45267 = n45266 ^ n15982 ^ 1'b0 ;
  assign n45268 = n7722 & ~n11102 ;
  assign n45269 = n18134 ^ n6643 ^ 1'b0 ;
  assign n45276 = n3666 & n17128 ;
  assign n45277 = n45276 ^ n25479 ^ 1'b0 ;
  assign n45270 = n3882 ^ n204 ^ 1'b0 ;
  assign n45271 = n16731 & ~n45270 ;
  assign n45272 = n15396 & ~n45271 ;
  assign n45273 = ~n15560 & n45272 ;
  assign n45274 = ( ~n1677 & n45128 ) | ( ~n1677 & n45273 ) | ( n45128 & n45273 ) ;
  assign n45275 = n7087 | n45274 ;
  assign n45278 = n45277 ^ n45275 ^ 1'b0 ;
  assign n45279 = ~n9416 & n14715 ;
  assign n45280 = n45279 ^ n19580 ^ 1'b0 ;
  assign n45281 = n8054 | n23930 ;
  assign n45282 = n45281 ^ n18556 ^ n9181 ;
  assign n45283 = n18601 & ~n45282 ;
  assign n45284 = ~n45280 & n45283 ;
  assign n45285 = n19258 ^ n14760 ^ n792 ;
  assign n45286 = n5335 | n15651 ;
  assign n45287 = n19654 & n30926 ;
  assign n45288 = n37067 ^ n16363 ^ n2532 ;
  assign n45289 = n45288 ^ n12225 ^ 1'b0 ;
  assign n45290 = n14740 & n45289 ;
  assign n45291 = n2196 & n10656 ;
  assign n45292 = n4110 & n45291 ;
  assign n45293 = ~n17473 & n45292 ;
  assign n45294 = n6711 | n14124 ;
  assign n45295 = n45294 ^ n6956 ^ 1'b0 ;
  assign n45296 = n9621 & n45295 ;
  assign n45297 = n30453 & n45296 ;
  assign n45298 = n33690 ^ n6199 ^ 1'b0 ;
  assign n45306 = n22903 ^ n5415 ^ 1'b0 ;
  assign n45300 = ~n5924 & n7505 ;
  assign n45301 = ~n18164 & n45300 ;
  assign n45302 = n45301 ^ n16047 ^ 1'b0 ;
  assign n45303 = n7228 ^ n4110 ^ 1'b0 ;
  assign n45304 = n45302 & ~n45303 ;
  assign n45299 = ~n18299 & n25902 ;
  assign n45305 = n45304 ^ n45299 ^ 1'b0 ;
  assign n45307 = n45306 ^ n45305 ^ 1'b0 ;
  assign n45308 = n5160 & ~n9162 ;
  assign n45309 = n45308 ^ n15815 ^ 1'b0 ;
  assign n45310 = n19147 & ~n28855 ;
  assign n45311 = ~n4427 & n45310 ;
  assign n45312 = n3961 & ~n34036 ;
  assign n45313 = n34345 & ~n45312 ;
  assign n45314 = ( n6578 & ~n26446 ) | ( n6578 & n45313 ) | ( ~n26446 & n45313 ) ;
  assign n45315 = n18730 ^ n17694 ^ n12167 ;
  assign n45316 = n10118 ^ n2721 ^ n499 ;
  assign n45317 = n45316 ^ n25933 ^ 1'b0 ;
  assign n45318 = n614 & n45317 ;
  assign n45319 = n8247 & ~n12670 ;
  assign n45320 = n45319 ^ n40674 ^ 1'b0 ;
  assign n45321 = n15064 | n44334 ;
  assign n45322 = n32743 & ~n45321 ;
  assign n45323 = n17798 & n27490 ;
  assign n45324 = n45323 ^ n2784 ^ 1'b0 ;
  assign n45325 = n9631 & n14572 ;
  assign n45326 = n1395 | n34884 ;
  assign n45327 = n45325 | n45326 ;
  assign n45328 = n30935 ^ n16075 ^ n249 ;
  assign n45329 = ( n31628 & n45327 ) | ( n31628 & ~n45328 ) | ( n45327 & ~n45328 ) ;
  assign n45331 = n31244 ^ n11032 ^ n3551 ;
  assign n45330 = n8371 & n19598 ;
  assign n45332 = n45331 ^ n45330 ^ 1'b0 ;
  assign n45333 = n11465 ^ n378 ^ 1'b0 ;
  assign n45334 = ( n8313 & n22055 ) | ( n8313 & ~n28476 ) | ( n22055 & ~n28476 ) ;
  assign n45335 = n45334 ^ n12779 ^ 1'b0 ;
  assign n45336 = ( n18421 & ~n21395 ) | ( n18421 & n42148 ) | ( ~n21395 & n42148 ) ;
  assign n45337 = n45336 ^ n756 ^ 1'b0 ;
  assign n45338 = ~n38188 & n45337 ;
  assign n45339 = n17440 & ~n19083 ;
  assign n45340 = ( n18998 & ~n28282 ) | ( n18998 & n34929 ) | ( ~n28282 & n34929 ) ;
  assign n45341 = n1097 ^ n350 ^ 1'b0 ;
  assign n45342 = n45341 ^ n19209 ^ n2049 ;
  assign n45343 = n45342 ^ n6496 ^ 1'b0 ;
  assign n45344 = n9633 | n45343 ;
  assign n45345 = n40703 ^ n5160 ^ 1'b0 ;
  assign n45346 = ~n25409 & n45345 ;
  assign n45347 = n31169 ^ n11256 ^ 1'b0 ;
  assign n45348 = ~n38437 & n45347 ;
  assign n45349 = n16223 ^ n2673 ^ 1'b0 ;
  assign n45350 = ~n6067 & n45349 ;
  assign n45351 = n9802 | n32447 ;
  assign n45352 = n45351 ^ n13316 ^ 1'b0 ;
  assign n45353 = n26043 ^ n5749 ^ 1'b0 ;
  assign n45354 = ~n19236 & n45353 ;
  assign n45355 = n17993 ^ n2955 ^ 1'b0 ;
  assign n45356 = n17994 & n45355 ;
  assign n45357 = n35103 & n45356 ;
  assign n45358 = n13201 ^ n8023 ^ 1'b0 ;
  assign n45359 = n12696 | n45358 ;
  assign n45360 = ( ~n5076 & n10211 ) | ( ~n5076 & n17290 ) | ( n10211 & n17290 ) ;
  assign n45361 = n9843 ^ n7862 ^ 1'b0 ;
  assign n45362 = ( ~n10707 & n31520 ) | ( ~n10707 & n45361 ) | ( n31520 & n45361 ) ;
  assign n45363 = n15084 ^ n7282 ^ 1'b0 ;
  assign n45365 = n3059 & n18587 ;
  assign n45364 = n1332 & n23463 ;
  assign n45366 = n45365 ^ n45364 ^ 1'b0 ;
  assign n45367 = n22941 ^ n13394 ^ 1'b0 ;
  assign n45368 = n15370 | n45367 ;
  assign n45369 = n19346 ^ n8400 ^ n925 ;
  assign n45370 = n45369 ^ n10733 ^ 1'b0 ;
  assign n45371 = n7325 | n45370 ;
  assign n45372 = ( n9050 & n14102 ) | ( n9050 & n42977 ) | ( n14102 & n42977 ) ;
  assign n45378 = n13469 | n37786 ;
  assign n45379 = n45378 ^ n24863 ^ 1'b0 ;
  assign n45375 = n15678 ^ n13991 ^ 1'b0 ;
  assign n45376 = ~n9130 & n45375 ;
  assign n45377 = n45376 ^ n13164 ^ 1'b0 ;
  assign n45373 = n43841 ^ n34899 ^ 1'b0 ;
  assign n45374 = n2544 & ~n45373 ;
  assign n45380 = n45379 ^ n45377 ^ n45374 ;
  assign n45381 = n567 & ~n23351 ;
  assign n45382 = n45381 ^ n3491 ^ 1'b0 ;
  assign n45383 = n3022 & n16841 ;
  assign n45384 = n45383 ^ n8676 ^ 1'b0 ;
  assign n45385 = n5132 | n44753 ;
  assign n45386 = n45384 & ~n45385 ;
  assign n45387 = ( n23193 & n45382 ) | ( n23193 & ~n45386 ) | ( n45382 & ~n45386 ) ;
  assign n45388 = n23726 & n29929 ;
  assign n45389 = n26175 ^ n8975 ^ 1'b0 ;
  assign n45390 = n5099 & ~n45389 ;
  assign n45391 = n22639 ^ n2105 ^ 1'b0 ;
  assign n45392 = n23500 ^ n19461 ^ n8655 ;
  assign n45393 = n45392 ^ n20096 ^ 1'b0 ;
  assign n45394 = n45393 ^ n33633 ^ n18509 ;
  assign n45395 = n45394 ^ n29049 ^ 1'b0 ;
  assign n45396 = n4126 & ~n36682 ;
  assign n45397 = n45396 ^ n6646 ^ 1'b0 ;
  assign n45398 = ~n1633 & n7975 ;
  assign n45399 = n3710 & n45398 ;
  assign n45400 = n41987 ^ n20743 ^ 1'b0 ;
  assign n45401 = n9952 & ~n35880 ;
  assign n45402 = n5803 & ~n39954 ;
  assign n45403 = ~n45401 & n45402 ;
  assign n45404 = n20336 & ~n30479 ;
  assign n45405 = n17499 & n45404 ;
  assign n45406 = n1186 & n21612 ;
  assign n45407 = ~n36656 & n45406 ;
  assign n45408 = n9570 & ~n45407 ;
  assign n45409 = n18509 ^ n10689 ^ n6746 ;
  assign n45410 = n26997 ^ n12991 ^ n5607 ;
  assign n45411 = ~n13548 & n29930 ;
  assign n45412 = n45411 ^ n983 ^ 1'b0 ;
  assign n45413 = n20570 ^ n17679 ^ 1'b0 ;
  assign n45414 = ~n18508 & n45413 ;
  assign n45415 = n45412 & n45414 ;
  assign n45416 = n14462 ^ n1656 ^ 1'b0 ;
  assign n45417 = n20252 | n24842 ;
  assign n45418 = n45417 ^ n44417 ^ 1'b0 ;
  assign n45419 = n6783 | n15172 ;
  assign n45420 = ~n24205 & n30938 ;
  assign n45421 = n45419 & n45420 ;
  assign n45422 = n43570 ^ n4872 ^ 1'b0 ;
  assign n45423 = n4827 & n14760 ;
  assign n45424 = n1972 & ~n5399 ;
  assign n45425 = n45423 | n45424 ;
  assign n45426 = n6030 & ~n28081 ;
  assign n45427 = n45426 ^ n34351 ^ 1'b0 ;
  assign n45428 = n3317 & ~n33399 ;
  assign n45429 = n42412 & ~n45428 ;
  assign n45430 = n21773 | n45429 ;
  assign n45431 = n2671 | n45430 ;
  assign n45432 = n4878 & n45431 ;
  assign n45433 = n23958 ^ n9061 ^ 1'b0 ;
  assign n45434 = ~n4202 & n11023 ;
  assign n45435 = n45434 ^ n2055 ^ 1'b0 ;
  assign n45436 = n45433 & n45435 ;
  assign n45437 = n19322 & n45436 ;
  assign n45438 = n33896 ^ n19267 ^ 1'b0 ;
  assign n45439 = ~n15108 & n23177 ;
  assign n45440 = ~n10176 & n45439 ;
  assign n45441 = n28511 ^ n14657 ^ 1'b0 ;
  assign n45442 = n37328 | n45441 ;
  assign n45443 = n45442 ^ n33507 ^ n18495 ;
  assign n45444 = ( n18826 & ~n34362 ) | ( n18826 & n38720 ) | ( ~n34362 & n38720 ) ;
  assign n45445 = n31157 ^ n5493 ^ 1'b0 ;
  assign n45446 = n23870 ^ n10185 ^ 1'b0 ;
  assign n45447 = n32100 & ~n45446 ;
  assign n45448 = n26773 & n39900 ;
  assign n45449 = ( ~n2115 & n14999 ) | ( ~n2115 & n45448 ) | ( n14999 & n45448 ) ;
  assign n45450 = n11172 & ~n45449 ;
  assign n45451 = n45450 ^ n21703 ^ 1'b0 ;
  assign n45452 = n45451 ^ n21681 ^ 1'b0 ;
  assign n45453 = n8878 ^ n1856 ^ 1'b0 ;
  assign n45454 = n3758 | n14409 ;
  assign n45455 = n34977 | n45454 ;
  assign n45456 = n45455 ^ n2689 ^ 1'b0 ;
  assign n45457 = n23831 & n45456 ;
  assign n45458 = n3934 & n21437 ;
  assign n45459 = ( ~n45453 & n45457 ) | ( ~n45453 & n45458 ) | ( n45457 & n45458 ) ;
  assign n45460 = n2004 | n3255 ;
  assign n45461 = n14282 & ~n45460 ;
  assign n45462 = n7624 ^ n1281 ^ n53 ;
  assign n45463 = n42217 ^ n25506 ^ 1'b0 ;
  assign n45464 = n45462 & ~n45463 ;
  assign n45465 = n1041 & n35356 ;
  assign n45466 = ~n13017 & n24386 ;
  assign n45467 = ~n45465 & n45466 ;
  assign n45468 = n19319 | n27938 ;
  assign n45469 = n26504 | n45468 ;
  assign n45470 = ( n1857 & ~n16168 ) | ( n1857 & n32465 ) | ( ~n16168 & n32465 ) ;
  assign n45471 = n45470 ^ n38244 ^ n26702 ;
  assign n45472 = n17721 ^ n732 ^ 1'b0 ;
  assign n45473 = n45472 ^ n30996 ^ 1'b0 ;
  assign n45474 = n6309 ^ n5212 ^ 1'b0 ;
  assign n45477 = n1279 | n45195 ;
  assign n45478 = n30196 | n45477 ;
  assign n45476 = n2177 & ~n42979 ;
  assign n45479 = n45478 ^ n45476 ^ 1'b0 ;
  assign n45475 = ~n15636 & n17140 ;
  assign n45480 = n45479 ^ n45475 ^ 1'b0 ;
  assign n45481 = ( n25921 & n30905 ) | ( n25921 & ~n37589 ) | ( n30905 & ~n37589 ) ;
  assign n45482 = ~n14076 & n40763 ;
  assign n45483 = ~n5263 & n45482 ;
  assign n45484 = ~n45481 & n45483 ;
  assign n45486 = ( n37 & ~n16419 ) | ( n37 & n21139 ) | ( ~n16419 & n21139 ) ;
  assign n45485 = n13206 ^ n2544 ^ 1'b0 ;
  assign n45487 = n45486 ^ n45485 ^ n14468 ;
  assign n45488 = n45487 ^ n9926 ^ n6430 ;
  assign n45489 = ~n287 & n1124 ;
  assign n45490 = n45489 ^ n19974 ^ 1'b0 ;
  assign n45491 = n34639 | n45490 ;
  assign n45492 = n24532 ^ n12694 ^ 1'b0 ;
  assign n45493 = n36600 | n45492 ;
  assign n45496 = n29611 ^ n22659 ^ 1'b0 ;
  assign n45494 = n5481 & n24196 ;
  assign n45495 = n30162 | n45494 ;
  assign n45497 = n45496 ^ n45495 ^ 1'b0 ;
  assign n45498 = n45497 ^ n42157 ^ n30389 ;
  assign n45499 = n19716 | n41898 ;
  assign n45500 = n6860 & ~n30188 ;
  assign n45501 = n13089 & n14925 ;
  assign n45502 = n45500 & n45501 ;
  assign n45503 = n7121 ^ n965 ^ 1'b0 ;
  assign n45504 = ( n7873 & ~n13693 ) | ( n7873 & n20713 ) | ( ~n13693 & n20713 ) ;
  assign n45505 = n29476 ^ n19108 ^ 1'b0 ;
  assign n45506 = n36973 ^ n36346 ^ n31216 ;
  assign n45507 = n26087 & n45506 ;
  assign n45508 = n45167 ^ n19869 ^ n12576 ;
  assign n45509 = n37741 ^ n6146 ^ 1'b0 ;
  assign n45510 = ~n6921 & n45509 ;
  assign n45511 = ~n26788 & n31130 ;
  assign n45512 = n45511 ^ n14493 ^ 1'b0 ;
  assign n45513 = n13899 ^ n6082 ^ 1'b0 ;
  assign n45514 = ~n934 & n45513 ;
  assign n45515 = n45514 ^ n17377 ^ 1'b0 ;
  assign n45516 = n4412 | n5641 ;
  assign n45517 = n2048 | n45516 ;
  assign n45518 = n1997 | n45517 ;
  assign n45519 = n16722 & ~n45518 ;
  assign n45520 = ~n5853 & n20882 ;
  assign n45521 = ( n842 & n10404 ) | ( n842 & n15685 ) | ( n10404 & n15685 ) ;
  assign n45522 = n45521 ^ n34370 ^ 1'b0 ;
  assign n45523 = ~n45520 & n45522 ;
  assign n45524 = n1752 | n42394 ;
  assign n45525 = n17122 & ~n45524 ;
  assign n45526 = n38726 ^ n34945 ^ 1'b0 ;
  assign n45527 = ( n5602 & n18093 ) | ( n5602 & ~n25358 ) | ( n18093 & ~n25358 ) ;
  assign n45528 = n13829 & n45527 ;
  assign n45529 = n624 & n18541 ;
  assign n45530 = n10563 & n40710 ;
  assign n45531 = n45530 ^ n33405 ^ n11487 ;
  assign n45532 = n9144 ^ n6804 ^ 1'b0 ;
  assign n45533 = ~n9426 & n36157 ;
  assign n45534 = n45533 ^ n13366 ^ 1'b0 ;
  assign n45535 = n5876 | n26351 ;
  assign n45536 = n9150 | n14832 ;
  assign n45537 = n45536 ^ n7216 ^ 1'b0 ;
  assign n45538 = n20366 | n41481 ;
  assign n45539 = n45538 ^ n7022 ^ 1'b0 ;
  assign n45540 = n2367 ^ n1308 ^ 1'b0 ;
  assign n45541 = n9858 | n45540 ;
  assign n45542 = n34028 ^ n697 ^ 1'b0 ;
  assign n45543 = n12909 | n45542 ;
  assign n45544 = n25253 ^ n7925 ^ 1'b0 ;
  assign n45545 = n45543 | n45544 ;
  assign n45546 = n26436 & ~n45545 ;
  assign n45547 = n45541 & n45546 ;
  assign n45548 = n18225 ^ n5285 ^ 1'b0 ;
  assign n45549 = n10920 ^ n2486 ^ 1'b0 ;
  assign n45550 = n45548 & ~n45549 ;
  assign n45551 = n45550 ^ n20580 ^ n4903 ;
  assign n45552 = n6888 & n42799 ;
  assign n45553 = n2969 & n18462 ;
  assign n45554 = ~n44872 & n45553 ;
  assign n45555 = n19605 ^ n18587 ^ 1'b0 ;
  assign n45556 = n9597 & n45555 ;
  assign n45557 = n45556 ^ n24164 ^ 1'b0 ;
  assign n45558 = n1603 & n25637 ;
  assign n45559 = n31200 ^ n12494 ^ 1'b0 ;
  assign n45560 = ( n15586 & n45558 ) | ( n15586 & ~n45559 ) | ( n45558 & ~n45559 ) ;
  assign n45561 = n45560 ^ n12966 ^ 1'b0 ;
  assign n45562 = ~n13153 & n45561 ;
  assign n45563 = n11921 ^ n4175 ^ 1'b0 ;
  assign n45564 = n45563 ^ n11382 ^ 1'b0 ;
  assign n45565 = n12073 | n45564 ;
  assign n45566 = n4573 & n45565 ;
  assign n45567 = n21688 & n45566 ;
  assign n45571 = n12395 | n26941 ;
  assign n45568 = n853 & ~n23047 ;
  assign n45569 = ~n17114 & n45568 ;
  assign n45570 = n45569 ^ n34774 ^ n10804 ;
  assign n45572 = n45571 ^ n45570 ^ n31688 ;
  assign n45573 = ~n132 & n20781 ;
  assign n45574 = n10978 & n45573 ;
  assign n45575 = n45574 ^ n33307 ^ 1'b0 ;
  assign n45576 = n41375 ^ n27560 ^ 1'b0 ;
  assign n45577 = n3018 & n45576 ;
  assign n45578 = ~n11692 & n45577 ;
  assign n45579 = n26171 & ~n35273 ;
  assign n45580 = ~n13123 & n41559 ;
  assign n45581 = n15017 & n39947 ;
  assign n45582 = n45581 ^ n30488 ^ 1'b0 ;
  assign n45583 = n16339 & n27308 ;
  assign n45584 = n11986 & n45583 ;
  assign n45585 = n7468 & n9495 ;
  assign n45586 = n20819 ^ n12525 ^ 1'b0 ;
  assign n45587 = n45585 | n45586 ;
  assign n45588 = ~n6008 & n26259 ;
  assign n45589 = n7478 ^ n1069 ^ 1'b0 ;
  assign n45595 = ( ~n8195 & n10773 ) | ( ~n8195 & n13368 ) | ( n10773 & n13368 ) ;
  assign n45590 = ~n5770 & n6169 ;
  assign n45591 = ~n8861 & n45590 ;
  assign n45592 = n10527 | n45591 ;
  assign n45593 = ( n8526 & n24505 ) | ( n8526 & n45592 ) | ( n24505 & n45592 ) ;
  assign n45594 = n45593 ^ n485 ^ 1'b0 ;
  assign n45596 = n45595 ^ n45594 ^ n2579 ;
  assign n45597 = ( n5077 & ~n16215 ) | ( n5077 & n19165 ) | ( ~n16215 & n19165 ) ;
  assign n45598 = n14440 ^ n11233 ^ n5897 ;
  assign n45599 = n37200 ^ n2612 ^ 1'b0 ;
  assign n45600 = n7144 & ~n45599 ;
  assign n45601 = n36546 ^ n11967 ^ 1'b0 ;
  assign n45602 = n45600 & n45601 ;
  assign n45603 = n25594 & n44820 ;
  assign n45604 = ~n12477 & n35457 ;
  assign n45605 = n45604 ^ n11345 ^ 1'b0 ;
  assign n45606 = n11609 & ~n45605 ;
  assign n45607 = ~n30068 & n45606 ;
  assign n45608 = n3165 & n45607 ;
  assign n45609 = n4447 | n29158 ;
  assign n45610 = n45609 ^ n38541 ^ 1'b0 ;
  assign n45611 = n17824 & n24173 ;
  assign n45612 = n45611 ^ n19592 ^ 1'b0 ;
  assign n45613 = n45610 & n45612 ;
  assign n45614 = n18716 ^ n17564 ^ 1'b0 ;
  assign n45615 = ~n621 & n6664 ;
  assign n45616 = n45615 ^ n5246 ^ 1'b0 ;
  assign n45617 = n5042 & ~n45616 ;
  assign n45618 = n5109 & n27956 ;
  assign n45619 = n29638 & n45618 ;
  assign n45620 = n25111 ^ n24835 ^ 1'b0 ;
  assign n45621 = n1807 & ~n6557 ;
  assign n45622 = n19472 & n45621 ;
  assign n45623 = n9837 & ~n45622 ;
  assign n45624 = ( n1368 & ~n1840 ) | ( n1368 & n13517 ) | ( ~n1840 & n13517 ) ;
  assign n45625 = n18783 ^ n2579 ^ 1'b0 ;
  assign n45626 = n8550 | n13159 ;
  assign n45627 = ( n2613 & ~n11044 ) | ( n2613 & n45626 ) | ( ~n11044 & n45626 ) ;
  assign n45628 = ( n14443 & ~n34527 ) | ( n14443 & n45627 ) | ( ~n34527 & n45627 ) ;
  assign n45629 = n2729 & n14710 ;
  assign n45630 = n45629 ^ n15856 ^ 1'b0 ;
  assign n45631 = n23950 & n33105 ;
  assign n45632 = n45631 ^ n27666 ^ 1'b0 ;
  assign n45634 = n28952 ^ n4529 ^ 1'b0 ;
  assign n45635 = n12149 & ~n45634 ;
  assign n45636 = n45635 ^ n15592 ^ 1'b0 ;
  assign n45633 = n5022 | n5657 ;
  assign n45637 = n45636 ^ n45633 ^ 1'b0 ;
  assign n45638 = ( ~n16851 & n39033 ) | ( ~n16851 & n41613 ) | ( n39033 & n41613 ) ;
  assign n45639 = n1376 & n8530 ;
  assign n45640 = n3096 & ~n42979 ;
  assign n45641 = ~n13388 & n45640 ;
  assign n45642 = n45641 ^ n11630 ^ 1'b0 ;
  assign n45643 = n20085 & ~n35080 ;
  assign n45644 = n2525 & n45643 ;
  assign n45647 = n8656 & ~n11409 ;
  assign n45645 = n696 & ~n18433 ;
  assign n45646 = n45645 ^ n2216 ^ n564 ;
  assign n45648 = n45647 ^ n45646 ^ n16473 ;
  assign n45649 = n38686 ^ n33207 ^ 1'b0 ;
  assign n45650 = n4064 | n45649 ;
  assign n45651 = ( n16406 & n20791 ) | ( n16406 & ~n21803 ) | ( n20791 & ~n21803 ) ;
  assign n45652 = n8619 & ~n45651 ;
  assign n45653 = n22324 | n45652 ;
  assign n45654 = ~n3679 & n21073 ;
  assign n45655 = n39314 ^ n10227 ^ 1'b0 ;
  assign n45656 = n27553 ^ n9993 ^ n9818 ;
  assign n45657 = n20110 ^ n4974 ^ 1'b0 ;
  assign n45658 = ~n45656 & n45657 ;
  assign n45659 = ( n3666 & n15220 ) | ( n3666 & n19060 ) | ( n15220 & n19060 ) ;
  assign n45660 = n25949 ^ n13534 ^ 1'b0 ;
  assign n45661 = n2776 | n45660 ;
  assign n45662 = ( n24904 & ~n40667 ) | ( n24904 & n45661 ) | ( ~n40667 & n45661 ) ;
  assign n45663 = n20378 | n45662 ;
  assign n45664 = ( n1154 & n2397 ) | ( n1154 & ~n20446 ) | ( n2397 & ~n20446 ) ;
  assign n45665 = n2650 | n19911 ;
  assign n45666 = n63 & ~n45665 ;
  assign n45667 = n45666 ^ n40349 ^ 1'b0 ;
  assign n45668 = ( ~n3189 & n4688 ) | ( ~n3189 & n45667 ) | ( n4688 & n45667 ) ;
  assign n45669 = n45668 ^ n5562 ^ 1'b0 ;
  assign n45670 = n32150 ^ n22951 ^ n15428 ;
  assign n45671 = ~n6929 & n45670 ;
  assign n45672 = n45671 ^ n15670 ^ 1'b0 ;
  assign n45673 = n1734 & ~n2810 ;
  assign n45674 = n25208 & n45673 ;
  assign n45675 = ~n11920 & n25551 ;
  assign n45676 = ~n461 & n26510 ;
  assign n45677 = n45675 | n45676 ;
  assign n45678 = n10411 & n15166 ;
  assign n45679 = n5304 ^ n2222 ^ 1'b0 ;
  assign n45680 = n45678 & ~n45679 ;
  assign n45681 = n19476 | n20005 ;
  assign n45682 = n6444 & ~n45681 ;
  assign n45683 = n3381 | n45682 ;
  assign n45686 = n8876 & ~n26977 ;
  assign n45687 = n17493 & n45686 ;
  assign n45688 = n12310 & n45687 ;
  assign n45684 = n11692 & ~n17803 ;
  assign n45685 = ~n1412 & n45684 ;
  assign n45689 = n45688 ^ n45685 ^ 1'b0 ;
  assign n45690 = ~n3866 & n16092 ;
  assign n45691 = ~n5262 & n45690 ;
  assign n45692 = n12961 & n37122 ;
  assign n45693 = n4440 & n8512 ;
  assign n45694 = n45693 ^ n2114 ^ 1'b0 ;
  assign n45695 = n4638 & ~n5732 ;
  assign n45696 = n45694 & n45695 ;
  assign n45697 = ( n9296 & n28191 ) | ( n9296 & n45696 ) | ( n28191 & n45696 ) ;
  assign n45698 = n19491 ^ n13459 ^ 1'b0 ;
  assign n45699 = n45698 ^ n29638 ^ n19968 ;
  assign n45700 = n5229 ^ n878 ^ 1'b0 ;
  assign n45701 = n24345 | n45700 ;
  assign n45702 = n4646 & ~n45701 ;
  assign n45703 = n24418 & n28983 ;
  assign n45704 = n35136 ^ n1426 ^ 1'b0 ;
  assign n45705 = ~n30221 & n39256 ;
  assign n45706 = n24028 & ~n42771 ;
  assign n45707 = n45706 ^ n28006 ^ 1'b0 ;
  assign n45708 = n28380 ^ n633 ^ 1'b0 ;
  assign n45709 = n40033 & ~n45708 ;
  assign n45710 = ~n5520 & n16712 ;
  assign n45711 = n30593 & ~n45710 ;
  assign n45712 = n33723 | n45711 ;
  assign n45713 = n15582 & ~n45712 ;
  assign n45714 = n31047 ^ n15999 ^ 1'b0 ;
  assign n45715 = n4105 & ~n45714 ;
  assign n45716 = n583 & n7373 ;
  assign n45717 = ~n583 & n45716 ;
  assign n45718 = n7041 & ~n45717 ;
  assign n45719 = ~n45715 & n45718 ;
  assign n45720 = n45719 ^ n16417 ^ 1'b0 ;
  assign n45721 = ( n11009 & ~n17064 ) | ( n11009 & n27525 ) | ( ~n17064 & n27525 ) ;
  assign n45722 = ( n569 & ~n9236 ) | ( n569 & n45721 ) | ( ~n9236 & n45721 ) ;
  assign n45723 = n34965 ^ n17595 ^ n4422 ;
  assign n45724 = ~n44323 & n45723 ;
  assign n45725 = ~n15504 & n45724 ;
  assign n45726 = n13151 | n19098 ;
  assign n45727 = n113 | n45726 ;
  assign n45728 = ~n28731 & n44910 ;
  assign n45729 = n45728 ^ n1922 ^ 1'b0 ;
  assign n45730 = n17932 ^ n3159 ^ 1'b0 ;
  assign n45731 = ~n11306 & n31696 ;
  assign n45732 = ~n34756 & n45731 ;
  assign n45733 = n12955 ^ n2665 ^ 1'b0 ;
  assign n45734 = ~n5239 & n15100 ;
  assign n45735 = ~n15269 & n45734 ;
  assign n45736 = n26262 ^ n4516 ^ 1'b0 ;
  assign n45737 = ~n22357 & n45736 ;
  assign n45738 = n13138 & n45737 ;
  assign n45739 = n45735 & n45738 ;
  assign n45740 = n34965 | n45739 ;
  assign n45741 = n2449 & n15690 ;
  assign n45742 = ~n1695 & n22788 ;
  assign n45743 = ~n27623 & n45742 ;
  assign n45746 = n11387 ^ n7536 ^ 1'b0 ;
  assign n45747 = n11879 & n45746 ;
  assign n45748 = n12418 & n45747 ;
  assign n45744 = n10479 ^ n5862 ^ 1'b0 ;
  assign n45745 = n9054 & n45744 ;
  assign n45749 = n45748 ^ n45745 ^ 1'b0 ;
  assign n45750 = ~n12439 & n25141 ;
  assign n45751 = n13983 | n24562 ;
  assign n45752 = n36847 & ~n45751 ;
  assign n45753 = n4977 | n25969 ;
  assign n45754 = n45752 | n45753 ;
  assign n45755 = n45750 & ~n45754 ;
  assign n45756 = n22224 & ~n40184 ;
  assign n45757 = n10845 | n11560 ;
  assign n45758 = n20693 & ~n29801 ;
  assign n45759 = ~n7471 & n45758 ;
  assign n45760 = n29448 ^ n1009 ^ 1'b0 ;
  assign n45761 = ~n4544 & n45760 ;
  assign n45762 = n2118 & n21323 ;
  assign n45764 = ~n7574 & n11593 ;
  assign n45765 = n45764 ^ n28742 ^ 1'b0 ;
  assign n45763 = ~n2843 & n30782 ;
  assign n45766 = n45765 ^ n45763 ^ 1'b0 ;
  assign n45767 = n23306 & ~n45766 ;
  assign n45768 = ~n45762 & n45767 ;
  assign n45769 = n42371 ^ n9454 ^ 1'b0 ;
  assign n45770 = n16852 & n20740 ;
  assign n45771 = ( n82 & n9918 ) | ( n82 & ~n45770 ) | ( n9918 & ~n45770 ) ;
  assign n45772 = ( n14508 & n30725 ) | ( n14508 & n45771 ) | ( n30725 & n45771 ) ;
  assign n45773 = n10822 & ~n30812 ;
  assign n45774 = n34525 & n45773 ;
  assign n45775 = ( ~n20350 & n22118 ) | ( ~n20350 & n34201 ) | ( n22118 & n34201 ) ;
  assign n45776 = n34705 ^ n29559 ^ n4140 ;
  assign n45777 = n2039 & ~n14385 ;
  assign n45778 = n150 & n45777 ;
  assign n45779 = n17936 & ~n45407 ;
  assign n45780 = ~n45778 & n45779 ;
  assign n45781 = n25192 ^ n17938 ^ 1'b0 ;
  assign n45782 = n25976 | n45781 ;
  assign n45783 = n993 & ~n45782 ;
  assign n45784 = n14624 & n45783 ;
  assign n45785 = n27595 ^ n23005 ^ n645 ;
  assign n45786 = n12418 | n45785 ;
  assign n45787 = n22013 & ~n45786 ;
  assign n45788 = n31715 ^ n8314 ^ 1'b0 ;
  assign n45789 = n45787 & ~n45788 ;
  assign n45797 = n4681 & n9314 ;
  assign n45790 = ~n2128 & n9758 ;
  assign n45791 = n45790 ^ n4810 ^ 1'b0 ;
  assign n45792 = n989 & n11904 ;
  assign n45793 = n45792 ^ n30904 ^ 1'b0 ;
  assign n45794 = n45791 | n45793 ;
  assign n45795 = n9286 | n45794 ;
  assign n45796 = n7188 | n45795 ;
  assign n45798 = n45797 ^ n45796 ^ 1'b0 ;
  assign n45799 = n45798 ^ n1718 ^ 1'b0 ;
  assign n45803 = n18025 & n28826 ;
  assign n45801 = n15562 ^ n5730 ^ 1'b0 ;
  assign n45800 = n1143 & ~n43558 ;
  assign n45802 = n45801 ^ n45800 ^ 1'b0 ;
  assign n45804 = n45803 ^ n45802 ^ n13256 ;
  assign n45805 = ( n7641 & n12323 ) | ( n7641 & ~n28090 ) | ( n12323 & ~n28090 ) ;
  assign n45806 = ( ~n18987 & n31459 ) | ( ~n18987 & n45805 ) | ( n31459 & n45805 ) ;
  assign n45807 = n24207 ^ n19909 ^ n5599 ;
  assign n45808 = n7848 | n11171 ;
  assign n45809 = n16550 & n45808 ;
  assign n45810 = ~n3736 & n45809 ;
  assign n45811 = n45807 & n45810 ;
  assign n45812 = n8236 & ~n16288 ;
  assign n45813 = n25545 ^ n24809 ^ n5754 ;
  assign n45814 = ( ~n4640 & n15263 ) | ( ~n4640 & n29107 ) | ( n15263 & n29107 ) ;
  assign n45815 = n45814 ^ n40602 ^ 1'b0 ;
  assign n45816 = n45813 & ~n45815 ;
  assign n45817 = n230 & n45816 ;
  assign n45818 = n24041 ^ n15516 ^ n903 ;
  assign n45819 = n45818 ^ n5266 ^ 1'b0 ;
  assign n45820 = ( ~n11827 & n18110 ) | ( ~n11827 & n31904 ) | ( n18110 & n31904 ) ;
  assign n45821 = n9309 & ~n18822 ;
  assign n45822 = n29488 ^ n23796 ^ 1'b0 ;
  assign n45823 = n20361 & n45822 ;
  assign n45824 = n12556 | n28839 ;
  assign n45825 = n45824 ^ n3441 ^ 1'b0 ;
  assign n45826 = n23718 | n45825 ;
  assign n45827 = ( n5891 & n7963 ) | ( n5891 & ~n13265 ) | ( n7963 & ~n13265 ) ;
  assign n45828 = n11769 ^ n628 ^ 1'b0 ;
  assign n45829 = n13513 & n45828 ;
  assign n45830 = n3040 & n45829 ;
  assign n45831 = ~n3111 & n25251 ;
  assign n45832 = n13161 ^ n5227 ^ 1'b0 ;
  assign n45833 = n1937 & ~n20033 ;
  assign n45834 = ~n45832 & n45833 ;
  assign n45835 = n16327 ^ n11880 ^ 1'b0 ;
  assign n45836 = n25296 ^ n18361 ^ 1'b0 ;
  assign n45837 = n30513 ^ n14054 ^ 1'b0 ;
  assign n45838 = n2395 & ~n26589 ;
  assign n45839 = n45838 ^ n364 ^ 1'b0 ;
  assign n45840 = n27697 ^ n20366 ^ 1'b0 ;
  assign n45841 = ~n12264 & n45840 ;
  assign n45842 = ~n33553 & n45841 ;
  assign n45843 = ~n9588 & n23106 ;
  assign n45844 = n18510 ^ n17334 ^ 1'b0 ;
  assign n45845 = n5220 | n7741 ;
  assign n45846 = n11057 & n45845 ;
  assign n45847 = n45846 ^ n19952 ^ 1'b0 ;
  assign n45848 = n45847 ^ n45341 ^ n42552 ;
  assign n45849 = n45848 ^ n17505 ^ 1'b0 ;
  assign n45850 = n33430 ^ n19210 ^ 1'b0 ;
  assign n45851 = n22085 & ~n45850 ;
  assign n45852 = n2752 | n20679 ;
  assign n45853 = n23392 ^ n6987 ^ 1'b0 ;
  assign n45854 = n15544 ^ n14698 ^ 1'b0 ;
  assign n45855 = ~n30723 & n45854 ;
  assign n45856 = n45855 ^ n11347 ^ 1'b0 ;
  assign n45857 = n26360 ^ n16327 ^ 1'b0 ;
  assign n45858 = n18373 & ~n45857 ;
  assign n45859 = n6357 ^ n6226 ^ 1'b0 ;
  assign n45860 = n698 | n45859 ;
  assign n45861 = n45860 ^ n18586 ^ 1'b0 ;
  assign n45862 = n4249 & n43889 ;
  assign n45863 = n27100 ^ n20513 ^ n17407 ;
  assign n45864 = n1214 & n14505 ;
  assign n45865 = ( n6759 & n8859 ) | ( n6759 & n45864 ) | ( n8859 & n45864 ) ;
  assign n45866 = n30072 ^ n1623 ^ 1'b0 ;
  assign n45867 = n28887 ^ n8849 ^ 1'b0 ;
  assign n45868 = n7440 | n21858 ;
  assign n45869 = n18711 ^ n4240 ^ 1'b0 ;
  assign n45870 = n12856 & n39546 ;
  assign n45871 = n2067 | n5955 ;
  assign n45872 = n45871 ^ n24395 ^ 1'b0 ;
  assign n45873 = n12328 & n45872 ;
  assign n45874 = n34129 & ~n45873 ;
  assign n45875 = ~n14452 & n43220 ;
  assign n45876 = n2443 & n12140 ;
  assign n45877 = n12558 & ~n13511 ;
  assign n45878 = ~n11143 & n28285 ;
  assign n45879 = n21297 ^ n6676 ^ 1'b0 ;
  assign n45880 = ~n38265 & n45879 ;
  assign n45881 = n29559 ^ n23149 ^ 1'b0 ;
  assign n45882 = ~n45880 & n45881 ;
  assign n45883 = n29448 ^ n21146 ^ n14715 ;
  assign n45884 = ~n21688 & n45883 ;
  assign n45885 = n32750 ^ n24234 ^ n216 ;
  assign n45886 = n6602 & ~n25676 ;
  assign n45887 = ~n7065 & n29426 ;
  assign n45888 = n45887 ^ n27285 ^ 1'b0 ;
  assign n45889 = n34734 ^ n31676 ^ 1'b0 ;
  assign n45890 = n27583 & ~n32324 ;
  assign n45891 = n8018 & n9894 ;
  assign n45892 = n45891 ^ n45829 ^ 1'b0 ;
  assign n45893 = n32237 & ~n45892 ;
  assign n45894 = n36037 ^ n9216 ^ 1'b0 ;
  assign n45895 = n39158 & ~n45894 ;
  assign n45896 = ~n9078 & n20517 ;
  assign n45897 = ~n8828 & n45896 ;
  assign n45898 = n4495 & n23959 ;
  assign n45899 = n45897 & n45898 ;
  assign n45900 = n10690 | n17640 ;
  assign n45901 = n45900 ^ n32262 ^ 1'b0 ;
  assign n45902 = n24889 ^ n9773 ^ 1'b0 ;
  assign n45903 = n19176 | n45902 ;
  assign n45904 = n1495 & n3645 ;
  assign n45905 = n45904 ^ n18555 ^ 1'b0 ;
  assign n45906 = ~n1105 & n23578 ;
  assign n45907 = n45905 & n45906 ;
  assign n45908 = n27024 ^ n13334 ^ 1'b0 ;
  assign n45910 = ~n3918 & n4888 ;
  assign n45911 = n45910 ^ n4122 ^ 1'b0 ;
  assign n45909 = n2561 | n15943 ;
  assign n45912 = n45911 ^ n45909 ^ 1'b0 ;
  assign n45913 = n21844 ^ n11247 ^ 1'b0 ;
  assign n45914 = n9417 ^ n2810 ^ 1'b0 ;
  assign n45915 = n4622 & ~n43496 ;
  assign n45916 = n951 | n4339 ;
  assign n45917 = n45916 ^ n31979 ^ n12366 ;
  assign n45918 = n45915 & ~n45917 ;
  assign n45919 = ~n4686 & n14010 ;
  assign n45922 = n24518 ^ n21865 ^ 1'b0 ;
  assign n45921 = n1082 & n24468 ;
  assign n45923 = n45922 ^ n45921 ^ 1'b0 ;
  assign n45924 = n12701 | n35447 ;
  assign n45925 = n45923 | n45924 ;
  assign n45926 = n35441 & n45925 ;
  assign n45927 = ~n16637 & n45926 ;
  assign n45920 = n879 | n40788 ;
  assign n45928 = n45927 ^ n45920 ^ 1'b0 ;
  assign n45929 = n32457 ^ n13169 ^ n9619 ;
  assign n45932 = n998 | n3971 ;
  assign n45930 = n19510 & n19778 ;
  assign n45931 = n38976 & ~n45930 ;
  assign n45933 = n45932 ^ n45931 ^ 1'b0 ;
  assign n45934 = ~n2176 & n4405 ;
  assign n45935 = n24936 ^ n21543 ^ 1'b0 ;
  assign n45936 = n45934 | n45935 ;
  assign n45937 = n600 & n12286 ;
  assign n45938 = n6996 & n45937 ;
  assign n45939 = n45938 ^ n3926 ^ 1'b0 ;
  assign n45940 = n18592 | n45939 ;
  assign n45941 = n3461 | n9430 ;
  assign n45942 = n26410 ^ n24131 ^ n1931 ;
  assign n45943 = n12668 | n45702 ;
  assign n45944 = n9033 & ~n45943 ;
  assign n45945 = n45944 ^ n42430 ^ n9832 ;
  assign n45946 = n40051 ^ n17951 ^ 1'b0 ;
  assign n45947 = ~n12330 & n29621 ;
  assign n45948 = n13846 & ~n41474 ;
  assign n45949 = n11716 | n25383 ;
  assign n45950 = n13113 & ~n45949 ;
  assign n45951 = n4138 & ~n17513 ;
  assign n45952 = ~n654 & n45951 ;
  assign n45953 = n31172 | n45952 ;
  assign n45954 = n45953 ^ n15459 ^ 1'b0 ;
  assign n45955 = ( ~n80 & n10490 ) | ( ~n80 & n37350 ) | ( n10490 & n37350 ) ;
  assign n45956 = n14790 & n45955 ;
  assign n45957 = n45956 ^ n31674 ^ 1'b0 ;
  assign n45958 = n38894 ^ n11729 ^ 1'b0 ;
  assign n45959 = n22355 & ~n45958 ;
  assign n45960 = n45959 ^ n23457 ^ 1'b0 ;
  assign n45961 = n45960 ^ n44580 ^ n14315 ;
  assign n45963 = n27851 ^ n23861 ^ 1'b0 ;
  assign n45962 = ( n870 & ~n5536 ) | ( n870 & n11229 ) | ( ~n5536 & n11229 ) ;
  assign n45964 = n45963 ^ n45962 ^ 1'b0 ;
  assign n45965 = n4186 & n7736 ;
  assign n45966 = ( n3578 & n25123 ) | ( n3578 & n30756 ) | ( n25123 & n30756 ) ;
  assign n45969 = n19237 | n25565 ;
  assign n45968 = n652 & ~n21718 ;
  assign n45970 = n45969 ^ n45968 ^ 1'b0 ;
  assign n45967 = n27340 ^ n4657 ^ 1'b0 ;
  assign n45971 = n45970 ^ n45967 ^ 1'b0 ;
  assign n45972 = n2218 | n45971 ;
  assign n45973 = ( ~n45965 & n45966 ) | ( ~n45965 & n45972 ) | ( n45966 & n45972 ) ;
  assign n45974 = n24831 ^ n14993 ^ 1'b0 ;
  assign n45975 = n17323 & n45974 ;
  assign n45976 = n8594 | n8678 ;
  assign n45977 = n22092 & ~n45976 ;
  assign n45978 = ~n45975 & n45977 ;
  assign n45979 = n27003 ^ n22380 ^ 1'b0 ;
  assign n45980 = n16807 & ~n45979 ;
  assign n45981 = n45980 ^ n12477 ^ 1'b0 ;
  assign n45982 = ~n24354 & n26775 ;
  assign n45983 = n28780 & ~n45982 ;
  assign n45984 = n45983 ^ n31984 ^ 1'b0 ;
  assign n45985 = n26243 ^ n9029 ^ 1'b0 ;
  assign n45986 = n2621 | n29685 ;
  assign n45987 = n4345 | n45986 ;
  assign n45988 = n13670 ^ n4508 ^ 1'b0 ;
  assign n45989 = ~n6008 & n45988 ;
  assign n45990 = n8115 & n45989 ;
  assign n45991 = n45990 ^ n3840 ^ 1'b0 ;
  assign n45992 = ( n4536 & n7153 ) | ( n4536 & ~n45991 ) | ( n7153 & ~n45991 ) ;
  assign n45993 = n7791 ^ n7261 ^ 1'b0 ;
  assign n45994 = n11442 & n45993 ;
  assign n45995 = ( n37 & ~n45992 ) | ( n37 & n45994 ) | ( ~n45992 & n45994 ) ;
  assign n45996 = n34627 ^ n25631 ^ n11844 ;
  assign n45997 = n11577 ^ n4071 ^ 1'b0 ;
  assign n45998 = n25690 & ~n45997 ;
  assign n45999 = n25829 & n45998 ;
  assign n46000 = n26910 & ~n38235 ;
  assign n46001 = n23479 & ~n33084 ;
  assign n46002 = n24432 ^ n15509 ^ n1944 ;
  assign n46003 = n11366 & n20649 ;
  assign n46004 = n11040 & n46003 ;
  assign n46008 = n30758 ^ n3446 ^ n780 ;
  assign n46009 = n35420 | n46008 ;
  assign n46010 = n46009 ^ n9892 ^ 1'b0 ;
  assign n46005 = ~n953 & n6384 ;
  assign n46006 = n20068 | n28627 ;
  assign n46007 = n46005 | n46006 ;
  assign n46011 = n46010 ^ n46007 ^ 1'b0 ;
  assign n46012 = n11076 & n43634 ;
  assign n46013 = n46012 ^ n40773 ^ 1'b0 ;
  assign n46014 = n9568 & ~n46013 ;
  assign n46015 = n46014 ^ n11295 ^ 1'b0 ;
  assign n46016 = n4216 ^ n2650 ^ n1316 ;
  assign n46017 = n8970 | n46016 ;
  assign n46018 = n2314 | n46017 ;
  assign n46019 = n9903 | n46018 ;
  assign n46020 = n21181 ^ n5123 ^ 1'b0 ;
  assign n46021 = n46019 & n46020 ;
  assign n46022 = n1435 | n7167 ;
  assign n46023 = ~n3259 & n6638 ;
  assign n46024 = ~n1565 & n46023 ;
  assign n46025 = n45792 ^ n7482 ^ 1'b0 ;
  assign n46026 = n46024 | n46025 ;
  assign n46027 = ( n976 & n23139 ) | ( n976 & ~n46026 ) | ( n23139 & ~n46026 ) ;
  assign n46028 = n46027 ^ n28924 ^ 1'b0 ;
  assign n46029 = n35868 ^ n9566 ^ 1'b0 ;
  assign n46030 = n12292 & n46029 ;
  assign n46031 = n19140 ^ n16710 ^ 1'b0 ;
  assign n46032 = n1245 & n46031 ;
  assign n46033 = n42701 ^ n7026 ^ 1'b0 ;
  assign n46034 = ~n26001 & n27533 ;
  assign n46035 = ~n6717 & n46034 ;
  assign n46036 = n44873 ^ n7289 ^ 1'b0 ;
  assign n46037 = ~n46035 & n46036 ;
  assign n46038 = n3460 & ~n11691 ;
  assign n46039 = n42817 ^ n28879 ^ 1'b0 ;
  assign n46040 = n34770 | n46039 ;
  assign n46041 = n2820 & n3246 ;
  assign n46042 = n13267 & ~n46041 ;
  assign n46043 = n46042 ^ n40673 ^ 1'b0 ;
  assign n46044 = n944 | n17801 ;
  assign n46045 = n46044 ^ n13220 ^ 1'b0 ;
  assign n46046 = ~n10053 & n46045 ;
  assign n46047 = n46046 ^ n25998 ^ 1'b0 ;
  assign n46048 = n23922 ^ n4704 ^ 1'b0 ;
  assign n46049 = n18571 & n46048 ;
  assign n46050 = n46049 ^ n26948 ^ n16745 ;
  assign n46051 = n25067 ^ n18514 ^ n14386 ;
  assign n46052 = n376 & n8043 ;
  assign n46053 = n32026 | n46052 ;
  assign n46054 = n3231 | n46053 ;
  assign n46055 = ( n4000 & ~n6473 ) | ( n4000 & n30483 ) | ( ~n6473 & n30483 ) ;
  assign n46056 = n19155 & ~n46055 ;
  assign n46057 = n19562 ^ n17110 ^ n10971 ;
  assign n46058 = n3441 ^ n713 ^ 1'b0 ;
  assign n46059 = n25406 | n46058 ;
  assign n46060 = ~n46057 & n46059 ;
  assign n46061 = n6842 & ~n15102 ;
  assign n46062 = n46061 ^ n1000 ^ 1'b0 ;
  assign n46063 = n9599 ^ n1805 ^ 1'b0 ;
  assign n46064 = n37495 & ~n46063 ;
  assign n46065 = n25100 ^ n12349 ^ n5098 ;
  assign n46066 = n46065 ^ n45428 ^ n24531 ;
  assign n46067 = ~n11355 & n18994 ;
  assign n46068 = ~n46066 & n46067 ;
  assign n46069 = ~n5396 & n8070 ;
  assign n46070 = ~n15123 & n24959 ;
  assign n46071 = n18679 ^ n2635 ^ 1'b0 ;
  assign n46072 = n46071 ^ n30862 ^ 1'b0 ;
  assign n46073 = n46072 ^ n22612 ^ n2813 ;
  assign n46074 = n42301 ^ n11633 ^ 1'b0 ;
  assign n46075 = n7255 & ~n29363 ;
  assign n46076 = n46075 ^ n12443 ^ 1'b0 ;
  assign n46077 = n24041 ^ n13579 ^ n11982 ;
  assign n46078 = ( ~n19305 & n38310 ) | ( ~n19305 & n46077 ) | ( n38310 & n46077 ) ;
  assign n46079 = ( n6181 & n13502 ) | ( n6181 & n42837 ) | ( n13502 & n42837 ) ;
  assign n46080 = ( n816 & n861 ) | ( n816 & ~n46079 ) | ( n861 & ~n46079 ) ;
  assign n46081 = n42273 | n46080 ;
  assign n46082 = ( n12277 & ~n13917 ) | ( n12277 & n46081 ) | ( ~n13917 & n46081 ) ;
  assign n46083 = n22528 ^ n8625 ^ n473 ;
  assign n46084 = n15426 & n22783 ;
  assign n46085 = n46084 ^ n3447 ^ 1'b0 ;
  assign n46086 = ~n8647 & n46085 ;
  assign n46087 = n24569 ^ n10459 ^ 1'b0 ;
  assign n46088 = n26409 & ~n46087 ;
  assign n46092 = ~n38479 & n40659 ;
  assign n46093 = n5256 & n46092 ;
  assign n46089 = n15470 & n45165 ;
  assign n46090 = ~n20772 & n46089 ;
  assign n46091 = n31507 | n46090 ;
  assign n46094 = n46093 ^ n46091 ^ 1'b0 ;
  assign n46095 = ~n4204 & n45861 ;
  assign n46096 = ~n8967 & n15970 ;
  assign n46097 = n31932 ^ n30357 ^ 1'b0 ;
  assign n46098 = n22292 & n46097 ;
  assign n46099 = n41316 ^ n19473 ^ 1'b0 ;
  assign n46100 = n20811 & n46099 ;
  assign n46101 = n7763 & n24277 ;
  assign n46102 = n21849 & n46101 ;
  assign n46103 = n3855 | n17913 ;
  assign n46104 = n46102 & ~n46103 ;
  assign n46105 = ( n9606 & n46100 ) | ( n9606 & ~n46104 ) | ( n46100 & ~n46104 ) ;
  assign n46106 = ( n24370 & ~n37997 ) | ( n24370 & n46105 ) | ( ~n37997 & n46105 ) ;
  assign n46107 = n3789 & ~n12499 ;
  assign n46108 = n7268 & ~n25560 ;
  assign n46109 = n46108 ^ n39038 ^ n14023 ;
  assign n46110 = n46107 & n46109 ;
  assign n46111 = ~n9346 & n45809 ;
  assign n46112 = n26929 ^ n11850 ^ 1'b0 ;
  assign n46113 = ~n3575 & n7434 ;
  assign n46114 = ( ~n25523 & n31455 ) | ( ~n25523 & n46113 ) | ( n31455 & n46113 ) ;
  assign n46115 = n46114 ^ n19383 ^ 1'b0 ;
  assign n46116 = n45271 ^ n41475 ^ n150 ;
  assign n46117 = n40425 | n44446 ;
  assign n46118 = n46117 ^ n20396 ^ 1'b0 ;
  assign n46119 = n25289 & ~n29841 ;
  assign n46120 = n6142 & n36300 ;
  assign n46121 = n46120 ^ n3209 ^ 1'b0 ;
  assign n46122 = n39572 ^ n1890 ^ 1'b0 ;
  assign n46123 = n39262 ^ n24278 ^ 1'b0 ;
  assign n46124 = n40181 & ~n44995 ;
  assign n46125 = ~n2461 & n46124 ;
  assign n46126 = n12578 & n13388 ;
  assign n46127 = n46126 ^ n24968 ^ 1'b0 ;
  assign n46128 = n13197 ^ n1279 ^ 1'b0 ;
  assign n46129 = n6687 | n10093 ;
  assign n46130 = n46129 ^ n34645 ^ 1'b0 ;
  assign n46131 = n42437 ^ n36112 ^ 1'b0 ;
  assign n46132 = n31712 ^ n18316 ^ 1'b0 ;
  assign n46133 = ~n46131 & n46132 ;
  assign n46134 = n28837 ^ n2952 ^ 1'b0 ;
  assign n46135 = ~n12249 & n46134 ;
  assign n46136 = n38467 ^ n3376 ^ 1'b0 ;
  assign n46137 = n31130 ^ n9275 ^ 1'b0 ;
  assign n46138 = n45569 ^ n221 ^ 1'b0 ;
  assign n46139 = n28670 ^ n11949 ^ 1'b0 ;
  assign n46140 = n6648 | n33154 ;
  assign n46141 = n1832 & n46140 ;
  assign n46142 = n46139 & n46141 ;
  assign n46143 = n38841 ^ n17820 ^ n4396 ;
  assign n46144 = ( n1979 & ~n6438 ) | ( n1979 & n9791 ) | ( ~n6438 & n9791 ) ;
  assign n46145 = n8077 ^ n3736 ^ 1'b0 ;
  assign n46146 = n20491 & ~n46145 ;
  assign n46147 = n46146 ^ n12569 ^ 1'b0 ;
  assign n46148 = n5637 | n20654 ;
  assign n46149 = n32982 ^ n948 ^ 1'b0 ;
  assign n46150 = n36508 & n46149 ;
  assign n46151 = n46150 ^ n7273 ^ 1'b0 ;
  assign n46152 = n19195 & ~n36417 ;
  assign n46153 = n32845 & n46152 ;
  assign n46154 = n6702 | n12710 ;
  assign n46155 = n18894 | n27347 ;
  assign n46156 = n46154 & ~n46155 ;
  assign n46157 = n24271 & ~n29448 ;
  assign n46158 = n46156 & n46157 ;
  assign n46159 = n46153 & ~n46158 ;
  assign n46160 = n4252 & ~n16130 ;
  assign n46161 = ( n628 & n37068 ) | ( n628 & n46160 ) | ( n37068 & n46160 ) ;
  assign n46162 = n46161 ^ n2609 ^ 1'b0 ;
  assign n46163 = n35254 ^ n12004 ^ 1'b0 ;
  assign n46164 = n44292 & ~n46163 ;
  assign n46165 = n46164 ^ n24819 ^ 1'b0 ;
  assign n46166 = n18463 & n46165 ;
  assign n46167 = n17854 ^ n12849 ^ n4217 ;
  assign n46168 = n46167 ^ n4088 ^ 1'b0 ;
  assign n46169 = ~n3696 & n34005 ;
  assign n46170 = n46169 ^ n16557 ^ 1'b0 ;
  assign n46171 = n46170 ^ n2278 ^ 1'b0 ;
  assign n46172 = n7049 & ~n41171 ;
  assign n46173 = ~n597 & n19523 ;
  assign n46174 = ~n23294 & n46173 ;
  assign n46175 = ~n14148 & n31360 ;
  assign n46176 = n4257 & n46175 ;
  assign n46177 = n11062 & ~n36562 ;
  assign n46178 = ~n18590 & n45972 ;
  assign n46179 = n25823 & n28301 ;
  assign n46180 = ~n2440 & n24453 ;
  assign n46181 = n46180 ^ n25477 ^ 1'b0 ;
  assign n46182 = n890 ^ n691 ^ 1'b0 ;
  assign n46183 = ~n7402 & n46182 ;
  assign n46184 = n32992 ^ n31343 ^ 1'b0 ;
  assign n46185 = ~n9770 & n46184 ;
  assign n46194 = n3614 & n3645 ;
  assign n46195 = ~n3645 & n46194 ;
  assign n46196 = n2283 | n46195 ;
  assign n46197 = n2283 & ~n46196 ;
  assign n46198 = n101 & ~n46197 ;
  assign n46199 = ~n101 & n46198 ;
  assign n46200 = n46199 ^ n8242 ^ 1'b0 ;
  assign n46188 = n8884 & n41296 ;
  assign n46189 = ~n41296 & n46188 ;
  assign n46190 = n772 & n3084 ;
  assign n46191 = ~n3084 & n46190 ;
  assign n46192 = n46191 ^ n16625 ^ 1'b0 ;
  assign n46193 = n46189 | n46192 ;
  assign n46186 = ~n8426 & n11137 ;
  assign n46187 = n46186 ^ n9685 ^ 1'b0 ;
  assign n46201 = n46200 ^ n46193 ^ n46187 ;
  assign n46202 = n45128 ^ n40776 ^ 1'b0 ;
  assign n46203 = n6683 ^ n6161 ^ 1'b0 ;
  assign n46204 = ~n46202 & n46203 ;
  assign n46205 = ~n7807 & n17768 ;
  assign n46206 = n32142 | n32809 ;
  assign n46207 = ~n14764 & n20681 ;
  assign n46208 = n8960 & n46207 ;
  assign n46209 = n2815 & n24348 ;
  assign n46210 = ( n46206 & ~n46208 ) | ( n46206 & n46209 ) | ( ~n46208 & n46209 ) ;
  assign n46211 = n11188 | n43858 ;
  assign n46212 = n15884 ^ n4216 ^ 1'b0 ;
  assign n46213 = n2412 & n33749 ;
  assign n46214 = n46213 ^ n3912 ^ 1'b0 ;
  assign n46215 = ( ~n4536 & n9787 ) | ( ~n4536 & n18522 ) | ( n9787 & n18522 ) ;
  assign n46216 = ( n5212 & n15142 ) | ( n5212 & n32886 ) | ( n15142 & n32886 ) ;
  assign n46217 = n46215 | n46216 ;
  assign n46218 = n46217 ^ n23302 ^ 1'b0 ;
  assign n46219 = ( n12346 & ~n22831 ) | ( n12346 & n30597 ) | ( ~n22831 & n30597 ) ;
  assign n46220 = ( n321 & n879 ) | ( n321 & ~n2449 ) | ( n879 & ~n2449 ) ;
  assign n46221 = ( n1249 & n17942 ) | ( n1249 & ~n46220 ) | ( n17942 & ~n46220 ) ;
  assign n46223 = ~n4446 & n35334 ;
  assign n46224 = n46223 ^ n14523 ^ 1'b0 ;
  assign n46225 = ( n17493 & n30450 ) | ( n17493 & ~n46224 ) | ( n30450 & ~n46224 ) ;
  assign n46222 = n7854 & n36613 ;
  assign n46226 = n46225 ^ n46222 ^ 1'b0 ;
  assign n46227 = ~n36011 & n43942 ;
  assign n46228 = n6657 & n16381 ;
  assign n46229 = n21856 | n31661 ;
  assign n46230 = n8467 | n46229 ;
  assign n46231 = ( n31351 & n32584 ) | ( n31351 & ~n46230 ) | ( n32584 & ~n46230 ) ;
  assign n46232 = n224 & n46017 ;
  assign n46233 = ~n608 & n27499 ;
  assign n46234 = n46233 ^ n10240 ^ 1'b0 ;
  assign n46235 = n32953 ^ n14189 ^ 1'b0 ;
  assign n46236 = ~n16791 & n46235 ;
  assign n46237 = n13694 | n20415 ;
  assign n46238 = n15020 & ~n44242 ;
  assign n46239 = n20876 & n46238 ;
  assign n46240 = ( n13356 & n15651 ) | ( n13356 & ~n27317 ) | ( n15651 & ~n27317 ) ;
  assign n46241 = ( n6528 & ~n10850 ) | ( n6528 & n46240 ) | ( ~n10850 & n46240 ) ;
  assign n46242 = n32565 ^ n7707 ^ n2794 ;
  assign n46243 = n28350 ^ n2579 ^ 1'b0 ;
  assign n46244 = n12282 & n46243 ;
  assign n46245 = n1230 & n46244 ;
  assign n46246 = n46245 ^ n12479 ^ 1'b0 ;
  assign n46247 = n17168 | n30141 ;
  assign n46248 = n46247 ^ n33582 ^ 1'b0 ;
  assign n46249 = n10012 & ~n46248 ;
  assign n46250 = ~n17180 & n43443 ;
  assign n46251 = n46249 & n46250 ;
  assign n46252 = n3985 | n20496 ;
  assign n46253 = ~n3054 & n46252 ;
  assign n46254 = n46251 & n46253 ;
  assign n46255 = n2885 | n29024 ;
  assign n46256 = n505 | n46255 ;
  assign n46257 = n19558 ^ n5315 ^ 1'b0 ;
  assign n46258 = n19497 ^ n15940 ^ 1'b0 ;
  assign n46259 = ( n1241 & ~n39267 ) | ( n1241 & n46258 ) | ( ~n39267 & n46258 ) ;
  assign n46260 = n17100 | n24703 ;
  assign n46261 = ~n23582 & n46260 ;
  assign n46262 = ~n29582 & n34476 ;
  assign n46263 = n46262 ^ n29321 ^ 1'b0 ;
  assign n46264 = n43133 & ~n46263 ;
  assign n46265 = n2704 & n27118 ;
  assign n46266 = n31159 ^ n6574 ^ 1'b0 ;
  assign n46267 = n4900 | n46266 ;
  assign n46268 = n19962 ^ n2802 ^ 1'b0 ;
  assign n46269 = ~n17173 & n46268 ;
  assign n46271 = n11534 & ~n43080 ;
  assign n46270 = n39235 ^ n19658 ^ 1'b0 ;
  assign n46272 = n46271 ^ n46270 ^ n6895 ;
  assign n46273 = n8476 & n22508 ;
  assign n46274 = n46273 ^ n3081 ^ 1'b0 ;
  assign n46275 = ~n11870 & n42121 ;
  assign n46276 = ~n14570 & n46275 ;
  assign n46279 = n2304 | n13444 ;
  assign n46280 = n4918 & ~n46279 ;
  assign n46277 = ( n9173 & ~n12234 ) | ( n9173 & n24794 ) | ( ~n12234 & n24794 ) ;
  assign n46278 = n46277 ^ n29363 ^ 1'b0 ;
  assign n46281 = n46280 ^ n46278 ^ 1'b0 ;
  assign n46282 = ~n18966 & n46281 ;
  assign n46283 = ~n8356 & n46282 ;
  assign n46284 = n46283 ^ n12369 ^ 1'b0 ;
  assign n46285 = n23836 ^ n2054 ^ 1'b0 ;
  assign n46286 = n15086 & n20686 ;
  assign n46287 = n46286 ^ n3125 ^ 1'b0 ;
  assign n46288 = n7154 | n12255 ;
  assign n46289 = ( n2617 & n6352 ) | ( n2617 & n17450 ) | ( n6352 & n17450 ) ;
  assign n46290 = n46289 ^ n15879 ^ 1'b0 ;
  assign n46291 = n46288 | n46290 ;
  assign n46292 = ~n26918 & n39271 ;
  assign n46293 = ( n177 & ~n8980 ) | ( n177 & n39380 ) | ( ~n8980 & n39380 ) ;
  assign n46294 = ( n3690 & ~n4969 ) | ( n3690 & n25885 ) | ( ~n4969 & n25885 ) ;
  assign n46295 = n46294 ^ n11880 ^ 1'b0 ;
  assign n46296 = n32643 | n46295 ;
  assign n46297 = n46293 | n46296 ;
  assign n46298 = n16093 & ~n41353 ;
  assign n46299 = n46298 ^ n10124 ^ 1'b0 ;
  assign n46300 = n5113 ^ n2720 ^ 1'b0 ;
  assign n46301 = n3656 & n46300 ;
  assign n46302 = ~n672 & n13754 ;
  assign n46303 = ~n7728 & n46302 ;
  assign n46304 = n3578 | n46303 ;
  assign n46305 = n25343 | n35457 ;
  assign n46306 = n24165 & n46305 ;
  assign n46310 = n33974 & ~n40694 ;
  assign n46311 = n1081 & n46310 ;
  assign n46307 = n35099 ^ n20191 ^ 1'b0 ;
  assign n46308 = n41599 ^ n3089 ^ 1'b0 ;
  assign n46309 = n46307 & n46308 ;
  assign n46312 = n46311 ^ n46309 ^ 1'b0 ;
  assign n46313 = n13679 | n46312 ;
  assign n46314 = n6296 | n18519 ;
  assign n46315 = n13960 & ~n46314 ;
  assign n46316 = n23359 ^ n10453 ^ 1'b0 ;
  assign n46317 = n14493 | n46316 ;
  assign n46318 = n36189 & ~n46317 ;
  assign n46319 = n46318 ^ n44175 ^ 1'b0 ;
  assign n46320 = n4104 & ~n46319 ;
  assign n46321 = n46320 ^ n26884 ^ 1'b0 ;
  assign n46322 = n7269 & n18539 ;
  assign n46323 = n46322 ^ n43756 ^ 1'b0 ;
  assign n46325 = ~n12442 & n15595 ;
  assign n46326 = n7610 & n46325 ;
  assign n46324 = n7240 ^ n5464 ^ 1'b0 ;
  assign n46327 = n46326 ^ n46324 ^ n242 ;
  assign n46328 = ( n16305 & ~n20950 ) | ( n16305 & n46327 ) | ( ~n20950 & n46327 ) ;
  assign n46329 = n46328 ^ n37068 ^ 1'b0 ;
  assign n46330 = n8030 | n19616 ;
  assign n46331 = ~n27556 & n39182 ;
  assign n46336 = ~n200 & n2888 ;
  assign n46337 = n46336 ^ n8950 ^ 1'b0 ;
  assign n46338 = ~n2857 & n46337 ;
  assign n46339 = n890 & n46338 ;
  assign n46334 = ( ~n6770 & n11594 ) | ( ~n6770 & n44251 ) | ( n11594 & n44251 ) ;
  assign n46333 = n13387 ^ n2470 ^ 1'b0 ;
  assign n46335 = n46334 ^ n46333 ^ n514 ;
  assign n46332 = n11231 ^ n7051 ^ 1'b0 ;
  assign n46340 = n46339 ^ n46335 ^ n46332 ;
  assign n46341 = ~n3730 & n13113 ;
  assign n46342 = n5915 & ~n46341 ;
  assign n46343 = n46342 ^ n10883 ^ n3791 ;
  assign n46344 = n8445 ^ n1159 ^ 1'b0 ;
  assign n46346 = n6988 ^ n108 ^ 1'b0 ;
  assign n46347 = n7434 & n46346 ;
  assign n46348 = n38136 ^ n22052 ^ 1'b0 ;
  assign n46349 = n46347 & ~n46348 ;
  assign n46345 = n1290 | n16407 ;
  assign n46350 = n46349 ^ n46345 ^ 1'b0 ;
  assign n46351 = n37309 & ~n41077 ;
  assign n46352 = n46351 ^ n8458 ^ 1'b0 ;
  assign n46353 = n9400 & n19354 ;
  assign n46354 = n46353 ^ n31682 ^ 1'b0 ;
  assign n46355 = n7144 & n32110 ;
  assign n46356 = n46355 ^ n36828 ^ n4417 ;
  assign n46357 = n245 | n36050 ;
  assign n46358 = n33750 | n46357 ;
  assign n46359 = ~n24675 & n46358 ;
  assign n46360 = ( n17034 & ~n17320 ) | ( n17034 & n36185 ) | ( ~n17320 & n36185 ) ;
  assign n46361 = ~n6247 & n46360 ;
  assign n46362 = n42512 & ~n46361 ;
  assign n46363 = n46362 ^ n287 ^ 1'b0 ;
  assign n46364 = n22900 ^ n5554 ^ 1'b0 ;
  assign n46365 = n46363 & n46364 ;
  assign n46366 = n41296 ^ n15886 ^ 1'b0 ;
  assign n46367 = n1209 & ~n25841 ;
  assign n46368 = n46367 ^ n705 ^ 1'b0 ;
  assign n46369 = n10428 & n30924 ;
  assign n46370 = n46369 ^ n18649 ^ 1'b0 ;
  assign n46371 = n1465 & ~n11769 ;
  assign n46372 = n2485 & ~n35176 ;
  assign n46373 = n6039 & n46372 ;
  assign n46374 = ( ~n6096 & n11961 ) | ( ~n6096 & n18118 ) | ( n11961 & n18118 ) ;
  assign n46375 = ( n6844 & ~n46373 ) | ( n6844 & n46374 ) | ( ~n46373 & n46374 ) ;
  assign n46376 = n46375 ^ n5477 ^ 1'b0 ;
  assign n46377 = n2076 & n13344 ;
  assign n46378 = ( ~n12878 & n46376 ) | ( ~n12878 & n46377 ) | ( n46376 & n46377 ) ;
  assign n46379 = n9680 ^ n8891 ^ 1'b0 ;
  assign n46380 = ~n7295 & n46379 ;
  assign n46381 = n46380 ^ n33399 ^ n1154 ;
  assign n46382 = n4066 | n5725 ;
  assign n46383 = ~n10795 & n24216 ;
  assign n46384 = ~n5641 & n46383 ;
  assign n46385 = ~n11693 & n46384 ;
  assign n46386 = n41678 ^ n38509 ^ 1'b0 ;
  assign n46387 = n37972 | n46386 ;
  assign n46388 = n33089 ^ n4222 ^ 1'b0 ;
  assign n46389 = n46388 ^ n24702 ^ 1'b0 ;
  assign n46390 = ~n36201 & n46389 ;
  assign n46391 = n3578 | n18867 ;
  assign n46392 = n1926 | n10320 ;
  assign n46393 = n46392 ^ n9908 ^ 1'b0 ;
  assign n46394 = ( n44754 & n45808 ) | ( n44754 & n46393 ) | ( n45808 & n46393 ) ;
  assign n46395 = n46394 ^ n20664 ^ 1'b0 ;
  assign n46396 = n46395 ^ n13610 ^ 1'b0 ;
  assign n46397 = ( n7171 & n32230 ) | ( n7171 & n32689 ) | ( n32230 & n32689 ) ;
  assign n46398 = n18316 & n21065 ;
  assign n46399 = n46398 ^ n43332 ^ 1'b0 ;
  assign n46400 = n863 & n11599 ;
  assign n46401 = ~n20845 & n46400 ;
  assign n46402 = n25771 ^ n3071 ^ 1'b0 ;
  assign n46403 = n13337 ^ n8871 ^ 1'b0 ;
  assign n46404 = ~n46402 & n46403 ;
  assign n46405 = n46404 ^ n33392 ^ 1'b0 ;
  assign n46406 = n22170 & n46405 ;
  assign n46408 = n8921 ^ n4851 ^ 1'b0 ;
  assign n46409 = n11727 | n46408 ;
  assign n46410 = n22182 | n46409 ;
  assign n46407 = n10551 & n43203 ;
  assign n46411 = n46410 ^ n46407 ^ 1'b0 ;
  assign n46412 = n13747 ^ n10227 ^ 1'b0 ;
  assign n46413 = n46412 ^ n30075 ^ n12474 ;
  assign n46414 = n3205 & n22369 ;
  assign n46415 = n46414 ^ n43015 ^ 1'b0 ;
  assign n46416 = n39205 ^ n14204 ^ 1'b0 ;
  assign n46417 = n5173 & ~n16762 ;
  assign n46419 = n7167 | n32611 ;
  assign n46418 = ~n13030 & n31609 ;
  assign n46420 = n46419 ^ n46418 ^ 1'b0 ;
  assign n46421 = ( n1773 & n1940 ) | ( n1773 & n19689 ) | ( n1940 & n19689 ) ;
  assign n46422 = n41156 ^ n6269 ^ 1'b0 ;
  assign n46423 = ~n46421 & n46422 ;
  assign n46424 = ~n10911 & n46423 ;
  assign n46425 = n38539 & n46424 ;
  assign n46426 = n46425 ^ n37746 ^ 1'b0 ;
  assign n46427 = n3686 | n17513 ;
  assign n46428 = ( n31087 & n42269 ) | ( n31087 & n46427 ) | ( n42269 & n46427 ) ;
  assign n46429 = n20849 | n37137 ;
  assign n46430 = n46429 ^ n44770 ^ 1'b0 ;
  assign n46432 = n4582 | n25200 ;
  assign n46433 = ( ~n999 & n1864 ) | ( ~n999 & n29761 ) | ( n1864 & n29761 ) ;
  assign n46434 = ~n46432 & n46433 ;
  assign n46431 = n4258 & n10812 ;
  assign n46435 = n46434 ^ n46431 ^ 1'b0 ;
  assign n46436 = n11432 ^ n3368 ^ 1'b0 ;
  assign n46437 = n29160 | n46436 ;
  assign n46438 = n7668 | n14100 ;
  assign n46439 = n46437 & ~n46438 ;
  assign n46440 = n30967 | n46439 ;
  assign n46441 = n13904 ^ n9947 ^ 1'b0 ;
  assign n46442 = n12251 | n46441 ;
  assign n46443 = n6437 & ~n46442 ;
  assign n46444 = n23904 | n25424 ;
  assign n46445 = n3923 | n46444 ;
  assign n46446 = n33078 ^ n1185 ^ 1'b0 ;
  assign n46447 = ( ~n6566 & n24086 ) | ( ~n6566 & n46446 ) | ( n24086 & n46446 ) ;
  assign n46448 = n1623 & n3398 ;
  assign n46449 = n46448 ^ n3214 ^ 1'b0 ;
  assign n46450 = n46449 ^ n31670 ^ n11035 ;
  assign n46451 = n5914 & n23499 ;
  assign n46452 = ~n20532 & n22760 ;
  assign n46453 = n46451 | n46452 ;
  assign n46454 = n43757 ^ n5315 ^ 1'b0 ;
  assign n46455 = ~n19985 & n46454 ;
  assign n46456 = n18667 ^ n1250 ^ 1'b0 ;
  assign n46457 = n5342 | n46456 ;
  assign n46458 = n12120 & n46457 ;
  assign n46459 = n28567 | n30870 ;
  assign n46460 = n26794 & n46459 ;
  assign n46461 = n46460 ^ n37081 ^ n10314 ;
  assign n46462 = n12077 & ~n13993 ;
  assign n46463 = n46462 ^ n7104 ^ 1'b0 ;
  assign n46464 = n12071 | n46463 ;
  assign n46465 = ~n989 & n46464 ;
  assign n46466 = n5648 | n18929 ;
  assign n46467 = n25621 ^ n1924 ^ 1'b0 ;
  assign n46468 = n35200 & n46467 ;
  assign n46469 = n19244 ^ n17685 ^ 1'b0 ;
  assign n46470 = n46469 ^ n37817 ^ 1'b0 ;
  assign n46471 = n10490 & n46470 ;
  assign n46472 = n34192 ^ n12668 ^ n8403 ;
  assign n46473 = n45431 ^ n25824 ^ n4681 ;
  assign n46474 = n6914 ^ n2725 ^ 1'b0 ;
  assign n46475 = n10371 | n46474 ;
  assign n46476 = ~n33180 & n41273 ;
  assign n46477 = ( n34589 & ~n46475 ) | ( n34589 & n46476 ) | ( ~n46475 & n46476 ) ;
  assign n46478 = n11269 & n20772 ;
  assign n46479 = n13215 & ~n29596 ;
  assign n46480 = ( n3102 & n9993 ) | ( n3102 & n19180 ) | ( n9993 & n19180 ) ;
  assign n46481 = n46480 ^ n46185 ^ 1'b0 ;
  assign n46482 = n29118 ^ n15601 ^ 1'b0 ;
  assign n46483 = n27226 & n46482 ;
  assign n46485 = n15026 ^ n5994 ^ 1'b0 ;
  assign n46484 = n13858 ^ n7280 ^ 1'b0 ;
  assign n46486 = n46485 ^ n46484 ^ 1'b0 ;
  assign n46487 = n46486 ^ n16657 ^ 1'b0 ;
  assign n46488 = ( n14395 & n21130 ) | ( n14395 & ~n26371 ) | ( n21130 & ~n26371 ) ;
  assign n46489 = n46488 ^ n14684 ^ 1'b0 ;
  assign n46490 = ~n25891 & n46489 ;
  assign n46491 = n3930 & n9564 ;
  assign n46492 = n12126 & n18729 ;
  assign n46493 = n2328 & n46492 ;
  assign n46494 = ( n7097 & n7215 ) | ( n7097 & ~n46493 ) | ( n7215 & ~n46493 ) ;
  assign n46495 = ( n17971 & ~n46491 ) | ( n17971 & n46494 ) | ( ~n46491 & n46494 ) ;
  assign n46496 = n46495 ^ n20903 ^ 1'b0 ;
  assign n46497 = n35515 ^ n7000 ^ 1'b0 ;
  assign n46498 = ~n1337 & n46497 ;
  assign n46499 = n46498 ^ n3573 ^ 1'b0 ;
  assign n46500 = n7534 | n24323 ;
  assign n46501 = ~n12369 & n39212 ;
  assign n46502 = n37438 ^ n12618 ^ 1'b0 ;
  assign n46503 = n27414 | n46502 ;
  assign n46504 = n4914 & ~n20314 ;
  assign n46505 = n1437 & n37236 ;
  assign n46506 = ( n46503 & n46504 ) | ( n46503 & n46505 ) | ( n46504 & n46505 ) ;
  assign n46507 = n611 & ~n5504 ;
  assign n46508 = n24061 & n46507 ;
  assign n46509 = n46508 ^ n7001 ^ n210 ;
  assign n46510 = n2949 & n6083 ;
  assign n46511 = n46510 ^ n1387 ^ 1'b0 ;
  assign n46512 = ( n7913 & n25391 ) | ( n7913 & ~n46511 ) | ( n25391 & ~n46511 ) ;
  assign n46513 = n46512 ^ n30553 ^ 1'b0 ;
  assign n46514 = n27087 & ~n33010 ;
  assign n46515 = n46514 ^ n4593 ^ 1'b0 ;
  assign n46516 = n3778 & ~n38100 ;
  assign n46517 = n46516 ^ n15868 ^ 1'b0 ;
  assign n46518 = n46517 ^ n9507 ^ 1'b0 ;
  assign n46519 = n20176 | n46518 ;
  assign n46520 = n29040 ^ n5483 ^ 1'b0 ;
  assign n46521 = n6415 & n43572 ;
  assign n46522 = n25526 ^ n9390 ^ 1'b0 ;
  assign n46524 = ~n27726 & n30718 ;
  assign n46523 = ~n6135 & n17359 ;
  assign n46525 = n46524 ^ n46523 ^ 1'b0 ;
  assign n46526 = n25579 ^ n980 ^ 1'b0 ;
  assign n46527 = ~n809 & n46526 ;
  assign n46528 = ~n5084 & n46527 ;
  assign n46529 = n12794 & n46528 ;
  assign n46530 = n22507 ^ n6219 ^ 1'b0 ;
  assign n46531 = n6191 | n10712 ;
  assign n46532 = n46531 ^ n32929 ^ 1'b0 ;
  assign n46533 = n45222 & ~n46532 ;
  assign n46534 = ( n16200 & n16682 ) | ( n16200 & ~n17842 ) | ( n16682 & ~n17842 ) ;
  assign n46535 = n17414 ^ n10781 ^ 1'b0 ;
  assign n46536 = n764 & ~n46535 ;
  assign n46537 = ~n3125 & n46536 ;
  assign n46538 = n772 & n46537 ;
  assign n46539 = n46534 & n46538 ;
  assign n46540 = ( n9532 & ~n15617 ) | ( n9532 & n17805 ) | ( ~n15617 & n17805 ) ;
  assign n46541 = n46540 ^ n29366 ^ n17969 ;
  assign n46542 = ( n310 & n5580 ) | ( n310 & ~n6659 ) | ( n5580 & ~n6659 ) ;
  assign n46543 = ~n4892 & n29200 ;
  assign n46544 = n6931 & n46543 ;
  assign n46546 = ~n19536 & n25655 ;
  assign n46547 = ~n10106 & n46546 ;
  assign n46545 = n21233 & n44940 ;
  assign n46548 = n46547 ^ n46545 ^ 1'b0 ;
  assign n46549 = n17094 | n46548 ;
  assign n46550 = n46549 ^ n24477 ^ 1'b0 ;
  assign n46551 = n5491 & ~n30934 ;
  assign n46552 = n46551 ^ n9860 ^ 1'b0 ;
  assign n46553 = n2859 | n44601 ;
  assign n46554 = n46553 ^ n22562 ^ 1'b0 ;
  assign n46555 = ( n12803 & n46552 ) | ( n12803 & n46554 ) | ( n46552 & n46554 ) ;
  assign n46556 = n25824 ^ n5397 ^ n2495 ;
  assign n46557 = n10936 ^ n4465 ^ 1'b0 ;
  assign n46558 = n24991 | n46557 ;
  assign n46559 = n10511 & n43494 ;
  assign n46560 = n46559 ^ n30553 ^ 1'b0 ;
  assign n46561 = n40014 ^ n13697 ^ n10098 ;
  assign n46562 = ~n4071 & n46561 ;
  assign n46563 = n46562 ^ n11065 ^ 1'b0 ;
  assign n46564 = n38895 ^ n32669 ^ 1'b0 ;
  assign n46565 = n20285 | n46564 ;
  assign n46566 = n46565 ^ n341 ^ 1'b0 ;
  assign n46567 = n4684 | n46566 ;
  assign n46568 = n11037 & ~n46567 ;
  assign n46569 = n46568 ^ n16761 ^ 1'b0 ;
  assign n46570 = n113 | n792 ;
  assign n46571 = n46570 ^ n37677 ^ 1'b0 ;
  assign n46572 = n16402 ^ n4477 ^ 1'b0 ;
  assign n46573 = n41099 & n46572 ;
  assign n46574 = n45245 ^ n361 ^ 1'b0 ;
  assign n46575 = ~n27845 & n34273 ;
  assign n46576 = n8746 & ~n15979 ;
  assign n46578 = ( n4618 & ~n8746 ) | ( n4618 & n14283 ) | ( ~n8746 & n14283 ) ;
  assign n46577 = n10346 | n33041 ;
  assign n46579 = n46578 ^ n46577 ^ 1'b0 ;
  assign n46580 = ( n7400 & n11019 ) | ( n7400 & ~n15943 ) | ( n11019 & ~n15943 ) ;
  assign n46581 = n1924 & n9351 ;
  assign n46582 = n46581 ^ n12645 ^ 1'b0 ;
  assign n46583 = ~n813 & n46582 ;
  assign n46584 = n21997 & n27273 ;
  assign n46585 = n36425 & ~n46584 ;
  assign n46586 = ~n42016 & n46585 ;
  assign n46594 = n13770 ^ n1789 ^ 1'b0 ;
  assign n46591 = n4799 ^ n4534 ^ 1'b0 ;
  assign n46592 = n628 | n46591 ;
  assign n46587 = n2775 & n16947 ;
  assign n46588 = n38247 & n46587 ;
  assign n46589 = n46588 ^ n3758 ^ 1'b0 ;
  assign n46590 = ~n576 & n46589 ;
  assign n46593 = n46592 ^ n46590 ^ 1'b0 ;
  assign n46595 = n46594 ^ n46593 ^ n42749 ;
  assign n46596 = n14849 | n22007 ;
  assign n46597 = n46596 ^ n2749 ^ 1'b0 ;
  assign n46598 = n38500 & n46597 ;
  assign n46599 = n46598 ^ n44457 ^ n3477 ;
  assign n46600 = n46599 ^ n6011 ^ 1'b0 ;
  assign n46601 = ~n6335 & n31180 ;
  assign n46602 = n46601 ^ n622 ^ 1'b0 ;
  assign n46605 = n33844 ^ n21858 ^ n4633 ;
  assign n46603 = n3982 ^ n3236 ^ n760 ;
  assign n46604 = n46603 ^ n17590 ^ n13531 ;
  assign n46606 = n46605 ^ n46604 ^ 1'b0 ;
  assign n46607 = n24237 | n30680 ;
  assign n46608 = n46607 ^ n17860 ^ 1'b0 ;
  assign n46609 = n1414 & ~n14379 ;
  assign n46610 = n46609 ^ n27316 ^ 1'b0 ;
  assign n46611 = n2516 & n46610 ;
  assign n46612 = ~n21434 & n32573 ;
  assign n46613 = n22068 & n38957 ;
  assign n46614 = n46613 ^ n3667 ^ 1'b0 ;
  assign n46615 = n498 | n2718 ;
  assign n46616 = n32909 | n42679 ;
  assign n46617 = n25973 & ~n46616 ;
  assign n46618 = n34066 ^ n31604 ^ 1'b0 ;
  assign n46619 = n8873 ^ n6027 ^ 1'b0 ;
  assign n46620 = n9659 & ~n46619 ;
  assign n46621 = n19245 ^ n11583 ^ 1'b0 ;
  assign n46622 = n12698 & ~n27032 ;
  assign n46623 = n46622 ^ n26976 ^ 1'b0 ;
  assign n46624 = n1094 & n22237 ;
  assign n46625 = ~n46623 & n46624 ;
  assign n46626 = n3650 & ~n37503 ;
  assign n46627 = n30055 & ~n46626 ;
  assign n46628 = n46625 & n46627 ;
  assign n46629 = n46628 ^ n42493 ^ 1'b0 ;
  assign n46630 = x3 | n18689 ;
  assign n46631 = n31012 & n46630 ;
  assign n46632 = n7884 & n46631 ;
  assign n46633 = n46632 ^ n9376 ^ 1'b0 ;
  assign n46634 = n14997 ^ n963 ^ 1'b0 ;
  assign n46635 = ( n2509 & ~n40008 ) | ( n2509 & n46634 ) | ( ~n40008 & n46634 ) ;
  assign n46636 = n13660 & n46635 ;
  assign n46637 = n46633 & n46636 ;
  assign n46638 = n32530 ^ n13678 ^ 1'b0 ;
  assign n46639 = n46638 ^ n11683 ^ 1'b0 ;
  assign n46640 = n582 | n694 ;
  assign n46641 = ~n10587 & n36388 ;
  assign n46642 = n46641 ^ n22290 ^ 1'b0 ;
  assign n46643 = n34018 ^ n791 ^ n200 ;
  assign n46644 = n30525 & ~n31689 ;
  assign n46645 = ~n46643 & n46644 ;
  assign n46646 = n112 | n3684 ;
  assign n46647 = n7267 & n8241 ;
  assign n46648 = n46646 & ~n46647 ;
  assign n46649 = n3901 & ~n9264 ;
  assign n46650 = ~n33795 & n46649 ;
  assign n46651 = n11498 | n34519 ;
  assign n46652 = ( n14487 & n30350 ) | ( n14487 & ~n46651 ) | ( n30350 & ~n46651 ) ;
  assign n46653 = ( n5844 & n7989 ) | ( n5844 & n27505 ) | ( n7989 & n27505 ) ;
  assign n46654 = n34596 & ~n42448 ;
  assign n46655 = n33433 ^ n11870 ^ 1'b0 ;
  assign n46656 = n46655 ^ n14288 ^ 1'b0 ;
  assign n46657 = n28709 | n46656 ;
  assign n46658 = n26921 | n34869 ;
  assign n46659 = n46658 ^ n5209 ^ 1'b0 ;
  assign n46660 = n14112 & n21352 ;
  assign n46661 = n46660 ^ n19597 ^ 1'b0 ;
  assign n46662 = n3898 & ~n46661 ;
  assign n46663 = ~n51 & n8120 ;
  assign n46664 = n46663 ^ n9117 ^ 1'b0 ;
  assign n46665 = n22373 | n46664 ;
  assign n46666 = n46665 ^ n33318 ^ 1'b0 ;
  assign n46667 = n36697 ^ n15182 ^ 1'b0 ;
  assign n46668 = n9416 | n19605 ;
  assign n46669 = n46668 ^ n33148 ^ n28564 ;
  assign n46671 = n31483 ^ n16409 ^ 1'b0 ;
  assign n46670 = n4004 & ~n11132 ;
  assign n46672 = n46671 ^ n46670 ^ 1'b0 ;
  assign n46673 = n38326 ^ n25767 ^ n14534 ;
  assign n46674 = n46170 | n46673 ;
  assign n46678 = n3772 | n8165 ;
  assign n46675 = ~n4307 & n41613 ;
  assign n46676 = n46675 ^ n25812 ^ 1'b0 ;
  assign n46677 = n4571 & ~n46676 ;
  assign n46679 = n46678 ^ n46677 ^ 1'b0 ;
  assign n46680 = n12507 & n28295 ;
  assign n46681 = n29641 ^ n1798 ^ 1'b0 ;
  assign n46682 = ~n2065 & n46681 ;
  assign n46683 = n2943 | n6635 ;
  assign n46684 = n46683 ^ n3498 ^ 1'b0 ;
  assign n46685 = n46684 ^ n14710 ^ 1'b0 ;
  assign n46686 = n7557 | n35920 ;
  assign n46687 = n46686 ^ n21366 ^ 1'b0 ;
  assign n46688 = n42663 ^ n18453 ^ n12940 ;
  assign n46689 = n46688 ^ n43111 ^ n16252 ;
  assign n46690 = n34853 ^ n26571 ^ n1311 ;
  assign n46691 = n12307 & ~n24380 ;
  assign n46692 = n46691 ^ n34768 ^ 1'b0 ;
  assign n46693 = n28081 ^ n3825 ^ 1'b0 ;
  assign n46694 = n46692 & ~n46693 ;
  assign n46695 = n23036 & n46694 ;
  assign n46696 = n22713 & n46695 ;
  assign n46697 = n12340 | n46696 ;
  assign n46698 = n11233 ^ n3754 ^ 1'b0 ;
  assign n46699 = n29424 | n42289 ;
  assign n46700 = n17887 ^ n9036 ^ 1'b0 ;
  assign n46701 = ~n13453 & n46700 ;
  assign n46702 = n23593 & n35051 ;
  assign n46703 = n46702 ^ n221 ^ 1'b0 ;
  assign n46704 = n7122 ^ n1176 ^ 1'b0 ;
  assign n46705 = n1279 | n46704 ;
  assign n46706 = n6827 | n46705 ;
  assign n46707 = n46706 ^ n3371 ^ 1'b0 ;
  assign n46708 = n6010 | n9005 ;
  assign n46709 = n13903 ^ n990 ^ 1'b0 ;
  assign n46710 = ~n46708 & n46709 ;
  assign n46711 = n12494 ^ n11871 ^ 1'b0 ;
  assign n46712 = n15787 & n46711 ;
  assign n46713 = n7312 | n16504 ;
  assign n46714 = n28775 & n46713 ;
  assign n46715 = n46714 ^ n14826 ^ n369 ;
  assign n46716 = n40649 ^ n33720 ^ 1'b0 ;
  assign n46718 = n1526 & n3382 ;
  assign n46719 = ~n12349 & n46718 ;
  assign n46717 = n2794 & n13854 ;
  assign n46720 = n46719 ^ n46717 ^ 1'b0 ;
  assign n46721 = n9033 & n15483 ;
  assign n46722 = n46721 ^ n6930 ^ 1'b0 ;
  assign n46723 = n12772 & n40467 ;
  assign n46724 = n46723 ^ n953 ^ 1'b0 ;
  assign n46725 = n46724 ^ n32244 ^ 1'b0 ;
  assign n46726 = n3762 & ~n46725 ;
  assign n46727 = n44912 ^ n24395 ^ n3180 ;
  assign n46728 = ( n22466 & ~n38910 ) | ( n22466 & n46727 ) | ( ~n38910 & n46727 ) ;
  assign n46729 = ~n16363 & n33231 ;
  assign n46730 = n14718 & ~n31648 ;
  assign n46731 = n9137 & n46730 ;
  assign n46732 = n20509 ^ n6351 ^ 1'b0 ;
  assign n46733 = ~n46731 & n46732 ;
  assign n46734 = n7612 | n18924 ;
  assign n46735 = n19328 | n46734 ;
  assign n46736 = ( n1036 & n4265 ) | ( n1036 & n38551 ) | ( n4265 & n38551 ) ;
  assign n46740 = n510 & ~n8215 ;
  assign n46737 = n16153 & ~n21734 ;
  assign n46738 = n46737 ^ n22745 ^ 1'b0 ;
  assign n46739 = n21664 & ~n46738 ;
  assign n46741 = n46740 ^ n46739 ^ 1'b0 ;
  assign n46742 = n30614 ^ n28620 ^ 1'b0 ;
  assign n46743 = n1064 & ~n32110 ;
  assign n46744 = n46743 ^ n14030 ^ 1'b0 ;
  assign n46745 = n134 & n28574 ;
  assign n46746 = n4460 & ~n46745 ;
  assign n46747 = n4023 & n46746 ;
  assign n46748 = n1160 ^ n757 ^ 1'b0 ;
  assign n46749 = ~n46747 & n46748 ;
  assign n46750 = n19099 & n19497 ;
  assign n46751 = n23404 & n39655 ;
  assign n46752 = n18570 & n46751 ;
  assign n46753 = ~n5816 & n21020 ;
  assign n46754 = n46753 ^ n6703 ^ 1'b0 ;
  assign n46755 = n989 | n6662 ;
  assign n46756 = n1531 & n10171 ;
  assign n46757 = ~n46755 & n46756 ;
  assign n46758 = ( n6716 & n11806 ) | ( n6716 & n46757 ) | ( n11806 & n46757 ) ;
  assign n46759 = ( n18246 & n40255 ) | ( n18246 & n44447 ) | ( n40255 & n44447 ) ;
  assign n46760 = ( ~n4862 & n12529 ) | ( ~n4862 & n46759 ) | ( n12529 & n46759 ) ;
  assign n46761 = n10909 ^ n485 ^ 1'b0 ;
  assign n46762 = n46761 ^ n28054 ^ n23675 ;
  assign n46763 = n30853 ^ n20692 ^ 1'b0 ;
  assign n46764 = n7319 | n46763 ;
  assign n46765 = n16719 & ~n18033 ;
  assign n46766 = n46765 ^ n25181 ^ 1'b0 ;
  assign n46767 = ~n922 & n46766 ;
  assign n46770 = n6013 | n33540 ;
  assign n46768 = n39526 & ~n46495 ;
  assign n46769 = n15537 & n46768 ;
  assign n46771 = n46770 ^ n46769 ^ 1'b0 ;
  assign n46772 = n16506 & n46614 ;
  assign n46773 = ~n27720 & n46772 ;
  assign n46774 = n9975 & ~n12033 ;
  assign n46775 = n46774 ^ n36299 ^ n10035 ;
  assign n46776 = n5791 & ~n13046 ;
  assign n46777 = n15317 ^ n8911 ^ 1'b0 ;
  assign n46778 = n7338 & n16722 ;
  assign n46779 = n4112 & ~n35900 ;
  assign n46780 = n46779 ^ n14247 ^ 1'b0 ;
  assign n46781 = n14183 & n27205 ;
  assign n46782 = n46781 ^ n42506 ^ n23588 ;
  assign n46783 = ( n27984 & n31764 ) | ( n27984 & ~n42996 ) | ( n31764 & ~n42996 ) ;
  assign n46784 = n27864 ^ n20812 ^ n2885 ;
  assign n46785 = n5461 & ~n19623 ;
  assign n46786 = n46785 ^ n1214 ^ 1'b0 ;
  assign n46787 = n46786 ^ n20220 ^ 1'b0 ;
  assign n46788 = n32589 | n46787 ;
  assign n46789 = n19198 ^ n15349 ^ 1'b0 ;
  assign n46790 = n21085 & n46789 ;
  assign n46791 = ~n6131 & n28398 ;
  assign n46792 = n471 | n13974 ;
  assign n46793 = n19483 & ~n46792 ;
  assign n46794 = ~n9548 & n19872 ;
  assign n46795 = n3260 & n13275 ;
  assign n46796 = n46795 ^ n6438 ^ 1'b0 ;
  assign n46797 = n46796 ^ n1698 ^ n1437 ;
  assign n46798 = n9656 & n46797 ;
  assign n46799 = n865 | n20470 ;
  assign n46800 = n15476 & ~n46799 ;
  assign n46801 = n46800 ^ n12046 ^ n11406 ;
  assign n46802 = n15807 ^ n9908 ^ 1'b0 ;
  assign n46803 = n13956 ^ n10108 ^ n2760 ;
  assign n46804 = n33416 ^ n2422 ^ 1'b0 ;
  assign n46805 = ~n14658 & n24934 ;
  assign n46807 = ~n12851 & n22018 ;
  assign n46808 = ~n9031 & n46807 ;
  assign n46806 = n23393 | n35328 ;
  assign n46809 = n46808 ^ n46806 ^ n20622 ;
  assign n46810 = n32216 ^ n15169 ^ n11082 ;
  assign n46811 = ~n17377 & n18904 ;
  assign n46812 = n38166 ^ n30269 ^ 1'b0 ;
  assign n46813 = n46812 ^ n12850 ^ 1'b0 ;
  assign n46814 = n27043 & n46813 ;
  assign n46815 = n46814 ^ n26114 ^ 1'b0 ;
  assign n46816 = n46811 & n46815 ;
  assign n46817 = n14074 ^ n8657 ^ 1'b0 ;
  assign n46818 = n29298 ^ n23590 ^ 1'b0 ;
  assign n46819 = ~n34450 & n46818 ;
  assign n46820 = ( n1296 & ~n2779 ) | ( n1296 & n29225 ) | ( ~n2779 & n29225 ) ;
  assign n46821 = ~n1326 & n28360 ;
  assign n46822 = n32576 ^ n9513 ^ n1910 ;
  assign n46824 = n26673 & n39526 ;
  assign n46823 = n7776 & n21183 ;
  assign n46825 = n46824 ^ n46823 ^ 1'b0 ;
  assign n46826 = n46825 ^ n36853 ^ 1'b0 ;
  assign n46827 = n27382 ^ n8305 ^ n2472 ;
  assign n46828 = n18611 ^ n2679 ^ 1'b0 ;
  assign n46829 = n46827 & ~n46828 ;
  assign n46830 = n26412 ^ n257 ^ 1'b0 ;
  assign n46831 = ~n1491 & n4262 ;
  assign n46832 = n46831 ^ n362 ^ 1'b0 ;
  assign n46833 = n46832 ^ n1348 ^ 1'b0 ;
  assign n46834 = n41670 ^ n30196 ^ 1'b0 ;
  assign n46835 = n12827 ^ n10423 ^ 1'b0 ;
  assign n46836 = n34274 & ~n46835 ;
  assign n46837 = ~n3446 & n12976 ;
  assign n46838 = ~n46836 & n46837 ;
  assign n46839 = n5443 & ~n34774 ;
  assign n46840 = ~n9151 & n28278 ;
  assign n46841 = n46840 ^ n27191 ^ 1'b0 ;
  assign n46842 = n3187 ^ n1387 ^ 1'b0 ;
  assign n46843 = ~n26373 & n46842 ;
  assign n46844 = n24374 & ~n29759 ;
  assign n46845 = ~n46843 & n46844 ;
  assign n46846 = n15920 & ~n39804 ;
  assign n46847 = n37466 ^ n33784 ^ n8919 ;
  assign n46848 = n20679 & n33784 ;
  assign n46849 = ( ~n12703 & n24801 ) | ( ~n12703 & n32211 ) | ( n24801 & n32211 ) ;
  assign n46850 = n27255 ^ n7483 ^ 1'b0 ;
  assign n46851 = n44642 ^ n383 ^ 1'b0 ;
  assign n46852 = n46850 & n46851 ;
  assign n46853 = n34974 ^ n2190 ^ 1'b0 ;
  assign n46854 = ~n7772 & n12812 ;
  assign n46855 = n46854 ^ n39377 ^ 1'b0 ;
  assign n46856 = n8993 & ~n46855 ;
  assign n46857 = ~n5978 & n46856 ;
  assign n46858 = n5312 & ~n6648 ;
  assign n46859 = ( ~n4908 & n10829 ) | ( ~n4908 & n13587 ) | ( n10829 & n13587 ) ;
  assign n46860 = ~n20896 & n46859 ;
  assign n46861 = n46860 ^ n2270 ^ 1'b0 ;
  assign n46862 = n11718 | n43035 ;
  assign n46863 = n46861 & ~n46862 ;
  assign n46864 = ( ~n3457 & n3802 ) | ( ~n3457 & n21640 ) | ( n3802 & n21640 ) ;
  assign n46865 = n29199 & n39235 ;
  assign n46866 = ( n10634 & n14141 ) | ( n10634 & n16816 ) | ( n14141 & n16816 ) ;
  assign n46867 = n46866 ^ n24108 ^ 1'b0 ;
  assign n46868 = n11207 | n46867 ;
  assign n46869 = n8830 & ~n46868 ;
  assign n46870 = n46869 ^ n7581 ^ 1'b0 ;
  assign n46872 = n12959 | n29333 ;
  assign n46873 = n46872 ^ n38175 ^ 1'b0 ;
  assign n46871 = n44412 ^ n20938 ^ 1'b0 ;
  assign n46874 = n46873 ^ n46871 ^ 1'b0 ;
  assign n46875 = n46870 & n46874 ;
  assign n46876 = n10729 ^ n2979 ^ 1'b0 ;
  assign n46877 = n27418 | n46876 ;
  assign n46878 = n19906 & ~n46877 ;
  assign n46879 = n6908 & n46878 ;
  assign n46880 = n34162 & n46879 ;
  assign n46881 = n18745 ^ n1022 ^ 1'b0 ;
  assign n46882 = n63 | n16086 ;
  assign n46883 = n46881 & ~n46882 ;
  assign n46884 = n21955 & ~n46883 ;
  assign n46885 = n32188 & n46884 ;
  assign n46886 = n22721 | n22744 ;
  assign n46887 = n4211 & ~n46886 ;
  assign n46888 = ~n2071 & n8821 ;
  assign n46889 = n46888 ^ n12527 ^ 1'b0 ;
  assign n46895 = n2798 & n14932 ;
  assign n46890 = ~n15716 & n21204 ;
  assign n46891 = ~n811 & n46890 ;
  assign n46892 = n1447 & n29567 ;
  assign n46893 = ~n11135 & n46892 ;
  assign n46894 = ~n46891 & n46893 ;
  assign n46896 = n46895 ^ n46894 ^ 1'b0 ;
  assign n46897 = n38292 & ~n46896 ;
  assign n46898 = n34922 | n37664 ;
  assign n46899 = n8821 | n24121 ;
  assign n46900 = n46899 ^ n26099 ^ 1'b0 ;
  assign n46901 = n43438 ^ n35719 ^ 1'b0 ;
  assign n46902 = ~n46900 & n46901 ;
  assign n46903 = n6875 ^ n6566 ^ 1'b0 ;
  assign n46904 = n46903 ^ n963 ^ 1'b0 ;
  assign n46905 = n210 | n11015 ;
  assign n46906 = n46905 ^ n3370 ^ 1'b0 ;
  assign n46909 = n1178 & ~n4799 ;
  assign n46907 = n22144 | n37112 ;
  assign n46908 = n46907 ^ n6128 ^ 1'b0 ;
  assign n46910 = n46909 ^ n46908 ^ 1'b0 ;
  assign n46911 = ~n46906 & n46910 ;
  assign n46912 = ~n15871 & n46911 ;
  assign n46913 = n6412 & n46912 ;
  assign n46914 = n18804 | n20031 ;
  assign n46915 = n46914 ^ n11601 ^ 1'b0 ;
  assign n46916 = n4475 & ~n21935 ;
  assign n46917 = n46916 ^ n12097 ^ 1'b0 ;
  assign n46918 = n18369 | n20142 ;
  assign n46919 = n34001 ^ n26916 ^ n19505 ;
  assign n46920 = n16620 & n46919 ;
  assign n46921 = n46920 ^ n3196 ^ 1'b0 ;
  assign n46922 = n39163 ^ n16278 ^ n6510 ;
  assign n46923 = n33843 | n46922 ;
  assign n46924 = n46923 ^ n11554 ^ 1'b0 ;
  assign n46925 = ~n14500 & n14820 ;
  assign n46926 = n27480 & n46925 ;
  assign n46927 = n10340 & n25622 ;
  assign n46928 = ~n334 & n46927 ;
  assign n46929 = ( n850 & n9202 ) | ( n850 & n45622 ) | ( n9202 & n45622 ) ;
  assign n46930 = ~n46928 & n46929 ;
  assign n46931 = ~n18681 & n45680 ;
  assign n46932 = n32853 ^ n87 ^ 1'b0 ;
  assign n46933 = ( n17086 & n24624 ) | ( n17086 & ~n46932 ) | ( n24624 & ~n46932 ) ;
  assign n46934 = n16352 ^ n2806 ^ n126 ;
  assign n46935 = ( n3308 & ~n27440 ) | ( n3308 & n34077 ) | ( ~n27440 & n34077 ) ;
  assign n46936 = n5809 & ~n10272 ;
  assign n46937 = n46936 ^ n15705 ^ 1'b0 ;
  assign n46938 = n36279 & n46937 ;
  assign n46939 = n46938 ^ n4316 ^ 1'b0 ;
  assign n46940 = n31639 | n46939 ;
  assign n46941 = n46940 ^ n22506 ^ 1'b0 ;
  assign n46942 = n13593 | n30036 ;
  assign n46943 = n23033 & ~n31180 ;
  assign n46944 = n46943 ^ n24072 ^ 1'b0 ;
  assign n46945 = n22240 ^ n7943 ^ n5581 ;
  assign n46946 = n46945 ^ n9286 ^ 1'b0 ;
  assign n46947 = ~n17828 & n19915 ;
  assign n46948 = n46947 ^ n4825 ^ 1'b0 ;
  assign n46949 = n23825 & n26465 ;
  assign n46950 = n17513 & n46949 ;
  assign n46951 = n46950 ^ n32218 ^ 1'b0 ;
  assign n46952 = n46948 & n46951 ;
  assign n46953 = n341 & n875 ;
  assign n46954 = n9132 & ~n11657 ;
  assign n46955 = n132 & n46954 ;
  assign n46956 = n31130 ^ n21568 ^ 1'b0 ;
  assign n46957 = n29319 | n34290 ;
  assign n46958 = n26344 ^ n5220 ^ 1'b0 ;
  assign n46959 = ~n18371 & n46958 ;
  assign n46960 = n46747 & n46959 ;
  assign n46961 = n350 & ~n18822 ;
  assign n46962 = n45595 ^ n14156 ^ 1'b0 ;
  assign n46963 = n13567 ^ n5128 ^ 1'b0 ;
  assign n46964 = n46963 ^ n44244 ^ 1'b0 ;
  assign n46965 = n11108 & ~n19808 ;
  assign n46966 = ( n1368 & ~n46964 ) | ( n1368 & n46965 ) | ( ~n46964 & n46965 ) ;
  assign n46967 = n17173 ^ n1538 ^ 1'b0 ;
  assign n46968 = n13159 | n46967 ;
  assign n46969 = n7261 & ~n46968 ;
  assign n46971 = n25702 | n26196 ;
  assign n46972 = n20638 & n46971 ;
  assign n46970 = ~n6866 & n16733 ;
  assign n46973 = n46972 ^ n46970 ^ 1'b0 ;
  assign n46974 = n20395 ^ n12091 ^ n11771 ;
  assign n46975 = n46974 ^ n11917 ^ 1'b0 ;
  assign n46976 = n32327 & n46975 ;
  assign n46977 = n46976 ^ n22466 ^ 1'b0 ;
  assign n46978 = n46973 & ~n46977 ;
  assign n46979 = n10291 & ~n29192 ;
  assign n46980 = n44 & n46979 ;
  assign n46981 = n20149 ^ n4977 ^ 1'b0 ;
  assign n46982 = n25301 | n31398 ;
  assign n46983 = n381 | n46982 ;
  assign n46984 = ~n44019 & n46983 ;
  assign n46985 = n4140 & n10072 ;
  assign n46986 = n26124 ^ n22057 ^ 1'b0 ;
  assign n46987 = n16271 & ~n46986 ;
  assign n46988 = n46987 ^ n10808 ^ 1'b0 ;
  assign n46989 = ( n6202 & n6460 ) | ( n6202 & n32623 ) | ( n6460 & n32623 ) ;
  assign n46990 = ~n7490 & n37200 ;
  assign n46991 = n4977 & ~n8071 ;
  assign n46993 = n23654 ^ n10617 ^ n1063 ;
  assign n46992 = n32308 ^ n17574 ^ 1'b0 ;
  assign n46994 = n46993 ^ n46992 ^ n24996 ;
  assign n46995 = n37274 ^ n10348 ^ 1'b0 ;
  assign n46996 = n20871 & n23938 ;
  assign n46997 = n46996 ^ n34959 ^ 1'b0 ;
  assign n46998 = n17016 & ~n46759 ;
  assign n46999 = n34935 ^ n16012 ^ 1'b0 ;
  assign n47000 = n3894 ^ n2986 ^ 1'b0 ;
  assign n47001 = ( n1435 & n16171 ) | ( n1435 & n47000 ) | ( n16171 & n47000 ) ;
  assign n47002 = n16389 & n47001 ;
  assign n47004 = n14231 ^ n5649 ^ 1'b0 ;
  assign n47003 = ~n3460 & n44222 ;
  assign n47005 = n47004 ^ n47003 ^ 1'b0 ;
  assign n47006 = ( n18568 & n26382 ) | ( n18568 & n27885 ) | ( n26382 & n27885 ) ;
  assign n47007 = n32692 ^ n4845 ^ 1'b0 ;
  assign n47008 = ( n28414 & n35411 ) | ( n28414 & n47007 ) | ( n35411 & n47007 ) ;
  assign n47009 = n14247 ^ n9357 ^ 1'b0 ;
  assign n47010 = n7561 ^ n3567 ^ 1'b0 ;
  assign n47011 = n11442 & ~n44137 ;
  assign n47012 = ~n47010 & n47011 ;
  assign n47013 = n827 & ~n32653 ;
  assign n47014 = n14517 & ~n18533 ;
  assign n47015 = n18782 & n20536 ;
  assign n47016 = n47015 ^ n5640 ^ 1'b0 ;
  assign n47018 = ~n2472 & n10038 ;
  assign n47017 = n34762 & ~n45369 ;
  assign n47019 = n47018 ^ n47017 ^ 1'b0 ;
  assign n47020 = ( ~n5337 & n29643 ) | ( ~n5337 & n47019 ) | ( n29643 & n47019 ) ;
  assign n47021 = n13644 ^ n672 ^ 1'b0 ;
  assign n47022 = n27231 ^ n12903 ^ n2139 ;
  assign n47023 = n47021 & ~n47022 ;
  assign n47024 = n18806 & n23215 ;
  assign n47025 = n5691 & n8424 ;
  assign n47026 = n929 & n2195 ;
  assign n47027 = n47026 ^ n2778 ^ 1'b0 ;
  assign n47028 = n47027 ^ n37471 ^ 1'b0 ;
  assign n47029 = n47025 & n47028 ;
  assign n47030 = n1006 & n47029 ;
  assign n47031 = n14801 & n20761 ;
  assign n47032 = n42433 & n47031 ;
  assign n47033 = ( ~n11524 & n12461 ) | ( ~n11524 & n15747 ) | ( n12461 & n15747 ) ;
  assign n47034 = n9176 & n47033 ;
  assign n47035 = n47034 ^ n29617 ^ 1'b0 ;
  assign n47036 = n448 | n5654 ;
  assign n47037 = n47036 ^ n827 ^ 1'b0 ;
  assign n47038 = ~n6100 & n47037 ;
  assign n47039 = n38402 ^ n35261 ^ 1'b0 ;
  assign n47040 = n47038 | n47039 ;
  assign n47041 = n2220 ^ n1718 ^ 1'b0 ;
  assign n47042 = ~n33028 & n47041 ;
  assign n47043 = ~n17146 & n47042 ;
  assign n47044 = n22720 & ~n35453 ;
  assign n47045 = ~n30248 & n47044 ;
  assign n47046 = ~n26938 & n42150 ;
  assign n47047 = n19884 | n20596 ;
  assign n47049 = n12854 ^ n934 ^ 1'b0 ;
  assign n47050 = ~n16644 & n47049 ;
  assign n47048 = n25148 & n28460 ;
  assign n47051 = n47050 ^ n47048 ^ 1'b0 ;
  assign n47053 = n15914 ^ n3812 ^ 1'b0 ;
  assign n47054 = n22450 | n47053 ;
  assign n47052 = ~n6206 & n29434 ;
  assign n47055 = n47054 ^ n47052 ^ 1'b0 ;
  assign n47056 = n34096 ^ n17094 ^ n659 ;
  assign n47057 = ( ~n2012 & n13587 ) | ( ~n2012 & n27959 ) | ( n13587 & n27959 ) ;
  assign n47058 = n47057 ^ n4810 ^ 1'b0 ;
  assign n47059 = n1350 & n13249 ;
  assign n47060 = n47059 ^ n24323 ^ n22363 ;
  assign n47061 = ~n41948 & n47060 ;
  assign n47062 = n2297 | n27148 ;
  assign n47063 = n28972 & ~n47062 ;
  assign n47064 = n27217 ^ n18768 ^ n2280 ;
  assign n47065 = n47064 ^ n26496 ^ n7399 ;
  assign n47066 = n47065 ^ n22546 ^ 1'b0 ;
  assign n47067 = ~n47063 & n47066 ;
  assign n47069 = n13737 ^ n6440 ^ n1656 ;
  assign n47070 = n47069 ^ n5617 ^ 1'b0 ;
  assign n47071 = n22649 ^ n11490 ^ 1'b0 ;
  assign n47072 = n47070 | n47071 ;
  assign n47068 = n2551 & ~n8682 ;
  assign n47073 = n47072 ^ n47068 ^ 1'b0 ;
  assign n47074 = n34791 & n47073 ;
  assign n47075 = n10382 ^ n7196 ^ 1'b0 ;
  assign n47076 = n7493 | n47075 ;
  assign n47077 = n33511 ^ n2106 ^ n1837 ;
  assign n47078 = ~n1945 & n24547 ;
  assign n47079 = n2697 | n6899 ;
  assign n47080 = ( n5388 & n6386 ) | ( n5388 & ~n37491 ) | ( n6386 & ~n37491 ) ;
  assign n47081 = n47080 ^ n6392 ^ 1'b0 ;
  assign n47082 = n22426 | n41575 ;
  assign n47083 = n5303 | n28651 ;
  assign n47084 = n47083 ^ n11892 ^ 1'b0 ;
  assign n47085 = n46270 ^ n43699 ^ n41874 ;
  assign n47086 = ~n16215 & n43595 ;
  assign n47087 = ~n17893 & n25313 ;
  assign n47088 = n397 & ~n1162 ;
  assign n47089 = ~n15389 & n47088 ;
  assign n47090 = n47089 ^ n46147 ^ 1'b0 ;
  assign n47091 = n32669 ^ n7404 ^ n5397 ;
  assign n47092 = n91 & n47091 ;
  assign n47093 = n47092 ^ n40675 ^ 1'b0 ;
  assign n47094 = n3076 & n8424 ;
  assign n47095 = n44286 & n47094 ;
  assign n47096 = n47095 ^ n21376 ^ 1'b0 ;
  assign n47097 = n35308 ^ n34246 ^ n7239 ;
  assign n47098 = ~n7807 & n17237 ;
  assign n47099 = n26459 | n47098 ;
  assign n47102 = n523 & ~n4498 ;
  assign n47100 = n5915 & n12941 ;
  assign n47101 = n15292 | n47100 ;
  assign n47103 = n47102 ^ n47101 ^ 1'b0 ;
  assign n47104 = n24908 ^ n842 ^ 1'b0 ;
  assign n47105 = n26693 ^ n23922 ^ 1'b0 ;
  assign n47107 = n7120 ^ n790 ^ 1'b0 ;
  assign n47108 = n28822 & ~n47107 ;
  assign n47109 = n47108 ^ n33905 ^ n855 ;
  assign n47106 = n4092 & n43498 ;
  assign n47110 = n47109 ^ n47106 ^ 1'b0 ;
  assign n47111 = n14796 | n35931 ;
  assign n47112 = ~n3080 & n29721 ;
  assign n47113 = n10140 ^ n3663 ^ 1'b0 ;
  assign n47114 = ~n22534 & n39192 ;
  assign n47115 = n47113 | n47114 ;
  assign n47116 = n1464 | n2177 ;
  assign n47117 = n47116 ^ n10211 ^ 1'b0 ;
  assign n47118 = n22196 | n22229 ;
  assign n47119 = n27316 & n47118 ;
  assign n47120 = ~n27535 & n47119 ;
  assign n47121 = n15064 | n15287 ;
  assign n47122 = n15534 | n44023 ;
  assign n47123 = n47121 & ~n47122 ;
  assign n47125 = n8414 ^ n7275 ^ 1'b0 ;
  assign n47126 = n47125 ^ n14646 ^ n710 ;
  assign n47127 = n31070 | n47126 ;
  assign n47124 = n24013 & n41931 ;
  assign n47128 = n47127 ^ n47124 ^ 1'b0 ;
  assign n47129 = n5290 & n26929 ;
  assign n47130 = n7774 & n19383 ;
  assign n47131 = n5022 | n10421 ;
  assign n47132 = x3 | n47131 ;
  assign n47133 = n1261 & ~n47132 ;
  assign n47134 = n7708 & n40596 ;
  assign n47135 = n47134 ^ n10339 ^ 1'b0 ;
  assign n47136 = n4072 | n18994 ;
  assign n47137 = ~n4275 & n13272 ;
  assign n47138 = ~n31937 & n47137 ;
  assign n47139 = n13784 & ~n47138 ;
  assign n47140 = n40823 ^ n28506 ^ 1'b0 ;
  assign n47141 = ( n5337 & n13540 ) | ( n5337 & ~n47140 ) | ( n13540 & ~n47140 ) ;
  assign n47142 = n30319 ^ n2609 ^ 1'b0 ;
  assign n47143 = n1450 | n22083 ;
  assign n47144 = n1791 | n34933 ;
  assign n47145 = ~n4988 & n22768 ;
  assign n47146 = n23933 ^ n15042 ^ 1'b0 ;
  assign n47147 = n34266 & n36343 ;
  assign n47148 = n47147 ^ n13064 ^ 1'b0 ;
  assign n47149 = n47146 & n47148 ;
  assign n47150 = n13954 | n28206 ;
  assign n47151 = n47150 ^ n36 ^ 1'b0 ;
  assign n47152 = n18150 & ~n32431 ;
  assign n47153 = ~n41475 & n47152 ;
  assign n47154 = n9039 ^ n8884 ^ 1'b0 ;
  assign n47155 = ~n35404 & n47154 ;
  assign n47156 = n47155 ^ n26642 ^ n5311 ;
  assign n47161 = ~n2657 & n5618 ;
  assign n47162 = n47161 ^ n15600 ^ 1'b0 ;
  assign n47157 = n25651 & ~n44812 ;
  assign n47158 = n47157 ^ n34891 ^ 1'b0 ;
  assign n47159 = n37246 & ~n47158 ;
  assign n47160 = n47159 ^ n8874 ^ 1'b0 ;
  assign n47163 = n47162 ^ n47160 ^ n6335 ;
  assign n47167 = ~n7617 & n38613 ;
  assign n47164 = n10810 ^ n2563 ^ 1'b0 ;
  assign n47165 = n25585 | n47164 ;
  assign n47166 = n19197 & ~n47165 ;
  assign n47168 = n47167 ^ n47166 ^ n43976 ;
  assign n47169 = n7650 & ~n10008 ;
  assign n47170 = n47169 ^ n10723 ^ 1'b0 ;
  assign n47171 = n11761 & n26499 ;
  assign n47172 = ~n39702 & n47171 ;
  assign n47173 = n17797 & ~n47172 ;
  assign n47174 = n13542 ^ n6743 ^ 1'b0 ;
  assign n47175 = ~n40914 & n47174 ;
  assign n47176 = n15335 & n23443 ;
  assign n47177 = n22427 ^ n7962 ^ 1'b0 ;
  assign n47178 = n1959 & ~n47177 ;
  assign n47179 = n24378 & n47178 ;
  assign n47180 = n3599 & n47179 ;
  assign n47181 = n47180 ^ n3081 ^ 1'b0 ;
  assign n47182 = ~n12975 & n20548 ;
  assign n47183 = n47182 ^ n26551 ^ 1'b0 ;
  assign n47184 = n47183 ^ n5527 ^ 1'b0 ;
  assign n47185 = n43855 ^ n14201 ^ 1'b0 ;
  assign n47186 = n8457 & n47185 ;
  assign n47187 = n47186 ^ n35618 ^ 1'b0 ;
  assign n47188 = ~n22479 & n47187 ;
  assign n47189 = n23607 & ~n47188 ;
  assign n47190 = n17251 ^ n3389 ^ n1527 ;
  assign n47191 = ~n17493 & n47190 ;
  assign n47192 = n14545 & n47191 ;
  assign n47193 = ~n16504 & n18462 ;
  assign n47194 = n47193 ^ n14037 ^ 1'b0 ;
  assign n47195 = n47194 ^ n38504 ^ 1'b0 ;
  assign n47196 = n21388 & n33056 ;
  assign n47197 = ~n6322 & n47109 ;
  assign n47198 = n47197 ^ n3375 ^ 1'b0 ;
  assign n47199 = ~n25159 & n47198 ;
  assign n47200 = ~n7941 & n44144 ;
  assign n47201 = n13376 & n47200 ;
  assign n47202 = n32684 ^ n25724 ^ 1'b0 ;
  assign n47203 = n25965 & ~n47202 ;
  assign n47204 = n47203 ^ n26770 ^ 1'b0 ;
  assign n47205 = n15610 ^ n9231 ^ 1'b0 ;
  assign n47206 = n27649 ^ n6925 ^ 1'b0 ;
  assign n47207 = ~n47205 & n47206 ;
  assign n47208 = n36708 ^ n10087 ^ 1'b0 ;
  assign n47209 = n7113 & ~n47208 ;
  assign n47210 = n41640 ^ n17252 ^ 1'b0 ;
  assign n47211 = n22110 & ~n47210 ;
  assign n47212 = n47211 ^ n30752 ^ n172 ;
  assign n47213 = n29174 & ~n34133 ;
  assign n47214 = n47213 ^ n38712 ^ 1'b0 ;
  assign n47215 = n40 | n28924 ;
  assign n47216 = n47215 ^ n36327 ^ 1'b0 ;
  assign n47217 = ( ~n1036 & n11170 ) | ( ~n1036 & n21461 ) | ( n11170 & n21461 ) ;
  assign n47218 = ~n3345 & n9576 ;
  assign n47219 = n47218 ^ n2922 ^ 1'b0 ;
  assign n47220 = n46451 ^ n36708 ^ 1'b0 ;
  assign n47221 = ~n47219 & n47220 ;
  assign n47222 = n356 & n47221 ;
  assign n47223 = n37911 ^ n30904 ^ 1'b0 ;
  assign n47224 = n18104 | n18490 ;
  assign n47225 = n47224 ^ n10705 ^ 1'b0 ;
  assign n47226 = n551 | n33979 ;
  assign n47227 = ( n181 & ~n3784 ) | ( n181 & n47226 ) | ( ~n3784 & n47226 ) ;
  assign n47228 = n32576 ^ n29113 ^ n19014 ;
  assign n47229 = n33526 & n41551 ;
  assign n47230 = n47229 ^ n5372 ^ 1'b0 ;
  assign n47231 = n2555 & n38955 ;
  assign n47232 = ~n11385 & n47231 ;
  assign n47233 = ~n36210 & n47232 ;
  assign n47234 = n14464 & ~n21220 ;
  assign n47235 = n30237 ^ n22269 ^ 1'b0 ;
  assign n47236 = n741 & ~n47235 ;
  assign n47237 = ~n47234 & n47236 ;
  assign n47238 = ~n941 & n25427 ;
  assign n47239 = ~n10506 & n47238 ;
  assign n47240 = n30464 ^ n4467 ^ 1'b0 ;
  assign n47241 = n20370 | n38089 ;
  assign n47243 = n23486 ^ n21325 ^ 1'b0 ;
  assign n47244 = n28020 & ~n47243 ;
  assign n47242 = n12703 ^ n3293 ^ n3033 ;
  assign n47245 = n47244 ^ n47242 ^ n9909 ;
  assign n47246 = n47241 | n47245 ;
  assign n47250 = n6186 & ~n28052 ;
  assign n47251 = n47250 ^ n17629 ^ 1'b0 ;
  assign n47252 = n9904 | n47251 ;
  assign n47247 = n40 | n18745 ;
  assign n47248 = n25296 & ~n47247 ;
  assign n47249 = ( n6948 & ~n8426 ) | ( n6948 & n47248 ) | ( ~n8426 & n47248 ) ;
  assign n47253 = n47252 ^ n47249 ^ 1'b0 ;
  assign n47254 = n27658 ^ n18063 ^ n17468 ;
  assign n47256 = n8296 ^ n7715 ^ n1801 ;
  assign n47255 = n514 & n8056 ;
  assign n47257 = n47256 ^ n47255 ^ 1'b0 ;
  assign n47258 = n47254 | n47257 ;
  assign n47259 = n28176 ^ n12782 ^ 1'b0 ;
  assign n47260 = ~n11706 & n16728 ;
  assign n47261 = n15009 ^ n4041 ^ 1'b0 ;
  assign n47262 = n47260 | n47261 ;
  assign n47263 = n25372 & ~n47262 ;
  assign n47264 = n2635 | n36052 ;
  assign n47265 = n2408 | n4074 ;
  assign n47266 = n2729 | n47265 ;
  assign n47267 = n47266 ^ n13791 ^ n589 ;
  assign n47268 = ~n4160 & n47267 ;
  assign n47269 = n47268 ^ n24762 ^ 1'b0 ;
  assign n47270 = n47269 ^ n37016 ^ n263 ;
  assign n47271 = ~n954 & n28342 ;
  assign n47272 = n19683 & n47271 ;
  assign n47273 = n33468 ^ n12536 ^ 1'b0 ;
  assign n47274 = n47272 | n47273 ;
  assign n47275 = n21740 & ~n47274 ;
  assign n47276 = n12874 & n42461 ;
  assign n47277 = n2174 & ~n47276 ;
  assign n47278 = n6339 | n41552 ;
  assign n47279 = n5706 & n47278 ;
  assign n47280 = n24716 ^ n1564 ^ 1'b0 ;
  assign n47281 = n47279 & ~n47280 ;
  assign n47282 = n4226 & n36885 ;
  assign n47283 = ~n29390 & n47282 ;
  assign n47284 = n6667 ^ n2466 ^ 1'b0 ;
  assign n47285 = ( n12789 & n28316 ) | ( n12789 & ~n47284 ) | ( n28316 & ~n47284 ) ;
  assign n47286 = n17296 ^ n12745 ^ n3221 ;
  assign n47287 = ( n7911 & n8032 ) | ( n7911 & n47286 ) | ( n8032 & n47286 ) ;
  assign n47288 = n46900 ^ n22281 ^ 1'b0 ;
  assign n47289 = n11706 & ~n20705 ;
  assign n47290 = n5535 & n47289 ;
  assign n47291 = n16865 & ~n34953 ;
  assign n47292 = n10040 & ~n47291 ;
  assign n47293 = n1801 & ~n24485 ;
  assign n47294 = n4772 & n47293 ;
  assign n47295 = ~n6759 & n47294 ;
  assign n47296 = ~n12443 & n17938 ;
  assign n47297 = n47295 & n47296 ;
  assign n47298 = n28388 ^ n51 ^ 1'b0 ;
  assign n47299 = n35137 | n47298 ;
  assign n47300 = n16094 ^ n5380 ^ 1'b0 ;
  assign n47301 = n26767 | n47300 ;
  assign n47302 = n6862 & n47301 ;
  assign n47303 = n17895 ^ n12413 ^ n3548 ;
  assign n47304 = n2414 & ~n7101 ;
  assign n47305 = n47304 ^ n5736 ^ 1'b0 ;
  assign n47306 = n8918 ^ n3342 ^ 1'b0 ;
  assign n47307 = n7761 & n47306 ;
  assign n47308 = n9785 & ~n30133 ;
  assign n47309 = ~n47307 & n47308 ;
  assign n47310 = n34825 ^ n11010 ^ n3351 ;
  assign n47311 = ( n24689 & ~n41253 ) | ( n24689 & n43638 ) | ( ~n41253 & n43638 ) ;
  assign n47312 = ( ~n5533 & n17576 ) | ( ~n5533 & n42565 ) | ( n17576 & n42565 ) ;
  assign n47313 = n22106 & n26849 ;
  assign n47314 = n47312 | n47313 ;
  assign n47315 = n19843 ^ n5484 ^ 1'b0 ;
  assign n47316 = n23200 & ~n47315 ;
  assign n47317 = n47314 | n47316 ;
  assign n47318 = n47317 ^ n33801 ^ 1'b0 ;
  assign n47319 = n27875 & n47318 ;
  assign n47320 = n28278 ^ n611 ^ 1'b0 ;
  assign n47321 = n25777 & n47320 ;
  assign n47322 = ~n16771 & n30292 ;
  assign n47323 = ~n1805 & n10902 ;
  assign n47324 = ~n8536 & n47323 ;
  assign n47325 = ( n16345 & ~n22315 ) | ( n16345 & n47000 ) | ( ~n22315 & n47000 ) ;
  assign n47326 = n11917 | n27632 ;
  assign n47327 = n47325 & ~n47326 ;
  assign n47328 = n5102 ^ n3420 ^ 1'b0 ;
  assign n47329 = n16476 & ~n47328 ;
  assign n47330 = n47329 ^ n1786 ^ 1'b0 ;
  assign n47331 = n47327 | n47330 ;
  assign n47332 = n14423 | n16801 ;
  assign n47333 = n47332 ^ n12082 ^ 1'b0 ;
  assign n47334 = n876 | n47333 ;
  assign n47335 = n14945 ^ n2794 ^ n280 ;
  assign n47336 = n47335 ^ n8247 ^ n2330 ;
  assign n47337 = n47 & ~n40473 ;
  assign n47338 = n47337 ^ n24463 ^ 1'b0 ;
  assign n47339 = n47338 ^ n31402 ^ 1'b0 ;
  assign n47340 = n40901 | n47339 ;
  assign n47341 = n18186 | n36320 ;
  assign n47342 = n23320 & ~n24658 ;
  assign n47343 = n47342 ^ n34601 ^ 1'b0 ;
  assign n47344 = n18071 | n47343 ;
  assign n47345 = n24105 ^ n18688 ^ n5185 ;
  assign n47346 = n5442 | n18473 ;
  assign n47347 = n1932 & ~n20961 ;
  assign n47348 = n47347 ^ n37716 ^ 1'b0 ;
  assign n47349 = n47348 ^ n21395 ^ 1'b0 ;
  assign n47350 = n1991 | n47349 ;
  assign n47351 = ~n102 & n47350 ;
  assign n47353 = n24365 ^ n23205 ^ 1'b0 ;
  assign n47352 = n26853 ^ n22721 ^ 1'b0 ;
  assign n47354 = n47353 ^ n47352 ^ n44601 ;
  assign n47355 = n17422 ^ n8615 ^ 1'b0 ;
  assign n47356 = n47355 ^ n40009 ^ n26872 ;
  assign n47357 = n42465 ^ n27097 ^ n9143 ;
  assign n47358 = n700 & n34901 ;
  assign n47359 = n34034 & n37582 ;
  assign n47360 = ~n40303 & n47359 ;
  assign n47361 = n16019 | n22909 ;
  assign n47362 = n47361 ^ n13361 ^ 1'b0 ;
  assign n47363 = n1817 & ~n26833 ;
  assign n47364 = n57 & n47363 ;
  assign n47365 = ~n21785 & n27586 ;
  assign n47366 = n25047 & n47365 ;
  assign n47367 = n47366 ^ n19197 ^ 1'b0 ;
  assign n47368 = n20494 ^ n7363 ^ n3856 ;
  assign n47369 = n8683 & ~n30391 ;
  assign n47370 = n11607 & ~n47369 ;
  assign n47371 = n47370 ^ n33844 ^ n16405 ;
  assign n47372 = n47368 & n47371 ;
  assign n47373 = n7607 ^ n2114 ^ 1'b0 ;
  assign n47374 = n8070 | n47373 ;
  assign n47375 = ( ~n1432 & n17890 ) | ( ~n1432 & n42534 ) | ( n17890 & n42534 ) ;
  assign n47376 = ~n59 & n17572 ;
  assign n47380 = n22315 & ~n24523 ;
  assign n47381 = n47380 ^ n16654 ^ 1'b0 ;
  assign n47382 = n38018 & ~n47381 ;
  assign n47383 = ( n8792 & n19372 ) | ( n8792 & n47382 ) | ( n19372 & n47382 ) ;
  assign n47377 = n14632 ^ n1661 ^ 1'b0 ;
  assign n47378 = n10764 | n47377 ;
  assign n47379 = n17121 | n47378 ;
  assign n47384 = n47383 ^ n47379 ^ 1'b0 ;
  assign n47385 = n18396 & n22360 ;
  assign n47386 = n10073 & ~n47385 ;
  assign n47387 = n2542 & ~n9667 ;
  assign n47388 = n47387 ^ n9849 ^ 1'b0 ;
  assign n47389 = n28430 | n42887 ;
  assign n47390 = n47389 ^ n8838 ^ 1'b0 ;
  assign n47391 = n47390 ^ n3971 ^ 1'b0 ;
  assign n47392 = ~n17171 & n29332 ;
  assign n47393 = n47391 & n47392 ;
  assign n47394 = n46285 ^ n18038 ^ 1'b0 ;
  assign n47395 = n23876 & ~n44987 ;
  assign n47396 = n47395 ^ n18681 ^ 1'b0 ;
  assign n47397 = n21532 | n47396 ;
  assign n47398 = ( ~n3087 & n39452 ) | ( ~n3087 & n47397 ) | ( n39452 & n47397 ) ;
  assign n47399 = ~n14030 & n40181 ;
  assign n47404 = n4633 & n5205 ;
  assign n47405 = n47404 ^ n4538 ^ 1'b0 ;
  assign n47402 = n20299 ^ n132 ^ 1'b0 ;
  assign n47403 = ~n4957 & n47402 ;
  assign n47406 = n47405 ^ n47403 ^ 1'b0 ;
  assign n47407 = n47406 ^ n45591 ^ n14290 ;
  assign n47400 = n7891 & n11700 ;
  assign n47401 = n47400 ^ n8209 ^ 1'b0 ;
  assign n47408 = n47407 ^ n47401 ^ 1'b0 ;
  assign n47409 = n38980 & n45997 ;
  assign n47410 = n9699 ^ n4445 ^ 1'b0 ;
  assign n47411 = ~n1604 & n5204 ;
  assign n47412 = n26132 ^ n17233 ^ 1'b0 ;
  assign n47413 = n35384 ^ n28333 ^ 1'b0 ;
  assign n47414 = n1577 & n47413 ;
  assign n47415 = n47414 ^ n2008 ^ 1'b0 ;
  assign n47416 = n40497 ^ n37864 ^ 1'b0 ;
  assign n47417 = ( ~n5793 & n6578 ) | ( ~n5793 & n47416 ) | ( n6578 & n47416 ) ;
  assign n47418 = n31399 ^ n10993 ^ 1'b0 ;
  assign n47419 = ( ~n27241 & n28634 ) | ( ~n27241 & n47418 ) | ( n28634 & n47418 ) ;
  assign n47420 = n22912 & n45075 ;
  assign n47421 = ~n30779 & n47420 ;
  assign n47422 = ~n13023 & n39378 ;
  assign n47423 = n7335 & n47422 ;
  assign n47424 = n20695 ^ n15022 ^ 1'b0 ;
  assign n47425 = n47423 | n47424 ;
  assign n47426 = n13737 & ~n22204 ;
  assign n47427 = n9314 & n47426 ;
  assign n47428 = ~n3170 & n47427 ;
  assign n47429 = n18371 & n47428 ;
  assign n47430 = n2646 | n15351 ;
  assign n47431 = n39860 & ~n47430 ;
  assign n47432 = n47431 ^ n9667 ^ 1'b0 ;
  assign n47433 = n23059 ^ n11433 ^ 1'b0 ;
  assign n47434 = ~n14576 & n15962 ;
  assign n47435 = n47433 & n47434 ;
  assign n47436 = n6365 | n20786 ;
  assign n47437 = n21881 & ~n30289 ;
  assign n47438 = n4563 & n47437 ;
  assign n47439 = n6614 ^ n1155 ^ 1'b0 ;
  assign n47440 = ~n42202 & n47439 ;
  assign n47441 = n4857 & n10411 ;
  assign n47442 = ( n15430 & n47440 ) | ( n15430 & n47441 ) | ( n47440 & n47441 ) ;
  assign n47444 = ( n624 & ~n1225 ) | ( n624 & n7446 ) | ( ~n1225 & n7446 ) ;
  assign n47443 = ~n14220 & n24771 ;
  assign n47445 = n47444 ^ n47443 ^ n4377 ;
  assign n47446 = n30812 ^ n15154 ^ 1'b0 ;
  assign n47447 = n47446 ^ n41588 ^ 1'b0 ;
  assign n47448 = n33566 ^ n21607 ^ n6895 ;
  assign n47449 = n32806 & n47448 ;
  assign n47450 = n18015 ^ n2667 ^ 1'b0 ;
  assign n47451 = n5768 & n22668 ;
  assign n47452 = n47451 ^ n20064 ^ 1'b0 ;
  assign n47453 = n47450 & ~n47452 ;
  assign n47454 = n14418 ^ n4588 ^ 1'b0 ;
  assign n47455 = n14013 & ~n47454 ;
  assign n47456 = n46694 ^ n18080 ^ 1'b0 ;
  assign n47457 = n28503 ^ n14851 ^ n7539 ;
  assign n47458 = n47457 ^ n47080 ^ n14826 ;
  assign n47459 = ~n2138 & n3898 ;
  assign n47460 = ~n3441 & n12787 ;
  assign n47462 = n46295 ^ n31663 ^ n3790 ;
  assign n47461 = n12112 | n42576 ;
  assign n47463 = n47462 ^ n47461 ^ 1'b0 ;
  assign n47464 = n11157 ^ n734 ^ 1'b0 ;
  assign n47465 = n31377 & n47464 ;
  assign n47466 = n19066 | n20798 ;
  assign n47467 = n47465 | n47466 ;
  assign n47468 = ~n496 & n18532 ;
  assign n47469 = n47468 ^ n34114 ^ 1'b0 ;
  assign n47470 = ( n310 & n25150 ) | ( n310 & n47469 ) | ( n25150 & n47469 ) ;
  assign n47471 = n47470 ^ n40390 ^ n3020 ;
  assign n47472 = ( ~n2076 & n19829 ) | ( ~n2076 & n33275 ) | ( n19829 & n33275 ) ;
  assign n47473 = n31788 ^ n10217 ^ 1'b0 ;
  assign n47474 = n47472 | n47473 ;
  assign n47475 = n7666 & n47474 ;
  assign n47476 = n8635 ^ n2858 ^ 1'b0 ;
  assign n47477 = n3636 | n32981 ;
  assign n47478 = n47477 ^ n43392 ^ 1'b0 ;
  assign n47479 = ~n8442 & n11529 ;
  assign n47480 = n47479 ^ n31469 ^ 1'b0 ;
  assign n47481 = n33342 ^ n20368 ^ 1'b0 ;
  assign n47482 = n15678 | n47481 ;
  assign n47483 = n47482 ^ n35413 ^ 1'b0 ;
  assign n47484 = n33773 ^ n25181 ^ 1'b0 ;
  assign n47485 = n47484 ^ n37442 ^ n32584 ;
  assign n47486 = n8504 ^ n969 ^ 1'b0 ;
  assign n47487 = ~n2759 & n47486 ;
  assign n47488 = n31687 ^ n28850 ^ n8707 ;
  assign n47489 = n31392 ^ n16415 ^ 1'b0 ;
  assign n47490 = ~n4823 & n29318 ;
  assign n47491 = ( n47488 & ~n47489 ) | ( n47488 & n47490 ) | ( ~n47489 & n47490 ) ;
  assign n47492 = n47487 | n47491 ;
  assign n47493 = ~n10215 & n25611 ;
  assign n47494 = n47493 ^ n26600 ^ 1'b0 ;
  assign n47495 = n22840 ^ n12675 ^ 1'b0 ;
  assign n47496 = n37861 & n47495 ;
  assign n47497 = ~n7756 & n9549 ;
  assign n47498 = ~n28339 & n47497 ;
  assign n47499 = n3776 | n47498 ;
  assign n47500 = n34498 | n47499 ;
  assign n47502 = n3410 & n17214 ;
  assign n47503 = n47502 ^ n40338 ^ 1'b0 ;
  assign n47501 = n25808 | n34689 ;
  assign n47504 = n47503 ^ n47501 ^ 1'b0 ;
  assign n47505 = n30032 ^ n18263 ^ 1'b0 ;
  assign n47506 = ( n30617 & ~n37562 ) | ( n30617 & n47505 ) | ( ~n37562 & n47505 ) ;
  assign n47507 = n8088 ^ n5199 ^ n1197 ;
  assign n47508 = n47507 ^ n473 ^ 1'b0 ;
  assign n47509 = ( n11901 & n15975 ) | ( n11901 & ~n47508 ) | ( n15975 & ~n47508 ) ;
  assign n47510 = n24193 ^ n8462 ^ 1'b0 ;
  assign n47511 = n26206 ^ n3949 ^ 1'b0 ;
  assign n47512 = n3750 & n47511 ;
  assign n47513 = n41066 ^ n20092 ^ 1'b0 ;
  assign n47514 = n27224 | n47513 ;
  assign n47515 = n3421 ^ n3043 ^ 1'b0 ;
  assign n47516 = ~n11488 & n47515 ;
  assign n47517 = ( n2830 & ~n16996 ) | ( n2830 & n23238 ) | ( ~n16996 & n23238 ) ;
  assign n47518 = n12747 & n13952 ;
  assign n47519 = ~n16297 & n33638 ;
  assign n47520 = ~n32419 & n47519 ;
  assign n47521 = n47520 ^ n21206 ^ 1'b0 ;
  assign n47522 = n1122 & n42022 ;
  assign n47523 = n11704 & ~n37016 ;
  assign n47524 = n47523 ^ n47455 ^ 1'b0 ;
  assign n47525 = n3241 | n34408 ;
  assign n47526 = ( n8790 & n25851 ) | ( n8790 & ~n42545 ) | ( n25851 & ~n42545 ) ;
  assign n47527 = ( n6262 & ~n19354 ) | ( n6262 & n47526 ) | ( ~n19354 & n47526 ) ;
  assign n47528 = n39232 & ~n47527 ;
  assign n47529 = n349 | n14566 ;
  assign n47530 = n26886 ^ n13316 ^ n12239 ;
  assign n47531 = n3979 & n22025 ;
  assign n47532 = n28285 & ~n47531 ;
  assign n47533 = n15249 & n22993 ;
  assign n47534 = n29341 & ~n39377 ;
  assign n47535 = n24262 & n47534 ;
  assign n47536 = ~n13958 & n15562 ;
  assign n47537 = n185 | n47536 ;
  assign n47538 = n47537 ^ n18257 ^ 1'b0 ;
  assign n47539 = n44085 ^ n21167 ^ 1'b0 ;
  assign n47540 = n47538 & n47539 ;
  assign n47541 = n19559 ^ n13502 ^ 1'b0 ;
  assign n47542 = ~n29746 & n36856 ;
  assign n47543 = n8740 & n17380 ;
  assign n47544 = n394 & ~n47543 ;
  assign n47545 = n18971 & n47544 ;
  assign n47546 = n431 | n18085 ;
  assign n47547 = ~n23992 & n47546 ;
  assign n47548 = n47547 ^ n27533 ^ 1'b0 ;
  assign n47549 = ( ~n14752 & n18299 ) | ( ~n14752 & n47548 ) | ( n18299 & n47548 ) ;
  assign n47550 = n37510 ^ n6096 ^ 1'b0 ;
  assign n47551 = n47550 ^ n39989 ^ 1'b0 ;
  assign n47552 = n14385 & n46630 ;
  assign n47553 = n47552 ^ n31786 ^ 1'b0 ;
  assign n47554 = ~n36539 & n47553 ;
  assign n47555 = n26994 ^ n10669 ^ n8483 ;
  assign n47556 = n2991 & n47555 ;
  assign n47557 = n29944 & n47556 ;
  assign n47558 = n6307 | n26540 ;
  assign n47559 = ( ~n15923 & n26850 ) | ( ~n15923 & n32820 ) | ( n26850 & n32820 ) ;
  assign n47560 = n17675 & n47559 ;
  assign n47561 = n27786 ^ n12682 ^ n11410 ;
  assign n47562 = ( ~n32148 & n39651 ) | ( ~n32148 & n47561 ) | ( n39651 & n47561 ) ;
  assign n47563 = ( n2650 & n33640 ) | ( n2650 & n37124 ) | ( n33640 & n37124 ) ;
  assign n47564 = n26152 ^ n10673 ^ 1'b0 ;
  assign n47565 = n47564 ^ n5323 ^ n2288 ;
  assign n47566 = n23900 | n42179 ;
  assign n47567 = n34521 ^ n226 ^ 1'b0 ;
  assign n47568 = n3428 & ~n47567 ;
  assign n47569 = n17800 ^ n14335 ^ 1'b0 ;
  assign n47570 = ~n19270 & n24934 ;
  assign n47571 = n47570 ^ n14032 ^ 1'b0 ;
  assign n47572 = n27912 ^ n3181 ^ n2463 ;
  assign n47573 = n47572 ^ n5678 ^ 1'b0 ;
  assign n47574 = ~n30105 & n47446 ;
  assign n47575 = n23015 ^ n7749 ^ 1'b0 ;
  assign n47576 = n19209 | n47575 ;
  assign n47577 = n24744 ^ n17698 ^ 1'b0 ;
  assign n47578 = n1364 & ~n47577 ;
  assign n47579 = n24869 & n28965 ;
  assign n47580 = n47358 | n47579 ;
  assign n47581 = n1212 & n18017 ;
  assign n47582 = ~n2230 & n47581 ;
  assign n47583 = n10670 & ~n47582 ;
  assign n47584 = ~n14363 & n47583 ;
  assign n47585 = n11698 & ~n43704 ;
  assign n47586 = n47585 ^ n46158 ^ 1'b0 ;
  assign n47587 = n8701 & n12748 ;
  assign n47588 = n23674 ^ n23662 ^ n22052 ;
  assign n47589 = n47555 ^ n20623 ^ 1'b0 ;
  assign n47590 = n38645 & ~n47589 ;
  assign n47592 = ~n3540 & n6235 ;
  assign n47591 = n6731 | n17837 ;
  assign n47593 = n47592 ^ n47591 ^ 1'b0 ;
  assign n47594 = n15608 | n47593 ;
  assign n47595 = n21212 | n47594 ;
  assign n47596 = n990 & n3413 ;
  assign n47597 = n20013 ^ n14227 ^ 1'b0 ;
  assign n47598 = n47596 & n47597 ;
  assign n47600 = n115 & ~n26572 ;
  assign n47599 = n46868 ^ n25672 ^ n19305 ;
  assign n47601 = n47600 ^ n47599 ^ 1'b0 ;
  assign n47602 = n10587 | n11891 ;
  assign n47603 = n9984 | n39838 ;
  assign n47604 = ~n4845 & n13533 ;
  assign n47605 = n47604 ^ n24397 ^ 1'b0 ;
  assign n47606 = n11648 & n45663 ;
  assign n47607 = n47606 ^ n30439 ^ 1'b0 ;
  assign n47608 = n6568 & ~n8427 ;
  assign n47609 = n47608 ^ n7150 ^ 1'b0 ;
  assign n47610 = n12175 & ~n26351 ;
  assign n47611 = n47610 ^ n4799 ^ 1'b0 ;
  assign n47612 = ~n11226 & n47611 ;
  assign n47613 = ~n5350 & n47612 ;
  assign n47614 = ~n594 & n2030 ;
  assign n47615 = n39318 ^ n5135 ^ 1'b0 ;
  assign n47616 = n8119 | n30035 ;
  assign n47617 = n47616 ^ n23520 ^ 1'b0 ;
  assign n47618 = n10962 & n47617 ;
  assign n47619 = ~n2553 & n14104 ;
  assign n47620 = n47619 ^ n15663 ^ 1'b0 ;
  assign n47621 = ~n22099 & n47620 ;
  assign n47622 = n6131 & n25711 ;
  assign n47623 = n47622 ^ n2735 ^ 1'b0 ;
  assign n47624 = ~n6377 & n31026 ;
  assign n47625 = n47624 ^ n1185 ^ 1'b0 ;
  assign n47626 = n30208 | n47625 ;
  assign n47627 = n1789 & ~n47626 ;
  assign n47628 = n24123 ^ n5357 ^ 1'b0 ;
  assign n47629 = n20693 & n22213 ;
  assign n47630 = ( n20343 & n47628 ) | ( n20343 & ~n47629 ) | ( n47628 & ~n47629 ) ;
  assign n47631 = n19837 ^ n11363 ^ 1'b0 ;
  assign n47632 = ~n1093 & n22723 ;
  assign n47633 = n47632 ^ n9674 ^ 1'b0 ;
  assign n47634 = n459 & ~n15647 ;
  assign n47635 = n242 & n47634 ;
  assign n47636 = ~n39227 & n47635 ;
  assign n47637 = n1209 & ~n22526 ;
  assign n47638 = ( n6613 & ~n15276 ) | ( n6613 & n19884 ) | ( ~n15276 & n19884 ) ;
  assign n47639 = n17825 & n19815 ;
  assign n47640 = n448 | n16459 ;
  assign n47641 = ( n9255 & n21706 ) | ( n9255 & ~n47640 ) | ( n21706 & ~n47640 ) ;
  assign n47642 = ( n403 & ~n47639 ) | ( n403 & n47641 ) | ( ~n47639 & n47641 ) ;
  assign n47643 = ( ~n9330 & n21228 ) | ( ~n9330 & n26453 ) | ( n21228 & n26453 ) ;
  assign n47644 = n2128 & n13943 ;
  assign n47645 = n25383 ^ n16766 ^ 1'b0 ;
  assign n47646 = ( n257 & n5873 ) | ( n257 & ~n10159 ) | ( n5873 & ~n10159 ) ;
  assign n47647 = n13275 & ~n34774 ;
  assign n47648 = n47646 & n47647 ;
  assign n47651 = ~n24670 & n42368 ;
  assign n47649 = n35269 ^ n16771 ^ 1'b0 ;
  assign n47650 = n21160 | n47649 ;
  assign n47652 = n47651 ^ n47650 ^ 1'b0 ;
  assign n47653 = ( n2231 & n4333 ) | ( n2231 & ~n10178 ) | ( n4333 & ~n10178 ) ;
  assign n47654 = n462 & n10308 ;
  assign n47655 = n5164 & n47654 ;
  assign n47656 = n47655 ^ n16697 ^ n14487 ;
  assign n47657 = ( n533 & ~n4948 ) | ( n533 & n47656 ) | ( ~n4948 & n47656 ) ;
  assign n47658 = ~n7583 & n23605 ;
  assign n47659 = n47658 ^ n11991 ^ 1'b0 ;
  assign n47660 = n7129 & n47659 ;
  assign n47661 = ( n26997 & n43195 ) | ( n26997 & ~n47660 ) | ( n43195 & ~n47660 ) ;
  assign n47662 = n14192 ^ n14049 ^ 1'b0 ;
  assign n47663 = n5655 | n47662 ;
  assign n47664 = n37234 & ~n47663 ;
  assign n47665 = n10329 | n24331 ;
  assign n47666 = n14228 | n47665 ;
  assign n47667 = n22707 ^ n20250 ^ n2710 ;
  assign n47668 = ~n1357 & n17656 ;
  assign n47669 = n47668 ^ n23189 ^ 1'b0 ;
  assign n47670 = n47667 & ~n47669 ;
  assign n47671 = ~n37990 & n47670 ;
  assign n47672 = ( n22524 & n29366 ) | ( n22524 & n45449 ) | ( n29366 & n45449 ) ;
  assign n47673 = n43549 & ~n47672 ;
  assign n47674 = ( n9996 & ~n21062 ) | ( n9996 & n45997 ) | ( ~n21062 & n45997 ) ;
  assign n47675 = n14744 ^ n13589 ^ 1'b0 ;
  assign n47676 = n8672 & ~n12530 ;
  assign n47677 = n43458 ^ n13082 ^ n5129 ;
  assign n47678 = n38655 & ~n47677 ;
  assign n47679 = n47678 ^ n3179 ^ 1'b0 ;
  assign n47680 = n5827 | n47679 ;
  assign n47681 = ~n1462 & n14520 ;
  assign n47682 = n30516 & ~n47681 ;
  assign n47683 = n10519 & n47682 ;
  assign n47684 = n5990 & ~n10167 ;
  assign n47685 = n47684 ^ n9191 ^ 1'b0 ;
  assign n47686 = n47685 ^ n12481 ^ 1'b0 ;
  assign n47687 = n30156 | n47686 ;
  assign n47691 = n16124 & ~n23780 ;
  assign n47690 = ~n10560 & n32554 ;
  assign n47692 = n47691 ^ n47690 ^ 1'b0 ;
  assign n47688 = n82 | n30970 ;
  assign n47689 = n37336 | n47688 ;
  assign n47693 = n47692 ^ n47689 ^ 1'b0 ;
  assign n47694 = n15420 ^ n14766 ^ n7080 ;
  assign n47695 = n8975 & n47694 ;
  assign n47696 = n10444 & ~n32845 ;
  assign n47697 = n12018 & n47696 ;
  assign n47698 = ~n18297 & n47697 ;
  assign n47699 = ( n10444 & n16966 ) | ( n10444 & ~n28743 ) | ( n16966 & ~n28743 ) ;
  assign n47700 = n42829 ^ n8157 ^ 1'b0 ;
  assign n47701 = n20220 & n47700 ;
  assign n47702 = n47701 ^ n7498 ^ 1'b0 ;
  assign n47703 = n6396 & ~n27816 ;
  assign n47704 = n27816 & n47703 ;
  assign n47705 = n19597 | n47704 ;
  assign n47706 = n47704 & ~n47705 ;
  assign n47707 = n35956 ^ n3932 ^ 1'b0 ;
  assign n47708 = n12826 & ~n19368 ;
  assign n47709 = n23132 & n47708 ;
  assign n47710 = n7904 | n23515 ;
  assign n47711 = n34938 | n47710 ;
  assign n47712 = n20726 ^ n14972 ^ 1'b0 ;
  assign n47713 = ( n12241 & n25540 ) | ( n12241 & n44846 ) | ( n25540 & n44846 ) ;
  assign n47714 = n684 | n46607 ;
  assign n47715 = n6104 ^ n3908 ^ 1'b0 ;
  assign n47716 = n38223 ^ n21868 ^ 1'b0 ;
  assign n47717 = ~n47715 & n47716 ;
  assign n47718 = n35080 ^ n17217 ^ 1'b0 ;
  assign n47719 = ~n5338 & n33253 ;
  assign n47720 = n17880 ^ n8494 ^ 1'b0 ;
  assign n47721 = n639 | n35195 ;
  assign n47722 = n27247 ^ n16375 ^ 1'b0 ;
  assign n47723 = n14213 & ~n47722 ;
  assign n47724 = n45865 ^ n180 ^ 1'b0 ;
  assign n47725 = ~n20079 & n47724 ;
  assign n47726 = ( n3856 & n18825 ) | ( n3856 & ~n30009 ) | ( n18825 & ~n30009 ) ;
  assign n47727 = n16935 | n47726 ;
  assign n47728 = n47727 ^ n16378 ^ 1'b0 ;
  assign n47729 = ( n965 & n9321 ) | ( n965 & n17147 ) | ( n9321 & n17147 ) ;
  assign n47730 = ( ~n5128 & n12664 ) | ( ~n5128 & n47729 ) | ( n12664 & n47729 ) ;
  assign n47731 = n47730 ^ n15240 ^ 1'b0 ;
  assign n47732 = n15651 | n28548 ;
  assign n47733 = n47732 ^ n6879 ^ 1'b0 ;
  assign n47734 = n47205 ^ n706 ^ 1'b0 ;
  assign n47735 = n25100 & n47734 ;
  assign n47736 = ~n47733 & n47735 ;
  assign n47737 = n47736 ^ n47416 ^ 1'b0 ;
  assign n47738 = n15904 ^ n1231 ^ 1'b0 ;
  assign n47739 = n11971 & ~n46812 ;
  assign n47740 = n47738 & n47739 ;
  assign n47741 = ~n15555 & n32060 ;
  assign n47742 = ~n12021 & n47741 ;
  assign n47743 = n47742 ^ n17753 ^ 1'b0 ;
  assign n47744 = n4023 | n5781 ;
  assign n47745 = n47744 ^ n27237 ^ 1'b0 ;
  assign n47746 = n47745 ^ n19237 ^ n536 ;
  assign n47747 = ( ~n732 & n4948 ) | ( ~n732 & n20339 ) | ( n4948 & n20339 ) ;
  assign n47748 = n47747 ^ n32470 ^ n6807 ;
  assign n47749 = n18444 & n31904 ;
  assign n47750 = n45207 | n47749 ;
  assign n47751 = n36288 | n47750 ;
  assign n47752 = ~n28520 & n47751 ;
  assign n47753 = n47752 ^ n13325 ^ 1'b0 ;
  assign n47754 = n14677 | n16005 ;
  assign n47755 = n21478 | n47754 ;
  assign n47756 = n18913 | n47755 ;
  assign n47758 = n7005 & n10568 ;
  assign n47757 = n11867 & n15166 ;
  assign n47759 = n47758 ^ n47757 ^ 1'b0 ;
  assign n47765 = n16305 ^ n926 ^ 1'b0 ;
  assign n47766 = n27917 & n47765 ;
  assign n47767 = ~n5793 & n47766 ;
  assign n47760 = n490 & n7193 ;
  assign n47761 = ~n1357 & n47760 ;
  assign n47762 = n3087 | n47761 ;
  assign n47763 = n19767 & ~n47762 ;
  assign n47764 = n9109 & ~n47763 ;
  assign n47768 = n47767 ^ n47764 ^ 1'b0 ;
  assign n47769 = n4072 ^ n490 ^ 1'b0 ;
  assign n47770 = n47769 ^ n10897 ^ 1'b0 ;
  assign n47771 = n43347 ^ n40088 ^ 1'b0 ;
  assign n47772 = n47770 | n47771 ;
  assign n47773 = n21815 | n31293 ;
  assign n47774 = ( n521 & n8811 ) | ( n521 & ~n47773 ) | ( n8811 & ~n47773 ) ;
  assign n47775 = n14033 ^ n8035 ^ n4318 ;
  assign n47776 = n14634 ^ n10501 ^ 1'b0 ;
  assign n47777 = n12477 | n47776 ;
  assign n47778 = ( n1155 & n15012 ) | ( n1155 & n47777 ) | ( n15012 & n47777 ) ;
  assign n47779 = n32429 & n47014 ;
  assign n47780 = ( ~n11209 & n12482 ) | ( ~n11209 & n16316 ) | ( n12482 & n16316 ) ;
  assign n47781 = n29663 ^ n18010 ^ 1'b0 ;
  assign n47782 = ~n47780 & n47781 ;
  assign n47783 = ( n11439 & ~n12866 ) | ( n11439 & n32790 ) | ( ~n12866 & n32790 ) ;
  assign n47784 = n44217 ^ n42968 ^ n25823 ;
  assign n47785 = n6978 & ~n13485 ;
  assign n47786 = ~n21007 & n47785 ;
  assign n47787 = n15984 ^ n15573 ^ 1'b0 ;
  assign n47788 = ~n15592 & n47787 ;
  assign n47789 = n15271 & ~n47788 ;
  assign n47790 = n18029 ^ n12181 ^ 1'b0 ;
  assign n47791 = n1775 | n47790 ;
  assign n47792 = n14510 ^ n2826 ^ 1'b0 ;
  assign n47793 = n11560 | n27285 ;
  assign n47794 = n47793 ^ n1983 ^ 1'b0 ;
  assign n47795 = n37149 ^ n19324 ^ n11473 ;
  assign n47796 = n22298 ^ n4336 ^ 1'b0 ;
  assign n47797 = n5825 | n47796 ;
  assign n47798 = n47797 ^ n4743 ^ n4010 ;
  assign n47799 = ~n2375 & n5436 ;
  assign n47800 = n8213 & n47799 ;
  assign n47801 = n16482 ^ n5331 ^ 1'b0 ;
  assign n47802 = n8532 ^ n6969 ^ 1'b0 ;
  assign n47803 = ~n15742 & n47802 ;
  assign n47804 = n47801 & ~n47803 ;
  assign n47805 = ~n47800 & n47804 ;
  assign n47806 = n17991 ^ n10387 ^ 1'b0 ;
  assign n47807 = n17450 & ~n47806 ;
  assign n47808 = n21254 ^ n20767 ^ 1'b0 ;
  assign n47809 = n33398 ^ n19510 ^ n2143 ;
  assign n47810 = n47809 ^ n15560 ^ 1'b0 ;
  assign n47811 = n35366 & ~n47810 ;
  assign n47812 = ( n24296 & ~n47808 ) | ( n24296 & n47811 ) | ( ~n47808 & n47811 ) ;
  assign n47813 = ~n21773 & n22277 ;
  assign n47814 = n47813 ^ n30944 ^ n10885 ;
  assign n47815 = n47814 ^ n1990 ^ 1'b0 ;
  assign n47816 = ( n8574 & n11025 ) | ( n8574 & n23317 ) | ( n11025 & n23317 ) ;
  assign n47819 = n4986 ^ n1154 ^ 1'b0 ;
  assign n47820 = ~n22084 & n47819 ;
  assign n47817 = n20836 & n37266 ;
  assign n47818 = n47817 ^ n14229 ^ 1'b0 ;
  assign n47821 = n47820 ^ n47818 ^ 1'b0 ;
  assign n47822 = n7996 ^ n2385 ^ 1'b0 ;
  assign n47823 = n4497 & ~n47822 ;
  assign n47824 = n5954 & ~n47823 ;
  assign n47825 = n47824 ^ n9923 ^ 1'b0 ;
  assign n47826 = n12252 & ~n13991 ;
  assign n47827 = n10597 & n47826 ;
  assign n47828 = n44362 & n47827 ;
  assign n47829 = n47828 ^ n36417 ^ 1'b0 ;
  assign n47830 = n47825 & ~n47829 ;
  assign n47831 = n24681 ^ n11346 ^ 1'b0 ;
  assign n47832 = n25622 & ~n47831 ;
  assign n47833 = ~n33304 & n45851 ;
  assign n47834 = n47833 ^ n36389 ^ 1'b0 ;
  assign n47835 = ~n10049 & n15372 ;
  assign n47836 = n30422 & n47835 ;
  assign n47837 = n6713 & n42503 ;
  assign n47838 = n46317 ^ n21898 ^ n11529 ;
  assign n47839 = n4795 | n11986 ;
  assign n47840 = n283 & ~n47839 ;
  assign n47841 = n47840 ^ n30636 ^ 1'b0 ;
  assign n47842 = ( n12588 & n36853 ) | ( n12588 & ~n47841 ) | ( n36853 & ~n47841 ) ;
  assign n47843 = n28146 ^ n5311 ^ 1'b0 ;
  assign n47844 = ~n18039 & n47843 ;
  assign n47845 = n2775 & n4845 ;
  assign n47846 = n47845 ^ n192 ^ 1'b0 ;
  assign n47847 = n47846 ^ n2718 ^ 1'b0 ;
  assign n47848 = n5617 & n47847 ;
  assign n47849 = n4803 & n38373 ;
  assign n47850 = n47849 ^ n38172 ^ 1'b0 ;
  assign n47851 = ~n2612 & n3580 ;
  assign n47852 = n47851 ^ n4703 ^ 1'b0 ;
  assign n47853 = n47852 ^ n44358 ^ 1'b0 ;
  assign n47854 = ~n28640 & n47853 ;
  assign n47855 = n42016 ^ n38380 ^ n27499 ;
  assign n47856 = ~n9901 & n25308 ;
  assign n47857 = n15849 & n47856 ;
  assign n47858 = n29962 ^ n29634 ^ 1'b0 ;
  assign n47859 = ~n9255 & n44649 ;
  assign n47860 = ~n47858 & n47859 ;
  assign n47861 = n4364 & n35527 ;
  assign n47862 = n26259 & n47861 ;
  assign n47863 = ( ~n859 & n12126 ) | ( ~n859 & n18866 ) | ( n12126 & n18866 ) ;
  assign n47864 = n36776 ^ n11567 ^ n9517 ;
  assign n47865 = n47863 & ~n47864 ;
  assign n47866 = n10383 & n12441 ;
  assign n47867 = ~n46599 & n47866 ;
  assign n47868 = ( n9838 & n19248 ) | ( n9838 & ~n43756 ) | ( n19248 & ~n43756 ) ;
  assign n47869 = n65 & n39831 ;
  assign n47870 = n47869 ^ n23032 ^ n2861 ;
  assign n47871 = n38393 ^ n10238 ^ 1'b0 ;
  assign n47872 = n28025 & ~n37661 ;
  assign n47873 = ( n3170 & n47871 ) | ( n3170 & n47872 ) | ( n47871 & n47872 ) ;
  assign n47874 = n39548 ^ n19344 ^ 1'b0 ;
  assign n47875 = n16497 & n31655 ;
  assign n47876 = ~n4804 & n47875 ;
  assign n47877 = n1666 | n47876 ;
  assign n47878 = n47877 ^ n8376 ^ 1'b0 ;
  assign n47879 = n7171 & ~n10745 ;
  assign n47880 = n47879 ^ n7550 ^ 1'b0 ;
  assign n47881 = ( ~n3581 & n18664 ) | ( ~n3581 & n47880 ) | ( n18664 & n47880 ) ;
  assign n47882 = ~n6827 & n47881 ;
  assign n47883 = n11871 & n13946 ;
  assign n47884 = n46202 ^ n36734 ^ 1'b0 ;
  assign n47885 = n11890 ^ n9860 ^ 1'b0 ;
  assign n47886 = n45198 ^ n24135 ^ 1'b0 ;
  assign n47887 = n7072 & ~n15909 ;
  assign n47888 = n23083 ^ n14403 ^ n4115 ;
  assign n47889 = n28255 | n47888 ;
  assign n47890 = n15140 & ~n22353 ;
  assign n47891 = n47890 ^ n33210 ^ 1'b0 ;
  assign n47892 = n5053 | n47891 ;
  assign n47893 = n47892 ^ n12468 ^ n10555 ;
  assign n47894 = n16863 & ~n24513 ;
  assign n47895 = ~n9160 & n47894 ;
  assign n47896 = n47895 ^ n29809 ^ n20795 ;
  assign n47897 = n11329 ^ n3833 ^ 1'b0 ;
  assign n47898 = ~n2596 & n28540 ;
  assign n47899 = ~n28029 & n28582 ;
  assign n47901 = n884 & n8403 ;
  assign n47900 = n17812 & ~n30996 ;
  assign n47902 = n47901 ^ n47900 ^ 1'b0 ;
  assign n47903 = ~n7399 & n12761 ;
  assign n47906 = n36144 ^ n27969 ^ 1'b0 ;
  assign n47907 = n39908 | n47906 ;
  assign n47904 = n41971 ^ n18052 ^ 1'b0 ;
  assign n47905 = ~n18351 & n47904 ;
  assign n47908 = n47907 ^ n47905 ^ 1'b0 ;
  assign n47909 = n8355 ^ n3526 ^ n2118 ;
  assign n47910 = n12353 ^ n3704 ^ 1'b0 ;
  assign n47911 = n47909 & n47910 ;
  assign n47912 = n47911 ^ n26794 ^ n3985 ;
  assign n47913 = ( n13677 & n47908 ) | ( n13677 & n47912 ) | ( n47908 & n47912 ) ;
  assign n47914 = ( ~n3140 & n23690 ) | ( ~n3140 & n34856 ) | ( n23690 & n34856 ) ;
  assign n47915 = ~n4114 & n47914 ;
  assign n47916 = n29991 ^ n10414 ^ 1'b0 ;
  assign n47917 = n26478 & n30520 ;
  assign n47918 = n30182 & n47917 ;
  assign n47919 = n37454 ^ n35437 ^ n420 ;
  assign n47920 = n47919 ^ n17440 ^ 1'b0 ;
  assign n47921 = ~n26148 & n47920 ;
  assign n47922 = n43592 ^ n15489 ^ 1'b0 ;
  assign n47923 = n31155 & ~n47922 ;
  assign n47924 = n12314 & n47923 ;
  assign n47925 = n14934 & ~n26126 ;
  assign n47926 = n42707 ^ n29778 ^ 1'b0 ;
  assign n47927 = n2784 | n6226 ;
  assign n47928 = n9117 | n47927 ;
  assign n47929 = n8736 & ~n34843 ;
  assign n47930 = n9717 | n47929 ;
  assign n47931 = n47928 | n47930 ;
  assign n47932 = ( ~n34891 & n35346 ) | ( ~n34891 & n47931 ) | ( n35346 & n47931 ) ;
  assign n47933 = ~n18945 & n38683 ;
  assign n47934 = n47933 ^ n9462 ^ 1'b0 ;
  assign n47935 = ( n11236 & ~n42989 ) | ( n11236 & n47934 ) | ( ~n42989 & n47934 ) ;
  assign n47936 = ~n19826 & n30470 ;
  assign n47937 = n6257 | n29117 ;
  assign n47938 = n6257 & ~n47937 ;
  assign n47939 = ( n27807 & n31634 ) | ( n27807 & ~n47938 ) | ( n31634 & ~n47938 ) ;
  assign n47940 = ( ~n1408 & n2580 ) | ( ~n1408 & n44068 ) | ( n2580 & n44068 ) ;
  assign n47941 = n5066 & ~n47940 ;
  assign n47942 = ~n47939 & n47941 ;
  assign n47943 = n15670 & ~n29648 ;
  assign n47944 = ~n20674 & n47943 ;
  assign n47945 = ~n44127 & n47944 ;
  assign n47946 = ~n14684 & n38271 ;
  assign n47947 = ~n1439 & n16288 ;
  assign n47951 = n16196 ^ n12113 ^ n8590 ;
  assign n47948 = n43223 ^ n16171 ^ 1'b0 ;
  assign n47949 = n47948 ^ n22104 ^ n11930 ;
  assign n47950 = ( n26360 & n45816 ) | ( n26360 & ~n47949 ) | ( n45816 & ~n47949 ) ;
  assign n47952 = n47951 ^ n47950 ^ 1'b0 ;
  assign n47953 = n36302 ^ n25671 ^ 1'b0 ;
  assign n47954 = n37309 ^ n27408 ^ 1'b0 ;
  assign n47955 = ( n2696 & n4545 ) | ( n2696 & n12317 ) | ( n4545 & n12317 ) ;
  assign n47956 = n1995 & n19727 ;
  assign n47957 = n7998 & n47956 ;
  assign n47958 = ( n31910 & n47955 ) | ( n31910 & n47957 ) | ( n47955 & n47957 ) ;
  assign n47963 = n7433 ^ n4701 ^ n1781 ;
  assign n47964 = n32861 & ~n47963 ;
  assign n47959 = n27805 ^ n8828 ^ 1'b0 ;
  assign n47960 = n11447 | n47959 ;
  assign n47961 = n19256 & ~n47960 ;
  assign n47962 = n44951 & n47961 ;
  assign n47965 = n47964 ^ n47962 ^ n17521 ;
  assign n47966 = n39341 ^ n33402 ^ n10002 ;
  assign n47967 = n25604 & n26669 ;
  assign n47968 = n19868 | n36019 ;
  assign n47969 = n37733 | n47968 ;
  assign n47970 = n39227 & n47056 ;
  assign n47974 = n12617 & n14296 ;
  assign n47971 = n29523 ^ n6139 ^ n2896 ;
  assign n47972 = n23067 ^ n3730 ^ 1'b0 ;
  assign n47973 = n47971 & ~n47972 ;
  assign n47975 = n47974 ^ n47973 ^ n13825 ;
  assign n47976 = n47975 ^ n12629 ^ 1'b0 ;
  assign n47977 = n2845 & ~n27641 ;
  assign n47978 = n22193 & n47977 ;
  assign n47979 = ~n1727 & n35004 ;
  assign n47980 = n34087 ^ n5994 ^ n1028 ;
  assign n47981 = n31717 & ~n35935 ;
  assign n47982 = n7873 | n30153 ;
  assign n47983 = ~n8523 & n47982 ;
  assign n47984 = n47983 ^ n19005 ^ 1'b0 ;
  assign n47985 = n1642 ^ n1355 ^ 1'b0 ;
  assign n47986 = n8128 & n47985 ;
  assign n47987 = n47986 ^ n38127 ^ n4769 ;
  assign n47988 = ~n14067 & n42669 ;
  assign n47989 = ~n18675 & n45222 ;
  assign n47990 = n22575 ^ n10318 ^ 1'b0 ;
  assign n47991 = n536 & n47990 ;
  assign n47992 = n2441 & n6537 ;
  assign n47993 = ( n13287 & ~n18236 ) | ( n13287 & n47992 ) | ( ~n18236 & n47992 ) ;
  assign n47994 = n19906 ^ n17100 ^ 1'b0 ;
  assign n47995 = ~n47993 & n47994 ;
  assign n47996 = n17473 ^ n5155 ^ 1'b0 ;
  assign n47997 = n36337 | n43803 ;
  assign n47998 = n32319 ^ n18113 ^ n1684 ;
  assign n47999 = n20664 ^ n5072 ^ 1'b0 ;
  assign n48000 = n10931 ^ n463 ^ 1'b0 ;
  assign n48001 = ~n41931 & n48000 ;
  assign n48002 = n20601 & n30063 ;
  assign n48003 = n48002 ^ n41697 ^ 1'b0 ;
  assign n48004 = n33445 ^ n16297 ^ 1'b0 ;
  assign n48005 = ( n4039 & n20676 ) | ( n4039 & n33300 ) | ( n20676 & n33300 ) ;
  assign n48006 = n411 & n2484 ;
  assign n48007 = n33843 ^ n31544 ^ 1'b0 ;
  assign n48008 = n6029 | n17245 ;
  assign n48009 = n48008 ^ n28468 ^ 1'b0 ;
  assign n48010 = n48009 ^ n10079 ^ 1'b0 ;
  assign n48011 = n19237 | n48010 ;
  assign n48012 = ~n23656 & n27638 ;
  assign n48013 = n48012 ^ n28674 ^ 1'b0 ;
  assign n48014 = n48013 ^ n31772 ^ n21935 ;
  assign n48015 = n48014 ^ n6098 ^ 1'b0 ;
  assign n48016 = n1875 | n9321 ;
  assign n48017 = n36916 ^ n17848 ^ 1'b0 ;
  assign n48018 = n19463 ^ n13141 ^ n1943 ;
  assign n48019 = n48018 ^ n15173 ^ n2140 ;
  assign n48020 = n21382 ^ n15665 ^ 1'b0 ;
  assign n48021 = ~n28002 & n48020 ;
  assign n48022 = ( n31753 & ~n41655 ) | ( n31753 & n48021 ) | ( ~n41655 & n48021 ) ;
  assign n48023 = ( n7406 & n19745 ) | ( n7406 & ~n30586 ) | ( n19745 & ~n30586 ) ;
  assign n48024 = n29379 ^ n9734 ^ 1'b0 ;
  assign n48025 = n2678 & ~n29774 ;
  assign n48026 = n48024 & n48025 ;
  assign n48027 = n9706 & n39020 ;
  assign n48028 = n25455 & n48027 ;
  assign n48029 = n41178 & n44933 ;
  assign n48030 = n15687 ^ n7754 ^ 1'b0 ;
  assign n48031 = ( ~n14878 & n23986 ) | ( ~n14878 & n24278 ) | ( n23986 & n24278 ) ;
  assign n48032 = ( n154 & n1616 ) | ( n154 & n4461 ) | ( n1616 & n4461 ) ;
  assign n48033 = ~n48031 & n48032 ;
  assign n48034 = ~n3717 & n25239 ;
  assign n48035 = ~n15735 & n42801 ;
  assign n48036 = n31338 & n48035 ;
  assign n48038 = ~n8287 & n16263 ;
  assign n48037 = ~n4608 & n13760 ;
  assign n48039 = n48038 ^ n48037 ^ 1'b0 ;
  assign n48040 = ~n18176 & n32808 ;
  assign n48041 = n19946 ^ n13110 ^ 1'b0 ;
  assign n48042 = n22694 & n48041 ;
  assign n48043 = n29541 & n48042 ;
  assign n48044 = n48040 & ~n48043 ;
  assign n48045 = ~n1426 & n4715 ;
  assign n48046 = n47821 & n48045 ;
  assign n48047 = n7991 & ~n36113 ;
  assign n48048 = ~n17919 & n21787 ;
  assign n48049 = n5210 & n30940 ;
  assign n48050 = n48049 ^ n24703 ^ 1'b0 ;
  assign n48051 = ( n3608 & n3823 ) | ( n3608 & ~n16883 ) | ( n3823 & ~n16883 ) ;
  assign n48052 = n7864 & n48051 ;
  assign n48053 = n10502 & n48052 ;
  assign n48054 = n48050 & ~n48053 ;
  assign n48057 = ~n2367 & n3376 ;
  assign n48058 = ~n13926 & n48057 ;
  assign n48059 = n48058 ^ n36273 ^ 1'b0 ;
  assign n48055 = n43987 ^ n22968 ^ 1'b0 ;
  assign n48056 = n12089 & n48055 ;
  assign n48060 = n48059 ^ n48056 ^ n31955 ;
  assign n48063 = n20021 | n24623 ;
  assign n48061 = n9618 | n31457 ;
  assign n48062 = n23114 & ~n48061 ;
  assign n48064 = n48063 ^ n48062 ^ 1'b0 ;
  assign n48065 = n28743 ^ n10392 ^ 1'b0 ;
  assign n48066 = n19240 | n48065 ;
  assign n48067 = n48066 ^ n19767 ^ 1'b0 ;
  assign n48068 = ~n11717 & n48067 ;
  assign n48070 = n19858 ^ n7847 ^ 1'b0 ;
  assign n48069 = n5836 | n42135 ;
  assign n48071 = n48070 ^ n48069 ^ 1'b0 ;
  assign n48072 = n5301 & ~n27233 ;
  assign n48073 = ( n473 & n5563 ) | ( n473 & n44491 ) | ( n5563 & n44491 ) ;
  assign n48074 = ( n550 & ~n6418 ) | ( n550 & n40130 ) | ( ~n6418 & n40130 ) ;
  assign n48075 = n2317 | n47503 ;
  assign n48076 = n9005 & ~n48075 ;
  assign n48077 = n2935 & ~n17233 ;
  assign n48078 = n48077 ^ n27971 ^ 1'b0 ;
  assign n48081 = n19683 ^ n14178 ^ 1'b0 ;
  assign n48082 = n35258 | n48081 ;
  assign n48079 = n26956 ^ n7535 ^ 1'b0 ;
  assign n48080 = n11395 | n48079 ;
  assign n48083 = n48082 ^ n48080 ^ 1'b0 ;
  assign n48084 = n17260 ^ n2519 ^ 1'b0 ;
  assign n48085 = n6788 & n48084 ;
  assign n48086 = n17920 ^ n13632 ^ 1'b0 ;
  assign n48087 = n44333 | n48086 ;
  assign n48088 = ( ~n9635 & n15907 ) | ( ~n9635 & n48087 ) | ( n15907 & n48087 ) ;
  assign n48089 = n1337 | n18855 ;
  assign n48090 = n4608 | n48089 ;
  assign n48091 = ( ~n11069 & n41657 ) | ( ~n11069 & n48090 ) | ( n41657 & n48090 ) ;
  assign n48092 = ( n42803 & ~n48088 ) | ( n42803 & n48091 ) | ( ~n48088 & n48091 ) ;
  assign n48093 = n32452 ^ n27791 ^ 1'b0 ;
  assign n48094 = n4553 & ~n16379 ;
  assign n48095 = n16585 ^ n722 ^ 1'b0 ;
  assign n48096 = ~n48094 & n48095 ;
  assign n48097 = n38912 ^ n29371 ^ 1'b0 ;
  assign n48098 = n45780 ^ n29780 ^ 1'b0 ;
  assign n48099 = n26982 & n48098 ;
  assign n48100 = n9296 & n18940 ;
  assign n48101 = n1712 & n2895 ;
  assign n48102 = ( n19562 & n48100 ) | ( n19562 & n48101 ) | ( n48100 & n48101 ) ;
  assign n48104 = ~n6737 & n21707 ;
  assign n48103 = ~n7468 & n38033 ;
  assign n48105 = n48104 ^ n48103 ^ 1'b0 ;
  assign n48106 = n46567 ^ n39160 ^ 1'b0 ;
  assign n48107 = n18420 & ~n26283 ;
  assign n48108 = n48107 ^ n32407 ^ 1'b0 ;
  assign n48109 = n14530 ^ n7025 ^ 1'b0 ;
  assign n48110 = n9621 & n48109 ;
  assign n48111 = n574 & ~n10512 ;
  assign n48112 = n48110 & n48111 ;
  assign n48113 = n26245 & n48112 ;
  assign n48114 = ~n12742 & n22358 ;
  assign n48115 = n3773 & n4181 ;
  assign n48116 = n48115 ^ n1894 ^ 1'b0 ;
  assign n48117 = ( n32106 & n46319 ) | ( n32106 & n48116 ) | ( n46319 & n48116 ) ;
  assign n48118 = n29458 & n31383 ;
  assign n48119 = n48118 ^ n26994 ^ 1'b0 ;
  assign n48120 = n37775 ^ n22698 ^ n3730 ;
  assign n48121 = n48120 ^ n12202 ^ 1'b0 ;
  assign n48122 = n46486 & ~n48121 ;
  assign n48123 = n772 & n48122 ;
  assign n48124 = n48123 ^ n30486 ^ 1'b0 ;
  assign n48125 = ~n29133 & n48124 ;
  assign n48126 = n7377 ^ n3548 ^ 1'b0 ;
  assign n48127 = n1933 & n5151 ;
  assign n48128 = n22967 & ~n23040 ;
  assign n48129 = n48128 ^ n44882 ^ n20494 ;
  assign n48130 = n21784 ^ n14526 ^ 1'b0 ;
  assign n48131 = n48130 ^ n40739 ^ n11603 ;
  assign n48132 = n2880 & n4422 ;
  assign n48133 = n48132 ^ n6447 ^ 1'b0 ;
  assign n48134 = n7516 & n48133 ;
  assign n48135 = n21664 ^ n4768 ^ 1'b0 ;
  assign n48136 = n4683 & ~n48135 ;
  assign n48137 = ~n3940 & n48136 ;
  assign n48138 = n48137 ^ n45792 ^ 1'b0 ;
  assign n48139 = n22502 | n48138 ;
  assign n48140 = n48139 ^ n14882 ^ 1'b0 ;
  assign n48141 = n20086 | n36906 ;
  assign n48142 = n48141 ^ n19453 ^ 1'b0 ;
  assign n48143 = n37621 & ~n48142 ;
  assign n48144 = n29604 ^ n7831 ^ n4104 ;
  assign n48145 = n27076 | n48144 ;
  assign n48146 = n48145 ^ n17578 ^ 1'b0 ;
  assign n48147 = n48143 & ~n48146 ;
  assign n48148 = n9832 | n16291 ;
  assign n48149 = n48148 ^ n29344 ^ n4930 ;
  assign n48150 = n39993 & ~n41882 ;
  assign n48151 = n5115 & n48150 ;
  assign n48152 = n48151 ^ n21232 ^ 1'b0 ;
  assign n48153 = ~n31753 & n48152 ;
  assign n48154 = n15645 & n45786 ;
  assign n48155 = n48153 & n48154 ;
  assign n48156 = n3225 | n5883 ;
  assign n48157 = ( n1311 & n4622 ) | ( n1311 & ~n48156 ) | ( n4622 & ~n48156 ) ;
  assign n48158 = ~n8311 & n42710 ;
  assign n48159 = n1238 | n37921 ;
  assign n48160 = n44103 | n48159 ;
  assign n48161 = ~n7345 & n11769 ;
  assign n48162 = ~n5573 & n31813 ;
  assign n48163 = n48162 ^ n7235 ^ 1'b0 ;
  assign n48164 = n47656 ^ n3693 ^ 1'b0 ;
  assign n48165 = ~n9866 & n48164 ;
  assign n48166 = n36108 ^ n2459 ^ 1'b0 ;
  assign n48167 = n8443 & ~n9283 ;
  assign n48168 = n18845 & n48167 ;
  assign n48169 = ~n15537 & n48168 ;
  assign n48170 = n16464 & ~n16873 ;
  assign n48171 = n48170 ^ n4785 ^ 1'b0 ;
  assign n48172 = ( ~n8371 & n48169 ) | ( ~n8371 & n48171 ) | ( n48169 & n48171 ) ;
  assign n48173 = n26977 ^ n17487 ^ n16467 ;
  assign n48174 = n6683 | n15498 ;
  assign n48175 = ~n23669 & n31488 ;
  assign n48176 = n44406 ^ n32150 ^ 1'b0 ;
  assign n48177 = n45635 ^ n25016 ^ 1'b0 ;
  assign n48178 = ~n12272 & n25762 ;
  assign n48179 = ~n29073 & n48178 ;
  assign n48180 = n42985 ^ n22466 ^ n20647 ;
  assign n48181 = n23676 ^ n16559 ^ 1'b0 ;
  assign n48182 = n45163 ^ n22907 ^ n3464 ;
  assign n48183 = n48182 ^ n26416 ^ n9699 ;
  assign n48184 = n48183 ^ n40596 ^ 1'b0 ;
  assign n48185 = n4175 | n5608 ;
  assign n48186 = n22729 & ~n48185 ;
  assign n48187 = n1389 ^ n1340 ^ 1'b0 ;
  assign n48188 = n48186 | n48187 ;
  assign n48189 = n26128 | n48188 ;
  assign n48190 = n9890 & ~n48189 ;
  assign n48191 = n42017 & ~n48190 ;
  assign n48192 = ~n13594 & n48191 ;
  assign n48193 = n22941 & ~n25681 ;
  assign n48194 = n47488 ^ n32452 ^ 1'b0 ;
  assign n48195 = n48193 & ~n48194 ;
  assign n48196 = n38532 ^ n22687 ^ 1'b0 ;
  assign n48197 = n25142 & ~n48196 ;
  assign n48198 = n4372 & ~n8593 ;
  assign n48199 = n8646 | n11531 ;
  assign n48200 = n48199 ^ n47198 ^ n4978 ;
  assign n48201 = n47639 ^ n17656 ^ n5529 ;
  assign n48202 = n1509 | n20636 ;
  assign n48203 = n20636 & ~n48202 ;
  assign n48204 = n48203 ^ n18522 ^ n8713 ;
  assign n48205 = n48204 ^ n33773 ^ 1'b0 ;
  assign n48206 = n12976 | n15373 ;
  assign n48207 = n2309 ^ n1168 ^ 1'b0 ;
  assign n48208 = n38477 & n48207 ;
  assign n48209 = n12324 ^ n3261 ^ 1'b0 ;
  assign n48210 = n48209 ^ n16507 ^ 1'b0 ;
  assign n48211 = n8829 & n48210 ;
  assign n48212 = n19562 & ~n20767 ;
  assign n48213 = n26036 ^ n2114 ^ 1'b0 ;
  assign n48214 = n48213 ^ n40728 ^ 1'b0 ;
  assign n48216 = ( n2528 & n12807 ) | ( n2528 & ~n29244 ) | ( n12807 & ~n29244 ) ;
  assign n48215 = n5166 & n15238 ;
  assign n48217 = n48216 ^ n48215 ^ 1'b0 ;
  assign n48218 = ( n6251 & ~n10385 ) | ( n6251 & n48058 ) | ( ~n10385 & n48058 ) ;
  assign n48219 = ( n2104 & n42482 ) | ( n2104 & ~n48218 ) | ( n42482 & ~n48218 ) ;
  assign n48220 = n29539 & n45449 ;
  assign n48225 = n7864 | n38679 ;
  assign n48226 = n48225 ^ n39394 ^ 1'b0 ;
  assign n48221 = n4410 ^ n2831 ^ 1'b0 ;
  assign n48222 = n18368 & ~n48221 ;
  assign n48223 = n28748 ^ n25556 ^ 1'b0 ;
  assign n48224 = ~n48222 & n48223 ;
  assign n48227 = n48226 ^ n48224 ^ n38916 ;
  assign n48228 = n20679 & n48227 ;
  assign n48229 = ~n5570 & n22716 ;
  assign n48230 = n43572 ^ n9265 ^ n2313 ;
  assign n48231 = ( ~n28864 & n47402 ) | ( ~n28864 & n48230 ) | ( n47402 & n48230 ) ;
  assign n48232 = n48231 ^ n863 ^ 1'b0 ;
  assign n48233 = n9101 & n48043 ;
  assign n48234 = n27865 & ~n39969 ;
  assign n48235 = n14977 | n15408 ;
  assign n48236 = ( n39314 & n44427 ) | ( n39314 & n48235 ) | ( n44427 & n48235 ) ;
  assign n48237 = ~n24109 & n24890 ;
  assign n48238 = n9072 | n26611 ;
  assign n48239 = n8491 & n48238 ;
  assign n48240 = n48239 ^ n30460 ^ 1'b0 ;
  assign n48241 = n48240 ^ n36219 ^ 1'b0 ;
  assign n48242 = n43464 | n48241 ;
  assign n48243 = n48242 ^ n16639 ^ 1'b0 ;
  assign n48244 = n7580 & n12885 ;
  assign n48245 = n2579 ^ n2177 ^ 1'b0 ;
  assign n48246 = n7069 & n48245 ;
  assign n48247 = ( n6166 & n37776 ) | ( n6166 & n48246 ) | ( n37776 & n48246 ) ;
  assign n48248 = n36393 ^ n17996 ^ 1'b0 ;
  assign n48249 = n31871 | n48248 ;
  assign n48250 = n431 | n597 ;
  assign n48251 = ~n18243 & n47733 ;
  assign n48252 = n7357 ^ n3464 ^ 1'b0 ;
  assign n48253 = ~n14900 & n48252 ;
  assign n48254 = n11585 ^ n3046 ^ 1'b0 ;
  assign n48255 = ( ~n15610 & n26563 ) | ( ~n15610 & n30924 ) | ( n26563 & n30924 ) ;
  assign n48256 = ~n3747 & n6700 ;
  assign n48257 = ( n14112 & n16719 ) | ( n14112 & n48256 ) | ( n16719 & n48256 ) ;
  assign n48258 = n5069 | n25111 ;
  assign n48259 = n25167 & ~n48258 ;
  assign n48260 = n18989 & n44093 ;
  assign n48261 = ~n21267 & n48260 ;
  assign n48262 = n48261 ^ n34490 ^ 1'b0 ;
  assign n48263 = n18045 ^ n922 ^ 1'b0 ;
  assign n48264 = n48263 ^ n24191 ^ n7111 ;
  assign n48265 = n48264 ^ n26214 ^ 1'b0 ;
  assign n48266 = n1118 & n48265 ;
  assign n48267 = n31070 ^ n4367 ^ 1'b0 ;
  assign n48268 = n48266 & ~n48267 ;
  assign n48269 = n1025 & n2070 ;
  assign n48270 = ~n4387 & n48269 ;
  assign n48271 = n19237 & ~n21628 ;
  assign n48272 = n4141 | n10524 ;
  assign n48273 = n48272 ^ n42664 ^ 1'b0 ;
  assign n48274 = n2746 & ~n5212 ;
  assign n48275 = ( n1378 & n48120 ) | ( n1378 & ~n48274 ) | ( n48120 & ~n48274 ) ;
  assign n48276 = n5702 & ~n11365 ;
  assign n48277 = n12658 | n13160 ;
  assign n48278 = n48277 ^ n29304 ^ 1'b0 ;
  assign n48279 = ~n48276 & n48278 ;
  assign n48280 = n2980 & n5781 ;
  assign n48281 = n2436 | n37410 ;
  assign n48282 = n48281 ^ n1288 ^ 1'b0 ;
  assign n48283 = n26138 | n27217 ;
  assign n48284 = n48283 ^ n21119 ^ 1'b0 ;
  assign n48285 = n48284 ^ n22096 ^ n6990 ;
  assign n48287 = n20312 ^ n8612 ^ 1'b0 ;
  assign n48286 = n2486 | n16780 ;
  assign n48288 = n48287 ^ n48286 ^ 1'b0 ;
  assign n48289 = ( n5878 & ~n9143 ) | ( n5878 & n48288 ) | ( ~n9143 & n48288 ) ;
  assign n48290 = ~n13730 & n47085 ;
  assign n48291 = n8912 ^ n6008 ^ n5284 ;
  assign n48292 = n4315 & n48291 ;
  assign n48293 = n48292 ^ n38960 ^ 1'b0 ;
  assign n48294 = n48293 ^ n12404 ^ n6966 ;
  assign n48295 = n16835 | n33756 ;
  assign n48296 = n48294 & ~n48295 ;
  assign n48297 = n6062 | n23106 ;
  assign n48298 = n48297 ^ n28438 ^ 1'b0 ;
  assign n48299 = ~n8547 & n21430 ;
  assign n48300 = n3542 & n48299 ;
  assign n48301 = n31268 & ~n42010 ;
  assign n48302 = n11503 ^ n8145 ^ n5740 ;
  assign n48303 = n39764 ^ n27472 ^ n659 ;
  assign n48304 = n15574 & n43024 ;
  assign n48305 = n10133 & n17556 ;
  assign n48306 = ~n16901 & n48305 ;
  assign n48307 = n490 & ~n5214 ;
  assign n48308 = n46508 | n48307 ;
  assign n48309 = n9944 | n27989 ;
  assign n48310 = n46916 ^ n11785 ^ 1'b0 ;
  assign n48313 = ~n2393 & n9996 ;
  assign n48314 = n48313 ^ n9424 ^ 1'b0 ;
  assign n48311 = n22057 ^ n19899 ^ n16573 ;
  assign n48312 = ~n5122 & n48311 ;
  assign n48315 = n48314 ^ n48312 ^ 1'b0 ;
  assign n48317 = n32979 ^ n12806 ^ n10453 ;
  assign n48316 = ~n36988 & n39127 ;
  assign n48318 = n48317 ^ n48316 ^ 1'b0 ;
  assign n48319 = ( n887 & ~n16224 ) | ( n887 & n43759 ) | ( ~n16224 & n43759 ) ;
  assign n48320 = n10245 & ~n19285 ;
  assign n48321 = ( n21548 & n26744 ) | ( n21548 & n48320 ) | ( n26744 & n48320 ) ;
  assign n48322 = n28308 ^ n17954 ^ n3544 ;
  assign n48323 = n21744 ^ n37 ^ 1'b0 ;
  assign n48324 = ~n18818 & n48323 ;
  assign n48325 = n45636 | n48324 ;
  assign n48326 = n4817 ^ n2071 ^ 1'b0 ;
  assign n48327 = ( n20751 & ~n27731 ) | ( n20751 & n48326 ) | ( ~n27731 & n48326 ) ;
  assign n48328 = n12053 | n48327 ;
  assign n48329 = n20838 & n35267 ;
  assign n48330 = n23344 | n48329 ;
  assign n48331 = n48328 | n48330 ;
  assign n48332 = n28767 | n40756 ;
  assign n48333 = n1768 & ~n48332 ;
  assign n48334 = n10296 & ~n30934 ;
  assign n48335 = ( n3702 & n18806 ) | ( n3702 & ~n39900 ) | ( n18806 & ~n39900 ) ;
  assign n48336 = ( ~n10314 & n31330 ) | ( ~n10314 & n48335 ) | ( n31330 & n48335 ) ;
  assign n48337 = n2904 ^ n753 ^ 1'b0 ;
  assign n48338 = n48337 ^ n7631 ^ 1'b0 ;
  assign n48339 = ~n8950 & n34946 ;
  assign n48340 = n1606 & ~n20752 ;
  assign n48341 = n48340 ^ n3624 ^ 1'b0 ;
  assign n48342 = n20161 ^ n18940 ^ 1'b0 ;
  assign n48343 = ~n22202 & n48342 ;
  assign n48344 = n29831 | n33289 ;
  assign n48345 = n36459 | n48344 ;
  assign n48346 = n24834 ^ n13261 ^ n1118 ;
  assign n48347 = n13942 & ~n48346 ;
  assign n48348 = n24110 & n48347 ;
  assign n48349 = ( ~n39124 & n41164 ) | ( ~n39124 & n48348 ) | ( n41164 & n48348 ) ;
  assign n48350 = ~n24802 & n33482 ;
  assign n48354 = n12495 & ~n13071 ;
  assign n48355 = n48354 ^ n22101 ^ 1'b0 ;
  assign n48351 = n16500 ^ n8482 ^ 1'b0 ;
  assign n48352 = n14641 | n48351 ;
  assign n48353 = n8703 & ~n48352 ;
  assign n48356 = n48355 ^ n48353 ^ 1'b0 ;
  assign n48357 = n8369 & n9263 ;
  assign n48358 = ~n1507 & n48357 ;
  assign n48359 = n11772 ^ n496 ^ 1'b0 ;
  assign n48360 = n13764 | n48359 ;
  assign n48361 = n48360 ^ n15503 ^ 1'b0 ;
  assign n48362 = ~n16398 & n21213 ;
  assign n48363 = n3630 | n43411 ;
  assign n48364 = n48362 | n48363 ;
  assign n48365 = n43650 ^ n20830 ^ 1'b0 ;
  assign n48366 = n48364 & ~n48365 ;
  assign n48367 = ~n45682 & n47685 ;
  assign n48368 = ( n1752 & n17951 ) | ( n1752 & ~n48367 ) | ( n17951 & ~n48367 ) ;
  assign n48369 = n8195 ^ n3567 ^ 1'b0 ;
  assign n48372 = n25242 & n36126 ;
  assign n48370 = n6197 | n11275 ;
  assign n48371 = ~n43976 & n48370 ;
  assign n48373 = n48372 ^ n48371 ^ 1'b0 ;
  assign n48374 = n32255 & ~n37146 ;
  assign n48376 = n19387 | n20129 ;
  assign n48377 = n48376 ^ n15667 ^ 1'b0 ;
  assign n48378 = n48377 ^ n12666 ^ n5724 ;
  assign n48379 = n44242 & ~n48378 ;
  assign n48375 = n2250 | n8312 ;
  assign n48380 = n48379 ^ n48375 ^ 1'b0 ;
  assign n48381 = n26007 ^ n5123 ^ 1'b0 ;
  assign n48382 = ~n16591 & n30228 ;
  assign n48383 = n7542 & ~n15890 ;
  assign n48384 = n19729 & n48383 ;
  assign n48385 = n13438 | n48384 ;
  assign n48386 = n12119 ^ n7502 ^ n7062 ;
  assign n48387 = n21567 | n25522 ;
  assign n48388 = n6199 & n18664 ;
  assign n48389 = ( ~n32583 & n48387 ) | ( ~n32583 & n48388 ) | ( n48387 & n48388 ) ;
  assign n48390 = ~n15044 & n45849 ;
  assign n48391 = n48390 ^ n5880 ^ 1'b0 ;
  assign n48393 = n5083 & ~n23114 ;
  assign n48392 = n2895 & ~n5657 ;
  assign n48394 = n48393 ^ n48392 ^ 1'b0 ;
  assign n48395 = n13215 | n44609 ;
  assign n48396 = n48395 ^ n17354 ^ 1'b0 ;
  assign n48397 = n48396 ^ n15709 ^ 1'b0 ;
  assign n48398 = n4819 & n48397 ;
  assign n48399 = n45128 & n48398 ;
  assign n48400 = n4686 & ~n6562 ;
  assign n48401 = n15488 ^ n13101 ^ n7622 ;
  assign n48402 = n14067 ^ n13378 ^ 1'b0 ;
  assign n48403 = ( n19055 & n28406 ) | ( n19055 & ~n48402 ) | ( n28406 & ~n48402 ) ;
  assign n48404 = n2201 & n18759 ;
  assign n48405 = n1351 & n48404 ;
  assign n48406 = n48405 ^ n22426 ^ 1'b0 ;
  assign n48407 = n12758 ^ n7471 ^ 1'b0 ;
  assign n48408 = n34856 & ~n48407 ;
  assign n48409 = ~n12357 & n15754 ;
  assign n48410 = n42503 & n48409 ;
  assign n48411 = ~n12143 & n48410 ;
  assign n48412 = ~n20713 & n33783 ;
  assign n48413 = n44017 | n47025 ;
  assign n48414 = n24739 ^ n16922 ^ 1'b0 ;
  assign n48415 = n43069 ^ n38498 ^ n34307 ;
  assign n48416 = n29634 ^ n29586 ^ 1'b0 ;
  assign n48417 = ~n771 & n48416 ;
  assign n48418 = n8173 & ~n43324 ;
  assign n48419 = ~n1488 & n48418 ;
  assign n48420 = n48419 ^ n6985 ^ 1'b0 ;
  assign n48421 = n267 & n48420 ;
  assign n48422 = n37860 ^ n23571 ^ 1'b0 ;
  assign n48423 = ( n10686 & ~n19169 ) | ( n10686 & n20392 ) | ( ~n19169 & n20392 ) ;
  assign n48424 = ( n39798 & n44279 ) | ( n39798 & ~n48423 ) | ( n44279 & ~n48423 ) ;
  assign n48425 = n41190 ^ n12095 ^ n3750 ;
  assign n48426 = ( n11288 & n43592 ) | ( n11288 & n48425 ) | ( n43592 & n48425 ) ;
  assign n48427 = n7399 ^ n3455 ^ 1'b0 ;
  assign n48428 = n9973 | n11529 ;
  assign n48429 = n31026 | n48428 ;
  assign n48430 = n2982 | n26596 ;
  assign n48431 = n48430 ^ n28063 ^ 1'b0 ;
  assign n48432 = n12850 ^ n1314 ^ 1'b0 ;
  assign n48433 = ( n2915 & n11177 ) | ( n2915 & ~n21848 ) | ( n11177 & ~n21848 ) ;
  assign n48434 = n48433 ^ n7443 ^ 1'b0 ;
  assign n48435 = n48432 | n48434 ;
  assign n48436 = n22494 & ~n48435 ;
  assign n48437 = n11009 | n25775 ;
  assign n48438 = n18044 ^ n9610 ^ 1'b0 ;
  assign n48439 = n18478 & ~n48438 ;
  assign n48440 = ~n356 & n2094 ;
  assign n48441 = n48440 ^ n13226 ^ 1'b0 ;
  assign n48442 = n7071 | n48441 ;
  assign n48443 = n4202 | n48442 ;
  assign n48444 = n31295 | n33128 ;
  assign n48445 = n22858 | n43803 ;
  assign n48446 = n48445 ^ n10850 ^ 1'b0 ;
  assign n48447 = n9060 & ~n29603 ;
  assign n48448 = ~n27314 & n48447 ;
  assign n48449 = n48448 ^ n2738 ^ 1'b0 ;
  assign n48450 = n9904 & n19871 ;
  assign n48451 = n35445 ^ n27000 ^ 1'b0 ;
  assign n48452 = n43881 ^ n15821 ^ n11433 ;
  assign n48453 = n9618 ^ n5994 ^ 1'b0 ;
  assign n48454 = ( n2556 & ~n6654 ) | ( n2556 & n21578 ) | ( ~n6654 & n21578 ) ;
  assign n48455 = n7210 ^ n7089 ^ 1'b0 ;
  assign n48456 = ( n14124 & n15734 ) | ( n14124 & ~n48455 ) | ( n15734 & ~n48455 ) ;
  assign n48457 = ( n11389 & ~n46803 ) | ( n11389 & n47484 ) | ( ~n46803 & n47484 ) ;
  assign n48458 = n38935 ^ n10551 ^ 1'b0 ;
  assign n48459 = ~n2445 & n48458 ;
  assign n48460 = n11269 & n48459 ;
  assign n48461 = n44336 ^ n40181 ^ 1'b0 ;
  assign n48462 = n15826 | n48461 ;
  assign n48463 = n8662 & ~n12761 ;
  assign n48464 = n48463 ^ n12159 ^ 1'b0 ;
  assign n48465 = ( n2752 & n23636 ) | ( n2752 & n48464 ) | ( n23636 & n48464 ) ;
  assign n48466 = n48465 ^ n23841 ^ n13650 ;
  assign n48467 = n24302 ^ n17257 ^ n2484 ;
  assign n48468 = n48467 ^ n44534 ^ 1'b0 ;
  assign n48469 = n18225 | n48468 ;
  assign n48470 = n6390 | n8848 ;
  assign n48471 = n48470 ^ n32339 ^ 1'b0 ;
  assign n48472 = ~n8017 & n48471 ;
  assign n48473 = ~n39528 & n48472 ;
  assign n48474 = n10504 ^ n216 ^ 1'b0 ;
  assign n48475 = n45564 ^ n15111 ^ 1'b0 ;
  assign n48476 = n13769 & ~n48475 ;
  assign n48477 = n21510 & n48476 ;
  assign n48478 = n33909 ^ n18368 ^ 1'b0 ;
  assign n48479 = n13228 & ~n48478 ;
  assign n48480 = n48479 ^ n36625 ^ 1'b0 ;
  assign n48481 = n25089 ^ n13710 ^ n3825 ;
  assign n48482 = n48481 ^ n1231 ^ 1'b0 ;
  assign n48483 = n12994 & ~n48482 ;
  assign n48484 = n37559 ^ n15159 ^ 1'b0 ;
  assign n48485 = n21752 ^ n14920 ^ 1'b0 ;
  assign n48486 = n48485 ^ n21849 ^ n16536 ;
  assign n48487 = ( n28582 & n46868 ) | ( n28582 & n47804 ) | ( n46868 & n47804 ) ;
  assign n48488 = n21381 ^ n11035 ^ 1'b0 ;
  assign n48489 = ~n9290 & n48488 ;
  assign n48490 = n26885 | n48465 ;
  assign n48491 = n1292 | n35770 ;
  assign n48492 = n8683 | n48491 ;
  assign n48493 = n23033 ^ n19952 ^ 1'b0 ;
  assign n48494 = ~n36377 & n48493 ;
  assign n48495 = n36982 ^ n29091 ^ n13928 ;
  assign n48496 = n48495 ^ n27555 ^ 1'b0 ;
  assign n48497 = n27541 & n45506 ;
  assign n48498 = n48497 ^ n23168 ^ 1'b0 ;
  assign n48499 = n895 | n9189 ;
  assign n48500 = n48499 ^ n13589 ^ 1'b0 ;
  assign n48501 = n7385 ^ n1647 ^ 1'b0 ;
  assign n48502 = n8697 & n48501 ;
  assign n48503 = n39937 ^ n25145 ^ n6991 ;
  assign n48504 = ( n5387 & n6316 ) | ( n5387 & n48503 ) | ( n6316 & n48503 ) ;
  assign n48505 = ( n15461 & n17114 ) | ( n15461 & n39391 ) | ( n17114 & n39391 ) ;
  assign n48506 = n45243 ^ n29905 ^ n352 ;
  assign n48507 = ~n13768 & n24776 ;
  assign n48508 = n28323 & n48507 ;
  assign n48509 = ~n2982 & n18916 ;
  assign n48510 = n48509 ^ n1796 ^ 1'b0 ;
  assign n48511 = n73 | n11946 ;
  assign n48512 = n12903 | n16231 ;
  assign n48513 = n48512 ^ n22340 ^ n10313 ;
  assign n48514 = n1412 & ~n38357 ;
  assign n48515 = n9798 & n19815 ;
  assign n48516 = n8027 | n30934 ;
  assign n48517 = n48515 | n48516 ;
  assign n48518 = n48517 ^ n35049 ^ 1'b0 ;
  assign n48519 = ~n11581 & n48518 ;
  assign n48520 = n48519 ^ n25976 ^ 1'b0 ;
  assign n48521 = n14321 ^ n7876 ^ 1'b0 ;
  assign n48522 = ~n5147 & n48521 ;
  assign n48523 = ~n5898 & n5906 ;
  assign n48524 = n48523 ^ n27319 ^ 1'b0 ;
  assign n48525 = n48522 & ~n48524 ;
  assign n48526 = n30058 ^ n706 ^ 1'b0 ;
  assign n48527 = n1956 & n46100 ;
  assign n48528 = n45925 ^ n33791 ^ n12054 ;
  assign n48529 = n13956 ^ n2190 ^ 1'b0 ;
  assign n48530 = n19845 & ~n48529 ;
  assign n48531 = n1851 ^ n879 ^ 1'b0 ;
  assign n48532 = ( ~n5204 & n7136 ) | ( ~n5204 & n10219 ) | ( n7136 & n10219 ) ;
  assign n48533 = n17821 ^ n543 ^ 1'b0 ;
  assign n48534 = n48532 | n48533 ;
  assign n48535 = n48534 ^ n13298 ^ 1'b0 ;
  assign n48536 = n17939 | n38127 ;
  assign n48537 = n5250 | n39996 ;
  assign n48538 = n166 & ~n23971 ;
  assign n48539 = n16393 & ~n42150 ;
  assign n48540 = n48539 ^ n30398 ^ 1'b0 ;
  assign n48541 = n20085 | n48540 ;
  assign n48542 = n10780 & ~n21770 ;
  assign n48543 = n10885 & n48542 ;
  assign n48544 = n48543 ^ n9484 ^ 1'b0 ;
  assign n48545 = ~n20438 & n48544 ;
  assign n48546 = ~n40259 & n43080 ;
  assign n48547 = n33490 ^ n17243 ^ 1'b0 ;
  assign n48548 = n28206 ^ n5738 ^ 1'b0 ;
  assign n48549 = n48547 | n48548 ;
  assign n48550 = ~n1772 & n29746 ;
  assign n48551 = n48550 ^ n2001 ^ 1'b0 ;
  assign n48552 = n46167 & ~n48551 ;
  assign n48553 = n48552 ^ n510 ^ 1'b0 ;
  assign n48554 = n12002 | n19850 ;
  assign n48555 = n48554 ^ n9050 ^ 1'b0 ;
  assign n48556 = n5873 ^ n4685 ^ 1'b0 ;
  assign n48557 = ~n3872 & n7287 ;
  assign n48558 = ( n18059 & ~n48485 ) | ( n18059 & n48557 ) | ( ~n48485 & n48557 ) ;
  assign n48559 = n6851 & ~n21997 ;
  assign n48560 = n27727 ^ n1444 ^ 1'b0 ;
  assign n48561 = n19038 | n48560 ;
  assign n48562 = n3593 ^ n54 ^ 1'b0 ;
  assign n48563 = n15087 | n48562 ;
  assign n48564 = n492 | n10830 ;
  assign n48565 = n48564 ^ n43344 ^ 1'b0 ;
  assign n48566 = n48565 ^ n2471 ^ n1167 ;
  assign n48567 = n26055 | n48566 ;
  assign n48568 = n2905 | n9765 ;
  assign n48569 = n2795 & ~n48568 ;
  assign n48570 = n48569 ^ n12271 ^ 1'b0 ;
  assign n48571 = n17788 | n48570 ;
  assign n48573 = n14758 & n23497 ;
  assign n48572 = n5212 & n7527 ;
  assign n48574 = n48573 ^ n48572 ^ 1'b0 ;
  assign n48575 = n48556 ^ n11219 ^ 1'b0 ;
  assign n48576 = n7913 & ~n15371 ;
  assign n48577 = ( n3568 & n47655 ) | ( n3568 & ~n48576 ) | ( n47655 & ~n48576 ) ;
  assign n48578 = n20560 | n48577 ;
  assign n48579 = n40904 ^ n25110 ^ 1'b0 ;
  assign n48580 = ~n4277 & n48579 ;
  assign n48581 = ( n13621 & n21429 ) | ( n13621 & n48580 ) | ( n21429 & n48580 ) ;
  assign n48582 = n13046 ^ n11592 ^ n1080 ;
  assign n48583 = n28602 | n46463 ;
  assign n48584 = n48583 ^ n6134 ^ 1'b0 ;
  assign n48585 = n7205 & n48584 ;
  assign n48586 = n7094 | n37302 ;
  assign n48587 = n37081 & ~n48586 ;
  assign n48588 = n21469 & n48587 ;
  assign n48589 = ~n221 & n4825 ;
  assign n48590 = n48589 ^ n43711 ^ n8586 ;
  assign n48591 = ~n48588 & n48590 ;
  assign n48592 = n41588 ^ n36625 ^ 1'b0 ;
  assign n48593 = n47176 & ~n48592 ;
  assign n48594 = n48593 ^ n14850 ^ 1'b0 ;
  assign n48595 = n31679 & ~n35773 ;
  assign n48596 = n1138 & ~n37385 ;
  assign n48597 = n48596 ^ n2826 ^ 1'b0 ;
  assign n48598 = n21632 | n26148 ;
  assign n48599 = ~n29249 & n48598 ;
  assign n48600 = ( n9292 & n42313 ) | ( n9292 & n48599 ) | ( n42313 & n48599 ) ;
  assign n48601 = n14120 ^ n12502 ^ 1'b0 ;
  assign n48602 = n13752 ^ n9357 ^ 1'b0 ;
  assign n48603 = n6343 & n48602 ;
  assign n48604 = n48603 ^ n23949 ^ n23018 ;
  assign n48605 = n13554 | n41931 ;
  assign n48606 = n25164 & ~n48605 ;
  assign n48607 = ( n11852 & n17413 ) | ( n11852 & n18998 ) | ( n17413 & n18998 ) ;
  assign n48608 = n44392 & n48607 ;
  assign n48609 = n10232 & ~n48608 ;
  assign n48614 = n1693 & n8601 ;
  assign n48612 = n21188 & n39675 ;
  assign n48613 = n29048 & n48612 ;
  assign n48615 = n48614 ^ n48613 ^ 1'b0 ;
  assign n48610 = ( n4949 & n19811 ) | ( n4949 & n36033 ) | ( n19811 & n36033 ) ;
  assign n48611 = n19407 & ~n48610 ;
  assign n48616 = n48615 ^ n48611 ^ 1'b0 ;
  assign n48617 = n21305 ^ n1607 ^ 1'b0 ;
  assign n48618 = n16106 | n20343 ;
  assign n48619 = n1704 & ~n48618 ;
  assign n48620 = n48619 ^ n36277 ^ 1'b0 ;
  assign n48621 = ( ~n10411 & n29650 ) | ( ~n10411 & n41434 ) | ( n29650 & n41434 ) ;
  assign n48622 = n33937 ^ n5542 ^ 1'b0 ;
  assign n48623 = n30249 & ~n48622 ;
  assign n48624 = ( ~n13198 & n35191 ) | ( ~n13198 & n48623 ) | ( n35191 & n48623 ) ;
  assign n48625 = ~n1930 & n24438 ;
  assign n48626 = n36109 ^ n11320 ^ 1'b0 ;
  assign n48627 = n27405 & ~n48626 ;
  assign n48628 = n48627 ^ n13078 ^ 1'b0 ;
  assign n48629 = n48625 & n48628 ;
  assign n48630 = n9230 & n11749 ;
  assign n48631 = ~n44353 & n48630 ;
  assign n48635 = n32686 ^ n2557 ^ 1'b0 ;
  assign n48636 = ~n22674 & n48635 ;
  assign n48632 = n33941 ^ n4375 ^ 1'b0 ;
  assign n48633 = n15833 & n48632 ;
  assign n48634 = n5470 & n48633 ;
  assign n48637 = n48636 ^ n48634 ^ 1'b0 ;
  assign n48638 = n7230 | n12880 ;
  assign n48639 = n2619 & ~n48638 ;
  assign n48640 = n48639 ^ n24815 ^ 1'b0 ;
  assign n48641 = n7795 & n13060 ;
  assign n48642 = n15859 ^ n10720 ^ 1'b0 ;
  assign n48643 = n4930 & ~n48642 ;
  assign n48644 = n3915 | n48643 ;
  assign n48645 = ~n48641 & n48644 ;
  assign n48646 = ~n1389 & n10284 ;
  assign n48647 = n27449 & n48646 ;
  assign n48648 = ~n11772 & n24943 ;
  assign n48649 = n19056 ^ n5684 ^ 1'b0 ;
  assign n48650 = n4725 | n48649 ;
  assign n48651 = n33429 ^ n25559 ^ n19234 ;
  assign n48652 = n11762 & n48651 ;
  assign n48653 = n46549 ^ n9852 ^ 1'b0 ;
  assign n48654 = ~n13226 & n37660 ;
  assign n48655 = n19320 | n42624 ;
  assign n48656 = n48655 ^ n42576 ^ n22099 ;
  assign n48657 = n6524 & n48656 ;
  assign n48658 = n48657 ^ n11561 ^ 1'b0 ;
  assign n48659 = n20951 ^ n17371 ^ 1'b0 ;
  assign n48660 = ~n35834 & n48659 ;
  assign n48661 = ( n6866 & n10715 ) | ( n6866 & n12779 ) | ( n10715 & n12779 ) ;
  assign n48662 = n6656 & n48661 ;
  assign n48663 = n25307 & n48662 ;
  assign n48664 = n7577 & n10650 ;
  assign n48665 = n2049 & ~n12532 ;
  assign n48666 = n48665 ^ n8854 ^ 1'b0 ;
  assign n48667 = n48666 ^ n24458 ^ n15964 ;
  assign n48670 = n2433 & ~n21875 ;
  assign n48669 = n16154 & n21624 ;
  assign n48668 = n23464 ^ n12915 ^ 1'b0 ;
  assign n48671 = n48670 ^ n48669 ^ n48668 ;
  assign n48672 = ~n17098 & n36656 ;
  assign n48673 = n48672 ^ n14881 ^ 1'b0 ;
  assign n48674 = n24834 ^ n12752 ^ 1'b0 ;
  assign n48675 = n4904 | n48674 ;
  assign n48676 = n732 | n8947 ;
  assign n48677 = n48676 ^ n16997 ^ 1'b0 ;
  assign n48678 = n7116 & n15392 ;
  assign n48679 = n1506 & n48678 ;
  assign n48680 = n35839 & ~n48679 ;
  assign n48681 = n178 | n7087 ;
  assign n48682 = ~n47878 & n48681 ;
  assign n48683 = ~n15605 & n24388 ;
  assign n48684 = ~n41699 & n48683 ;
  assign n48685 = n16798 | n48684 ;
  assign n48686 = n28895 ^ n1318 ^ 1'b0 ;
  assign n48687 = ( n962 & n1064 ) | ( n962 & ~n9832 ) | ( n1064 & ~n9832 ) ;
  assign n48688 = n18504 | n48687 ;
  assign n48689 = ( n18454 & n25535 ) | ( n18454 & n48688 ) | ( n25535 & n48688 ) ;
  assign n48690 = ~n4681 & n44294 ;
  assign n48691 = n16828 & n27222 ;
  assign n48692 = n45942 ^ n34921 ^ 1'b0 ;
  assign n48693 = n48691 & n48692 ;
  assign n48694 = n21747 | n40338 ;
  assign n48695 = n28319 & n48694 ;
  assign n48696 = n28375 & n48695 ;
  assign n48697 = ~n2933 & n27875 ;
  assign n48698 = n48697 ^ n31325 ^ 1'b0 ;
  assign n48699 = n3035 & ~n10884 ;
  assign n48700 = n26206 & n48699 ;
  assign n48702 = n4717 & ~n14450 ;
  assign n48703 = n48702 ^ n533 ^ 1'b0 ;
  assign n48704 = n3985 & ~n48703 ;
  assign n48705 = n12796 & n48704 ;
  assign n48701 = n1771 & n13002 ;
  assign n48706 = n48705 ^ n48701 ^ 1'b0 ;
  assign n48708 = ( n11927 & n20356 ) | ( n11927 & ~n40641 ) | ( n20356 & ~n40641 ) ;
  assign n48709 = n48708 ^ n48031 ^ n17102 ;
  assign n48707 = n14275 ^ n5418 ^ 1'b0 ;
  assign n48710 = n48709 ^ n48707 ^ 1'b0 ;
  assign n48711 = n7980 | n36420 ;
  assign n48712 = n28428 & ~n48711 ;
  assign n48713 = n6716 | n33821 ;
  assign n48714 = n48713 ^ n26929 ^ 1'b0 ;
  assign n48715 = n14509 ^ n9894 ^ 1'b0 ;
  assign n48716 = n650 & n48715 ;
  assign n48717 = n10020 | n48716 ;
  assign n48718 = n14639 & n48717 ;
  assign n48719 = n7046 | n23143 ;
  assign n48720 = n48719 ^ n48661 ^ 1'b0 ;
  assign n48721 = n21674 ^ n5866 ^ n2302 ;
  assign n48722 = n6498 & ~n7128 ;
  assign n48723 = n48722 ^ n31572 ^ n11936 ;
  assign n48724 = ( n34958 & n48721 ) | ( n34958 & n48723 ) | ( n48721 & n48723 ) ;
  assign n48725 = n11716 ^ n6554 ^ 1'b0 ;
  assign n48726 = n48725 ^ n48305 ^ n6541 ;
  assign n48727 = n30099 ^ n3571 ^ 1'b0 ;
  assign n48728 = n19203 ^ n8745 ^ 1'b0 ;
  assign n48729 = n656 | n19897 ;
  assign n48730 = n48729 ^ n1457 ^ 1'b0 ;
  assign n48731 = ~n25331 & n48730 ;
  assign n48732 = n9914 & n14151 ;
  assign n48733 = n48732 ^ n20110 ^ 1'b0 ;
  assign n48734 = n48733 ^ n20855 ^ 1'b0 ;
  assign n48735 = ~n9656 & n25214 ;
  assign n48736 = ~n34910 & n48735 ;
  assign n48737 = ( n7663 & n16212 ) | ( n7663 & ~n48736 ) | ( n16212 & ~n48736 ) ;
  assign n48738 = n811 | n4454 ;
  assign n48739 = ( n2446 & n40076 ) | ( n2446 & n48738 ) | ( n40076 & n48738 ) ;
  assign n48741 = n17202 ^ n1746 ^ 1'b0 ;
  assign n48742 = n6451 | n48741 ;
  assign n48740 = n3575 & ~n18299 ;
  assign n48743 = n48742 ^ n48740 ^ 1'b0 ;
  assign n48744 = n3776 & ~n42280 ;
  assign n48745 = ~n863 & n44730 ;
  assign n48746 = n48745 ^ n43243 ^ 1'b0 ;
  assign n48747 = n68 & n41247 ;
  assign n48748 = n38610 & n48747 ;
  assign n48750 = n10279 & n32131 ;
  assign n48749 = n4713 | n44668 ;
  assign n48751 = n48750 ^ n48749 ^ 1'b0 ;
  assign n48752 = n26719 & n27095 ;
  assign n48753 = n27339 & n48752 ;
  assign n48754 = n45248 ^ n21837 ^ 1'b0 ;
  assign n48755 = n39810 ^ n17439 ^ 1'b0 ;
  assign n48756 = n929 & n11405 ;
  assign n48757 = n23229 & n48756 ;
  assign n48758 = n18319 & ~n23615 ;
  assign n48759 = ( ~n35329 & n48757 ) | ( ~n35329 & n48758 ) | ( n48757 & n48758 ) ;
  assign n48760 = ~n4385 & n18642 ;
  assign n48761 = ~n17698 & n48760 ;
  assign n48762 = n36928 ^ n16080 ^ 1'b0 ;
  assign n48763 = n48761 | n48762 ;
  assign n48764 = n19289 | n48763 ;
  assign n48765 = n39964 | n45281 ;
  assign n48766 = n16245 ^ n8159 ^ 1'b0 ;
  assign n48768 = n16806 & ~n22690 ;
  assign n48769 = n25966 & n48768 ;
  assign n48767 = n5791 | n13316 ;
  assign n48770 = n48769 ^ n48767 ^ 1'b0 ;
  assign n48771 = n48766 & ~n48770 ;
  assign n48773 = n46620 ^ n14329 ^ n563 ;
  assign n48772 = ~n576 & n30258 ;
  assign n48774 = n48773 ^ n48772 ^ 1'b0 ;
  assign n48775 = n13246 & n48774 ;
  assign n48777 = n30049 ^ n26253 ^ 1'b0 ;
  assign n48778 = n2249 & n48777 ;
  assign n48776 = n21339 & n23363 ;
  assign n48779 = n48778 ^ n48776 ^ 1'b0 ;
  assign n48780 = n7633 & n7722 ;
  assign n48781 = n22900 | n23554 ;
  assign n48782 = n11155 | n48781 ;
  assign n48783 = n5481 & n31770 ;
  assign n48784 = ~n1876 & n48783 ;
  assign n48785 = n2048 & n48784 ;
  assign n48787 = n9027 & n13844 ;
  assign n48788 = ~n3584 & n48787 ;
  assign n48789 = ( n6093 & n22495 ) | ( n6093 & ~n48788 ) | ( n22495 & ~n48788 ) ;
  assign n48786 = n5101 | n38339 ;
  assign n48790 = n48789 ^ n48786 ^ n34000 ;
  assign n48791 = n1578 & n17264 ;
  assign n48792 = n48791 ^ n25054 ^ 1'b0 ;
  assign n48793 = n8544 & n48792 ;
  assign n48794 = ~n5419 & n48793 ;
  assign n48795 = n9143 ^ n4454 ^ 1'b0 ;
  assign n48796 = n6860 & ~n20829 ;
  assign n48797 = n48796 ^ n42121 ^ 1'b0 ;
  assign n48798 = ~n31445 & n48797 ;
  assign n48799 = n4644 | n15993 ;
  assign n48800 = n31621 ^ n14951 ^ n13040 ;
  assign n48801 = n15325 ^ n11150 ^ 1'b0 ;
  assign n48802 = n27924 & n48801 ;
  assign n48803 = n33298 & n48802 ;
  assign n48804 = n13112 ^ n10333 ^ n696 ;
  assign n48805 = n5433 | n45880 ;
  assign n48806 = n45970 ^ n13907 ^ 1'b0 ;
  assign n48807 = n7881 & ~n30487 ;
  assign n48808 = n48807 ^ n23128 ^ 1'b0 ;
  assign n48809 = n6616 & n13780 ;
  assign n48810 = n48809 ^ n18237 ^ 1'b0 ;
  assign n48811 = n2280 & ~n7500 ;
  assign n48812 = ~n9469 & n11302 ;
  assign n48813 = n14154 & n48812 ;
  assign n48814 = n115 | n13969 ;
  assign n48815 = n48814 ^ n11664 ^ 1'b0 ;
  assign n48816 = n27655 ^ n16298 ^ 1'b0 ;
  assign n48817 = n48815 | n48816 ;
  assign n48818 = n9209 & n18228 ;
  assign n48819 = ~n1767 & n14512 ;
  assign n48820 = n25341 ^ n5377 ^ 1'b0 ;
  assign n48821 = n7489 & ~n25885 ;
  assign n48822 = n48821 ^ n41041 ^ n1036 ;
  assign n48823 = n16707 & ~n33629 ;
  assign n48824 = n37727 ^ n13047 ^ 1'b0 ;
  assign n48825 = ~n48823 & n48824 ;
  assign n48826 = ( n11570 & n48822 ) | ( n11570 & ~n48825 ) | ( n48822 & ~n48825 ) ;
  assign n48827 = ~n10830 & n37168 ;
  assign n48828 = n31161 ^ n27105 ^ 1'b0 ;
  assign n48829 = n11599 & ~n48828 ;
  assign n48834 = ( n177 & n4057 ) | ( n177 & ~n34956 ) | ( n4057 & ~n34956 ) ;
  assign n48835 = n48834 ^ n8555 ^ n5563 ;
  assign n48830 = n22733 ^ n14423 ^ n8767 ;
  assign n48831 = n225 & n48830 ;
  assign n48832 = n48831 ^ n153 ^ 1'b0 ;
  assign n48833 = ~n11941 & n48832 ;
  assign n48836 = n48835 ^ n48833 ^ 1'b0 ;
  assign n48837 = ~n27657 & n43739 ;
  assign n48838 = ~n39281 & n48837 ;
  assign n48839 = n17271 ^ n10001 ^ 1'b0 ;
  assign n48840 = n48838 & n48839 ;
  assign n48841 = n4711 ^ n3548 ^ 1'b0 ;
  assign n48843 = n17304 ^ n1623 ^ 1'b0 ;
  assign n48844 = ~n8902 & n48843 ;
  assign n48845 = ~n48843 & n48844 ;
  assign n48842 = n14071 | n19759 ;
  assign n48846 = n48845 ^ n48842 ^ 1'b0 ;
  assign n48847 = n26441 | n48846 ;
  assign n48848 = n6671 & n11533 ;
  assign n48849 = n48848 ^ n24133 ^ 1'b0 ;
  assign n48850 = n23443 & n32874 ;
  assign n48851 = n48849 & n48850 ;
  assign n48852 = n14373 & n25325 ;
  assign n48853 = ~n3039 & n31457 ;
  assign n48854 = n15420 & n48853 ;
  assign n48855 = n22323 ^ n18683 ^ 1'b0 ;
  assign n48856 = n41526 & n48855 ;
  assign n48858 = n8816 | n15138 ;
  assign n48859 = n48858 ^ n5311 ^ 1'b0 ;
  assign n48857 = n16175 & n37124 ;
  assign n48860 = n48859 ^ n48857 ^ 1'b0 ;
  assign n48861 = ~n2346 & n34150 ;
  assign n48862 = n48860 & n48861 ;
  assign n48863 = ~n838 & n13442 ;
  assign n48864 = n48863 ^ n11642 ^ 1'b0 ;
  assign n48867 = ~n228 & n23221 ;
  assign n48865 = n10995 & ~n21651 ;
  assign n48866 = ~n30553 & n48865 ;
  assign n48868 = n48867 ^ n48866 ^ n34720 ;
  assign n48869 = n48864 & n48868 ;
  assign n48870 = ~n1409 & n11295 ;
  assign n48871 = ~n48869 & n48870 ;
  assign n48872 = n3039 & ~n5658 ;
  assign n48873 = ~n9066 & n48872 ;
  assign n48874 = n48873 ^ n13532 ^ 1'b0 ;
  assign n48875 = n48874 ^ n44993 ^ 1'b0 ;
  assign n48876 = n13145 & n27720 ;
  assign n48877 = n34730 & n48876 ;
  assign n48878 = ~n32075 & n44838 ;
  assign n48879 = n48878 ^ n16517 ^ 1'b0 ;
  assign n48880 = n10500 ^ n8380 ^ 1'b0 ;
  assign n48881 = ~n48879 & n48880 ;
  assign n48882 = n48881 ^ n321 ^ 1'b0 ;
  assign n48883 = n11607 | n48882 ;
  assign n48884 = ( n26719 & n27074 ) | ( n26719 & n45073 ) | ( n27074 & n45073 ) ;
  assign n48885 = n27374 | n42016 ;
  assign n48886 = n9241 | n48885 ;
  assign n48887 = n48886 ^ n19025 ^ 1'b0 ;
  assign n48888 = n172 | n652 ;
  assign n48889 = n48888 ^ n23652 ^ 1'b0 ;
  assign n48890 = n34282 ^ n9369 ^ n1876 ;
  assign n48891 = n9345 & n48890 ;
  assign n48892 = ~n14964 & n48891 ;
  assign n48893 = n9139 & n36041 ;
  assign n48894 = n27273 ^ n3840 ^ 1'b0 ;
  assign n48895 = n48893 & n48894 ;
  assign n48896 = ( n12102 & n37661 ) | ( n12102 & n44053 ) | ( n37661 & n44053 ) ;
  assign n48897 = n34935 ^ n20605 ^ 1'b0 ;
  assign n48898 = n4656 ^ n2148 ^ 1'b0 ;
  assign n48899 = n48898 ^ n20240 ^ 1'b0 ;
  assign n48900 = n41049 & n48899 ;
  assign n48901 = n9975 | n22970 ;
  assign n48902 = n48901 ^ n25700 ^ 1'b0 ;
  assign n48903 = ~n10469 & n48902 ;
  assign n48904 = n23378 ^ n15654 ^ n2374 ;
  assign n48905 = n48904 ^ n31232 ^ 1'b0 ;
  assign n48906 = ~n4706 & n48905 ;
  assign n48907 = n14565 ^ n9549 ^ 1'b0 ;
  assign n48908 = n43699 & n48907 ;
  assign n48909 = ~n214 & n6195 ;
  assign n48910 = ~n15235 & n48909 ;
  assign n48911 = n20031 ^ n8536 ^ 1'b0 ;
  assign n48912 = n48910 | n48911 ;
  assign n48913 = n14002 & ~n18351 ;
  assign n48914 = n48913 ^ n645 ^ 1'b0 ;
  assign n48915 = ~n20335 & n29898 ;
  assign n48916 = n48915 ^ n20664 ^ n11519 ;
  assign n48917 = n545 & n44609 ;
  assign n48918 = n953 & n26491 ;
  assign n48919 = n13905 & n48918 ;
  assign n48920 = n6842 & ~n48919 ;
  assign n48921 = n2259 & n16185 ;
  assign n48922 = n1021 & n48921 ;
  assign n48923 = n14674 | n48922 ;
  assign n48927 = n13617 & ~n38141 ;
  assign n48928 = n48927 ^ n20009 ^ 1'b0 ;
  assign n48924 = ~n3898 & n37669 ;
  assign n48925 = n99 & n48924 ;
  assign n48926 = n17168 | n48925 ;
  assign n48929 = n48928 ^ n48926 ^ 1'b0 ;
  assign n48930 = ~n8647 & n21968 ;
  assign n48931 = n8804 | n48930 ;
  assign n48932 = n18820 & n47278 ;
  assign n48933 = n8989 & ~n45608 ;
  assign n48935 = n14499 ^ n13477 ^ 1'b0 ;
  assign n48934 = n47366 ^ n15714 ^ 1'b0 ;
  assign n48936 = n48935 ^ n48934 ^ n34954 ;
  assign n48937 = n43857 ^ n42 ^ 1'b0 ;
  assign n48938 = n23104 & n48937 ;
  assign n48939 = n25396 ^ n20664 ^ 1'b0 ;
  assign n48940 = ~n8414 & n19988 ;
  assign n48941 = n29511 ^ n16106 ^ 1'b0 ;
  assign n48942 = n8452 | n31613 ;
  assign n48943 = ~n7276 & n20100 ;
  assign n48944 = n48942 & n48943 ;
  assign n48945 = n48941 & ~n48944 ;
  assign n48946 = n982 & n17551 ;
  assign n48947 = n48946 ^ n20617 ^ 1'b0 ;
  assign n48948 = n48947 ^ n18399 ^ 1'b0 ;
  assign n48949 = n33468 & n48948 ;
  assign n48950 = n48949 ^ n38642 ^ n8631 ;
  assign n48951 = n23567 ^ n13911 ^ 1'b0 ;
  assign n48952 = n8471 ^ n521 ^ 1'b0 ;
  assign n48953 = n23081 & ~n48952 ;
  assign n48954 = n22771 & n48953 ;
  assign n48955 = n9926 | n14881 ;
  assign n48956 = n24266 | n48955 ;
  assign n48957 = n20185 ^ n4906 ^ 1'b0 ;
  assign n48958 = n48956 & ~n48957 ;
  assign n48959 = n37119 ^ n29376 ^ 1'b0 ;
  assign n48960 = n26459 | n48959 ;
  assign n48961 = n48960 ^ n34647 ^ 1'b0 ;
  assign n48962 = n37112 ^ n8901 ^ 1'b0 ;
  assign n48963 = n48962 ^ n47715 ^ n3191 ;
  assign n48965 = n5673 | n18344 ;
  assign n48964 = n30400 ^ n8028 ^ 1'b0 ;
  assign n48966 = n48965 ^ n48964 ^ n44838 ;
  assign n48967 = n572 & ~n21202 ;
  assign n48968 = n48967 ^ n11593 ^ 1'b0 ;
  assign n48969 = ~n2084 & n17081 ;
  assign n48970 = ( ~n4019 & n48968 ) | ( ~n4019 & n48969 ) | ( n48968 & n48969 ) ;
  assign n48971 = n33852 ^ n9457 ^ 1'b0 ;
  assign n48972 = n4259 | n36278 ;
  assign n48974 = n1081 | n42947 ;
  assign n48975 = n2278 & ~n48974 ;
  assign n48973 = n19361 & ~n29259 ;
  assign n48976 = n48975 ^ n48973 ^ 1'b0 ;
  assign n48977 = n35836 ^ n27340 ^ 1'b0 ;
  assign n48978 = n14910 & n24161 ;
  assign n48979 = n48978 ^ n3079 ^ 1'b0 ;
  assign n48980 = n48979 ^ n24863 ^ 1'b0 ;
  assign n48981 = n20623 | n34695 ;
  assign n48982 = n14158 & ~n48981 ;
  assign n48983 = n42949 ^ n9996 ^ n8294 ;
  assign n48984 = n15405 & ~n23211 ;
  assign n48985 = n3397 ^ n1717 ^ 1'b0 ;
  assign n48986 = n9452 ^ n41 ^ 1'b0 ;
  assign n48987 = ( ~n24302 & n48985 ) | ( ~n24302 & n48986 ) | ( n48985 & n48986 ) ;
  assign n48988 = n1188 & ~n6451 ;
  assign n48989 = n48988 ^ n17130 ^ 1'b0 ;
  assign n48990 = n5708 ^ n1000 ^ 1'b0 ;
  assign n48991 = ~n18699 & n48990 ;
  assign n48992 = n221 & ~n22540 ;
  assign n48993 = n48992 ^ n44550 ^ 1'b0 ;
  assign n48994 = ( n9036 & n20501 ) | ( n9036 & ~n22208 ) | ( n20501 & ~n22208 ) ;
  assign n48995 = ~n10222 & n41667 ;
  assign n48996 = n48995 ^ n38566 ^ 1'b0 ;
  assign n48997 = ~n5876 & n7646 ;
  assign n48998 = ~n23309 & n48997 ;
  assign n48999 = n2571 & n48998 ;
  assign n49000 = n12079 ^ n3614 ^ 1'b0 ;
  assign n49001 = n48999 & ~n49000 ;
  assign n49002 = n49001 ^ n6403 ^ 1'b0 ;
  assign n49003 = n44366 ^ n720 ^ 1'b0 ;
  assign n49004 = ( ~n1885 & n2546 ) | ( ~n1885 & n35339 ) | ( n2546 & n35339 ) ;
  assign n49005 = n184 & n15226 ;
  assign n49006 = ~n49004 & n49005 ;
  assign n49007 = n4469 & ~n4768 ;
  assign n49008 = ~n6197 & n49007 ;
  assign n49009 = ( n91 & ~n41748 ) | ( n91 & n49008 ) | ( ~n41748 & n49008 ) ;
  assign n49010 = n21984 & ~n32709 ;
  assign n49011 = ( ~n4345 & n28301 ) | ( ~n4345 & n41598 ) | ( n28301 & n41598 ) ;
  assign n49012 = n27171 ^ n17335 ^ 1'b0 ;
  assign n49013 = n13899 | n49012 ;
  assign n49014 = n34337 | n49013 ;
  assign n49015 = n49014 ^ n20116 ^ 1'b0 ;
  assign n49016 = ~n21382 & n39075 ;
  assign n49017 = ~n13594 & n49016 ;
  assign n49018 = n24715 | n49017 ;
  assign n49019 = n19739 | n29795 ;
  assign n49020 = n3607 | n49019 ;
  assign n49021 = n49020 ^ n32339 ^ 1'b0 ;
  assign n49025 = n14732 | n15718 ;
  assign n49026 = n49025 ^ n31863 ^ 1'b0 ;
  assign n49022 = n16802 ^ n11121 ^ 1'b0 ;
  assign n49023 = n49022 ^ n37127 ^ 1'b0 ;
  assign n49024 = n740 & n49023 ;
  assign n49027 = n49026 ^ n49024 ^ 1'b0 ;
  assign n49028 = n32186 ^ n4308 ^ 1'b0 ;
  assign n49029 = n2939 & ~n23706 ;
  assign n49030 = ~n7215 & n49029 ;
  assign n49031 = n13169 & n43564 ;
  assign n49032 = ~n5615 & n6654 ;
  assign n49033 = n49032 ^ n27853 ^ 1'b0 ;
  assign n49034 = n12385 & ~n13684 ;
  assign n49035 = n16035 ^ n10689 ^ 1'b0 ;
  assign n49036 = ~n720 & n5754 ;
  assign n49037 = ~n36380 & n49036 ;
  assign n49038 = ~n14559 & n49037 ;
  assign n49039 = n26941 ^ n8534 ^ 1'b0 ;
  assign n49040 = n32669 | n49039 ;
  assign n49041 = n3387 | n49040 ;
  assign n49042 = n29078 ^ n3446 ^ 1'b0 ;
  assign n49043 = n6027 & ~n13896 ;
  assign n49044 = n24777 & n49043 ;
  assign n49045 = n22361 ^ n4351 ^ 1'b0 ;
  assign n49046 = n39823 & ~n49045 ;
  assign n49047 = n49046 ^ n47104 ^ 1'b0 ;
  assign n49048 = ~n24482 & n49047 ;
  assign n49049 = n16582 & ~n18154 ;
  assign n49050 = n17830 & n26793 ;
  assign n49051 = n19434 & ~n49050 ;
  assign n49052 = n6564 & ~n15903 ;
  assign n49053 = n2078 & n49052 ;
  assign n49054 = ( n10178 & ~n40506 ) | ( n10178 & n49053 ) | ( ~n40506 & n49053 ) ;
  assign n49055 = n29654 ^ n11245 ^ 1'b0 ;
  assign n49056 = ( n4319 & ~n5311 ) | ( n4319 & n49055 ) | ( ~n5311 & n49055 ) ;
  assign n49057 = n17556 & ~n25879 ;
  assign n49058 = ~n28130 & n49057 ;
  assign n49059 = ( ~n32227 & n35341 ) | ( ~n32227 & n49058 ) | ( n35341 & n49058 ) ;
  assign n49060 = ~n12149 & n27868 ;
  assign n49061 = n49060 ^ n31724 ^ 1'b0 ;
  assign n49062 = n7383 ^ n6370 ^ 1'b0 ;
  assign n49063 = n24525 ^ n21260 ^ 1'b0 ;
  assign n49064 = n1540 & ~n2528 ;
  assign n49065 = n49064 ^ n20491 ^ 1'b0 ;
  assign n49066 = n1773 & ~n49065 ;
  assign n49067 = ~n49063 & n49066 ;
  assign n49068 = n3288 & ~n5395 ;
  assign n49069 = n36234 & n49068 ;
  assign n49070 = ~n13747 & n48238 ;
  assign n49071 = n22712 & n49070 ;
  assign n49072 = n1295 & n13680 ;
  assign n49073 = ( n22673 & ~n46041 ) | ( n22673 & n47095 ) | ( ~n46041 & n47095 ) ;
  assign n49074 = ( n15213 & n32621 ) | ( n15213 & n46684 ) | ( n32621 & n46684 ) ;
  assign n49075 = n4751 ^ n729 ^ 1'b0 ;
  assign n49076 = n17717 & n49075 ;
  assign n49077 = n617 & ~n48423 ;
  assign n49078 = n34184 ^ n31550 ^ 1'b0 ;
  assign n49079 = ~n4140 & n5978 ;
  assign n49080 = n21238 & n49079 ;
  assign n49081 = n29381 ^ n609 ^ 1'b0 ;
  assign n49082 = ~n49080 & n49081 ;
  assign n49083 = ( ~n34836 & n35308 ) | ( ~n34836 & n37570 ) | ( n35308 & n37570 ) ;
  assign n49084 = n49083 ^ n30926 ^ 1'b0 ;
  assign n49085 = n29041 & ~n49084 ;
  assign n49086 = n16536 ^ n6991 ^ 1'b0 ;
  assign n49087 = ( ~n20439 & n24756 ) | ( ~n20439 & n49086 ) | ( n24756 & n49086 ) ;
  assign n49088 = ( n37358 & n49085 ) | ( n37358 & ~n49087 ) | ( n49085 & ~n49087 ) ;
  assign n49089 = ( ~n2124 & n32358 ) | ( ~n2124 & n49088 ) | ( n32358 & n49088 ) ;
  assign n49090 = ( n7949 & n16620 ) | ( n7949 & n26786 ) | ( n16620 & n26786 ) ;
  assign n49091 = n10895 & ~n11456 ;
  assign n49092 = n49091 ^ n5590 ^ 1'b0 ;
  assign n49093 = ~n44759 & n49092 ;
  assign n49094 = ~n4985 & n12874 ;
  assign n49095 = n49094 ^ n38605 ^ 1'b0 ;
  assign n49096 = n17885 & n43377 ;
  assign n49097 = n4567 & ~n34556 ;
  assign n49098 = n24530 | n49097 ;
  assign n49099 = n49098 ^ n30538 ^ 1'b0 ;
  assign n49100 = ~n2502 & n10772 ;
  assign n49101 = n6520 & ~n24984 ;
  assign n49102 = ~n49100 & n49101 ;
  assign n49103 = n41796 & ~n49102 ;
  assign n49104 = n17991 ^ n15105 ^ n10445 ;
  assign n49105 = n11967 ^ n11341 ^ n1926 ;
  assign n49106 = n2784 & n49105 ;
  assign n49107 = n28143 ^ n22925 ^ n14741 ;
  assign n49108 = ~n47880 & n49107 ;
  assign n49109 = n37376 ^ n10452 ^ 1'b0 ;
  assign n49110 = ~n49108 & n49109 ;
  assign n49111 = n32276 & n49110 ;
  assign n49112 = ~n12543 & n37256 ;
  assign n49113 = n49112 ^ n32782 ^ 1'b0 ;
  assign n49114 = n16679 ^ n2784 ^ 1'b0 ;
  assign n49115 = n39363 ^ n38614 ^ n2885 ;
  assign n49116 = n37749 ^ n33498 ^ 1'b0 ;
  assign n49117 = n12849 ^ n11381 ^ 1'b0 ;
  assign n49118 = n21644 | n49117 ;
  assign n49119 = n49118 ^ n43881 ^ 1'b0 ;
  assign n49120 = ~n48998 & n49119 ;
  assign n49121 = n17864 | n22376 ;
  assign n49122 = n20288 & ~n49121 ;
  assign n49123 = n5418 & ~n20213 ;
  assign n49124 = n8600 | n23802 ;
  assign n49125 = n30673 & ~n49124 ;
  assign n49126 = n20464 | n49125 ;
  assign n49127 = n10523 & ~n10843 ;
  assign n49128 = n4156 ^ n2804 ^ 1'b0 ;
  assign n49129 = ( n10975 & n44084 ) | ( n10975 & ~n49128 ) | ( n44084 & ~n49128 ) ;
  assign n49130 = n49129 ^ n29962 ^ 1'b0 ;
  assign n49131 = n49127 & n49130 ;
  assign n49132 = n49131 ^ n12969 ^ 1'b0 ;
  assign n49133 = n6399 ^ n2886 ^ 1'b0 ;
  assign n49134 = n13448 | n49133 ;
  assign n49135 = n16712 & ~n49134 ;
  assign n49136 = ~n34805 & n49135 ;
  assign n49137 = n11003 & ~n31533 ;
  assign n49138 = n8894 & ~n13800 ;
  assign n49141 = ~n7158 & n11090 ;
  assign n49142 = n49141 ^ n2470 ^ 1'b0 ;
  assign n49139 = n41971 ^ n9060 ^ 1'b0 ;
  assign n49140 = ~n5139 & n49139 ;
  assign n49143 = n49142 ^ n49140 ^ n34525 ;
  assign n49144 = n27351 ^ n19277 ^ 1'b0 ;
  assign n49145 = n19976 & n49144 ;
  assign n49146 = n49145 ^ n35190 ^ n25606 ;
  assign n49147 = ~n8303 & n12400 ;
  assign n49148 = n49147 ^ n25199 ^ 1'b0 ;
  assign n49149 = n2695 & ~n49134 ;
  assign n49150 = n7503 & n20024 ;
  assign n49151 = n7383 & ~n28215 ;
  assign n49152 = ~n15283 & n49151 ;
  assign n49153 = n49152 ^ n47050 ^ n867 ;
  assign n49154 = ~n3579 & n18966 ;
  assign n49155 = n33584 ^ n32911 ^ 1'b0 ;
  assign n49156 = n21331 | n49155 ;
  assign n49157 = n16620 & n38023 ;
  assign n49158 = ~n29585 & n49157 ;
  assign n49159 = n29746 ^ n18380 ^ 1'b0 ;
  assign n49160 = n44344 ^ n4123 ^ 1'b0 ;
  assign n49161 = ~n49159 & n49160 ;
  assign n49163 = n750 & n27540 ;
  assign n49164 = n49163 ^ n32553 ^ 1'b0 ;
  assign n49162 = n37251 ^ n31445 ^ n14342 ;
  assign n49165 = n49164 ^ n49162 ^ 1'b0 ;
  assign n49166 = n11029 & ~n37393 ;
  assign n49167 = n49166 ^ n11890 ^ 1'b0 ;
  assign n49168 = ~n4132 & n49167 ;
  assign n49169 = n14471 ^ n891 ^ 1'b0 ;
  assign n49170 = ( n14243 & ~n23312 ) | ( n14243 & n24923 ) | ( ~n23312 & n24923 ) ;
  assign n49172 = ( ~n3523 & n37270 ) | ( ~n3523 & n45574 ) | ( n37270 & n45574 ) ;
  assign n49173 = ~n34969 & n49172 ;
  assign n49171 = n3858 & n13449 ;
  assign n49174 = n49173 ^ n49171 ^ n21564 ;
  assign n49175 = ~n49170 & n49174 ;
  assign n49176 = n6147 & ~n9538 ;
  assign n49177 = n49176 ^ n9347 ^ 1'b0 ;
  assign n49178 = n1803 & n49177 ;
  assign n49179 = n49178 ^ n20588 ^ n7847 ;
  assign n49180 = n37719 & n49179 ;
  assign n49181 = n35584 & n49180 ;
  assign n49182 = n10811 & n30158 ;
  assign n49183 = n13909 & n49182 ;
  assign n49184 = ~n9097 & n11769 ;
  assign n49185 = n19491 | n49184 ;
  assign n49186 = n2905 | n7975 ;
  assign n49187 = n49186 ^ n16426 ^ n6648 ;
  assign n49188 = ( n2216 & n22645 ) | ( n2216 & ~n33025 ) | ( n22645 & ~n33025 ) ;
  assign n49189 = n10187 | n16727 ;
  assign n49190 = n4848 | n49189 ;
  assign n49191 = ( ~n1913 & n11374 ) | ( ~n1913 & n16582 ) | ( n11374 & n16582 ) ;
  assign n49192 = n49191 ^ n19371 ^ 1'b0 ;
  assign n49193 = ~n12805 & n17528 ;
  assign n49194 = n49193 ^ n39094 ^ 1'b0 ;
  assign n49195 = ~n32649 & n42810 ;
  assign n49196 = n49195 ^ n27020 ^ 1'b0 ;
  assign n49197 = n49196 ^ n35093 ^ n3093 ;
  assign n49198 = n12618 ^ n1328 ^ 1'b0 ;
  assign n49199 = n10002 | n49198 ;
  assign n49200 = n7804 ^ n2636 ^ n1992 ;
  assign n49201 = ~n23035 & n49200 ;
  assign n49202 = n49201 ^ n23339 ^ 1'b0 ;
  assign n49203 = ~n733 & n5822 ;
  assign n49204 = n49203 ^ n27867 ^ 1'b0 ;
  assign n49205 = n49179 & ~n49204 ;
  assign n49206 = n49205 ^ n15732 ^ 1'b0 ;
  assign n49207 = n23831 & ~n25063 ;
  assign n49208 = n49207 ^ n30847 ^ 1'b0 ;
  assign n49209 = n11356 & ~n45141 ;
  assign n49210 = n49209 ^ n4188 ^ 1'b0 ;
  assign n49211 = n18044 ^ n9914 ^ 1'b0 ;
  assign n49212 = n43918 ^ n36837 ^ n10991 ;
  assign n49213 = n39045 ^ n38435 ^ 1'b0 ;
  assign n49214 = n43341 ^ n40165 ^ 1'b0 ;
  assign n49215 = n29319 ^ n21347 ^ 1'b0 ;
  assign n49216 = n3370 & ~n10227 ;
  assign n49217 = ( n23042 & ~n41206 ) | ( n23042 & n49039 ) | ( ~n41206 & n49039 ) ;
  assign n49218 = n23342 & ~n25067 ;
  assign n49219 = n4142 & n43641 ;
  assign n49220 = n49219 ^ n9376 ^ 1'b0 ;
  assign n49221 = n3341 | n49220 ;
  assign n49222 = n24863 | n37252 ;
  assign n49223 = n23540 ^ n14286 ^ 1'b0 ;
  assign n49224 = n13608 | n49223 ;
  assign n49225 = ~n15555 & n33056 ;
  assign n49226 = n17932 & n49225 ;
  assign n49227 = n49226 ^ n13516 ^ n11638 ;
  assign n49228 = n1565 & ~n49227 ;
  assign n49229 = n49224 & n49228 ;
  assign n49231 = n24665 | n29721 ;
  assign n49230 = n34485 ^ n17034 ^ 1'b0 ;
  assign n49232 = n49231 ^ n49230 ^ 1'b0 ;
  assign n49233 = n21628 ^ n2556 ^ 1'b0 ;
  assign n49234 = n401 & ~n49233 ;
  assign n49235 = n45287 ^ n24207 ^ 1'b0 ;
  assign n49236 = n9760 & n49235 ;
  assign n49237 = n7594 ^ n4936 ^ n826 ;
  assign n49238 = ~n43298 & n49237 ;
  assign n49241 = n36221 ^ n22561 ^ n299 ;
  assign n49242 = ~n21411 & n49241 ;
  assign n49239 = ( n38838 & n41759 ) | ( n38838 & ~n48985 ) | ( n41759 & ~n48985 ) ;
  assign n49240 = n38476 | n49239 ;
  assign n49243 = n49242 ^ n49240 ^ 1'b0 ;
  assign n49244 = ( n7977 & n30357 ) | ( n7977 & ~n31015 ) | ( n30357 & ~n31015 ) ;
  assign n49245 = n2147 & ~n3805 ;
  assign n49246 = ~n49244 & n49245 ;
  assign n49247 = n47553 ^ n23341 ^ 1'b0 ;
  assign n49248 = n46307 & ~n49247 ;
  assign n49249 = ~n3460 & n12332 ;
  assign n49250 = n49249 ^ n29192 ^ n818 ;
  assign n49251 = n49250 ^ n44133 ^ n24375 ;
  assign n49252 = ( n10745 & n35215 ) | ( n10745 & n45808 ) | ( n35215 & n45808 ) ;
  assign n49253 = n36683 ^ n17740 ^ 1'b0 ;
  assign n49255 = n13846 ^ n8530 ^ n8496 ;
  assign n49256 = ~n16627 & n49255 ;
  assign n49254 = n6288 & ~n18090 ;
  assign n49257 = n49256 ^ n49254 ^ 1'b0 ;
  assign n49258 = n11872 | n49257 ;
  assign n49259 = n35355 ^ n6877 ^ 1'b0 ;
  assign n49260 = n36027 & n49259 ;
  assign n49261 = n962 & ~n30197 ;
  assign n49262 = ~n9265 & n49261 ;
  assign n49263 = n33213 ^ n14414 ^ 1'b0 ;
  assign n49264 = n3218 | n14718 ;
  assign n49265 = ~n10178 & n20959 ;
  assign n49266 = n49265 ^ n47050 ^ n18381 ;
  assign n49267 = n25639 ^ n1450 ^ 1'b0 ;
  assign n49268 = n2060 | n49267 ;
  assign n49269 = n49268 ^ n1426 ^ n1175 ;
  assign n49270 = n37160 ^ n6676 ^ 1'b0 ;
  assign n49271 = n46140 & n49270 ;
  assign n49272 = n13849 & n49271 ;
  assign n49273 = n24618 & ~n41845 ;
  assign n49274 = n31650 ^ n6616 ^ 1'b0 ;
  assign n49275 = ~n38912 & n49274 ;
  assign n49276 = ~n3308 & n49275 ;
  assign n49277 = n1487 & ~n48890 ;
  assign n49278 = n49277 ^ n77 ^ 1'b0 ;
  assign n49279 = n769 | n10360 ;
  assign n49280 = n34677 | n49279 ;
  assign n49281 = n137 & ~n46871 ;
  assign n49282 = n18373 & n49281 ;
  assign n49283 = n6750 | n44361 ;
  assign n49284 = n49283 ^ n43124 ^ n4812 ;
  assign n49285 = n3205 & ~n15715 ;
  assign n49286 = n49285 ^ n563 ^ 1'b0 ;
  assign n49287 = n9857 & n10544 ;
  assign n49288 = n8740 | n17109 ;
  assign n49289 = n28825 & ~n49288 ;
  assign n49290 = n15349 & ~n49289 ;
  assign n49291 = n49290 ^ n16738 ^ 1'b0 ;
  assign n49292 = n9395 & n9614 ;
  assign n49293 = n5240 & ~n26759 ;
  assign n49294 = n18339 & n49293 ;
  assign n49295 = n38683 ^ n9419 ^ 1'b0 ;
  assign n49296 = n5381 & n49295 ;
  assign n49297 = n2873 | n18324 ;
  assign n49298 = n49296 | n49297 ;
  assign n49299 = n17060 | n41494 ;
  assign n49300 = ( n4486 & n8319 ) | ( n4486 & n35571 ) | ( n8319 & n35571 ) ;
  assign n49301 = n13102 ^ n5159 ^ 1'b0 ;
  assign n49302 = ~n2944 & n4391 ;
  assign n49303 = n49302 ^ n57 ^ 1'b0 ;
  assign n49304 = n12698 & ~n18950 ;
  assign n49305 = n49304 ^ n30746 ^ 1'b0 ;
  assign n49306 = n37068 ^ n15338 ^ 1'b0 ;
  assign n49307 = ~n6041 & n49306 ;
  assign n49308 = n13819 | n31908 ;
  assign n49309 = n49308 ^ n6433 ^ 1'b0 ;
  assign n49310 = n11356 & ~n37048 ;
  assign n49311 = ( n25843 & n45647 ) | ( n25843 & n49310 ) | ( n45647 & n49310 ) ;
  assign n49312 = n17608 & ~n49311 ;
  assign n49314 = n16979 ^ n2776 ^ 1'b0 ;
  assign n49315 = n24169 | n49314 ;
  assign n49313 = n28533 & ~n38738 ;
  assign n49316 = n49315 ^ n49313 ^ 1'b0 ;
  assign n49317 = n2546 & n49316 ;
  assign n49318 = n49317 ^ n17854 ^ 1'b0 ;
  assign n49319 = n12966 & ~n29837 ;
  assign n49320 = n49319 ^ n3644 ^ 1'b0 ;
  assign n49321 = n45755 & ~n49320 ;
  assign n49322 = n24090 | n37995 ;
  assign n49323 = n49322 ^ n16168 ^ 1'b0 ;
  assign n49324 = n41474 ^ n4978 ^ 1'b0 ;
  assign n49325 = n11371 & n49324 ;
  assign n49326 = ~n7734 & n33646 ;
  assign n49327 = n9840 & n49326 ;
  assign n49328 = n26480 | n33664 ;
  assign n49329 = n49328 ^ n27622 ^ 1'b0 ;
  assign n49331 = ~n254 & n7144 ;
  assign n49330 = ~n11038 & n17371 ;
  assign n49332 = n49331 ^ n49330 ^ 1'b0 ;
  assign n49333 = ~n8166 & n8693 ;
  assign n49334 = n49333 ^ n28185 ^ 1'b0 ;
  assign n49335 = n8581 | n49334 ;
  assign n49336 = n49335 ^ n9186 ^ 1'b0 ;
  assign n49337 = n23016 ^ n3864 ^ 1'b0 ;
  assign n49338 = n452 & ~n49337 ;
  assign n49339 = ~n49336 & n49338 ;
  assign n49340 = ~n25121 & n25556 ;
  assign n49341 = ( n45766 & n46651 ) | ( n45766 & n49340 ) | ( n46651 & n49340 ) ;
  assign n49342 = n35724 ^ n6353 ^ 1'b0 ;
  assign n49343 = n18768 | n42040 ;
  assign n49344 = n49343 ^ n39455 ^ 1'b0 ;
  assign n49346 = n9557 & n22024 ;
  assign n49347 = n49346 ^ n48013 ^ 1'b0 ;
  assign n49345 = n39034 & ~n48726 ;
  assign n49348 = n49347 ^ n49345 ^ 1'b0 ;
  assign n49349 = n6903 & ~n27738 ;
  assign n49350 = n49349 ^ n47572 ^ 1'b0 ;
  assign n49352 = n18780 ^ n7670 ^ n852 ;
  assign n49351 = n8302 & n42883 ;
  assign n49353 = n49352 ^ n49351 ^ 1'b0 ;
  assign n49354 = n23994 & ~n49353 ;
  assign n49355 = n16269 & ~n44720 ;
  assign n49356 = n49355 ^ n36491 ^ 1'b0 ;
  assign n49357 = n26802 ^ n10163 ^ 1'b0 ;
  assign n49358 = n49357 ^ n20157 ^ n10348 ;
  assign n49359 = ~n15682 & n34665 ;
  assign n49360 = n14145 & ~n23553 ;
  assign n49361 = n49360 ^ n5564 ^ 1'b0 ;
  assign n49362 = n49361 ^ n29736 ^ 1'b0 ;
  assign n49363 = n4085 & n49362 ;
  assign n49364 = n11323 & ~n14666 ;
  assign n49365 = ~n25388 & n49364 ;
  assign n49366 = n22912 ^ n6805 ^ 1'b0 ;
  assign n49367 = n36897 ^ n398 ^ 1'b0 ;
  assign n49368 = n15066 & ~n49367 ;
  assign n49369 = n3304 & n30898 ;
  assign n49370 = ( n432 & n31344 ) | ( n432 & n43837 ) | ( n31344 & n43837 ) ;
  assign n49371 = n33464 ^ n12136 ^ 1'b0 ;
  assign n49372 = n18555 & ~n18836 ;
  assign n49373 = n14175 & n25350 ;
  assign n49374 = ~n29657 & n49373 ;
  assign n49375 = n1781 & ~n11276 ;
  assign n49376 = n1395 | n49375 ;
  assign n49377 = n49376 ^ n31268 ^ 1'b0 ;
  assign n49378 = n19453 & n49377 ;
  assign n49379 = n49378 ^ n43919 ^ 1'b0 ;
  assign n49380 = n49379 ^ n403 ^ 1'b0 ;
  assign n49381 = ~n49374 & n49380 ;
  assign n49382 = n22004 & n23019 ;
  assign n49383 = n9759 | n13787 ;
  assign n49384 = n11567 & n44939 ;
  assign n49385 = n9284 | n49384 ;
  assign n49390 = n35635 ^ n29785 ^ 1'b0 ;
  assign n49391 = ~n3222 & n49390 ;
  assign n49386 = n27758 ^ n14898 ^ 1'b0 ;
  assign n49387 = n27289 & ~n49386 ;
  assign n49388 = ( n11829 & n25521 ) | ( n11829 & ~n49387 ) | ( n25521 & ~n49387 ) ;
  assign n49389 = n49388 ^ n6312 ^ 1'b0 ;
  assign n49392 = n49391 ^ n49389 ^ 1'b0 ;
  assign n49395 = n28301 ^ n2314 ^ 1'b0 ;
  assign n49393 = n32196 ^ n19047 ^ 1'b0 ;
  assign n49394 = n44921 & n49393 ;
  assign n49396 = n49395 ^ n49394 ^ 1'b0 ;
  assign n49397 = n26210 & ~n49396 ;
  assign n49398 = ~n3140 & n14386 ;
  assign n49399 = n13566 & n49398 ;
  assign n49400 = n35755 & n49399 ;
  assign n49401 = n47696 ^ n44902 ^ 1'b0 ;
  assign n49404 = n19525 ^ n11234 ^ n3281 ;
  assign n49402 = n8896 ^ n6700 ^ 1'b0 ;
  assign n49403 = ~n25523 & n49402 ;
  assign n49405 = n49404 ^ n49403 ^ n6186 ;
  assign n49406 = n25472 & n25682 ;
  assign n49407 = n49406 ^ n4712 ^ 1'b0 ;
  assign n49408 = n49407 ^ n36258 ^ 1'b0 ;
  assign n49409 = n49408 ^ n5099 ^ 1'b0 ;
  assign n49410 = n8431 ^ n5204 ^ 1'b0 ;
  assign n49411 = n49410 ^ n23914 ^ 1'b0 ;
  assign n49412 = n43103 ^ n928 ^ 1'b0 ;
  assign n49413 = ( ~n839 & n17062 ) | ( ~n839 & n43142 ) | ( n17062 & n43142 ) ;
  assign n49414 = n9601 ^ n8247 ^ 1'b0 ;
  assign n49415 = n33887 ^ n9716 ^ 1'b0 ;
  assign n49416 = n28259 | n49415 ;
  assign n49417 = n9251 | n49416 ;
  assign n49418 = ~n13330 & n24333 ;
  assign n49419 = ~n2580 & n11715 ;
  assign n49420 = n2571 & ~n26300 ;
  assign n49421 = n49420 ^ n36269 ^ 1'b0 ;
  assign n49422 = n20733 | n49421 ;
  assign n49423 = n9550 & n16756 ;
  assign n49424 = n49423 ^ n4361 ^ 1'b0 ;
  assign n49425 = ~n21027 & n49424 ;
  assign n49426 = n23528 ^ n22970 ^ 1'b0 ;
  assign n49427 = ~n22202 & n29903 ;
  assign n49428 = ~n38393 & n49427 ;
  assign n49429 = ~n6181 & n47780 ;
  assign n49430 = n15645 ^ n10707 ^ n989 ;
  assign n49431 = n4141 | n49430 ;
  assign n49432 = n49429 | n49431 ;
  assign n49433 = ( ~n7017 & n17828 ) | ( ~n7017 & n49432 ) | ( n17828 & n49432 ) ;
  assign n49434 = n37187 ^ n5376 ^ 1'b0 ;
  assign n49435 = n39083 ^ n15660 ^ 1'b0 ;
  assign n49436 = n2350 | n49435 ;
  assign n49437 = n47929 | n49436 ;
  assign n49438 = n49437 ^ n23294 ^ 1'b0 ;
  assign n49439 = n23755 ^ n2568 ^ 1'b0 ;
  assign n49440 = n603 | n49439 ;
  assign n49441 = n7943 & n11084 ;
  assign n49442 = n28428 & n49441 ;
  assign n49443 = n38779 ^ n10042 ^ 1'b0 ;
  assign n49444 = n7818 & n49443 ;
  assign n49445 = ~n12460 & n15408 ;
  assign n49446 = ( ~n5816 & n17389 ) | ( ~n5816 & n43074 ) | ( n17389 & n43074 ) ;
  assign n49447 = n10868 & n14833 ;
  assign n49448 = n49447 ^ n46423 ^ 1'b0 ;
  assign n49449 = n159 | n49448 ;
  assign n49450 = ~n4932 & n35360 ;
  assign n49451 = ( n5373 & n11896 ) | ( n5373 & n18251 ) | ( n11896 & n18251 ) ;
  assign n49452 = n22542 ^ n1866 ^ 1'b0 ;
  assign n49453 = n3082 | n17935 ;
  assign n49454 = ( n14052 & n49452 ) | ( n14052 & n49453 ) | ( n49452 & n49453 ) ;
  assign n49455 = n1512 | n19558 ;
  assign n49456 = n49455 ^ n835 ^ 1'b0 ;
  assign n49457 = n21469 | n49456 ;
  assign n49458 = n16880 & ~n49457 ;
  assign n49459 = n39954 ^ n25269 ^ 1'b0 ;
  assign n49460 = n17643 ^ n8926 ^ 1'b0 ;
  assign n49461 = ~n28453 & n49460 ;
  assign n49462 = n28143 ^ n24825 ^ 1'b0 ;
  assign n49463 = n49461 & ~n49462 ;
  assign n49464 = n12237 & ~n31575 ;
  assign n49465 = ~n40707 & n49464 ;
  assign n49466 = ~n8913 & n29767 ;
  assign n49467 = n49466 ^ n45845 ^ 1'b0 ;
  assign n49468 = n12283 | n49467 ;
  assign n49469 = n49468 ^ n32425 ^ 1'b0 ;
  assign n49470 = n1105 | n11859 ;
  assign n49471 = n49470 ^ n304 ^ 1'b0 ;
  assign n49472 = ~n10838 & n49471 ;
  assign n49473 = ~n35133 & n44001 ;
  assign n49474 = n49473 ^ n5333 ^ 1'b0 ;
  assign n49475 = n24577 ^ n6292 ^ n4847 ;
  assign n49476 = ~n14437 & n29017 ;
  assign n49477 = ( n41433 & n41870 ) | ( n41433 & n49476 ) | ( n41870 & n49476 ) ;
  assign n49478 = n11644 ^ n8096 ^ 1'b0 ;
  assign n49479 = n8355 | n49478 ;
  assign n49480 = n49479 ^ n6272 ^ 1'b0 ;
  assign n49481 = ~n30427 & n49480 ;
  assign n49482 = n7035 & n10003 ;
  assign n49483 = ( n937 & ~n1787 ) | ( n937 & n3170 ) | ( ~n1787 & n3170 ) ;
  assign n49484 = n49483 ^ n20000 ^ 1'b0 ;
  assign n49485 = ~n26185 & n49484 ;
  assign n49486 = n13962 & n49485 ;
  assign n49487 = n49482 & n49486 ;
  assign n49488 = n23340 ^ n172 ^ 1'b0 ;
  assign n49489 = n25372 & ~n49488 ;
  assign n49490 = n35515 ^ n9785 ^ 1'b0 ;
  assign n49491 = n1876 & n2239 ;
  assign n49492 = ( ~n4226 & n17424 ) | ( ~n4226 & n49491 ) | ( n17424 & n49491 ) ;
  assign n49493 = n49492 ^ n177 ^ 1'b0 ;
  assign n49494 = n40042 & ~n49493 ;
  assign n49495 = n45306 ^ n2330 ^ 1'b0 ;
  assign n49496 = n20798 ^ n20649 ^ n8577 ;
  assign n49497 = n18265 | n49496 ;
  assign n49498 = n8759 & ~n49497 ;
  assign n49499 = n7219 & n7728 ;
  assign n49500 = n49499 ^ n35209 ^ 1'b0 ;
  assign n49501 = n17936 & n49500 ;
  assign n49502 = n18544 & n24743 ;
  assign n49503 = n49502 ^ n44804 ^ 1'b0 ;
  assign n49504 = n4231 | n13151 ;
  assign n49505 = n19083 ^ n10325 ^ 1'b0 ;
  assign n49506 = ~n49504 & n49505 ;
  assign n49507 = n7818 & ~n28100 ;
  assign n49508 = n49507 ^ n29948 ^ 1'b0 ;
  assign n49511 = n15170 & ~n20077 ;
  assign n49512 = n6294 & n49511 ;
  assign n49509 = n34114 ^ n19317 ^ 1'b0 ;
  assign n49510 = n25893 & n49509 ;
  assign n49513 = n49512 ^ n49510 ^ 1'b0 ;
  assign n49514 = n21556 & ~n49513 ;
  assign n49515 = ~n39824 & n49514 ;
  assign n49516 = n14487 ^ n8465 ^ 1'b0 ;
  assign n49517 = n29523 ^ n24897 ^ n12530 ;
  assign n49518 = n49517 ^ n19433 ^ 1'b0 ;
  assign n49519 = ~n49516 & n49518 ;
  assign n49520 = n49519 ^ n35666 ^ 1'b0 ;
  assign n49521 = ( n3855 & n5722 ) | ( n3855 & n45059 ) | ( n5722 & n45059 ) ;
  assign n49522 = n45335 | n49521 ;
  assign n49523 = n1796 & ~n49522 ;
  assign n49525 = n12603 ^ n2284 ^ n1256 ;
  assign n49524 = n3662 & n38199 ;
  assign n49526 = n49525 ^ n49524 ^ 1'b0 ;
  assign n49527 = n21525 ^ n5718 ^ 1'b0 ;
  assign n49528 = ~n5311 & n37100 ;
  assign n49529 = n49528 ^ n3274 ^ 1'b0 ;
  assign n49530 = ~n4099 & n9737 ;
  assign n49531 = n5113 ^ n4371 ^ 1'b0 ;
  assign n49532 = n49531 ^ n22711 ^ 1'b0 ;
  assign n49533 = n17153 | n49532 ;
  assign n49534 = n5778 | n49533 ;
  assign n49535 = n49530 | n49534 ;
  assign n49536 = n1083 & ~n42987 ;
  assign n49537 = n37438 ^ n21611 ^ n12292 ;
  assign n49538 = n47550 | n49537 ;
  assign n49539 = ( n8480 & n20679 ) | ( n8480 & n26073 ) | ( n20679 & n26073 ) ;
  assign n49540 = n19708 & n20053 ;
  assign n49541 = n49540 ^ n13503 ^ 1'b0 ;
  assign n49543 = n12103 ^ n4992 ^ 1'b0 ;
  assign n49542 = n4626 & ~n33476 ;
  assign n49544 = n49543 ^ n49542 ^ 1'b0 ;
  assign n49545 = ~n2655 & n19765 ;
  assign n49546 = ~n10705 & n49545 ;
  assign n49547 = n49546 ^ n20678 ^ 1'b0 ;
  assign n49548 = n9958 & n13099 ;
  assign n49549 = n49548 ^ n32850 ^ 1'b0 ;
  assign n49550 = n9620 ^ n1997 ^ 1'b0 ;
  assign n49551 = n2671 & ~n27755 ;
  assign n49552 = n49551 ^ n11330 ^ 1'b0 ;
  assign n49553 = n172 & n40473 ;
  assign n49554 = n44606 ^ n13289 ^ 1'b0 ;
  assign n49555 = n49554 ^ n43562 ^ n36729 ;
  assign n49556 = ~n13472 & n22135 ;
  assign n49557 = ~n7532 & n21957 ;
  assign n49558 = ( n405 & n436 ) | ( n405 & ~n12671 ) | ( n436 & ~n12671 ) ;
  assign n49559 = ~n19265 & n49558 ;
  assign n49560 = n20993 & n49559 ;
  assign n49561 = n5662 & n20560 ;
  assign n49562 = ~n27592 & n49561 ;
  assign n49563 = n38435 ^ n28955 ^ 1'b0 ;
  assign n49564 = n29746 & ~n49563 ;
  assign n49565 = n49564 ^ n4378 ^ 1'b0 ;
  assign n49566 = n18213 ^ n12146 ^ n2769 ;
  assign n49567 = n48501 ^ n32129 ^ 1'b0 ;
  assign n49568 = n26831 ^ n14037 ^ 1'b0 ;
  assign n49569 = n11560 | n49568 ;
  assign n49570 = n15800 & n32382 ;
  assign n49571 = n2408 | n48826 ;
  assign n49572 = n19991 ^ n19271 ^ n12439 ;
  assign n49573 = ( n700 & ~n22177 ) | ( n700 & n49572 ) | ( ~n22177 & n49572 ) ;
  assign n49574 = n49573 ^ n6531 ^ 1'b0 ;
  assign n49575 = n1400 & n9226 ;
  assign n49576 = n169 & n534 ;
  assign n49577 = ~n534 & n49576 ;
  assign n49578 = n257 | n2302 ;
  assign n49579 = n49577 & ~n49578 ;
  assign n49580 = n49579 ^ n442 ^ 1'b0 ;
  assign n49581 = n8721 & ~n49580 ;
  assign n49582 = n16010 & n49581 ;
  assign n49583 = n6309 | n19698 ;
  assign n49584 = n49582 & ~n49583 ;
  assign n49585 = n44061 ^ n23610 ^ 1'b0 ;
  assign n49586 = n424 & n49585 ;
  assign n49587 = n28740 ^ n9286 ^ 1'b0 ;
  assign n49588 = ~n20714 & n49587 ;
  assign n49593 = n3723 ^ n1691 ^ 1'b0 ;
  assign n49594 = n10512 | n49593 ;
  assign n49595 = n14244 & ~n49594 ;
  assign n49589 = n12454 ^ n11811 ^ 1'b0 ;
  assign n49590 = ~n48 & n33401 ;
  assign n49591 = n49590 ^ n29731 ^ 1'b0 ;
  assign n49592 = n49589 & ~n49591 ;
  assign n49596 = n49595 ^ n49592 ^ 1'b0 ;
  assign n49597 = n47729 ^ n9995 ^ 1'b0 ;
  assign n49598 = n26464 ^ n4972 ^ 1'b0 ;
  assign n49599 = ~n49597 & n49598 ;
  assign n49600 = n49599 ^ n34320 ^ 1'b0 ;
  assign n49601 = n6316 | n37147 ;
  assign n49602 = n49601 ^ n36753 ^ 1'b0 ;
  assign n49603 = n43304 ^ n16663 ^ 1'b0 ;
  assign n49604 = n49602 | n49603 ;
  assign n49605 = n29587 ^ n25922 ^ 1'b0 ;
  assign n49606 = n17938 ^ n191 ^ 1'b0 ;
  assign n49607 = n7831 & n23411 ;
  assign n49608 = n49606 & n49607 ;
  assign n49609 = n3713 & ~n49608 ;
  assign n49612 = n3286 | n33743 ;
  assign n49613 = n767 | n49612 ;
  assign n49610 = n9284 | n38821 ;
  assign n49611 = n16887 & ~n49610 ;
  assign n49614 = n49613 ^ n49611 ^ 1'b0 ;
  assign n49615 = n13109 ^ n10679 ^ 1'b0 ;
  assign n49616 = n6157 ^ n2821 ^ 1'b0 ;
  assign n49617 = n4281 & ~n11824 ;
  assign n49618 = ~n49616 & n49617 ;
  assign n49619 = ~n6501 & n11247 ;
  assign n49620 = ( n976 & n42813 ) | ( n976 & ~n49619 ) | ( n42813 & ~n49619 ) ;
  assign n49621 = n49618 & n49620 ;
  assign n49622 = ~n4138 & n27057 ;
  assign n49623 = n11350 ^ n10295 ^ n4296 ;
  assign n49624 = n42777 ^ n3592 ^ 1'b0 ;
  assign n49625 = n9796 & ~n30326 ;
  assign n49628 = n23440 ^ n4276 ^ n576 ;
  assign n49626 = n39470 ^ n34317 ^ 1'b0 ;
  assign n49627 = n25949 & n49626 ;
  assign n49629 = n49628 ^ n49627 ^ n7320 ;
  assign n49630 = n49629 ^ n12754 ^ 1'b0 ;
  assign n49631 = n12317 ^ n9457 ^ 1'b0 ;
  assign n49632 = n16557 ^ n4803 ^ 1'b0 ;
  assign n49633 = ~n33172 & n49632 ;
  assign n49634 = ( n31732 & ~n41613 ) | ( n31732 & n49633 ) | ( ~n41613 & n49633 ) ;
  assign n49635 = n12947 ^ n3217 ^ 1'b0 ;
  assign n49636 = n49635 ^ n13627 ^ 1'b0 ;
  assign n49637 = n32492 ^ n3245 ^ 1'b0 ;
  assign n49638 = n48788 | n49637 ;
  assign n49639 = ( ~n91 & n6933 ) | ( ~n91 & n49638 ) | ( n6933 & n49638 ) ;
  assign n49640 = n17876 & ~n36547 ;
  assign n49641 = n49640 ^ n9852 ^ 1'b0 ;
  assign n49642 = ~n1435 & n17629 ;
  assign n49643 = n49642 ^ n3346 ^ 1'b0 ;
  assign n49644 = n34151 & n49643 ;
  assign n49645 = n28495 ^ n24968 ^ n102 ;
  assign n49646 = n42233 & ~n49645 ;
  assign n49647 = n9941 & n23956 ;
  assign n49648 = n49647 ^ n31619 ^ 1'b0 ;
  assign n49649 = n38445 ^ n22866 ^ 1'b0 ;
  assign n49650 = n33976 ^ n28886 ^ 1'b0 ;
  assign n49651 = n30876 & n49650 ;
  assign n49652 = n49651 ^ n19465 ^ 1'b0 ;
  assign n49653 = n22224 ^ n8267 ^ 1'b0 ;
  assign n49654 = ~n3574 & n49653 ;
  assign n49655 = ( n8750 & n28087 ) | ( n8750 & n49654 ) | ( n28087 & n49654 ) ;
  assign n49656 = n21895 ^ n11447 ^ n3056 ;
  assign n49657 = n49655 & n49656 ;
  assign n49658 = ( n10895 & n32070 ) | ( n10895 & ~n49657 ) | ( n32070 & ~n49657 ) ;
  assign n49659 = ~n12459 & n12630 ;
  assign n49660 = n2538 & n49659 ;
  assign n49661 = ( n9120 & n12951 ) | ( n9120 & n49660 ) | ( n12951 & n49660 ) ;
  assign n49662 = ( n4231 & n47396 ) | ( n4231 & ~n49661 ) | ( n47396 & ~n49661 ) ;
  assign n49663 = n10533 ^ n10339 ^ 1'b0 ;
  assign n49664 = ~n10679 & n49663 ;
  assign n49665 = n3256 & ~n23665 ;
  assign n49666 = ~n49664 & n49665 ;
  assign n49667 = n2502 | n37674 ;
  assign n49668 = n49667 ^ n11768 ^ 1'b0 ;
  assign n49669 = n8170 & ~n49668 ;
  assign n49673 = n15897 & ~n35165 ;
  assign n49670 = n3120 & ~n37285 ;
  assign n49671 = n49670 ^ n16527 ^ 1'b0 ;
  assign n49672 = n1418 & n49671 ;
  assign n49674 = n49673 ^ n49672 ^ 1'b0 ;
  assign n49675 = n46271 ^ n7144 ^ 1'b0 ;
  assign n49676 = n14026 ^ n2787 ^ 1'b0 ;
  assign n49677 = ~n40987 & n49676 ;
  assign n49678 = ~n20274 & n49677 ;
  assign n49679 = n2300 & ~n2588 ;
  assign n49680 = n49679 ^ n19002 ^ 1'b0 ;
  assign n49681 = n5285 ^ n2868 ^ 1'b0 ;
  assign n49682 = n49681 ^ n20815 ^ n3650 ;
  assign n49683 = n24222 ^ n1933 ^ 1'b0 ;
  assign n49684 = ~n6156 & n6758 ;
  assign n49686 = n15683 ^ n15412 ^ n11958 ;
  assign n49687 = ( ~n6791 & n10594 ) | ( ~n6791 & n49686 ) | ( n10594 & n49686 ) ;
  assign n49685 = ~n16810 & n23449 ;
  assign n49688 = n49687 ^ n49685 ^ 1'b0 ;
  assign n49689 = ~n19551 & n33994 ;
  assign n49690 = n49689 ^ n7633 ^ 1'b0 ;
  assign n49691 = n1138 & ~n34000 ;
  assign n49692 = n27516 ^ n19377 ^ 1'b0 ;
  assign n49693 = ( n16666 & n22103 ) | ( n16666 & n49692 ) | ( n22103 & n49692 ) ;
  assign n49694 = ~n3581 & n10484 ;
  assign n49695 = n49694 ^ n8838 ^ 1'b0 ;
  assign n49696 = n16301 ^ n222 ^ 1'b0 ;
  assign n49697 = n6254 & ~n13395 ;
  assign n49698 = ( ~n49695 & n49696 ) | ( ~n49695 & n49697 ) | ( n49696 & n49697 ) ;
  assign n49699 = n13253 & ~n19298 ;
  assign n49700 = n49699 ^ n181 ^ 1'b0 ;
  assign n49701 = n31874 ^ n20026 ^ 1'b0 ;
  assign n49702 = ~n45622 & n49701 ;
  assign n49703 = n8941 & n13609 ;
  assign n49704 = ~n12591 & n49703 ;
  assign n49705 = n10952 | n30483 ;
  assign n49706 = n49705 ^ n23134 ^ n10105 ;
  assign n49707 = n14690 ^ n8421 ^ 1'b0 ;
  assign n49708 = n9105 & n49707 ;
  assign n49709 = n1010 & n49708 ;
  assign n49710 = n49709 ^ n34414 ^ 1'b0 ;
  assign n49711 = n9789 | n49710 ;
  assign n49712 = n49711 ^ n7129 ^ 1'b0 ;
  assign n49713 = n31603 ^ n28966 ^ 1'b0 ;
  assign n49714 = ~n11971 & n42852 ;
  assign n49715 = ~n22988 & n32372 ;
  assign n49716 = n17401 ^ n7728 ^ 1'b0 ;
  assign n49717 = ( ~n15005 & n49715 ) | ( ~n15005 & n49716 ) | ( n49715 & n49716 ) ;
  assign n49718 = n179 | n15356 ;
  assign n49719 = n179 & ~n49718 ;
  assign n49720 = ~n1820 & n8619 ;
  assign n49721 = ~n8619 & n49720 ;
  assign n49722 = n49719 | n49721 ;
  assign n49723 = n49717 | n49722 ;
  assign n49724 = n46827 ^ n42540 ^ 1'b0 ;
  assign n49725 = n27572 | n49724 ;
  assign n49726 = n3288 & n15336 ;
  assign n49727 = n49725 & n49726 ;
  assign n49728 = n3149 | n38118 ;
  assign n49729 = n49727 & ~n49728 ;
  assign n49730 = ~n3574 & n20433 ;
  assign n49731 = n49730 ^ n1009 ^ 1'b0 ;
  assign n49732 = n4394 ^ n1585 ^ 1'b0 ;
  assign n49733 = n49731 & ~n49732 ;
  assign n49734 = n126 | n26940 ;
  assign n49735 = ~n17763 & n19402 ;
  assign n49736 = n43778 & n49735 ;
  assign n49737 = ( n13250 & n49734 ) | ( n13250 & n49736 ) | ( n49734 & n49736 ) ;
  assign n49738 = n7713 & ~n49737 ;
  assign n49739 = ~n940 & n49738 ;
  assign n49740 = n37388 ^ n4715 ^ 1'b0 ;
  assign n49741 = n9711 & n49740 ;
  assign n49742 = ( n12088 & n12932 ) | ( n12088 & n18611 ) | ( n12932 & n18611 ) ;
  assign n49743 = ( n10284 & ~n26827 ) | ( n10284 & n49742 ) | ( ~n26827 & n49742 ) ;
  assign n49746 = n16497 & n19105 ;
  assign n49744 = n14208 ^ n11982 ^ 1'b0 ;
  assign n49745 = n7776 & ~n49744 ;
  assign n49747 = n49746 ^ n49745 ^ n5380 ;
  assign n49748 = n49747 ^ n37457 ^ n6180 ;
  assign n49749 = n15960 ^ n4681 ^ 1'b0 ;
  assign n49750 = n17053 & ~n49749 ;
  assign n49751 = n49750 ^ n43153 ^ n3018 ;
  assign n49752 = n10218 & n49751 ;
  assign n49753 = n7404 & n22205 ;
  assign n49754 = ( n12619 & n39087 ) | ( n12619 & ~n49753 ) | ( n39087 & ~n49753 ) ;
  assign n49755 = n2004 & n25472 ;
  assign n49756 = n49755 ^ n12387 ^ 1'b0 ;
  assign n49757 = n7454 & n9469 ;
  assign n49758 = ( n1628 & n6343 ) | ( n1628 & ~n6521 ) | ( n6343 & ~n6521 ) ;
  assign n49759 = n48999 ^ n15497 ^ 1'b0 ;
  assign n49760 = n49758 & ~n49759 ;
  assign n49761 = n49760 ^ n45302 ^ 1'b0 ;
  assign n49762 = ~n62 & n7404 ;
  assign n49763 = n49762 ^ n26426 ^ 1'b0 ;
  assign n49764 = n10457 | n16802 ;
  assign n49765 = n13719 | n49764 ;
  assign n49766 = n7400 & n49765 ;
  assign n49767 = n16424 ^ n10703 ^ n446 ;
  assign n49768 = ~n12186 & n49767 ;
  assign n49769 = n18683 | n49768 ;
  assign n49770 = n49769 ^ n16462 ^ 1'b0 ;
  assign n49771 = n14943 ^ n4531 ^ 1'b0 ;
  assign n49772 = ~n15564 & n49771 ;
  assign n49773 = n49772 ^ n1412 ^ 1'b0 ;
  assign n49774 = ~n14878 & n30339 ;
  assign n49775 = n32052 & n49774 ;
  assign n49776 = n3574 | n29054 ;
  assign n49777 = n3660 | n49776 ;
  assign n49778 = n34085 & n49777 ;
  assign n49779 = n49778 ^ n23831 ^ 1'b0 ;
  assign n49780 = n49775 | n49779 ;
  assign n49781 = ~n1167 & n21837 ;
  assign n49782 = n37030 & n43621 ;
  assign n49783 = n2904 & ~n18594 ;
  assign n49784 = n49783 ^ n279 ^ 1'b0 ;
  assign n49785 = ~n9928 & n49784 ;
  assign n49786 = n33381 ^ n13408 ^ 1'b0 ;
  assign n49787 = n38828 ^ n18969 ^ 1'b0 ;
  assign n49788 = n49271 ^ n29437 ^ 1'b0 ;
  assign n49789 = n21958 | n22612 ;
  assign n49790 = n35817 | n49789 ;
  assign n49791 = n49790 ^ n23603 ^ 1'b0 ;
  assign n49792 = n49791 ^ n250 ^ 1'b0 ;
  assign n49793 = n17062 | n49792 ;
  assign n49794 = n3906 & n46796 ;
  assign n49795 = n32873 & n49794 ;
  assign n49796 = n33503 ^ n28691 ^ 1'b0 ;
  assign n49797 = n46400 ^ n33115 ^ n6564 ;
  assign n49798 = n6888 & n43053 ;
  assign n49799 = ~n18539 & n49798 ;
  assign n49800 = ~n49797 & n49799 ;
  assign n49801 = n23856 | n47348 ;
  assign n49802 = n13815 & n24749 ;
  assign n49803 = n18174 & n37507 ;
  assign n49804 = n28764 ^ n1661 ^ 1'b0 ;
  assign n49805 = ~n11266 & n49804 ;
  assign n49806 = n3652 | n26845 ;
  assign n49809 = n194 & ~n15373 ;
  assign n49810 = n49809 ^ n21667 ^ 1'b0 ;
  assign n49807 = n2696 | n28414 ;
  assign n49808 = n8380 | n49807 ;
  assign n49811 = n49810 ^ n49808 ^ 1'b0 ;
  assign n49812 = ~n16232 & n29852 ;
  assign n49813 = ~n5322 & n49812 ;
  assign n49814 = n5769 & n49813 ;
  assign n49815 = n39299 ^ n16117 ^ 1'b0 ;
  assign n49816 = n46209 & ~n49815 ;
  assign n49817 = ( n10537 & ~n16101 ) | ( n10537 & n42448 ) | ( ~n16101 & n42448 ) ;
  assign n49818 = ( n24744 & n26628 ) | ( n24744 & ~n45316 ) | ( n26628 & ~n45316 ) ;
  assign n49819 = n49818 ^ n17339 ^ n3581 ;
  assign n49820 = ( n9411 & n23810 ) | ( n9411 & n39598 ) | ( n23810 & n39598 ) ;
  assign n49821 = ~n23524 & n49820 ;
  assign n49822 = ( n9246 & n23970 ) | ( n9246 & ~n29720 ) | ( n23970 & ~n29720 ) ;
  assign n49823 = ~n38660 & n49822 ;
  assign n49824 = n35747 & n49823 ;
  assign n49825 = n49824 ^ n42461 ^ 1'b0 ;
  assign n49826 = n34754 ^ n15554 ^ 1'b0 ;
  assign n49827 = ~n9519 & n49826 ;
  assign n49828 = n4954 ^ n1507 ^ 1'b0 ;
  assign n49829 = ~n4165 & n49828 ;
  assign n49830 = n9667 ^ n5172 ^ 1'b0 ;
  assign n49831 = n8355 | n49830 ;
  assign n49832 = n49831 ^ n12183 ^ 1'b0 ;
  assign n49833 = n49829 & ~n49832 ;
  assign n49834 = n43828 ^ n16939 ^ 1'b0 ;
  assign n49835 = n49811 | n49834 ;
  assign n49841 = n524 & ~n19113 ;
  assign n49842 = ~n524 & n49841 ;
  assign n49843 = n342 | n3198 ;
  assign n49844 = n49842 & ~n49843 ;
  assign n49845 = n490 & ~n49844 ;
  assign n49846 = n49844 & n49845 ;
  assign n49839 = n1290 & ~n12075 ;
  assign n49840 = ~n1290 & n49839 ;
  assign n49836 = n5660 & ~n29105 ;
  assign n49837 = n29105 & n49836 ;
  assign n49838 = n49837 ^ n38317 ^ 1'b0 ;
  assign n49847 = n49846 ^ n49840 ^ n49838 ;
  assign n49848 = ( n15562 & ~n19770 ) | ( n15562 & n49847 ) | ( ~n19770 & n49847 ) ;
  assign n49849 = n887 & n31663 ;
  assign n49850 = n49849 ^ n1490 ^ 1'b0 ;
  assign n49851 = n174 & ~n29227 ;
  assign n49852 = n49850 & n49851 ;
  assign n49853 = n9498 & ~n31928 ;
  assign n49854 = n17966 & ~n37738 ;
  assign n49855 = n49854 ^ n12892 ^ 1'b0 ;
  assign n49856 = n49855 ^ n34509 ^ n27387 ;
  assign n49860 = n33580 ^ n16132 ^ 1'b0 ;
  assign n49857 = ~n11077 & n12202 ;
  assign n49858 = n16546 | n49857 ;
  assign n49859 = n57 | n49858 ;
  assign n49861 = n49860 ^ n49859 ^ n1602 ;
  assign n49862 = n38514 ^ n1642 ^ 1'b0 ;
  assign n49863 = n27107 & ~n49862 ;
  assign n49864 = n24032 & n38827 ;
  assign n49866 = ~n12049 & n20543 ;
  assign n49867 = n49866 ^ n4084 ^ 1'b0 ;
  assign n49865 = n15912 & ~n25594 ;
  assign n49868 = n49867 ^ n49865 ^ 1'b0 ;
  assign n49869 = n457 | n46244 ;
  assign n49870 = n30377 ^ n24865 ^ n3784 ;
  assign n49871 = ~n31795 & n45685 ;
  assign n49872 = n2550 & n32506 ;
  assign n49873 = n47996 ^ n38009 ^ 1'b0 ;
  assign n49874 = n2431 & n49873 ;
  assign n49875 = n12323 | n39943 ;
  assign n49876 = n15367 & ~n27902 ;
  assign n49877 = ~n12750 & n49876 ;
  assign n49878 = n49877 ^ n4647 ^ 1'b0 ;
  assign n49879 = n14890 | n31348 ;
  assign n49880 = n49879 ^ n21163 ^ 1'b0 ;
  assign n49881 = n34582 | n49880 ;
  assign n49883 = n28485 ^ n9273 ^ n4957 ;
  assign n49884 = n15097 | n49883 ;
  assign n49885 = n49884 ^ n37170 ^ n27429 ;
  assign n49882 = n12856 & n22658 ;
  assign n49886 = n49885 ^ n49882 ^ 1'b0 ;
  assign n49887 = n41437 ^ n41077 ^ 1'b0 ;
  assign n49888 = ~n15328 & n49887 ;
  assign n49889 = ~n21419 & n27138 ;
  assign n49890 = n49889 ^ n2382 ^ 1'b0 ;
  assign n49891 = ( n4077 & n18919 ) | ( n4077 & ~n41455 ) | ( n18919 & ~n41455 ) ;
  assign n49892 = n24755 ^ n2858 ^ 1'b0 ;
  assign n49893 = n14172 & ~n49892 ;
  assign n49894 = n27029 ^ n17720 ^ 1'b0 ;
  assign n49895 = ( n26845 & n49893 ) | ( n26845 & n49894 ) | ( n49893 & n49894 ) ;
  assign n49896 = n30422 | n40575 ;
  assign n49897 = n49896 ^ n37911 ^ 1'b0 ;
  assign n49898 = n49897 ^ n14278 ^ 1'b0 ;
  assign n49899 = n9621 & n49898 ;
  assign n49900 = n49899 ^ n38312 ^ 1'b0 ;
  assign n49901 = n25120 ^ n771 ^ 1'b0 ;
  assign n49902 = n10827 ^ n10040 ^ 1'b0 ;
  assign n49903 = n39947 ^ n31532 ^ 1'b0 ;
  assign n49906 = ~n5113 & n26226 ;
  assign n49907 = n49906 ^ n17996 ^ 1'b0 ;
  assign n49904 = n20316 ^ n3151 ^ 1'b0 ;
  assign n49905 = n8962 & n49904 ;
  assign n49908 = n49907 ^ n49905 ^ n2946 ;
  assign n49909 = n16005 ^ n12901 ^ n8451 ;
  assign n49910 = n11205 | n27041 ;
  assign n49911 = n1350 & ~n12090 ;
  assign n49912 = n36166 ^ n18132 ^ 1'b0 ;
  assign n49913 = n49911 & n49912 ;
  assign n49914 = n3837 & n7558 ;
  assign n49915 = n43305 ^ n4986 ^ 1'b0 ;
  assign n49916 = ~n44756 & n49915 ;
  assign n49917 = n44257 ^ n19404 ^ 1'b0 ;
  assign n49918 = n11519 | n17873 ;
  assign n49919 = n49918 ^ n42709 ^ 1'b0 ;
  assign n49920 = ( ~n19755 & n49917 ) | ( ~n19755 & n49919 ) | ( n49917 & n49919 ) ;
  assign n49921 = ~n14831 & n36622 ;
  assign n49922 = n9377 & n49921 ;
  assign n49923 = n49922 ^ n23786 ^ 1'b0 ;
  assign n49924 = n11628 | n15600 ;
  assign n49925 = ( n16602 & n38770 ) | ( n16602 & n49924 ) | ( n38770 & n49924 ) ;
  assign n49926 = n27840 ^ n26169 ^ n18193 ;
  assign n49927 = n38012 | n49926 ;
  assign n49928 = n49927 ^ n16419 ^ 1'b0 ;
  assign n49929 = ~n35724 & n49928 ;
  assign n49930 = n17078 & n48175 ;
  assign n49931 = n49930 ^ n47190 ^ 1'b0 ;
  assign n49932 = n10598 ^ n115 ^ 1'b0 ;
  assign n49933 = ~n3092 & n49932 ;
  assign n49934 = ~n38317 & n43258 ;
  assign n49935 = ~n49933 & n49934 ;
  assign n49936 = n3294 ^ n2596 ^ 1'b0 ;
  assign n49937 = n49936 ^ n7183 ^ 1'b0 ;
  assign n49938 = n22942 | n49937 ;
  assign n49939 = n28161 ^ n10342 ^ 1'b0 ;
  assign n49940 = ~n49938 & n49939 ;
  assign n49941 = n7260 & n24117 ;
  assign n49942 = ~n5372 & n49941 ;
  assign n49943 = ( ~n3936 & n8640 ) | ( ~n3936 & n49942 ) | ( n8640 & n49942 ) ;
  assign n49944 = n16284 & ~n38115 ;
  assign n49945 = n9770 & ~n45530 ;
  assign n49946 = n33472 & n36965 ;
  assign n49947 = n38835 ^ n18541 ^ 1'b0 ;
  assign n49950 = n4208 & n28101 ;
  assign n49951 = n49950 ^ n12696 ^ 1'b0 ;
  assign n49948 = n44036 ^ n43412 ^ n2339 ;
  assign n49949 = n49948 ^ n31118 ^ 1'b0 ;
  assign n49952 = n49951 ^ n49949 ^ n33489 ;
  assign n49953 = n34903 ^ n16187 ^ 1'b0 ;
  assign n49954 = n12969 | n31276 ;
  assign n49955 = n7291 & ~n49954 ;
  assign n49956 = n49955 ^ n36178 ^ n9352 ;
  assign n49957 = n23393 ^ n19090 ^ 1'b0 ;
  assign n49958 = n30898 ^ n7523 ^ n1088 ;
  assign n49959 = n49958 ^ n12898 ^ 1'b0 ;
  assign n49960 = ~n17128 & n49959 ;
  assign n49961 = n24288 ^ n23456 ^ 1'b0 ;
  assign n49962 = ~n6533 & n49961 ;
  assign n49963 = n12554 | n32880 ;
  assign n49964 = n26501 & ~n49963 ;
  assign n49965 = n37398 | n49964 ;
  assign n49966 = n36009 ^ n18103 ^ 1'b0 ;
  assign n49967 = n20210 & ~n42887 ;
  assign n49968 = n49967 ^ n9765 ^ 1'b0 ;
  assign n49969 = n19894 ^ n14760 ^ 1'b0 ;
  assign n49970 = ~n10456 & n24101 ;
  assign n49971 = n49970 ^ n16369 ^ 1'b0 ;
  assign n49972 = n39202 ^ n7417 ^ 1'b0 ;
  assign n49973 = n14534 | n49972 ;
  assign n49974 = n40212 ^ n30961 ^ 1'b0 ;
  assign n49975 = n1815 | n12143 ;
  assign n49976 = ~n3040 & n35079 ;
  assign n49977 = n8920 & ~n30733 ;
  assign n49978 = ~n9452 & n49977 ;
  assign n49979 = n40399 ^ n6204 ^ 1'b0 ;
  assign n49980 = ~n49978 & n49979 ;
  assign n49981 = n23354 ^ n12573 ^ 1'b0 ;
  assign n49982 = n14791 & ~n41931 ;
  assign n49983 = n49982 ^ n29694 ^ 1'b0 ;
  assign n49984 = n49981 & ~n49983 ;
  assign n49985 = n2449 | n38967 ;
  assign n49986 = ~n49984 & n49985 ;
  assign n49987 = n12454 ^ n7275 ^ 1'b0 ;
  assign n49988 = n2652 & n49987 ;
  assign n49989 = ~n22255 & n49988 ;
  assign n49990 = n49989 ^ n16405 ^ 1'b0 ;
  assign n49991 = n33578 & ~n49990 ;
  assign n49992 = n4060 | n40210 ;
  assign n49993 = n15794 ^ n8001 ^ 1'b0 ;
  assign n49994 = ~n1103 & n49993 ;
  assign n49995 = ~n23833 & n49994 ;
  assign n49996 = n398 & n49995 ;
  assign n49997 = ( n11949 & ~n16403 ) | ( n11949 & n49996 ) | ( ~n16403 & n49996 ) ;
  assign n49998 = n4412 | n7460 ;
  assign n49999 = n49998 ^ n47808 ^ n12763 ;
  assign n50000 = n34506 ^ n342 ^ 1'b0 ;
  assign n50001 = n26715 & n32758 ;
  assign n50002 = n46280 & n50001 ;
  assign n50003 = n11931 & n29903 ;
  assign n50004 = n44401 & n50003 ;
  assign n50005 = n26683 | n29534 ;
  assign n50008 = n14497 | n19212 ;
  assign n50006 = n17558 ^ n13903 ^ 1'b0 ;
  assign n50007 = n19565 | n50006 ;
  assign n50009 = n50008 ^ n50007 ^ 1'b0 ;
  assign n50010 = n4981 & ~n50009 ;
  assign n50011 = n50010 ^ n42441 ^ 1'b0 ;
  assign n50012 = n20061 ^ n2073 ^ 1'b0 ;
  assign n50013 = ~n6528 & n25625 ;
  assign n50014 = n7756 | n25251 ;
  assign n50015 = n45923 ^ n21652 ^ 1'b0 ;
  assign n50016 = n48708 ^ n13122 ^ 1'b0 ;
  assign n50017 = n14047 & ~n31362 ;
  assign n50018 = n18000 | n44616 ;
  assign n50019 = n50018 ^ n12945 ^ 1'b0 ;
  assign n50020 = n29604 ^ n23211 ^ 1'b0 ;
  assign n50021 = n37385 & ~n41516 ;
  assign n50022 = n3812 & n50021 ;
  assign n50023 = n30742 ^ n21212 ^ n5908 ;
  assign n50026 = ( n10893 & n18107 ) | ( n10893 & n36824 ) | ( n18107 & n36824 ) ;
  assign n50024 = n676 ^ n547 ^ 1'b0 ;
  assign n50025 = ~n19483 & n50024 ;
  assign n50027 = n50026 ^ n50025 ^ 1'b0 ;
  assign n50028 = n50027 ^ n39699 ^ 1'b0 ;
  assign n50029 = n45408 ^ n29117 ^ 1'b0 ;
  assign n50030 = n25164 & n25702 ;
  assign n50031 = n42264 ^ n6616 ^ n3127 ;
  assign n50032 = ~n923 & n9474 ;
  assign n50033 = n48063 | n50032 ;
  assign n50034 = n50033 ^ n40415 ^ n13113 ;
  assign n50035 = n28472 ^ n8472 ^ 1'b0 ;
  assign n50036 = n24092 & n50035 ;
  assign n50037 = n32581 ^ n7328 ^ 1'b0 ;
  assign n50038 = n3795 & n14475 ;
  assign n50039 = n50038 ^ n15246 ^ 1'b0 ;
  assign n50043 = n10829 | n19038 ;
  assign n50040 = n289 & ~n11207 ;
  assign n50041 = n50040 ^ n28259 ^ 1'b0 ;
  assign n50042 = ~n29363 & n50041 ;
  assign n50044 = n50043 ^ n50042 ^ 1'b0 ;
  assign n50045 = ~n33099 & n50044 ;
  assign n50046 = n50045 ^ n18641 ^ 1'b0 ;
  assign n50047 = n17053 & n40708 ;
  assign n50048 = ~n18024 & n50047 ;
  assign n50049 = ( n4520 & n6343 ) | ( n4520 & ~n11440 ) | ( n6343 & ~n11440 ) ;
  assign n50050 = n50049 ^ n2203 ^ 1'b0 ;
  assign n50051 = ( n2245 & ~n2583 ) | ( n2245 & n35552 ) | ( ~n2583 & n35552 ) ;
  assign n50052 = n395 & n42308 ;
  assign n50053 = n20486 ^ n18409 ^ n1525 ;
  assign n50054 = n14218 & ~n50053 ;
  assign n50055 = n21366 ^ n18879 ^ n7760 ;
  assign n50056 = n22874 ^ n9105 ^ n1832 ;
  assign n50057 = n46326 ^ n9021 ^ 1'b0 ;
  assign n50058 = n9045 & n21654 ;
  assign n50059 = n30460 ^ n11143 ^ n10335 ;
  assign n50060 = n50059 ^ n9439 ^ 1'b0 ;
  assign n50061 = ~n33436 & n37404 ;
  assign n50062 = n50060 & n50061 ;
  assign n50063 = n3087 | n36477 ;
  assign n50064 = n603 & ~n33520 ;
  assign n50065 = n39059 ^ n22576 ^ 1'b0 ;
  assign n50066 = n43919 & ~n50065 ;
  assign n50067 = n10291 & ~n50066 ;
  assign n50068 = n23047 ^ n21495 ^ n18754 ;
  assign n50069 = n26800 & n50068 ;
  assign n50070 = n50069 ^ n32327 ^ 1'b0 ;
  assign n50071 = n50070 ^ n35129 ^ n24998 ;
  assign n50072 = ~n7493 & n21259 ;
  assign n50073 = n22139 ^ n790 ^ 1'b0 ;
  assign n50074 = n19000 & ~n50073 ;
  assign n50075 = n20186 & n30523 ;
  assign n50076 = n13183 & n50075 ;
  assign n50077 = n43287 & ~n46154 ;
  assign n50078 = n50077 ^ n6866 ^ 1'b0 ;
  assign n50079 = n40867 | n50078 ;
  assign n50080 = n3354 & n50079 ;
  assign n50081 = n44912 & n50080 ;
  assign n50082 = n39145 ^ n544 ^ 1'b0 ;
  assign n50083 = n32527 & ~n50082 ;
  assign n50084 = n17754 ^ n11670 ^ n162 ;
  assign n50085 = n37267 ^ n28378 ^ n22677 ;
  assign n50086 = ~n2706 & n33743 ;
  assign n50087 = n29298 & ~n39234 ;
  assign n50088 = n50087 ^ n13242 ^ 1'b0 ;
  assign n50089 = ~n17489 & n50088 ;
  assign n50090 = n8369 & ~n31148 ;
  assign n50091 = n12553 & ~n50090 ;
  assign n50092 = n38199 ^ n5131 ^ 1'b0 ;
  assign n50093 = n1506 & n19034 ;
  assign n50094 = n50093 ^ n18935 ^ 1'b0 ;
  assign n50095 = n19465 | n50094 ;
  assign n50096 = n14298 & ~n16513 ;
  assign n50097 = n50096 ^ n20534 ^ 1'b0 ;
  assign n50098 = n50097 ^ n25108 ^ 1'b0 ;
  assign n50099 = ~n102 & n23958 ;
  assign n50100 = n50099 ^ n44208 ^ n3866 ;
  assign n50101 = n8061 | n50100 ;
  assign n50102 = n50101 ^ n31944 ^ 1'b0 ;
  assign n50103 = n15029 & ~n49196 ;
  assign n50105 = n18877 ^ n2946 ^ 1'b0 ;
  assign n50106 = n19407 & n50105 ;
  assign n50104 = ~n7106 & n14821 ;
  assign n50107 = n50106 ^ n50104 ^ 1'b0 ;
  assign n50108 = n44207 ^ n23128 ^ 1'b0 ;
  assign n50109 = n22437 ^ n17383 ^ 1'b0 ;
  assign n50110 = ~n41550 & n50109 ;
  assign n50111 = ( ~n5656 & n26382 ) | ( ~n5656 & n30191 ) | ( n26382 & n30191 ) ;
  assign n50112 = ( n10481 & n18600 ) | ( n10481 & ~n30610 ) | ( n18600 & ~n30610 ) ;
  assign n50115 = n46578 ^ n20666 ^ 1'b0 ;
  assign n50113 = ~n33736 & n46326 ;
  assign n50114 = n2557 & n50113 ;
  assign n50116 = n50115 ^ n50114 ^ 1'b0 ;
  assign n50117 = n38866 ^ n201 ^ 1'b0 ;
  assign n50118 = n9125 & ~n37426 ;
  assign n50119 = n50117 & n50118 ;
  assign n50120 = ~n2933 & n23652 ;
  assign n50121 = n9748 & ~n26636 ;
  assign n50122 = n20517 | n21009 ;
  assign n50123 = n12980 | n34358 ;
  assign n50124 = n8174 & ~n40862 ;
  assign n50125 = ~n12472 & n50124 ;
  assign n50126 = n50125 ^ n5468 ^ 1'b0 ;
  assign n50130 = n1258 & ~n21718 ;
  assign n50131 = n50130 ^ n48167 ^ 1'b0 ;
  assign n50127 = n15936 ^ n1512 ^ 1'b0 ;
  assign n50128 = n50127 ^ n3801 ^ 1'b0 ;
  assign n50129 = ~n42077 & n50128 ;
  assign n50132 = n50131 ^ n50129 ^ 1'b0 ;
  assign n50133 = n12209 ^ n3060 ^ 1'b0 ;
  assign n50134 = n46995 & n50133 ;
  assign n50135 = n10531 & n50134 ;
  assign n50136 = n9528 ^ n2194 ^ 1'b0 ;
  assign n50137 = n45073 ^ n23332 ^ 1'b0 ;
  assign n50138 = n24512 ^ n7363 ^ 1'b0 ;
  assign n50139 = n4173 | n50138 ;
  assign n50140 = n17805 & ~n42927 ;
  assign n50141 = n2552 & n24237 ;
  assign n50142 = n50141 ^ n20705 ^ 1'b0 ;
  assign n50143 = ~n19237 & n50142 ;
  assign n50144 = n24973 & ~n36303 ;
  assign n50145 = n21307 | n42265 ;
  assign n50146 = n42864 ^ n19256 ^ n7795 ;
  assign n50147 = ~n15951 & n19140 ;
  assign n50148 = ~n38343 & n50147 ;
  assign n50149 = ~n12612 & n15386 ;
  assign n50150 = n50149 ^ n16346 ^ 1'b0 ;
  assign n50151 = n28410 ^ n18032 ^ 1'b0 ;
  assign n50152 = n49188 & n50151 ;
  assign n50153 = n50150 & n50152 ;
  assign n50154 = n885 ^ n676 ^ 1'b0 ;
  assign n50155 = n7767 & ~n50154 ;
  assign n50156 = ~n13279 & n50155 ;
  assign n50157 = n22929 & ~n50156 ;
  assign n50158 = ~n26984 & n50157 ;
  assign n50159 = n9217 ^ n7661 ^ n5102 ;
  assign n50160 = n16581 & n50159 ;
  assign n50161 = n18702 & ~n50160 ;
  assign n50162 = n43111 & n50161 ;
  assign n50163 = ~n14234 & n33179 ;
  assign n50164 = n6839 & n46596 ;
  assign n50165 = ~n50163 & n50164 ;
  assign n50166 = n32146 ^ n25966 ^ 1'b0 ;
  assign n50167 = ~n29259 & n50166 ;
  assign n50168 = ~n31667 & n50167 ;
  assign n50169 = n50165 & n50168 ;
  assign n50170 = n33597 & n50169 ;
  assign n50171 = ( ~n4852 & n15923 ) | ( ~n4852 & n18019 ) | ( n15923 & n18019 ) ;
  assign n50172 = n1636 | n3663 ;
  assign n50173 = n50172 ^ n25565 ^ 1'b0 ;
  assign n50174 = n50173 ^ n13958 ^ n13287 ;
  assign n50175 = n35444 ^ n1095 ^ 1'b0 ;
  assign n50176 = n17653 & n50175 ;
  assign n50177 = n38079 & n50176 ;
  assign n50178 = ~n10930 & n43360 ;
  assign n50179 = ~n10960 & n50178 ;
  assign n50180 = n36851 & ~n50179 ;
  assign n50181 = n17617 ^ n11548 ^ 1'b0 ;
  assign n50182 = n22247 | n50181 ;
  assign n50183 = n31635 ^ n10943 ^ 1'b0 ;
  assign n50184 = n18380 | n50183 ;
  assign n50186 = n6603 & ~n17034 ;
  assign n50185 = ~n1581 & n12087 ;
  assign n50187 = n50186 ^ n50185 ^ n6585 ;
  assign n50189 = n27382 ^ n20008 ^ 1'b0 ;
  assign n50188 = ~n2449 & n43740 ;
  assign n50190 = n50189 ^ n50188 ^ 1'b0 ;
  assign n50191 = n46 | n50190 ;
  assign n50192 = n16075 & n47329 ;
  assign n50193 = n34145 & n50192 ;
  assign n50194 = n6243 ^ n3558 ^ 1'b0 ;
  assign n50195 = ~n211 & n50194 ;
  assign n50196 = n16658 & n50195 ;
  assign n50197 = n50196 ^ n19753 ^ 1'b0 ;
  assign n50198 = n34040 ^ n9260 ^ 1'b0 ;
  assign n50199 = n30344 & n50198 ;
  assign n50200 = n26210 & n50199 ;
  assign n50203 = n4126 ^ n3730 ^ n811 ;
  assign n50202 = n1812 & ~n12277 ;
  assign n50204 = n50203 ^ n50202 ^ 1'b0 ;
  assign n50201 = n517 & n12169 ;
  assign n50205 = n50204 ^ n50201 ^ 1'b0 ;
  assign n50206 = ~n18223 & n25479 ;
  assign n50207 = ~n50205 & n50206 ;
  assign n50208 = n49179 ^ n5037 ^ 1'b0 ;
  assign n50209 = n18401 | n50208 ;
  assign n50210 = n36980 & ~n50209 ;
  assign n50211 = ~n21954 & n50210 ;
  assign n50212 = n18498 & ~n32547 ;
  assign n50213 = ~n19087 & n50212 ;
  assign n50214 = n38353 ^ n21859 ^ n1368 ;
  assign n50215 = n122 & ~n24670 ;
  assign n50216 = n50215 ^ n22450 ^ 1'b0 ;
  assign n50217 = n4251 & ~n23592 ;
  assign n50218 = n8816 & n50217 ;
  assign n50219 = n17280 & ~n27660 ;
  assign n50220 = n9217 | n47535 ;
  assign n50221 = n17378 | n50220 ;
  assign n50222 = n43823 ^ n20001 ^ n5466 ;
  assign n50223 = n46355 ^ n11612 ^ 1'b0 ;
  assign n50224 = n45225 | n50223 ;
  assign n50225 = n25468 ^ n19639 ^ n10273 ;
  assign n50226 = ~n50224 & n50225 ;
  assign n50227 = ~n17416 & n38965 ;
  assign n50228 = n17244 ^ n4845 ^ 1'b0 ;
  assign n50229 = n13882 | n50228 ;
  assign n50230 = n20713 ^ n10450 ^ 1'b0 ;
  assign n50231 = ~n15292 & n50230 ;
  assign n50232 = n50231 ^ n49984 ^ 1'b0 ;
  assign n50233 = n10316 & ~n13712 ;
  assign n50234 = n50233 ^ n4136 ^ 1'b0 ;
  assign n50235 = n20183 ^ n10950 ^ 1'b0 ;
  assign n50236 = ~n50234 & n50235 ;
  assign n50237 = n1344 | n11488 ;
  assign n50238 = n50237 ^ n34085 ^ 1'b0 ;
  assign n50239 = n2844 | n2858 ;
  assign n50240 = n711 | n44419 ;
  assign n50241 = n24182 & ~n33247 ;
  assign n50242 = n50241 ^ n46170 ^ 1'b0 ;
  assign n50243 = n1332 | n4228 ;
  assign n50244 = n4263 | n7798 ;
  assign n50245 = n6062 & ~n50244 ;
  assign n50246 = n44863 ^ n18451 ^ 1'b0 ;
  assign n50247 = n40770 & n50246 ;
  assign n50248 = ~n819 & n33072 ;
  assign n50249 = ~n27319 & n50248 ;
  assign n50250 = n3080 & ~n50249 ;
  assign n50251 = n50250 ^ n19698 ^ 1'b0 ;
  assign n50252 = ( n30870 & n41344 ) | ( n30870 & ~n50251 ) | ( n41344 & ~n50251 ) ;
  assign n50253 = ( n13896 & ~n14280 ) | ( n13896 & n30377 ) | ( ~n14280 & n30377 ) ;
  assign n50256 = ~n11796 & n16221 ;
  assign n50257 = n13602 & n50256 ;
  assign n50254 = n49065 ^ n26930 ^ 1'b0 ;
  assign n50255 = n39712 | n50254 ;
  assign n50258 = n50257 ^ n50255 ^ n25526 ;
  assign n50259 = n11620 | n11915 ;
  assign n50260 = n50259 ^ n33298 ^ 1'b0 ;
  assign n50261 = n38614 ^ n37136 ^ 1'b0 ;
  assign n50262 = n28881 & n50261 ;
  assign n50263 = n1169 | n23962 ;
  assign n50264 = n50263 ^ n11741 ^ 1'b0 ;
  assign n50265 = n31928 ^ n17477 ^ n8398 ;
  assign n50266 = n22139 ^ n19893 ^ n13011 ;
  assign n50267 = n4992 & ~n13346 ;
  assign n50268 = n20443 & n50267 ;
  assign n50269 = n48337 ^ n1391 ^ 1'b0 ;
  assign n50270 = ~n50268 & n50269 ;
  assign n50271 = n291 & n50270 ;
  assign n50272 = n50271 ^ n1622 ^ 1'b0 ;
  assign n50273 = n2561 & n17031 ;
  assign n50274 = n14057 & n50273 ;
  assign n50276 = n26317 ^ n6555 ^ 1'b0 ;
  assign n50277 = n8490 & n50276 ;
  assign n50275 = n4925 & n48417 ;
  assign n50278 = n50277 ^ n50275 ^ 1'b0 ;
  assign n50279 = n30338 ^ n24141 ^ 1'b0 ;
  assign n50280 = n18638 & ~n25296 ;
  assign n50281 = ( ~n2447 & n6753 ) | ( ~n2447 & n47582 ) | ( n6753 & n47582 ) ;
  assign n50282 = n50281 ^ n29415 ^ 1'b0 ;
  assign n50283 = n50280 & n50282 ;
  assign n50284 = n29316 | n36548 ;
  assign n50285 = n50284 ^ n9996 ^ 1'b0 ;
  assign n50287 = n14277 ^ n5113 ^ n1345 ;
  assign n50288 = n11082 & ~n50287 ;
  assign n50286 = ~n5057 & n6345 ;
  assign n50289 = n50288 ^ n50286 ^ 1'b0 ;
  assign n50290 = n25981 & n27379 ;
  assign n50291 = ~n12739 & n50290 ;
  assign n50292 = n2541 | n50291 ;
  assign n50293 = n16419 ^ n7227 ^ 1'b0 ;
  assign n50294 = n40795 ^ n33732 ^ n6365 ;
  assign n50295 = n50293 & ~n50294 ;
  assign n50296 = n3140 ^ n2464 ^ n1176 ;
  assign n50297 = ~n2041 & n50296 ;
  assign n50298 = ( n44 & n3119 ) | ( n44 & ~n50297 ) | ( n3119 & ~n50297 ) ;
  assign n50299 = n27729 | n36379 ;
  assign n50300 = n18061 & n25739 ;
  assign n50301 = ~n12554 & n34165 ;
  assign n50302 = n50301 ^ n16776 ^ 1'b0 ;
  assign n50303 = n5592 & n15930 ;
  assign n50304 = ~n32702 & n50303 ;
  assign n50305 = n19060 & ~n43324 ;
  assign n50306 = n98 | n1177 ;
  assign n50307 = n5481 ^ n1001 ^ 1'b0 ;
  assign n50308 = n50307 ^ n44977 ^ n1069 ;
  assign n50309 = n18200 & n23664 ;
  assign n50310 = n4646 | n50309 ;
  assign n50311 = n5312 & ~n50310 ;
  assign n50312 = ~n18490 & n23299 ;
  assign n50313 = n50312 ^ n6217 ^ 1'b0 ;
  assign n50314 = ( n48402 & ~n50311 ) | ( n48402 & n50313 ) | ( ~n50311 & n50313 ) ;
  assign n50315 = n8822 & n23997 ;
  assign n50316 = n30570 | n50315 ;
  assign n50317 = n1201 & n36266 ;
  assign n50318 = n14890 | n28721 ;
  assign n50319 = n42065 & ~n50318 ;
  assign n50321 = n1015 | n26412 ;
  assign n50320 = n24374 ^ n16291 ^ n8427 ;
  assign n50322 = n50321 ^ n50320 ^ 1'b0 ;
  assign n50323 = ( n3057 & n42960 ) | ( n3057 & ~n50322 ) | ( n42960 & ~n50322 ) ;
  assign n50324 = n16546 ^ n14039 ^ 1'b0 ;
  assign n50325 = n50323 & n50324 ;
  assign n50326 = n5692 | n35101 ;
  assign n50327 = n46128 ^ n3076 ^ 1'b0 ;
  assign n50328 = n15190 & ~n50327 ;
  assign n50332 = n23110 ^ n15944 ^ 1'b0 ;
  assign n50330 = n8129 ^ n3953 ^ 1'b0 ;
  assign n50331 = n29650 & ~n50330 ;
  assign n50329 = n20059 ^ n3741 ^ 1'b0 ;
  assign n50333 = n50332 ^ n50331 ^ n50329 ;
  assign n50334 = n10950 & n23126 ;
  assign n50335 = ( n10353 & n24998 ) | ( n10353 & n50334 ) | ( n24998 & n50334 ) ;
  assign n50336 = ~n9789 & n48639 ;
  assign n50337 = n50336 ^ n15350 ^ 1'b0 ;
  assign n50338 = n17042 | n21419 ;
  assign n50339 = n50338 ^ n30831 ^ 1'b0 ;
  assign n50340 = n15407 ^ n14277 ^ 1'b0 ;
  assign n50341 = ~n2750 & n50340 ;
  assign n50342 = ~n9201 & n16278 ;
  assign n50343 = ~n16680 & n43024 ;
  assign n50344 = n23645 & ~n50343 ;
  assign n50345 = n39221 ^ n12162 ^ 1'b0 ;
  assign n50346 = n32198 & ~n50345 ;
  assign n50347 = n50346 ^ n10443 ^ 1'b0 ;
  assign n50348 = n50344 & n50347 ;
  assign n50349 = n50209 & ~n50348 ;
  assign n50350 = n16118 & n50349 ;
  assign n50351 = n13020 & n50350 ;
  assign n50352 = n962 | n50351 ;
  assign n50353 = n7832 & n35847 ;
  assign n50354 = n2687 & n50353 ;
  assign n50355 = ( n16686 & n25218 ) | ( n16686 & n50354 ) | ( n25218 & n50354 ) ;
  assign n50361 = n10250 | n47810 ;
  assign n50362 = n50361 ^ n45559 ^ n39177 ;
  assign n50363 = ~n42431 & n50362 ;
  assign n50360 = n23443 ^ n3993 ^ 1'b0 ;
  assign n50356 = n11508 ^ n9711 ^ 1'b0 ;
  assign n50357 = n14440 & n50356 ;
  assign n50358 = n48964 & n50357 ;
  assign n50359 = n50358 ^ n20815 ^ 1'b0 ;
  assign n50364 = n50363 ^ n50360 ^ n50359 ;
  assign n50365 = n14013 & ~n23156 ;
  assign n50366 = n50365 ^ n4142 ^ 1'b0 ;
  assign n50367 = n10684 & ~n10708 ;
  assign n50368 = n12934 & n50367 ;
  assign n50369 = ( n10001 & n36338 ) | ( n10001 & n50368 ) | ( n36338 & n50368 ) ;
  assign n50370 = n7338 & ~n50369 ;
  assign n50371 = n6369 | n50370 ;
  assign n50372 = n42224 & ~n42495 ;
  assign n50373 = n50372 ^ n27522 ^ 1'b0 ;
  assign n50374 = ~n12578 & n31678 ;
  assign n50375 = n50374 ^ n44019 ^ 1'b0 ;
  assign n50376 = n42808 ^ n5591 ^ 1'b0 ;
  assign n50377 = ~n17838 & n32672 ;
  assign n50378 = n7335 & n20679 ;
  assign n50379 = n50378 ^ n34012 ^ 1'b0 ;
  assign n50380 = n28971 & n50379 ;
  assign n50381 = ( n19731 & n50377 ) | ( n19731 & ~n50380 ) | ( n50377 & ~n50380 ) ;
  assign n50382 = n34137 ^ n16120 ^ 1'b0 ;
  assign n50383 = n13285 ^ n2196 ^ 1'b0 ;
  assign n50384 = n50383 ^ n12923 ^ n1267 ;
  assign n50385 = n2064 & n50384 ;
  assign n50386 = n50385 ^ n10088 ^ 1'b0 ;
  assign n50387 = ~n38266 & n50386 ;
  assign n50388 = n6264 | n45576 ;
  assign n50389 = n41812 ^ n25164 ^ 1'b0 ;
  assign n50390 = n50388 & n50389 ;
  assign n50391 = n741 & ~n2671 ;
  assign n50392 = ~n3745 & n14361 ;
  assign n50393 = ~n7260 & n50392 ;
  assign n50394 = n50393 ^ n49705 ^ n8942 ;
  assign n50395 = n7243 ^ n801 ^ 1'b0 ;
  assign n50396 = n8625 & ~n50395 ;
  assign n50397 = n50396 ^ n1100 ^ 1'b0 ;
  assign n50399 = ~n1267 & n16303 ;
  assign n50400 = n3299 & n50399 ;
  assign n50398 = n1898 & n45692 ;
  assign n50401 = n50400 ^ n50398 ^ 1'b0 ;
  assign n50402 = ( n3377 & n6856 ) | ( n3377 & ~n6899 ) | ( n6856 & ~n6899 ) ;
  assign n50403 = n5073 & ~n50402 ;
  assign n50404 = ~n879 & n50403 ;
  assign n50405 = n50404 ^ n42327 ^ 1'b0 ;
  assign n50406 = ~n9409 & n46737 ;
  assign n50407 = n50406 ^ n10859 ^ 1'b0 ;
  assign n50408 = n178 & ~n18248 ;
  assign n50409 = n43193 ^ n23270 ^ n17346 ;
  assign n50410 = n50409 ^ n17866 ^ 1'b0 ;
  assign n50411 = n1264 & ~n50410 ;
  assign n50412 = ~n21307 & n50411 ;
  assign n50413 = ( ~n6052 & n7169 ) | ( ~n6052 & n35198 ) | ( n7169 & n35198 ) ;
  assign n50414 = n50413 ^ n11922 ^ 1'b0 ;
  assign n50415 = n47000 ^ n29138 ^ 1'b0 ;
  assign n50416 = n4932 & ~n50415 ;
  assign n50417 = ~n6034 & n19936 ;
  assign n50418 = n7460 | n30096 ;
  assign n50419 = n22848 ^ n18598 ^ 1'b0 ;
  assign n50420 = n41217 | n50419 ;
  assign n50421 = n31317 ^ n25482 ^ 1'b0 ;
  assign n50422 = ~n30706 & n50421 ;
  assign n50423 = n23873 | n50422 ;
  assign n50424 = n9770 ^ n6129 ^ 1'b0 ;
  assign n50425 = n50423 & n50424 ;
  assign n50426 = n49978 ^ n41746 ^ 1'b0 ;
  assign n50427 = ( n8411 & n23648 ) | ( n8411 & n33145 ) | ( n23648 & n33145 ) ;
  assign n50428 = n17656 ^ n11129 ^ 1'b0 ;
  assign n50429 = n17736 & n50428 ;
  assign n50430 = n49677 ^ n29889 ^ 1'b0 ;
  assign n50431 = ~n824 & n9571 ;
  assign n50432 = n50431 ^ n37 ^ 1'b0 ;
  assign n50433 = n50432 ^ n3777 ^ 1'b0 ;
  assign n50434 = n50430 | n50433 ;
  assign n50435 = n20548 & ~n21518 ;
  assign n50436 = n23813 ^ n317 ^ 1'b0 ;
  assign n50437 = n31359 & n50436 ;
  assign n50438 = ( n6320 & ~n50435 ) | ( n6320 & n50437 ) | ( ~n50435 & n50437 ) ;
  assign n50439 = n25539 ^ n16809 ^ 1'b0 ;
  assign n50440 = n10775 & ~n50439 ;
  assign n50441 = n49679 ^ n4372 ^ 1'b0 ;
  assign n50442 = n3330 & n50441 ;
  assign n50443 = n33863 ^ n14880 ^ 1'b0 ;
  assign n50447 = n50163 ^ n28397 ^ 1'b0 ;
  assign n50448 = n8355 & ~n50447 ;
  assign n50444 = n19959 ^ n153 ^ 1'b0 ;
  assign n50445 = ~n28991 & n50444 ;
  assign n50446 = n12275 & n50445 ;
  assign n50449 = n50448 ^ n50446 ^ n23723 ;
  assign n50450 = n13729 & ~n50449 ;
  assign n50451 = ~n8514 & n23492 ;
  assign n50452 = n47256 & ~n50451 ;
  assign n50453 = ~n30919 & n50452 ;
  assign n50454 = n1889 | n6618 ;
  assign n50455 = n33834 | n50454 ;
  assign n50456 = n13496 & n13640 ;
  assign n50457 = n50456 ^ n24072 ^ 1'b0 ;
  assign n50458 = n3214 & n27735 ;
  assign n50459 = n50458 ^ n19833 ^ 1'b0 ;
  assign n50460 = n4471 & ~n50459 ;
  assign n50461 = n50460 ^ n1845 ^ 1'b0 ;
  assign n50462 = n50461 ^ n21541 ^ 1'b0 ;
  assign n50463 = n16403 | n50462 ;
  assign n50464 = n19996 ^ n4877 ^ 1'b0 ;
  assign n50465 = n25377 ^ n9707 ^ 1'b0 ;
  assign n50466 = n9759 ^ n8493 ^ 1'b0 ;
  assign n50467 = n48111 & n50466 ;
  assign n50468 = n21781 ^ n6071 ^ 1'b0 ;
  assign n50469 = n50468 ^ n35284 ^ n16362 ;
  assign n50470 = n3652 & n22528 ;
  assign n50471 = n45061 ^ n34021 ^ n32135 ;
  assign n50472 = n23188 & n32425 ;
  assign n50473 = n30295 & n50472 ;
  assign n50474 = n25531 ^ n12590 ^ 1'b0 ;
  assign n50475 = n14857 ^ n9506 ^ 1'b0 ;
  assign n50476 = n9265 & ~n50475 ;
  assign n50477 = n12377 ^ n6230 ^ 1'b0 ;
  assign n50478 = n21946 & ~n50477 ;
  assign n50479 = n50478 ^ n50090 ^ n13275 ;
  assign n50480 = n4344 | n5734 ;
  assign n50481 = n26243 | n50480 ;
  assign n50482 = ~n9868 & n50481 ;
  assign n50484 = n6821 ^ n5373 ^ 1'b0 ;
  assign n50485 = n25216 & n50484 ;
  assign n50483 = n7601 & ~n23556 ;
  assign n50486 = n50485 ^ n50483 ^ 1'b0 ;
  assign n50487 = n7276 | n36604 ;
  assign n50488 = n12548 | n50487 ;
  assign n50489 = n36686 ^ n14185 ^ n9377 ;
  assign n50490 = n50489 ^ n16235 ^ 1'b0 ;
  assign n50491 = ~n77 & n46419 ;
  assign n50492 = n16540 ^ n2106 ^ 1'b0 ;
  assign n50493 = ~n14962 & n50492 ;
  assign n50494 = n25338 & n31436 ;
  assign n50495 = n6856 & n50494 ;
  assign n50496 = ( n13712 & ~n50493 ) | ( n13712 & n50495 ) | ( ~n50493 & n50495 ) ;
  assign n50497 = ~n4977 & n24627 ;
  assign n50498 = ~n8023 & n50497 ;
  assign n50499 = n50498 ^ n27619 ^ n523 ;
  assign n50500 = n1153 | n50499 ;
  assign n50501 = n4301 & ~n5925 ;
  assign n50502 = n45445 | n50501 ;
  assign n50503 = n50502 ^ n27563 ^ 1'b0 ;
  assign n50504 = ~n15563 & n17771 ;
  assign n50505 = n1105 & n21561 ;
  assign n50506 = n50505 ^ n15972 ^ 1'b0 ;
  assign n50507 = n50506 ^ n19795 ^ 1'b0 ;
  assign n50508 = n40054 & ~n50507 ;
  assign n50509 = n41211 ^ n10777 ^ 1'b0 ;
  assign n50510 = n20343 ^ n17204 ^ n15076 ;
  assign n50511 = n1729 & n50510 ;
  assign n50512 = n15347 | n31415 ;
  assign n50513 = n621 | n50512 ;
  assign n50514 = n18129 | n44895 ;
  assign n50515 = n39603 & ~n50514 ;
  assign n50516 = ( ~n33225 & n50513 ) | ( ~n33225 & n50515 ) | ( n50513 & n50515 ) ;
  assign n50517 = n19630 ^ n601 ^ 1'b0 ;
  assign n50518 = n2851 | n50517 ;
  assign n50520 = ~n25672 & n46388 ;
  assign n50521 = ~n2106 & n50520 ;
  assign n50519 = n5012 & ~n42849 ;
  assign n50522 = n50521 ^ n50519 ^ 1'b0 ;
  assign n50523 = ~n20399 & n28204 ;
  assign n50524 = n50523 ^ n49153 ^ 1'b0 ;
  assign n50525 = n9996 & n24642 ;
  assign n50526 = n50525 ^ n18503 ^ n10230 ;
  assign n50527 = n14243 ^ n2421 ^ 1'b0 ;
  assign n50528 = n7707 & n50527 ;
  assign n50529 = ~n6025 & n50528 ;
  assign n50530 = n22597 ^ n4491 ^ 1'b0 ;
  assign n50531 = n26671 ^ n14460 ^ 1'b0 ;
  assign n50532 = n50530 & ~n50531 ;
  assign n50533 = n40563 ^ n362 ^ 1'b0 ;
  assign n50535 = n3402 | n13340 ;
  assign n50536 = ~n21875 & n50535 ;
  assign n50534 = n5053 | n35471 ;
  assign n50537 = n50536 ^ n50534 ^ 1'b0 ;
  assign n50538 = n29571 ^ n8184 ^ 1'b0 ;
  assign n50539 = n33081 ^ n1407 ^ 1'b0 ;
  assign n50540 = n45346 ^ n39067 ^ n2140 ;
  assign n50541 = ~n10339 & n15308 ;
  assign n50542 = n40227 ^ n8832 ^ 1'b0 ;
  assign n50543 = n14635 ^ n6732 ^ 1'b0 ;
  assign n50544 = ~n45798 & n50543 ;
  assign n50545 = n11833 & n50544 ;
  assign n50546 = n32853 & n48143 ;
  assign n50547 = n50546 ^ n24877 ^ 1'b0 ;
  assign n50548 = n2418 | n26702 ;
  assign n50549 = n31276 ^ n17455 ^ n7482 ;
  assign n50550 = n17362 ^ n6852 ^ 1'b0 ;
  assign n50551 = ~n8911 & n50550 ;
  assign n50552 = n50551 ^ n2037 ^ 1'b0 ;
  assign n50553 = ~n50549 & n50552 ;
  assign n50554 = n2823 & ~n20469 ;
  assign n50555 = ~n11540 & n50554 ;
  assign n50556 = n50555 ^ n17371 ^ 1'b0 ;
  assign n50557 = ~n8952 & n21686 ;
  assign n50558 = n4497 ^ n4116 ^ 1'b0 ;
  assign n50559 = n50558 ^ n26392 ^ 1'b0 ;
  assign n50560 = ~n8356 & n31063 ;
  assign n50561 = n49673 & ~n50560 ;
  assign n50562 = n21893 & ~n39682 ;
  assign n50563 = n7377 & ~n33089 ;
  assign n50564 = n12959 & ~n50563 ;
  assign n50565 = n3866 ^ n2620 ^ 1'b0 ;
  assign n50566 = n37669 ^ n18248 ^ 1'b0 ;
  assign n50567 = n15396 ^ n12260 ^ n9923 ;
  assign n50568 = n33337 & n50567 ;
  assign n50569 = n50568 ^ n21205 ^ 1'b0 ;
  assign n50570 = ~n17763 & n28471 ;
  assign n50571 = n50526 | n50570 ;
  assign n50572 = n50571 ^ n23123 ^ 1'b0 ;
  assign n50573 = n35595 ^ n28885 ^ 1'b0 ;
  assign n50574 = ( n12875 & ~n43708 ) | ( n12875 & n50573 ) | ( ~n43708 & n50573 ) ;
  assign n50575 = n23227 ^ n11898 ^ 1'b0 ;
  assign n50576 = ~n6042 & n16572 ;
  assign n50577 = n26859 & n50576 ;
  assign n50578 = ( ~n47763 & n50575 ) | ( ~n47763 & n50577 ) | ( n50575 & n50577 ) ;
  assign n50579 = n24807 & ~n26395 ;
  assign n50580 = n25004 & ~n47348 ;
  assign n50581 = n50580 ^ n12875 ^ 1'b0 ;
  assign n50582 = n8346 | n50581 ;
  assign n50583 = n3420 & ~n18613 ;
  assign n50584 = ~n19903 & n50583 ;
  assign n50585 = n3038 & n10617 ;
  assign n50586 = n50585 ^ n31879 ^ 1'b0 ;
  assign n50587 = n10404 ^ n4775 ^ 1'b0 ;
  assign n50588 = n50586 & ~n50587 ;
  assign n50589 = n12879 & ~n19875 ;
  assign n50590 = n10579 & n36627 ;
  assign n50591 = n50590 ^ n6060 ^ 1'b0 ;
  assign n50592 = n39309 ^ n25662 ^ n6490 ;
  assign n50593 = n50592 ^ n15190 ^ 1'b0 ;
  assign n50594 = n13909 | n50593 ;
  assign n50595 = n156 & ~n47444 ;
  assign n50598 = n1330 | n6833 ;
  assign n50599 = n31220 & ~n50598 ;
  assign n50596 = n19741 & ~n29585 ;
  assign n50597 = n50596 ^ n37474 ^ n10741 ;
  assign n50600 = n50599 ^ n50597 ^ 1'b0 ;
  assign n50601 = n5776 ^ n4959 ^ x3 ;
  assign n50602 = n35505 & n39678 ;
  assign n50603 = n50601 & n50602 ;
  assign n50604 = n17150 | n33585 ;
  assign n50605 = ~n50603 & n50604 ;
  assign n50606 = n2897 & n31700 ;
  assign n50607 = n23605 & n30196 ;
  assign n50608 = n50607 ^ n11372 ^ 1'b0 ;
  assign n50609 = n15514 ^ n15490 ^ 1'b0 ;
  assign n50610 = n15332 & n50609 ;
  assign n50611 = ~n8282 & n50610 ;
  assign n50612 = ~n13002 & n34095 ;
  assign n50613 = n17220 & n37108 ;
  assign n50614 = n50613 ^ n563 ^ 1'b0 ;
  assign n50615 = ~n5995 & n8891 ;
  assign n50616 = n50615 ^ n11103 ^ 1'b0 ;
  assign n50617 = n6045 & n50616 ;
  assign n50618 = n11795 | n14801 ;
  assign n50619 = ( n2944 & n16647 ) | ( n2944 & n50618 ) | ( n16647 & n50618 ) ;
  assign n50620 = n50004 ^ n26566 ^ 1'b0 ;
  assign n50621 = n6247 & ~n50620 ;
  assign n50622 = n3941 & ~n38660 ;
  assign n50623 = n50622 ^ n36488 ^ n12671 ;
  assign n50624 = n50623 ^ n2922 ^ 1'b0 ;
  assign n50625 = ~n13938 & n29840 ;
  assign n50626 = ~n35378 & n50625 ;
  assign n50627 = n33923 ^ n13306 ^ 1'b0 ;
  assign n50628 = ~n12685 & n50627 ;
  assign n50629 = ( n1979 & ~n9912 ) | ( n1979 & n21896 ) | ( ~n9912 & n21896 ) ;
  assign n50630 = n9606 ^ n5724 ^ 1'b0 ;
  assign n50631 = n50630 ^ n18855 ^ n14766 ;
  assign n50632 = ~n2452 & n21119 ;
  assign n50633 = n8402 & ~n31189 ;
  assign n50634 = n21787 | n22185 ;
  assign n50635 = n50634 ^ n17042 ^ 1'b0 ;
  assign n50636 = n20919 ^ n1393 ^ 1'b0 ;
  assign n50637 = n50635 | n50636 ;
  assign n50638 = n1777 | n22835 ;
  assign n50639 = ( n398 & ~n23722 ) | ( n398 & n50638 ) | ( ~n23722 & n50638 ) ;
  assign n50640 = n5099 ^ n1118 ^ 1'b0 ;
  assign n50641 = ( n5890 & n50639 ) | ( n5890 & ~n50640 ) | ( n50639 & ~n50640 ) ;
  assign n50642 = n35121 ^ n20779 ^ 1'b0 ;
  assign n50643 = ( n20475 & ~n23458 ) | ( n20475 & n41722 ) | ( ~n23458 & n41722 ) ;
  assign n50644 = ~n14943 & n43721 ;
  assign n50645 = n40723 & n50644 ;
  assign n50646 = n22403 ^ n1154 ^ 1'b0 ;
  assign n50647 = n18779 & n50646 ;
  assign n50648 = n50647 ^ n47773 ^ 1'b0 ;
  assign n50649 = ~n1712 & n4457 ;
  assign n50650 = ~n4457 & n50649 ;
  assign n50651 = n36 & n442 ;
  assign n50652 = ~n36 & n50651 ;
  assign n50653 = n156 & ~n50652 ;
  assign n50654 = n50653 ^ n21743 ^ 1'b0 ;
  assign n50655 = ~n50650 & n50654 ;
  assign n50661 = n452 & ~n581 ;
  assign n50662 = ~n452 & n50661 ;
  assign n50663 = n50662 ^ n2728 ^ 1'b0 ;
  assign n50656 = n2787 & ~n11642 ;
  assign n50657 = n11642 & n50656 ;
  assign n50658 = ~n7655 & n50657 ;
  assign n50659 = n4177 & n50658 ;
  assign n50660 = n50659 ^ n16041 ^ 1'b0 ;
  assign n50664 = n50663 ^ n50660 ^ 1'b0 ;
  assign n50665 = n50655 & ~n50664 ;
  assign n50666 = n20436 ^ n10305 ^ n4884 ;
  assign n50667 = n16833 ^ n3003 ^ 1'b0 ;
  assign n50668 = n4815 | n50667 ;
  assign n50669 = n50668 ^ n1639 ^ 1'b0 ;
  assign n50670 = n5713 & ~n8519 ;
  assign n50671 = n50670 ^ n2823 ^ 1'b0 ;
  assign n50672 = n14595 | n19944 ;
  assign n50673 = ( ~n26228 & n50671 ) | ( ~n26228 & n50672 ) | ( n50671 & n50672 ) ;
  assign n50674 = n50673 ^ n7839 ^ n7062 ;
  assign n50675 = n37398 ^ n26360 ^ n8414 ;
  assign n50676 = n777 & ~n17567 ;
  assign n50677 = n12224 & ~n13524 ;
  assign n50678 = n50677 ^ n7749 ^ 1'b0 ;
  assign n50679 = n50678 ^ n381 ^ 1'b0 ;
  assign n50680 = ~n50676 & n50679 ;
  assign n50681 = n2059 & n25941 ;
  assign n50682 = n12878 & ~n40865 ;
  assign n50683 = n22550 | n23718 ;
  assign n50684 = n44046 ^ n30395 ^ n14760 ;
  assign n50685 = n12500 & n41791 ;
  assign n50686 = n50685 ^ n4858 ^ 1'b0 ;
  assign n50687 = n50686 ^ n19766 ^ n7553 ;
  assign n50688 = n4612 | n43652 ;
  assign n50689 = n32421 ^ n22815 ^ 1'b0 ;
  assign n50691 = n27270 ^ n19844 ^ 1'b0 ;
  assign n50690 = n740 | n36244 ;
  assign n50692 = n50691 ^ n50690 ^ 1'b0 ;
  assign n50693 = n37404 | n38155 ;
  assign n50694 = n863 & n20967 ;
  assign n50695 = ~n22063 & n50694 ;
  assign n50698 = ( n6934 & n14064 ) | ( n6934 & ~n33571 ) | ( n14064 & ~n33571 ) ;
  assign n50696 = n45447 ^ n40523 ^ 1'b0 ;
  assign n50697 = ~n6358 & n50696 ;
  assign n50699 = n50698 ^ n50697 ^ 1'b0 ;
  assign n50700 = ( n647 & n6996 ) | ( n647 & ~n34488 ) | ( n6996 & ~n34488 ) ;
  assign n50701 = ( n2086 & n2107 ) | ( n2086 & ~n18998 ) | ( n2107 & ~n18998 ) ;
  assign n50702 = n1013 & n5392 ;
  assign n50703 = n50701 | n50702 ;
  assign n50704 = ~n996 & n1204 ;
  assign n50705 = n44380 & n50704 ;
  assign n50706 = ~n878 & n12695 ;
  assign n50707 = n38639 ^ n8655 ^ 1'b0 ;
  assign n50708 = n50706 & ~n50707 ;
  assign n50709 = n20706 ^ n3505 ^ 1'b0 ;
  assign n50710 = n50709 ^ n46971 ^ n4131 ;
  assign n50711 = n3299 & n50710 ;
  assign n50712 = ~n8616 & n18935 ;
  assign n50713 = n43287 ^ n7310 ^ 1'b0 ;
  assign n50714 = n10754 & n35369 ;
  assign n50715 = n18036 ^ n16627 ^ n1906 ;
  assign n50716 = n22617 & n50715 ;
  assign n50717 = n32913 ^ n17170 ^ 1'b0 ;
  assign n50718 = n7055 & n50717 ;
  assign n50719 = n34798 ^ n14719 ^ 1'b0 ;
  assign n50720 = n35242 & n50719 ;
  assign n50721 = n50720 ^ n26843 ^ 1'b0 ;
  assign n50722 = n42929 ^ n11009 ^ n2513 ;
  assign n50723 = n11121 & n13586 ;
  assign n50724 = n50723 ^ n31329 ^ 1'b0 ;
  assign n50725 = n49470 & ~n50724 ;
  assign n50726 = n28278 & n34724 ;
  assign n50727 = n50726 ^ n48576 ^ 1'b0 ;
  assign n50728 = ~n11734 & n29593 ;
  assign n50729 = n50728 ^ n16719 ^ 1'b0 ;
  assign n50730 = n6079 & n18096 ;
  assign n50731 = ~n49988 & n50730 ;
  assign n50732 = n29579 & ~n47810 ;
  assign n50733 = n1332 | n15866 ;
  assign n50734 = n50733 ^ n3826 ^ 1'b0 ;
  assign n50735 = n4804 & ~n30188 ;
  assign n50736 = n50735 ^ n36035 ^ 1'b0 ;
  assign n50737 = n13631 & ~n33933 ;
  assign n50738 = n50737 ^ n40073 ^ n28091 ;
  assign n50739 = n28406 ^ n2935 ^ 1'b0 ;
  assign n50740 = n38957 ^ n27903 ^ n5535 ;
  assign n50741 = n4780 ^ n4288 ^ 1'b0 ;
  assign n50742 = n18912 ^ n15250 ^ 1'b0 ;
  assign n50743 = ~n3425 & n28125 ;
  assign n50744 = n50742 & n50743 ;
  assign n50745 = n25549 ^ n4789 ^ 1'b0 ;
  assign n50746 = n8099 & n50745 ;
  assign n50747 = n47816 ^ n3534 ^ 1'b0 ;
  assign n50748 = ~n24652 & n50747 ;
  assign n50752 = n38458 ^ n28206 ^ 1'b0 ;
  assign n50749 = ~n1525 & n1623 ;
  assign n50750 = n4845 & n50749 ;
  assign n50751 = n1766 | n50750 ;
  assign n50753 = n50752 ^ n50751 ^ 1'b0 ;
  assign n50754 = n8427 & ~n18458 ;
  assign n50755 = n48227 & n50754 ;
  assign n50756 = n47269 ^ n640 ^ 1'b0 ;
  assign n50757 = ( n3171 & n8148 ) | ( n3171 & n24477 ) | ( n8148 & n24477 ) ;
  assign n50758 = n22702 ^ n17109 ^ n11508 ;
  assign n50759 = n40486 ^ n9379 ^ 1'b0 ;
  assign n50760 = n13608 | n29242 ;
  assign n50761 = n50760 ^ n17110 ^ 1'b0 ;
  assign n50762 = n5895 | n23900 ;
  assign n50763 = n2485 | n50762 ;
  assign n50764 = n10392 & n46349 ;
  assign n50765 = ~n50763 & n50764 ;
  assign n50766 = n16829 | n36316 ;
  assign n50767 = n8958 & ~n50766 ;
  assign n50768 = n37632 & n50767 ;
  assign n50769 = n3751 | n5135 ;
  assign n50770 = n23905 | n50769 ;
  assign n50771 = n50770 ^ n20356 ^ 1'b0 ;
  assign n50772 = ( ~n11724 & n16521 ) | ( ~n11724 & n48378 ) | ( n16521 & n48378 ) ;
  assign n50773 = n3566 & ~n6071 ;
  assign n50774 = ~n6503 & n50773 ;
  assign n50775 = n44154 ^ n23550 ^ n12030 ;
  assign n50776 = n7945 | n27783 ;
  assign n50777 = n3284 & ~n50776 ;
  assign n50778 = ( n25724 & n50775 ) | ( n25724 & ~n50777 ) | ( n50775 & ~n50777 ) ;
  assign n50779 = n50774 | n50778 ;
  assign n50780 = n50779 ^ n7869 ^ n5156 ;
  assign n50781 = n50592 ^ n13208 ^ 1'b0 ;
  assign n50782 = n6678 | n50781 ;
  assign n50784 = n3606 & ~n15142 ;
  assign n50783 = n10406 | n13703 ;
  assign n50785 = n50784 ^ n50783 ^ 1'b0 ;
  assign n50786 = n45627 ^ n14071 ^ n10313 ;
  assign n50787 = n38023 ^ n1135 ^ 1'b0 ;
  assign n50788 = n25120 & n44358 ;
  assign n50789 = n37457 ^ n24998 ^ n13223 ;
  assign n50790 = ~n34570 & n50789 ;
  assign n50791 = n50790 ^ n9549 ^ 1'b0 ;
  assign n50792 = n16554 & n34496 ;
  assign n50793 = n24246 ^ n390 ^ 1'b0 ;
  assign n50794 = ~n12539 & n27605 ;
  assign n50795 = n42880 ^ n9634 ^ 1'b0 ;
  assign n50796 = ~n41436 & n50795 ;
  assign n50797 = n28333 ^ n18162 ^ n1529 ;
  assign n50798 = n50797 ^ n26094 ^ 1'b0 ;
  assign n50799 = n23108 ^ n6690 ^ 1'b0 ;
  assign n50800 = n3988 | n12459 ;
  assign n50801 = n50800 ^ n26233 ^ 1'b0 ;
  assign n50802 = n34648 & ~n34921 ;
  assign n50803 = n50801 & n50802 ;
  assign n50804 = n13620 | n23211 ;
  assign n50805 = ~n1371 & n4647 ;
  assign n50806 = n5716 & n50805 ;
  assign n50807 = ~n18849 & n25148 ;
  assign n50808 = n28333 & n50807 ;
  assign n50809 = n32587 ^ n12969 ^ 1'b0 ;
  assign n50811 = ~n16132 & n38057 ;
  assign n50810 = ( n4972 & ~n6440 ) | ( n4972 & n7188 ) | ( ~n6440 & n7188 ) ;
  assign n50812 = n50811 ^ n50810 ^ 1'b0 ;
  assign n50813 = ~n7886 & n8389 ;
  assign n50814 = n47085 ^ n26533 ^ 1'b0 ;
  assign n50815 = n10393 | n20524 ;
  assign n50816 = n17865 | n50815 ;
  assign n50817 = n50816 ^ n1435 ^ 1'b0 ;
  assign n50818 = n21823 & ~n50817 ;
  assign n50819 = n30192 ^ n19799 ^ 1'b0 ;
  assign n50820 = n27095 & ~n47846 ;
  assign n50821 = ~n28767 & n47136 ;
  assign n50822 = n50821 ^ n20155 ^ 1'b0 ;
  assign n50823 = ( n12940 & n16832 ) | ( n12940 & ~n23928 ) | ( n16832 & ~n23928 ) ;
  assign n50824 = n50823 ^ n44701 ^ n32029 ;
  assign n50825 = ( n12882 & n35164 ) | ( n12882 & n41384 ) | ( n35164 & n41384 ) ;
  assign n50826 = ( n9263 & ~n17078 ) | ( n9263 & n50825 ) | ( ~n17078 & n50825 ) ;
  assign n50827 = n13140 ^ n5397 ^ 1'b0 ;
  assign n50828 = n8466 & n50827 ;
  assign n50829 = n50828 ^ n8009 ^ n5102 ;
  assign n50830 = n32103 | n40212 ;
  assign n50831 = n6574 | n6816 ;
  assign n50832 = n12384 | n50831 ;
  assign n50833 = n28390 ^ n3174 ^ 1'b0 ;
  assign n50834 = n50832 & n50833 ;
  assign n50835 = n1767 & ~n7316 ;
  assign n50836 = n20311 & n50835 ;
  assign n50837 = n35961 & ~n50836 ;
  assign n50838 = n7792 | n14146 ;
  assign n50839 = ( n2375 & n30398 ) | ( n2375 & n50838 ) | ( n30398 & n50838 ) ;
  assign n50840 = n18495 & n50839 ;
  assign n50841 = ~n47734 & n50840 ;
  assign n50842 = n46531 ^ n34408 ^ n13298 ;
  assign n50843 = n21321 & n30791 ;
  assign n50844 = ( n1361 & n14677 ) | ( n1361 & ~n50843 ) | ( n14677 & ~n50843 ) ;
  assign n50845 = ~n9692 & n25313 ;
  assign n50846 = n19689 | n29683 ;
  assign n50847 = n50846 ^ n2399 ^ 1'b0 ;
  assign n50848 = n17769 & ~n50847 ;
  assign n50849 = n34428 & n50848 ;
  assign n50850 = n9816 | n26081 ;
  assign n50851 = n37559 & ~n50850 ;
  assign n50852 = n19084 & ~n50851 ;
  assign n50853 = n6278 & n50852 ;
  assign n50854 = n24320 & n25526 ;
  assign n50855 = n31901 ^ n8220 ^ 1'b0 ;
  assign n50856 = n49765 | n50855 ;
  assign n50857 = n30002 ^ x10 ^ 1'b0 ;
  assign n50858 = n27529 | n35900 ;
  assign n50859 = n50858 ^ n40563 ^ 1'b0 ;
  assign n50860 = ~n24196 & n50859 ;
  assign n50861 = ~n5132 & n20827 ;
  assign n50862 = ( n4283 & n10825 ) | ( n4283 & n21443 ) | ( n10825 & n21443 ) ;
  assign n50863 = n50862 ^ n38353 ^ n27391 ;
  assign n50864 = ( n24759 & n29515 ) | ( n24759 & ~n44685 ) | ( n29515 & ~n44685 ) ;
  assign n50865 = n11609 & ~n43254 ;
  assign n50866 = n4782 ^ n2234 ^ 1'b0 ;
  assign n50867 = n19915 ^ n3207 ^ 1'b0 ;
  assign n50868 = ~n50866 & n50867 ;
  assign n50869 = n11019 | n14482 ;
  assign n50870 = n24270 & ~n37454 ;
  assign n50871 = n3959 & ~n37554 ;
  assign n50872 = n14287 & ~n50871 ;
  assign n50873 = ~n46252 & n50872 ;
  assign n50874 = n19596 ^ n9605 ^ 1'b0 ;
  assign n50875 = n1045 | n50874 ;
  assign n50876 = ( n8498 & n24101 ) | ( n8498 & n50875 ) | ( n24101 & n50875 ) ;
  assign n50877 = ( ~n5722 & n20771 ) | ( ~n5722 & n38275 ) | ( n20771 & n38275 ) ;
  assign n50878 = n50877 ^ n21521 ^ 1'b0 ;
  assign n50879 = ( n1751 & n3799 ) | ( n1751 & n14373 ) | ( n3799 & n14373 ) ;
  assign n50880 = n29927 & n48928 ;
  assign n50881 = n48959 & n50880 ;
  assign n50882 = n48670 ^ n22450 ^ 1'b0 ;
  assign n50883 = n35147 ^ n7053 ^ n5478 ;
  assign n50884 = ~n8010 & n37497 ;
  assign n50885 = n1952 & n50884 ;
  assign n50889 = ~n8201 & n23739 ;
  assign n50886 = n7981 ^ n2751 ^ 1'b0 ;
  assign n50887 = n25766 | n50886 ;
  assign n50888 = n50887 ^ n38660 ^ 1'b0 ;
  assign n50890 = n50889 ^ n50888 ^ 1'b0 ;
  assign n50891 = n50885 | n50890 ;
  assign n50892 = n37004 ^ n9191 ^ n6778 ;
  assign n50893 = n2317 & n50892 ;
  assign n50894 = n18148 | n50893 ;
  assign n50895 = n26124 & ~n32283 ;
  assign n50896 = n50895 ^ n37403 ^ 1'b0 ;
  assign n50897 = n47774 ^ n45855 ^ 1'b0 ;
  assign n50900 = ~n13139 & n17827 ;
  assign n50898 = ( n13023 & n34496 ) | ( n13023 & ~n46041 ) | ( n34496 & ~n46041 ) ;
  assign n50899 = n5533 & n50898 ;
  assign n50901 = n50900 ^ n50899 ^ 1'b0 ;
  assign n50902 = ( ~n1575 & n26717 ) | ( ~n1575 & n50901 ) | ( n26717 & n50901 ) ;
  assign n50903 = ~n13478 & n16075 ;
  assign n50904 = ~n27851 & n50903 ;
  assign n50905 = n12387 | n16711 ;
  assign n50906 = n50904 & ~n50905 ;
  assign n50907 = ~n37376 & n46952 ;
  assign n50908 = n15066 & ~n50907 ;
  assign n50909 = n37946 ^ n20648 ^ 1'b0 ;
  assign n50910 = n34819 & n43830 ;
  assign n50911 = n15237 | n43660 ;
  assign n50912 = n16883 & ~n50911 ;
  assign n50913 = n14236 ^ n2511 ^ 1'b0 ;
  assign n50914 = n50913 ^ n34806 ^ n27272 ;
  assign n50915 = ~n11419 & n23046 ;
  assign n50916 = ~n50914 & n50915 ;
  assign n50917 = n27742 ^ n5841 ^ 1'b0 ;
  assign n50918 = ( n19527 & n48719 ) | ( n19527 & ~n50917 ) | ( n48719 & ~n50917 ) ;
  assign n50919 = n11798 & n22674 ;
  assign n50920 = n25120 ^ n5483 ^ 1'b0 ;
  assign n50921 = ~n50919 & n50920 ;
  assign n50922 = n50921 ^ n27686 ^ n10962 ;
  assign n50923 = n24537 | n27342 ;
  assign n50924 = n50923 ^ n4235 ^ 1'b0 ;
  assign n50925 = ~n33833 & n50924 ;
  assign n50926 = n26971 & n50925 ;
  assign n50927 = n6623 | n33514 ;
  assign n50928 = n21772 & n50927 ;
  assign n50929 = n13218 & ~n39750 ;
  assign n50930 = ~n1575 & n50929 ;
  assign n50931 = n1228 & n13110 ;
  assign n50932 = n43436 & n50931 ;
  assign n50933 = n12051 & ~n27414 ;
  assign n50934 = ( n1722 & n9766 ) | ( n1722 & ~n17480 ) | ( n9766 & ~n17480 ) ;
  assign n50935 = n25194 & ~n50934 ;
  assign n50936 = ( n31513 & n33148 ) | ( n31513 & ~n37652 ) | ( n33148 & ~n37652 ) ;
  assign n50937 = n16294 | n18242 ;
  assign n50938 = ~n11226 & n36265 ;
  assign n50939 = n14252 | n16786 ;
  assign n50940 = n28662 & ~n50939 ;
  assign n50941 = ~n50938 & n50940 ;
  assign n50942 = n16192 ^ n5219 ^ 1'b0 ;
  assign n50943 = n50942 ^ n10748 ^ n3861 ;
  assign n50944 = n22473 ^ n22451 ^ 1'b0 ;
  assign n50945 = ~n42972 & n50944 ;
  assign n50946 = ( n2124 & ~n37762 ) | ( n2124 & n50945 ) | ( ~n37762 & n50945 ) ;
  assign n50947 = ~n8177 & n30461 ;
  assign n50952 = n16373 ^ n6998 ^ 1'b0 ;
  assign n50953 = ~n5640 & n50952 ;
  assign n50948 = n15315 ^ n1391 ^ 1'b0 ;
  assign n50949 = n38769 & ~n45965 ;
  assign n50950 = n50948 & n50949 ;
  assign n50951 = n45339 & ~n50950 ;
  assign n50954 = n50953 ^ n50951 ^ 1'b0 ;
  assign n50955 = ~n13249 & n29693 ;
  assign n50956 = ( n21090 & ~n22353 ) | ( n21090 & n48526 ) | ( ~n22353 & n48526 ) ;
  assign n50957 = ~n8654 & n50956 ;
  assign n50958 = ~n50955 & n50957 ;
  assign n50959 = n28252 ^ n18863 ^ n18210 ;
  assign n50960 = ~n26029 & n50959 ;
  assign n50961 = n2747 & ~n20927 ;
  assign n50962 = n20158 ^ n17020 ^ n7470 ;
  assign n50963 = n32652 & n47094 ;
  assign n50964 = n50963 ^ n14843 ^ 1'b0 ;
  assign n50965 = n50962 & n50964 ;
  assign n50966 = ( n29559 & n31299 ) | ( n29559 & ~n42619 ) | ( n31299 & ~n42619 ) ;
  assign n50967 = n34887 ^ n20734 ^ n8504 ;
  assign n50968 = ~n24962 & n30211 ;
  assign n50969 = n10830 & n50968 ;
  assign n50970 = ~n1290 & n32766 ;
  assign n50971 = n50970 ^ n12337 ^ 1'b0 ;
  assign n50972 = n15776 ^ n4216 ^ 1'b0 ;
  assign n50973 = n4596 & n50972 ;
  assign n50976 = ~n7251 & n8241 ;
  assign n50977 = n1961 & n50976 ;
  assign n50978 = n12697 & ~n50977 ;
  assign n50979 = n50978 ^ n25635 ^ 1'b0 ;
  assign n50974 = n26794 ^ n8057 ^ 1'b0 ;
  assign n50975 = n33217 & ~n50974 ;
  assign n50980 = n50979 ^ n50975 ^ 1'b0 ;
  assign n50981 = n8955 ^ n209 ^ 1'b0 ;
  assign n50982 = n13062 & ~n50981 ;
  assign n50983 = n1176 & n14792 ;
  assign n50984 = ~n25095 & n28241 ;
  assign n50985 = n38481 ^ n26192 ^ n17900 ;
  assign n50986 = ~n26729 & n43721 ;
  assign n50987 = ~n50985 & n50986 ;
  assign n50988 = n7795 & ~n34378 ;
  assign n50989 = n1599 | n19453 ;
  assign n50990 = n40410 ^ n6417 ^ 1'b0 ;
  assign n50991 = n13429 & n50990 ;
  assign n50996 = n30028 ^ n16805 ^ 1'b0 ;
  assign n50997 = ~n34887 & n50996 ;
  assign n50998 = n1475 & n29678 ;
  assign n50999 = ~n50997 & n50998 ;
  assign n50992 = n8802 & ~n8891 ;
  assign n50993 = ~n16628 & n50992 ;
  assign n50994 = n16388 ^ n937 ^ 1'b0 ;
  assign n50995 = ~n50993 & n50994 ;
  assign n51000 = n50999 ^ n50995 ^ n816 ;
  assign n51001 = n18751 ^ n16049 ^ 1'b0 ;
  assign n51002 = n51000 | n51001 ;
  assign n51003 = n1462 | n51002 ;
  assign n51004 = n51003 ^ n2651 ^ 1'b0 ;
  assign n51007 = n43515 ^ n28320 ^ 1'b0 ;
  assign n51008 = n16794 & n51007 ;
  assign n51005 = n12481 ^ n8480 ^ 1'b0 ;
  assign n51006 = n40593 & n51005 ;
  assign n51009 = n51008 ^ n51006 ^ n7707 ;
  assign n51011 = n1791 & ~n37646 ;
  assign n51012 = n14872 & ~n27450 ;
  assign n51013 = ~n51011 & n51012 ;
  assign n51014 = n45207 & ~n51013 ;
  assign n51010 = n14867 | n40425 ;
  assign n51015 = n51014 ^ n51010 ^ 1'b0 ;
  assign n51016 = ( ~n30276 & n34874 ) | ( ~n30276 & n51015 ) | ( n34874 & n51015 ) ;
  assign n51017 = ( n15389 & ~n31757 ) | ( n15389 & n46361 ) | ( ~n31757 & n46361 ) ;
  assign n51018 = n9479 | n22052 ;
  assign n51019 = ~n16580 & n18236 ;
  assign n51020 = n2733 & n20874 ;
  assign n51023 = n8641 & ~n15730 ;
  assign n51024 = n8522 & n51023 ;
  assign n51022 = n46120 ^ n18084 ^ n12272 ;
  assign n51021 = n23628 | n29599 ;
  assign n51025 = n51024 ^ n51022 ^ n51021 ;
  assign n51026 = n25701 ^ n13640 ^ 1'b0 ;
  assign n51027 = n25340 | n50927 ;
  assign n51028 = n37828 & n39182 ;
  assign n51029 = n51028 ^ n3985 ^ 1'b0 ;
  assign n51030 = n47678 & ~n51029 ;
  assign n51031 = ~n878 & n24168 ;
  assign n51032 = n51031 ^ n6369 ^ 1'b0 ;
  assign n51033 = n16299 & ~n51032 ;
  assign n51034 = n25881 & n51033 ;
  assign n51035 = n12266 ^ n401 ^ 1'b0 ;
  assign n51036 = n38562 ^ n112 ^ 1'b0 ;
  assign n51037 = n34589 ^ n17229 ^ 1'b0 ;
  assign n51038 = n19312 ^ n11759 ^ n5563 ;
  assign n51039 = n25149 & n51038 ;
  assign n51040 = n51039 ^ n7729 ^ 1'b0 ;
  assign n51041 = ~n20705 & n51040 ;
  assign n51042 = n51041 ^ n31099 ^ 1'b0 ;
  assign n51043 = n19570 | n50405 ;
  assign n51044 = n19056 & n19700 ;
  assign n51045 = n25101 & n51044 ;
  assign n51046 = n14285 ^ n13056 ^ 1'b0 ;
  assign n51047 = ~n2640 & n51046 ;
  assign n51048 = n20884 | n51047 ;
  assign n51049 = n20370 | n42153 ;
  assign n51050 = n51049 ^ n34606 ^ 1'b0 ;
  assign n51051 = n3523 ^ n169 ^ 1'b0 ;
  assign n51052 = n3303 & n51051 ;
  assign n51053 = n10588 ^ n9151 ^ n1066 ;
  assign n51054 = n51053 ^ n28918 ^ 1'b0 ;
  assign n51055 = n51052 | n51054 ;
  assign n51056 = n3882 & ~n9078 ;
  assign n51057 = ~n4115 & n51056 ;
  assign n51058 = ~n3066 & n15271 ;
  assign n51059 = n51057 & n51058 ;
  assign n51060 = ( n6646 & ~n31723 ) | ( n6646 & n50789 ) | ( ~n31723 & n50789 ) ;
  assign n51061 = n51060 ^ n7300 ^ 1'b0 ;
  assign n51062 = n9858 | n29133 ;
  assign n51063 = ~n126 & n51062 ;
  assign n51064 = n21655 ^ n16846 ^ n3691 ;
  assign n51065 = ~n7726 & n19810 ;
  assign n51066 = n51065 ^ n26064 ^ 1'b0 ;
  assign n51067 = n5855 | n19787 ;
  assign n51068 = ~n20970 & n51067 ;
  assign n51069 = n46955 | n51068 ;
  assign n51070 = n1281 & ~n7250 ;
  assign n51071 = ~n16554 & n51070 ;
  assign n51072 = n51071 ^ n12500 ^ 1'b0 ;
  assign n51073 = n15166 ^ n104 ^ 1'b0 ;
  assign n51074 = n49635 | n51073 ;
  assign n51075 = n25728 | n51074 ;
  assign n51076 = ( n1533 & n9967 ) | ( n1533 & ~n42273 ) | ( n9967 & ~n42273 ) ;
  assign n51077 = ~n31653 & n48379 ;
  assign n51078 = n51077 ^ n26759 ^ 1'b0 ;
  assign n51079 = n31908 & n51078 ;
  assign n51080 = ( n3067 & n20729 ) | ( n3067 & n48821 ) | ( n20729 & n48821 ) ;
  assign n51081 = n9360 & n51080 ;
  assign n51082 = n4267 | n41408 ;
  assign n51083 = n30079 & ~n51082 ;
  assign n51084 = ~n34881 & n50918 ;
  assign n51087 = n4471 | n10820 ;
  assign n51085 = ( n2827 & n22839 ) | ( n2827 & ~n27916 ) | ( n22839 & ~n27916 ) ;
  assign n51086 = n51085 ^ n3574 ^ 1'b0 ;
  assign n51088 = n51087 ^ n51086 ^ 1'b0 ;
  assign n51089 = n11283 | n13663 ;
  assign n51090 = n9847 | n51089 ;
  assign n51091 = ~n906 & n25210 ;
  assign n51092 = ( n28622 & ~n51008 ) | ( n28622 & n51091 ) | ( ~n51008 & n51091 ) ;
  assign n51093 = n28114 & ~n34661 ;
  assign n51094 = ~n24370 & n51093 ;
  assign n51095 = n51094 ^ n45514 ^ 1'b0 ;
  assign n51096 = ( n6118 & n8382 ) | ( n6118 & n12838 ) | ( n8382 & n12838 ) ;
  assign n51097 = n21343 ^ n67 ^ 1'b0 ;
  assign n51098 = n51096 | n51097 ;
  assign n51099 = ~n5441 & n15431 ;
  assign n51100 = n3456 ^ n3324 ^ 1'b0 ;
  assign n51101 = n13079 & ~n21518 ;
  assign n51102 = n51100 & n51101 ;
  assign n51103 = n19778 | n49982 ;
  assign n51104 = n15353 | n51103 ;
  assign n51105 = ( n7040 & ~n13602 ) | ( n7040 & n51104 ) | ( ~n13602 & n51104 ) ;
  assign n51106 = n777 & ~n1308 ;
  assign n51107 = n9255 | n51106 ;
  assign n51108 = n10350 | n51107 ;
  assign n51109 = ( ~n10983 & n21597 ) | ( ~n10983 & n51108 ) | ( n21597 & n51108 ) ;
  assign n51110 = n43398 ^ n28506 ^ n9732 ;
  assign n51111 = n19795 ^ n5010 ^ 1'b0 ;
  assign n51112 = n20049 | n51111 ;
  assign n51113 = n30113 | n35896 ;
  assign n51114 = ( n2966 & ~n7935 ) | ( n2966 & n37877 ) | ( ~n7935 & n37877 ) ;
  assign n51118 = n3850 ^ n181 ^ 1'b0 ;
  assign n51119 = n48515 & n51118 ;
  assign n51120 = n8226 & n34319 ;
  assign n51121 = ~n51119 & n51120 ;
  assign n51115 = n19200 ^ n978 ^ 1'b0 ;
  assign n51116 = ~n11542 & n51115 ;
  assign n51117 = n43971 & n51116 ;
  assign n51122 = n51121 ^ n51117 ^ n43288 ;
  assign n51123 = n20112 & ~n38548 ;
  assign n51124 = ~n32446 & n42224 ;
  assign n51125 = n11403 & n51124 ;
  assign n51126 = n6286 & ~n19288 ;
  assign n51127 = n4725 & n51126 ;
  assign n51128 = n18299 ^ n13742 ^ 1'b0 ;
  assign n51129 = n50638 | n51128 ;
  assign n51130 = n7165 | n37502 ;
  assign n51131 = n40116 & ~n51130 ;
  assign n51132 = n5836 ^ n1348 ^ 1'b0 ;
  assign n51133 = n51132 ^ n6197 ^ n1969 ;
  assign n51134 = n25839 ^ n11877 ^ 1'b0 ;
  assign n51135 = n51133 & ~n51134 ;
  assign n51136 = ~n18060 & n51135 ;
  assign n51137 = n4417 & n16462 ;
  assign n51138 = n51137 ^ n79 ^ 1'b0 ;
  assign n51139 = ( n6333 & n29387 ) | ( n6333 & n30182 ) | ( n29387 & n30182 ) ;
  assign n51140 = ( n36209 & n51138 ) | ( n36209 & ~n51139 ) | ( n51138 & ~n51139 ) ;
  assign n51141 = n51136 & ~n51140 ;
  assign n51142 = ~n16269 & n26090 ;
  assign n51143 = n51142 ^ n91 ^ 1'b0 ;
  assign n51144 = n8215 | n51143 ;
  assign n51145 = n4243 & ~n30509 ;
  assign n51146 = ~n7869 & n30664 ;
  assign n51147 = ~n2118 & n51146 ;
  assign n51148 = n32495 & ~n45108 ;
  assign n51149 = ( n17957 & n33006 ) | ( n17957 & n51148 ) | ( n33006 & n51148 ) ;
  assign n51150 = ~n34969 & n51149 ;
  assign n51152 = ( ~n3377 & n5919 ) | ( ~n3377 & n39367 ) | ( n5919 & n39367 ) ;
  assign n51151 = ~n27105 & n35350 ;
  assign n51153 = n51152 ^ n51151 ^ 1'b0 ;
  assign n51154 = n32334 ^ n8882 ^ 1'b0 ;
  assign n51155 = n41564 | n51154 ;
  assign n51156 = n28301 | n28714 ;
  assign n51157 = n51156 ^ n42797 ^ 1'b0 ;
  assign n51158 = n21378 ^ n13174 ^ n10660 ;
  assign n51159 = n1851 & ~n51158 ;
  assign n51160 = n51159 ^ n48372 ^ n34684 ;
  assign n51161 = ( n324 & n1848 ) | ( n324 & n15310 ) | ( n1848 & n15310 ) ;
  assign n51162 = n51161 ^ n23456 ^ 1'b0 ;
  assign n51163 = ~n40040 & n51162 ;
  assign n51164 = n51163 ^ n48864 ^ n46638 ;
  assign n51165 = n10760 & n51164 ;
  assign n51166 = n6460 | n7943 ;
  assign n51167 = n51166 ^ n19281 ^ n12578 ;
  assign n51168 = ~n37670 & n51167 ;
  assign n51169 = n30961 ^ n14332 ^ n10340 ;
  assign n51170 = ~n23259 & n51169 ;
  assign n51171 = n43857 ^ n3526 ^ 1'b0 ;
  assign n51172 = n6173 & ~n24792 ;
  assign n51173 = n37562 | n51172 ;
  assign n51174 = n45883 ^ n16666 ^ 1'b0 ;
  assign n51175 = n15138 | n17134 ;
  assign n51176 = n51175 ^ n8119 ^ 1'b0 ;
  assign n51177 = n45595 ^ n36128 ^ 1'b0 ;
  assign n51178 = n3188 | n51177 ;
  assign n51179 = ~n1964 & n4686 ;
  assign n51180 = n51178 & n51179 ;
  assign n51181 = n45205 & ~n51180 ;
  assign n51182 = n51176 & n51181 ;
  assign n51183 = n12895 ^ n4364 ^ 1'b0 ;
  assign n51184 = ~n30332 & n51183 ;
  assign n51185 = n51184 ^ n13917 ^ 1'b0 ;
  assign n51186 = n51185 ^ n18592 ^ 1'b0 ;
  assign n51187 = n45787 ^ n34779 ^ 1'b0 ;
  assign n51188 = n51187 ^ n39235 ^ n1213 ;
  assign n51189 = n1616 & ~n5612 ;
  assign n51190 = n51189 ^ n1336 ^ 1'b0 ;
  assign n51191 = ( n2140 & n4199 ) | ( n2140 & n51190 ) | ( n4199 & n51190 ) ;
  assign n51192 = n22520 & n29919 ;
  assign n51193 = n51192 ^ n19164 ^ 1'b0 ;
  assign n51194 = n29995 ^ n14438 ^ 1'b0 ;
  assign n51195 = ~n23662 & n51194 ;
  assign n51196 = ( n50156 & ~n51193 ) | ( n50156 & n51195 ) | ( ~n51193 & n51195 ) ;
  assign n51197 = n12248 & ~n42803 ;
  assign n51198 = n51197 ^ n35427 ^ 1'b0 ;
  assign n51199 = n2760 & n45479 ;
  assign n51200 = ( n1188 & n1932 ) | ( n1188 & ~n13857 ) | ( n1932 & ~n13857 ) ;
  assign n51201 = ( n18926 & n32742 ) | ( n18926 & n51200 ) | ( n32742 & n51200 ) ;
  assign n51202 = n9986 | n12969 ;
  assign n51203 = n51201 | n51202 ;
  assign n51204 = ~n18330 & n45002 ;
  assign n51205 = n25167 & n51204 ;
  assign n51206 = n41895 ^ n38266 ^ 1'b0 ;
  assign n51207 = n14882 & ~n34569 ;
  assign n51208 = n10239 & n48853 ;
  assign n51209 = n51208 ^ n11258 ^ 1'b0 ;
  assign n51210 = ~n10915 & n29726 ;
  assign n51211 = n51210 ^ n30347 ^ n21484 ;
  assign n51212 = n37929 | n51211 ;
  assign n51213 = n3523 & ~n39175 ;
  assign n51214 = ~n45037 & n51213 ;
  assign n51215 = n41031 | n47572 ;
  assign n51216 = n31634 ^ n8274 ^ 1'b0 ;
  assign n51217 = n19755 & n51216 ;
  assign n51218 = n45243 ^ n11521 ^ 1'b0 ;
  assign n51219 = n49681 & ~n51218 ;
  assign n51220 = n32992 & n51219 ;
  assign n51222 = n4067 ^ n1182 ^ 1'b0 ;
  assign n51223 = n51222 ^ n31213 ^ n192 ;
  assign n51221 = ~n3168 & n14343 ;
  assign n51224 = n51223 ^ n51221 ^ 1'b0 ;
  assign n51225 = n7722 | n25740 ;
  assign n51226 = ~n40491 & n46113 ;
  assign n51227 = n51226 ^ n7962 ^ 1'b0 ;
  assign n51228 = ( n1311 & n17422 ) | ( n1311 & ~n41483 ) | ( n17422 & ~n41483 ) ;
  assign n51229 = ( n15302 & n38793 ) | ( n15302 & ~n51228 ) | ( n38793 & ~n51228 ) ;
  assign n51230 = ~n26936 & n30244 ;
  assign n51231 = ~n51229 & n51230 ;
  assign n51232 = ( n4064 & ~n11750 ) | ( n4064 & n14246 ) | ( ~n11750 & n14246 ) ;
  assign n51233 = ~n16414 & n51232 ;
  assign n51234 = ~n16051 & n51233 ;
  assign n51235 = n51234 ^ n40374 ^ n5197 ;
  assign n51236 = n50297 ^ n45680 ^ 1'b0 ;
  assign n51237 = ~n9514 & n51236 ;
  assign n51238 = n51237 ^ n7694 ^ 1'b0 ;
  assign n51240 = n276 & n22012 ;
  assign n51239 = ~n13465 & n43237 ;
  assign n51241 = n51240 ^ n51239 ^ 1'b0 ;
  assign n51242 = n1096 & ~n3885 ;
  assign n51243 = ~n21552 & n51242 ;
  assign n51244 = n51243 ^ n2211 ^ 1'b0 ;
  assign n51245 = n5509 & ~n51244 ;
  assign n51246 = n3040 & ~n27258 ;
  assign n51247 = n23341 | n51246 ;
  assign n51248 = n51247 ^ n293 ^ 1'b0 ;
  assign n51249 = n21037 & ~n35145 ;
  assign n51250 = ~n17259 & n31678 ;
  assign n51251 = n43895 ^ n20033 ^ 1'b0 ;
  assign n51252 = n35926 & ~n51251 ;
  assign n51253 = ~n1249 & n51252 ;
  assign n51254 = n3508 & ~n14338 ;
  assign n51255 = n34521 ^ n5675 ^ 1'b0 ;
  assign n51256 = n5176 | n51255 ;
  assign n51257 = n30310 & n50945 ;
  assign n51258 = ~n962 & n51257 ;
  assign n51259 = ( n19351 & ~n51256 ) | ( n19351 & n51258 ) | ( ~n51256 & n51258 ) ;
  assign n51260 = n24633 ^ n17799 ^ n949 ;
  assign n51261 = n21714 | n51260 ;
  assign n51262 = n51261 ^ n20068 ^ 1'b0 ;
  assign n51263 = n17622 | n21997 ;
  assign n51264 = n49746 ^ n43324 ^ n8248 ;
  assign n51265 = n51264 ^ n39095 ^ n3659 ;
  assign n51266 = n51265 ^ n45172 ^ 1'b0 ;
  assign n51267 = n9428 | n51266 ;
  assign n51268 = n17554 ^ n13331 ^ 1'b0 ;
  assign n51269 = ~n42714 & n51268 ;
  assign n51270 = n16782 & n51269 ;
  assign n51271 = n33172 ^ n15306 ^ 1'b0 ;
  assign n51272 = n1071 & n51271 ;
  assign n51273 = n46707 ^ n5160 ^ 1'b0 ;
  assign n51274 = n13226 & ~n51273 ;
  assign n51275 = n42773 & ~n43500 ;
  assign n51276 = n12498 & n20344 ;
  assign n51277 = ( ~n12510 & n29898 ) | ( ~n12510 & n51276 ) | ( n29898 & n51276 ) ;
  assign n51278 = n30079 ^ n14297 ^ n6197 ;
  assign n51279 = n51278 ^ n37691 ^ 1'b0 ;
  assign n51280 = n14958 & ~n17754 ;
  assign n51281 = n51280 ^ n23731 ^ 1'b0 ;
  assign n51282 = n26561 ^ n16 ^ 1'b0 ;
  assign n51283 = ~n26176 & n51282 ;
  assign n51284 = ~n20358 & n32403 ;
  assign n51285 = n14046 & n51284 ;
  assign n51286 = ( n25232 & n30574 ) | ( n25232 & n51285 ) | ( n30574 & n51285 ) ;
  assign n51287 = n44062 & n44125 ;
  assign n51288 = n35609 ^ n8285 ^ 1'b0 ;
  assign n51289 = n24601 & ~n33287 ;
  assign n51290 = n51289 ^ n32533 ^ 1'b0 ;
  assign n51291 = n31722 ^ n17183 ^ 1'b0 ;
  assign n51292 = n17487 ^ n12461 ^ 1'b0 ;
  assign n51293 = n23364 & ~n51292 ;
  assign n51294 = n51293 ^ n15986 ^ 1'b0 ;
  assign n51295 = n51294 ^ n3588 ^ 1'b0 ;
  assign n51296 = n51295 ^ n50843 ^ n953 ;
  assign n51297 = n18928 & ~n29192 ;
  assign n51298 = n51297 ^ n23053 ^ 1'b0 ;
  assign n51299 = n51298 ^ n42308 ^ 1'b0 ;
  assign n51300 = n48505 ^ n23283 ^ 1'b0 ;
  assign n51301 = n49143 ^ n3985 ^ 1'b0 ;
  assign n51302 = n12554 | n32009 ;
  assign n51303 = n51302 ^ n8655 ^ 1'b0 ;
  assign n51304 = n8988 ^ n6845 ^ 1'b0 ;
  assign n51305 = n51304 ^ n24168 ^ n65 ;
  assign n51308 = n45384 ^ n23900 ^ n3782 ;
  assign n51309 = ( n4796 & ~n40209 ) | ( n4796 & n51308 ) | ( ~n40209 & n51308 ) ;
  assign n51306 = n44613 ^ n14453 ^ 1'b0 ;
  assign n51307 = n27361 | n51306 ;
  assign n51310 = n51309 ^ n51307 ^ 1'b0 ;
  assign n51311 = ~n28683 & n49695 ;
  assign n51312 = n51311 ^ n13356 ^ 1'b0 ;
  assign n51313 = n31772 ^ n27003 ^ 1'b0 ;
  assign n51314 = n4041 & ~n9813 ;
  assign n51315 = ( n99 & n1395 ) | ( n99 & ~n3890 ) | ( n1395 & ~n3890 ) ;
  assign n51316 = n50980 & ~n51315 ;
  assign n51317 = n51316 ^ n18150 ^ 1'b0 ;
  assign n51318 = n10217 & ~n23354 ;
  assign n51319 = n27159 & n51318 ;
  assign n51320 = n19357 ^ n5276 ^ 1'b0 ;
  assign n51321 = n5872 ^ n3105 ^ 1'b0 ;
  assign n51322 = ~n26669 & n41502 ;
  assign n51323 = n51321 | n51322 ;
  assign n51324 = n2662 & n46072 ;
  assign n51325 = n177 & n51324 ;
  assign n51326 = n14009 ^ n7418 ^ 1'b0 ;
  assign n51327 = n37178 & n51326 ;
  assign n51328 = n12560 ^ n9580 ^ n7106 ;
  assign n51329 = n51328 ^ n6135 ^ 1'b0 ;
  assign n51330 = n51329 ^ n30832 ^ 1'b0 ;
  assign n51331 = n51087 ^ n23567 ^ 1'b0 ;
  assign n51332 = n51331 ^ n42462 ^ n41525 ;
  assign n51333 = n39937 ^ n5120 ^ 1'b0 ;
  assign n51334 = n1200 & n51333 ;
  assign n51335 = ~n9323 & n43793 ;
  assign n51336 = n51335 ^ n29265 ^ 1'b0 ;
  assign n51337 = ( ~n26805 & n51334 ) | ( ~n26805 & n51336 ) | ( n51334 & n51336 ) ;
  assign n51338 = n9795 | n29485 ;
  assign n51339 = n23379 ^ n515 ^ 1'b0 ;
  assign n51340 = n43816 & ~n51339 ;
  assign n51341 = n3137 & n5016 ;
  assign n51342 = n51341 ^ n32216 ^ 1'b0 ;
  assign n51343 = n26261 & ~n51342 ;
  assign n51344 = ( n13821 & n15702 ) | ( n13821 & ~n21706 ) | ( n15702 & ~n21706 ) ;
  assign n51345 = n51344 ^ n14635 ^ 1'b0 ;
  assign n51346 = n48041 & n51345 ;
  assign n51347 = n44807 ^ n29109 ^ 1'b0 ;
  assign n51348 = ~n6181 & n15643 ;
  assign n51349 = n51348 ^ n11374 ^ 1'b0 ;
  assign n51350 = n10167 | n20557 ;
  assign n51351 = ~n5113 & n21848 ;
  assign n51352 = n51351 ^ n44436 ^ 1'b0 ;
  assign n51353 = n10118 ^ n5241 ^ 1'b0 ;
  assign n51354 = n50417 & ~n51353 ;
  assign n51355 = n51354 ^ n48566 ^ 1'b0 ;
  assign n51356 = n15560 ^ n13413 ^ 1'b0 ;
  assign n51357 = ~n1487 & n51356 ;
  assign n51358 = n51357 ^ n4826 ^ 1'b0 ;
  assign n51359 = n22275 & n51358 ;
  assign n51360 = n37511 ^ n24438 ^ 1'b0 ;
  assign n51361 = n46373 ^ n29270 ^ 1'b0 ;
  assign n51362 = n51360 & ~n51361 ;
  assign n51363 = n1186 & ~n42797 ;
  assign n51364 = n1036 & n33045 ;
  assign n51365 = ~n4812 & n51364 ;
  assign n51366 = n51365 ^ n40892 ^ 1'b0 ;
  assign n51367 = n51366 ^ n43788 ^ n10412 ;
  assign n51368 = n2180 | n40259 ;
  assign n51369 = n17331 | n42403 ;
  assign n51370 = n8713 & ~n51369 ;
  assign n51371 = n51370 ^ n6116 ^ 1'b0 ;
  assign n51372 = n7096 ^ n2281 ^ 1'b0 ;
  assign n51373 = n51371 & ~n51372 ;
  assign n51374 = ~n7737 & n36265 ;
  assign n51375 = n48708 & n51374 ;
  assign n51376 = n39321 | n51375 ;
  assign n51377 = n51376 ^ n17814 ^ 1'b0 ;
  assign n51378 = n7244 & ~n48009 ;
  assign n51379 = n10973 | n30334 ;
  assign n51380 = n51379 ^ n27452 ^ 1'b0 ;
  assign n51381 = n26567 ^ n12562 ^ 1'b0 ;
  assign n51382 = n4825 & n36312 ;
  assign n51383 = ~n17625 & n51382 ;
  assign n51384 = n51383 ^ n23148 ^ 1'b0 ;
  assign n51385 = n23776 & ~n51384 ;
  assign n51386 = ~n27656 & n51385 ;
  assign n51387 = n51386 ^ n47370 ^ 1'b0 ;
  assign n51388 = n18935 ^ n16067 ^ 1'b0 ;
  assign n51389 = n1877 & ~n2064 ;
  assign n51390 = n51389 ^ n27671 ^ 1'b0 ;
  assign n51391 = n51388 | n51390 ;
  assign n51392 = n3342 & ~n4390 ;
  assign n51393 = n51392 ^ n43191 ^ n41159 ;
  assign n51394 = n36547 | n41293 ;
  assign n51395 = n18522 | n51394 ;
  assign n51396 = ( n19834 & ~n50188 ) | ( n19834 & n51395 ) | ( ~n50188 & n51395 ) ;
  assign n51397 = n13905 ^ n5771 ^ 1'b0 ;
  assign n51398 = n3387 | n18083 ;
  assign n51399 = ~n5301 & n10479 ;
  assign n51400 = ~n6040 & n51399 ;
  assign n51401 = n17139 | n51400 ;
  assign n51402 = ( n51397 & n51398 ) | ( n51397 & ~n51401 ) | ( n51398 & ~n51401 ) ;
  assign n51403 = n40367 ^ n17910 ^ 1'b0 ;
  assign n51404 = ~n27652 & n36663 ;
  assign n51405 = n51404 ^ n8043 ^ 1'b0 ;
  assign n51406 = n51403 & ~n51405 ;
  assign n51408 = n1082 & ~n20087 ;
  assign n51409 = n16836 & n51408 ;
  assign n51407 = n57 & ~n50765 ;
  assign n51410 = n51409 ^ n51407 ^ 1'b0 ;
  assign n51411 = n4156 | n11459 ;
  assign n51414 = n4004 & n24667 ;
  assign n51412 = n13743 | n22906 ;
  assign n51413 = n7916 | n51412 ;
  assign n51415 = n51414 ^ n51413 ^ 1'b0 ;
  assign n51416 = n35328 ^ n7318 ^ n723 ;
  assign n51417 = n51415 & n51416 ;
  assign n51418 = n9224 ^ n8631 ^ 1'b0 ;
  assign n51419 = n22942 | n51418 ;
  assign n51420 = n28775 ^ n4789 ^ 1'b0 ;
  assign n51421 = n51419 | n51420 ;
  assign n51422 = n14385 ^ n5307 ^ 1'b0 ;
  assign n51423 = n1727 & ~n51422 ;
  assign n51424 = ( n14032 & n42897 ) | ( n14032 & ~n51423 ) | ( n42897 & ~n51423 ) ;
  assign n51425 = ( n129 & n17785 ) | ( n129 & ~n42084 ) | ( n17785 & ~n42084 ) ;
  assign n51426 = n2119 | n21021 ;
  assign n51428 = n3755 & n17301 ;
  assign n51429 = n51428 ^ n19553 ^ 1'b0 ;
  assign n51427 = ~n18688 & n43355 ;
  assign n51430 = n51429 ^ n51427 ^ 1'b0 ;
  assign n51431 = n7004 & n29024 ;
  assign n51432 = n23165 & n51431 ;
  assign n51433 = n5932 & n11777 ;
  assign n51434 = n8082 | n25067 ;
  assign n51435 = n45748 ^ n23193 ^ 1'b0 ;
  assign n51436 = ( n221 & n51434 ) | ( n221 & n51435 ) | ( n51434 & n51435 ) ;
  assign n51437 = n5256 | n51436 ;
  assign n51438 = ~n19429 & n41713 ;
  assign n51439 = n48887 ^ n20964 ^ 1'b0 ;
  assign n51440 = n19621 & ~n25402 ;
  assign n51441 = n51440 ^ n29943 ^ 1'b0 ;
  assign n51442 = ~n51439 & n51441 ;
  assign n51443 = ~n11306 & n49643 ;
  assign n51444 = ~n44 & n3428 ;
  assign n51445 = ~n51443 & n51444 ;
  assign n51446 = n2983 | n50150 ;
  assign n51447 = n31148 | n51446 ;
  assign n51448 = n11147 & n51447 ;
  assign n51449 = n51448 ^ n47503 ^ 1'b0 ;
  assign n51450 = ( n21434 & ~n23456 ) | ( n21434 & n32554 ) | ( ~n23456 & n32554 ) ;
  assign n51451 = n12791 & ~n35544 ;
  assign n51452 = n1315 & ~n40192 ;
  assign n51453 = n28714 ^ n12053 ^ 1'b0 ;
  assign n51454 = n6036 | n45664 ;
  assign n51455 = n34764 | n51454 ;
  assign n51456 = n11051 | n26586 ;
  assign n51457 = n19246 & ~n51456 ;
  assign n51458 = n51457 ^ n17708 ^ 1'b0 ;
  assign n51459 = ~n29451 & n51458 ;
  assign n51460 = n37588 | n51459 ;
  assign n51461 = n41436 ^ n9068 ^ 1'b0 ;
  assign n51462 = n51461 ^ n42198 ^ n16832 ;
  assign n51464 = n32124 ^ n15380 ^ 1'b0 ;
  assign n51465 = ~n4002 & n51464 ;
  assign n51463 = n13496 & ~n30313 ;
  assign n51466 = n51465 ^ n51463 ^ 1'b0 ;
  assign n51467 = n24885 ^ n48 ^ 1'b0 ;
  assign n51468 = n1206 | n51467 ;
  assign n51469 = n1348 & ~n31350 ;
  assign n51470 = n5164 & n51469 ;
  assign n51471 = n27534 ^ n7544 ^ 1'b0 ;
  assign n51472 = n1962 & n51471 ;
  assign n51473 = n21061 & n51472 ;
  assign n51474 = ~n1890 & n16389 ;
  assign n51475 = ( n4062 & ~n6493 ) | ( n4062 & n8179 ) | ( ~n6493 & n8179 ) ;
  assign n51476 = n50580 ^ n48958 ^ n22034 ;
  assign n51477 = ( ~n3855 & n5120 ) | ( ~n3855 & n10204 ) | ( n5120 & n10204 ) ;
  assign n51478 = n44041 & ~n51477 ;
  assign n51479 = ~n28828 & n51478 ;
  assign n51480 = n15061 & ~n23580 ;
  assign n51481 = n9336 & ~n48199 ;
  assign n51482 = n51481 ^ n7540 ^ n3167 ;
  assign n51483 = ~n2387 & n51482 ;
  assign n51484 = n8297 & ~n41166 ;
  assign n51485 = n14650 | n50076 ;
  assign n51486 = n51485 ^ n36802 ^ 1'b0 ;
  assign n51487 = n41789 & ~n51486 ;
  assign n51488 = n7500 | n30182 ;
  assign n51489 = ~n3141 & n6173 ;
  assign n51490 = n46431 | n51489 ;
  assign n51491 = n45652 ^ n12695 ^ 1'b0 ;
  assign n51492 = n7227 & n16196 ;
  assign n51493 = n51492 ^ n38080 ^ 1'b0 ;
  assign n51494 = n1099 & n24121 ;
  assign n51495 = n16021 | n47876 ;
  assign n51496 = n30756 ^ n5745 ^ 1'b0 ;
  assign n51497 = ~n938 & n51496 ;
  assign n51498 = n51497 ^ n7208 ^ 1'b0 ;
  assign n51499 = n2732 ^ n1518 ^ 1'b0 ;
  assign n51500 = n51499 ^ n15075 ^ n12476 ;
  assign n51501 = n49524 ^ n44361 ^ n30124 ;
  assign n51502 = n25569 ^ n7579 ^ 1'b0 ;
  assign n51503 = n10625 | n26845 ;
  assign n51504 = n926 | n15748 ;
  assign n51505 = n34665 & n51504 ;
  assign n51506 = n51505 ^ n3642 ^ 1'b0 ;
  assign n51507 = n38338 ^ n856 ^ 1'b0 ;
  assign n51508 = ( n2760 & n9778 ) | ( n2760 & ~n34903 ) | ( n9778 & ~n34903 ) ;
  assign n51509 = n13844 & n24283 ;
  assign n51510 = ~n37733 & n51509 ;
  assign n51511 = ~n2365 & n23974 ;
  assign n51512 = n14051 | n37931 ;
  assign n51513 = n20652 | n51512 ;
  assign n51514 = n8661 & ~n51513 ;
  assign n51515 = ~n32229 & n51514 ;
  assign n51516 = n26430 ^ n15310 ^ 1'b0 ;
  assign n51517 = n11120 & ~n22211 ;
  assign n51518 = ~n1893 & n51517 ;
  assign n51519 = n51518 ^ n21435 ^ n9162 ;
  assign n51520 = ( ~n10189 & n30124 ) | ( ~n10189 & n35139 ) | ( n30124 & n35139 ) ;
  assign n51521 = n51355 ^ n40784 ^ 1'b0 ;
  assign n51522 = n8985 ^ n3740 ^ 1'b0 ;
  assign n51523 = n33003 | n51522 ;
  assign n51524 = n14042 & n18520 ;
  assign n51525 = n11599 | n51524 ;
  assign n51526 = ~n15886 & n49933 ;
  assign n51527 = ~n51525 & n51526 ;
  assign n51528 = n5982 & n37559 ;
  assign n51530 = ~n427 & n32958 ;
  assign n51531 = n51530 ^ n31799 ^ 1'b0 ;
  assign n51529 = n1109 | n16017 ;
  assign n51532 = n51531 ^ n51529 ^ n18657 ;
  assign n51533 = n13559 ^ n7680 ^ 1'b0 ;
  assign n51534 = ~n13376 & n51533 ;
  assign n51535 = n51534 ^ n27345 ^ 1'b0 ;
  assign n51536 = n666 & n22698 ;
  assign n51537 = ~n16261 & n51536 ;
  assign n51538 = n51537 ^ n9592 ^ 1'b0 ;
  assign n51543 = n22726 ^ n12519 ^ 1'b0 ;
  assign n51539 = n44103 ^ n17916 ^ 1'b0 ;
  assign n51540 = n39148 & n40749 ;
  assign n51541 = ~n51539 & n51540 ;
  assign n51542 = n3416 & ~n51541 ;
  assign n51544 = n51543 ^ n51542 ^ 1'b0 ;
  assign n51545 = n39457 ^ n29467 ^ 1'b0 ;
  assign n51546 = ~n38451 & n51545 ;
  assign n51547 = n299 & ~n1045 ;
  assign n51548 = n39329 ^ n10832 ^ n28 ;
  assign n51549 = n11875 ^ n9400 ^ n4471 ;
  assign n51550 = n51549 ^ n7404 ^ 1'b0 ;
  assign n51551 = n51548 & n51550 ;
  assign n51552 = ( n10919 & ~n17336 ) | ( n10919 & n36656 ) | ( ~n17336 & n36656 ) ;
  assign n51553 = n32079 ^ n13277 ^ 1'b0 ;
  assign n51554 = n22561 ^ n21913 ^ 1'b0 ;
  assign n51555 = n20470 ^ n13516 ^ 1'b0 ;
  assign n51556 = n40954 | n51555 ;
  assign n51557 = n30248 & n39336 ;
  assign n51558 = n51556 & n51557 ;
  assign n51559 = ~n5727 & n17996 ;
  assign n51560 = n22465 & ~n42996 ;
  assign n51561 = n51559 | n51560 ;
  assign n51562 = ~n10017 & n34314 ;
  assign n51567 = n4480 & n5466 ;
  assign n51568 = n51567 ^ n4100 ^ 1'b0 ;
  assign n51563 = ( ~n3175 & n4686 ) | ( ~n3175 & n23156 ) | ( n4686 & n23156 ) ;
  assign n51564 = ~n22037 & n51563 ;
  assign n51565 = ~n43390 & n51564 ;
  assign n51566 = n51565 ^ n18254 ^ 1'b0 ;
  assign n51569 = n51568 ^ n51566 ^ n37374 ;
  assign n51570 = n3876 & ~n51569 ;
  assign n51571 = n51570 ^ n7144 ^ 1'b0 ;
  assign n51572 = n18110 & ~n25321 ;
  assign n51573 = n51572 ^ n30908 ^ n498 ;
  assign n51577 = n9857 ^ n9060 ^ 1'b0 ;
  assign n51574 = ~n773 & n11503 ;
  assign n51575 = n51574 ^ n9098 ^ 1'b0 ;
  assign n51576 = ~n12396 & n51575 ;
  assign n51578 = n51577 ^ n51576 ^ 1'b0 ;
  assign n51579 = n51578 ^ n42711 ^ n475 ;
  assign n51580 = n19294 & n43391 ;
  assign n51581 = n2377 & n51580 ;
  assign n51582 = n51581 ^ n6850 ^ 1'b0 ;
  assign n51583 = ~n21667 & n22777 ;
  assign n51584 = n28359 & n51583 ;
  assign n51585 = n51584 ^ n18872 ^ 1'b0 ;
  assign n51586 = n25452 & n51585 ;
  assign n51587 = n47746 ^ n7586 ^ 1'b0 ;
  assign n51588 = n9887 & ~n51587 ;
  assign n51589 = n10950 ^ n8614 ^ 1'b0 ;
  assign n51590 = ~n42752 & n51589 ;
  assign n51591 = n1940 & ~n13197 ;
  assign n51592 = n51591 ^ n4253 ^ 1'b0 ;
  assign n51593 = n30107 | n51592 ;
  assign n51595 = n4416 & n46755 ;
  assign n51594 = n16559 & ~n20799 ;
  assign n51596 = n51595 ^ n51594 ^ 1'b0 ;
  assign n51597 = n51596 ^ n39124 ^ n22648 ;
  assign n51598 = n8440 | n14281 ;
  assign n51599 = n25000 & n51598 ;
  assign n51600 = n13524 ^ n4518 ^ 1'b0 ;
  assign n51601 = ~n25437 & n51600 ;
  assign n51602 = n5595 & ~n26192 ;
  assign n51603 = ~n51397 & n51602 ;
  assign n51604 = n14766 & ~n25786 ;
  assign n51605 = n11523 | n24302 ;
  assign n51606 = n2979 | n51605 ;
  assign n51607 = n51606 ^ n12713 ^ 1'b0 ;
  assign n51608 = n51604 & n51607 ;
  assign n51609 = n15037 ^ n10265 ^ 1'b0 ;
  assign n51610 = ~n13969 & n15420 ;
  assign n51611 = ~n51609 & n51610 ;
  assign n51612 = n837 | n1437 ;
  assign n51613 = n47640 ^ n12828 ^ 1'b0 ;
  assign n51614 = n51612 | n51613 ;
  assign n51615 = ~n922 & n51614 ;
  assign n51616 = ~n11325 & n21244 ;
  assign n51617 = ~n51615 & n51616 ;
  assign n51619 = n41789 ^ n22104 ^ n13057 ;
  assign n51618 = n24266 & n29525 ;
  assign n51620 = n51619 ^ n51618 ^ 1'b0 ;
  assign n51621 = n13429 & n18639 ;
  assign n51622 = ( n132 & n13546 ) | ( n132 & n16187 ) | ( n13546 & n16187 ) ;
  assign n51623 = ( n12493 & n14386 ) | ( n12493 & ~n33093 ) | ( n14386 & ~n33093 ) ;
  assign n51624 = n5933 | n25072 ;
  assign n51625 = ~n18387 & n28145 ;
  assign n51626 = n29844 & n51625 ;
  assign n51627 = n38421 | n39711 ;
  assign n51628 = n51584 & ~n51627 ;
  assign n51629 = n10976 & ~n11210 ;
  assign n51630 = ~n31344 & n51629 ;
  assign n51631 = n51630 ^ n2997 ^ 1'b0 ;
  assign n51632 = n2040 | n7189 ;
  assign n51633 = n13916 | n37991 ;
  assign n51634 = n1439 & n51633 ;
  assign n51635 = n8515 | n28246 ;
  assign n51636 = n37163 ^ n9821 ^ 1'b0 ;
  assign n51637 = n20759 | n51636 ;
  assign n51638 = ~n4948 & n14912 ;
  assign n51639 = n24672 & n48633 ;
  assign n51640 = n11311 | n25318 ;
  assign n51641 = n9418 | n51640 ;
  assign n51642 = n42500 ^ n10085 ^ 1'b0 ;
  assign n51643 = n51641 & ~n51642 ;
  assign n51644 = n22426 | n51643 ;
  assign n51645 = n51436 ^ n44097 ^ 1'b0 ;
  assign n51646 = n12037 & ~n51645 ;
  assign n51647 = n569 & n22223 ;
  assign n51648 = ~n14799 & n48053 ;
  assign n51649 = n9282 & n51648 ;
  assign n51650 = n51649 ^ n6901 ^ 1'b0 ;
  assign n51651 = n15609 & n28568 ;
  assign n51652 = ( n1395 & n1888 ) | ( n1395 & n5086 ) | ( n1888 & n5086 ) ;
  assign n51653 = n51652 ^ n51210 ^ 1'b0 ;
  assign n51654 = ~n890 & n12058 ;
  assign n51655 = n51654 ^ n15203 ^ 1'b0 ;
  assign n51656 = n897 & ~n51655 ;
  assign n51657 = ~n1511 & n28761 ;
  assign n51658 = n51657 ^ n40748 ^ 1'b0 ;
  assign n51659 = n20386 | n51658 ;
  assign n51660 = n17070 ^ n5210 ^ 1'b0 ;
  assign n51661 = n6601 & n47004 ;
  assign n51662 = ~n51660 & n51661 ;
  assign n51663 = n5183 & n12159 ;
  assign n51664 = ~n14175 & n51663 ;
  assign n51665 = n51329 ^ n5338 ^ 1'b0 ;
  assign n51666 = n24797 ^ n23452 ^ 1'b0 ;
  assign n51667 = n29821 ^ n11902 ^ n7286 ;
  assign n51668 = n3135 | n4187 ;
  assign n51669 = n51668 ^ n2686 ^ 1'b0 ;
  assign n51670 = n7836 ^ n2311 ^ 1'b0 ;
  assign n51671 = n51670 ^ n28090 ^ 1'b0 ;
  assign n51672 = n7740 & ~n51671 ;
  assign n51673 = n35571 | n51672 ;
  assign n51674 = n11867 & n14564 ;
  assign n51675 = n51674 ^ n23254 ^ 1'b0 ;
  assign n51676 = ( n23832 & n42591 ) | ( n23832 & ~n51675 ) | ( n42591 & ~n51675 ) ;
  assign n51677 = n42686 ^ n28662 ^ 1'b0 ;
  assign n51678 = ( n14983 & ~n39618 ) | ( n14983 & n51677 ) | ( ~n39618 & n51677 ) ;
  assign n51679 = ( n6856 & ~n9103 ) | ( n6856 & n17236 ) | ( ~n9103 & n17236 ) ;
  assign n51680 = n38841 | n51679 ;
  assign n51681 = n17405 | n51680 ;
  assign n51682 = ~n26349 & n51681 ;
  assign n51683 = n16414 & n51682 ;
  assign n51684 = n45917 ^ n8907 ^ 1'b0 ;
  assign n51685 = n19409 | n44251 ;
  assign n51686 = n6462 | n51685 ;
  assign n51687 = ~n15940 & n22357 ;
  assign n51688 = n51687 ^ n22410 ^ 1'b0 ;
  assign n51689 = n33643 ^ n21778 ^ 1'b0 ;
  assign n51690 = n17836 ^ n9105 ^ n4393 ;
  assign n51691 = n11549 | n20786 ;
  assign n51692 = n29395 & n32428 ;
  assign n51693 = ( n51690 & ~n51691 ) | ( n51690 & n51692 ) | ( ~n51691 & n51692 ) ;
  assign n51694 = n39049 ^ n29605 ^ 1'b0 ;
  assign n51695 = n30060 | n30431 ;
  assign n51696 = n51695 ^ n1800 ^ 1'b0 ;
  assign n51697 = n20320 ^ n10999 ^ 1'b0 ;
  assign n51698 = n11137 & n51697 ;
  assign n51699 = n50090 ^ n12291 ^ x2 ;
  assign n51700 = ( n3137 & n4226 ) | ( n3137 & n34513 ) | ( n4226 & n34513 ) ;
  assign n51701 = n51700 ^ n6368 ^ n5459 ;
  assign n51702 = n51701 ^ n18324 ^ 1'b0 ;
  assign n51703 = n26759 ^ n9357 ^ 1'b0 ;
  assign n51704 = n30597 | n45172 ;
  assign n51705 = n36251 & ~n51704 ;
  assign n51706 = n26717 & n36424 ;
  assign n51707 = n51706 ^ n3973 ^ 1'b0 ;
  assign n51708 = ~n20473 & n22847 ;
  assign n51709 = n51708 ^ n38105 ^ 1'b0 ;
  assign n51710 = n13632 | n15972 ;
  assign n51711 = n51710 ^ n28025 ^ 1'b0 ;
  assign n51712 = n39551 | n51711 ;
  assign n51713 = n41918 & ~n51712 ;
  assign n51714 = n3263 & ~n51713 ;
  assign n51715 = n44208 ^ n9156 ^ 1'b0 ;
  assign n51716 = n51714 & n51715 ;
  assign n51717 = n51716 ^ n17185 ^ 1'b0 ;
  assign n51718 = n32892 ^ n17865 ^ 1'b0 ;
  assign n51719 = n14443 | n51718 ;
  assign n51720 = n51719 ^ n31406 ^ 1'b0 ;
  assign n51721 = ( n14964 & n43753 ) | ( n14964 & n51720 ) | ( n43753 & n51720 ) ;
  assign n51722 = n28540 ^ n13372 ^ 1'b0 ;
  assign n51723 = n30192 & n51722 ;
  assign n51724 = ~n5289 & n29373 ;
  assign n51725 = n51724 ^ n22660 ^ 1'b0 ;
  assign n51726 = n24488 & n51725 ;
  assign n51727 = ~n51723 & n51726 ;
  assign n51728 = n51727 ^ n21485 ^ n5143 ;
  assign n51730 = n3635 & n4533 ;
  assign n51731 = ~n4533 & n51730 ;
  assign n51732 = ( n890 & n6457 ) | ( n890 & ~n20199 ) | ( n6457 & ~n20199 ) ;
  assign n51733 = n3144 & n51732 ;
  assign n51734 = n51731 & n51733 ;
  assign n51735 = ( n25585 & ~n28002 ) | ( n25585 & n51734 ) | ( ~n28002 & n51734 ) ;
  assign n51736 = n16971 & ~n51735 ;
  assign n51737 = n51736 ^ n12949 ^ 1'b0 ;
  assign n51729 = n3284 ^ n177 ^ 1'b0 ;
  assign n51738 = n51737 ^ n51729 ^ n16349 ;
  assign n51739 = n8458 | n25506 ;
  assign n51740 = n18447 & ~n51739 ;
  assign n51741 = ~n43478 & n51740 ;
  assign n51742 = n8017 & n31854 ;
  assign n51743 = n16906 & n43772 ;
  assign n51745 = n2186 & ~n24644 ;
  assign n51746 = ~n7076 & n51745 ;
  assign n51744 = ~n13567 & n19055 ;
  assign n51747 = n51746 ^ n51744 ^ 1'b0 ;
  assign n51748 = n47615 ^ n8338 ^ 1'b0 ;
  assign n51749 = n16067 & ~n47001 ;
  assign n51750 = n4845 | n18440 ;
  assign n51751 = n45015 ^ n37614 ^ 1'b0 ;
  assign n51752 = ( n35659 & n51750 ) | ( n35659 & n51751 ) | ( n51750 & n51751 ) ;
  assign n51753 = ~n3254 & n30553 ;
  assign n51754 = n51753 ^ n15449 ^ n14769 ;
  assign n51755 = n926 | n9246 ;
  assign n51756 = n51755 ^ n25472 ^ 1'b0 ;
  assign n51757 = n31263 & ~n51756 ;
  assign n51758 = n17766 ^ n5844 ^ 1'b0 ;
  assign n51759 = n51757 & n51758 ;
  assign n51760 = n22640 & n34327 ;
  assign n51761 = n14624 & n51760 ;
  assign n51762 = n7864 & ~n23166 ;
  assign n51763 = n11459 ^ n8753 ^ 1'b0 ;
  assign n51764 = n39432 & ~n47740 ;
  assign n51765 = n51764 ^ n23954 ^ 1'b0 ;
  assign n51766 = n5311 & n51140 ;
  assign n51767 = n44408 ^ n4488 ^ 1'b0 ;
  assign n51768 = n5571 | n10974 ;
  assign n51769 = n51768 ^ n30712 ^ 1'b0 ;
  assign n51770 = n13866 | n51769 ;
  assign n51771 = ( n13721 & n33043 ) | ( n13721 & ~n51770 ) | ( n33043 & ~n51770 ) ;
  assign n51772 = n2980 & ~n13931 ;
  assign n51773 = n13207 & n51772 ;
  assign n51774 = n51773 ^ n8055 ^ 1'b0 ;
  assign n51775 = n1773 & ~n42420 ;
  assign n51776 = n51775 ^ n27069 ^ 1'b0 ;
  assign n51777 = n10950 | n45297 ;
  assign n51778 = ~n2449 & n51777 ;
  assign n51779 = n51778 ^ n42458 ^ 1'b0 ;
  assign n51780 = n49745 ^ n6167 ^ 1'b0 ;
  assign n51781 = n25769 ^ n6561 ^ n1686 ;
  assign n51782 = ~n51780 & n51781 ;
  assign n51783 = n6673 & ~n10212 ;
  assign n51784 = n8480 | n39929 ;
  assign n51785 = ( ~n15287 & n15638 ) | ( ~n15287 & n22426 ) | ( n15638 & n22426 ) ;
  assign n51786 = n24235 & n25990 ;
  assign n51787 = n51786 ^ n11069 ^ 1'b0 ;
  assign n51788 = ~n5898 & n15821 ;
  assign n51789 = n4093 & n10247 ;
  assign n51790 = n2734 & n51789 ;
  assign n51791 = n33243 & n34001 ;
  assign n51792 = n51791 ^ n37354 ^ 1'b0 ;
  assign n51793 = n14974 ^ n5895 ^ 1'b0 ;
  assign n51794 = n51792 & n51793 ;
  assign n51795 = n4967 & ~n5578 ;
  assign n51796 = n8654 & n51795 ;
  assign n51797 = n35235 ^ n11736 ^ 1'b0 ;
  assign n51798 = n18482 ^ n9862 ^ 1'b0 ;
  assign n51799 = n34671 & ~n51798 ;
  assign n51800 = ~n8703 & n51799 ;
  assign n51801 = n50268 ^ n6098 ^ 1'b0 ;
  assign n51802 = n35907 ^ n16684 ^ n4750 ;
  assign n51803 = n30297 & ~n33881 ;
  assign n51804 = n15861 & ~n24807 ;
  assign n51805 = n5047 & ~n8452 ;
  assign n51806 = n31495 & n51805 ;
  assign n51807 = n17151 | n22243 ;
  assign n51808 = n51806 & ~n51807 ;
  assign n51809 = n7197 & ~n19097 ;
  assign n51810 = n14706 & n25457 ;
  assign n51811 = n4102 & n51810 ;
  assign n51812 = ~n1642 & n4421 ;
  assign n51813 = n51812 ^ n12995 ^ 1'b0 ;
  assign n51814 = n14719 | n48475 ;
  assign n51815 = n51814 ^ n26226 ^ 1'b0 ;
  assign n51816 = n12551 & n51815 ;
  assign n51817 = n31097 & ~n50160 ;
  assign n51818 = ~n11560 & n31249 ;
  assign n51819 = n23207 & n51818 ;
  assign n51820 = ( n16948 & ~n43413 ) | ( n16948 & n51819 ) | ( ~n43413 & n51819 ) ;
  assign n51821 = n11178 & ~n14118 ;
  assign n51822 = n51821 ^ n10420 ^ 1'b0 ;
  assign n51823 = n3415 & n51822 ;
  assign n51824 = ( n5713 & n31861 ) | ( n5713 & ~n51823 ) | ( n31861 & ~n51823 ) ;
  assign n51825 = n51824 ^ n4060 ^ 1'b0 ;
  assign n51826 = n10849 & ~n26643 ;
  assign n51827 = n51826 ^ n20628 ^ 1'b0 ;
  assign n51828 = n30636 & ~n51827 ;
  assign n51829 = n24902 ^ n3506 ^ 1'b0 ;
  assign n51830 = n5376 & ~n51829 ;
  assign n51831 = n40665 & n51830 ;
  assign n51832 = n5339 ^ n741 ^ 1'b0 ;
  assign n51833 = n40648 ^ n2126 ^ n1177 ;
  assign n51834 = n10077 | n32691 ;
  assign n51835 = n983 & n51834 ;
  assign n51836 = n36377 ^ n6231 ^ 1'b0 ;
  assign n51837 = n11956 & ~n51836 ;
  assign n51838 = n195 & ~n41190 ;
  assign n51839 = ~n10543 & n51838 ;
  assign n51840 = n51839 ^ n18330 ^ 1'b0 ;
  assign n51841 = n1295 & n51840 ;
  assign n51842 = ( n25678 & n39231 ) | ( n25678 & ~n51841 ) | ( n39231 & ~n51841 ) ;
  assign n51843 = n14375 & n27305 ;
  assign n51844 = ~n10893 & n51843 ;
  assign n51845 = n51844 ^ n36626 ^ n29217 ;
  assign n51846 = n6523 & n51845 ;
  assign n51847 = n51846 ^ n16092 ^ 1'b0 ;
  assign n51848 = n22335 | n29314 ;
  assign n51849 = n15248 & n15933 ;
  assign n51850 = ( n11962 & ~n15630 ) | ( n11962 & n25549 ) | ( ~n15630 & n25549 ) ;
  assign n51851 = n5182 & ~n33711 ;
  assign n51852 = ~n26809 & n51851 ;
  assign n51853 = ( ~n1426 & n4226 ) | ( ~n1426 & n51852 ) | ( n4226 & n51852 ) ;
  assign n51855 = n26210 ^ n7906 ^ 1'b0 ;
  assign n51856 = n6173 & n51855 ;
  assign n51854 = ~n4847 & n5904 ;
  assign n51857 = n51856 ^ n51854 ^ 1'b0 ;
  assign n51858 = ( n21985 & ~n50640 ) | ( n21985 & n51857 ) | ( ~n50640 & n51857 ) ;
  assign n51861 = n1482 & n1974 ;
  assign n51859 = n35658 ^ n16382 ^ 1'b0 ;
  assign n51860 = ~n18458 & n51859 ;
  assign n51862 = n51861 ^ n51860 ^ n2271 ;
  assign n51863 = n43350 & ~n51862 ;
  assign n51864 = ~n39096 & n51863 ;
  assign n51865 = n48083 ^ n28255 ^ 1'b0 ;
  assign n51866 = n46107 & ~n51865 ;
  assign n51867 = n26887 | n45965 ;
  assign n51868 = n51867 ^ n10491 ^ 1'b0 ;
  assign n51869 = n2735 & n34467 ;
  assign n51870 = n15142 ^ n928 ^ 1'b0 ;
  assign n51871 = n51869 & n51870 ;
  assign n51872 = n35125 ^ n22164 ^ 1'b0 ;
  assign n51873 = n43992 | n51872 ;
  assign n51874 = n8091 & ~n10393 ;
  assign n51875 = n51874 ^ n30898 ^ n29474 ;
  assign n51876 = n1443 ^ n664 ^ 1'b0 ;
  assign n51877 = n1000 & n51876 ;
  assign n51878 = n23563 | n51877 ;
  assign n51879 = ( n31443 & n35350 ) | ( n31443 & ~n51878 ) | ( n35350 & ~n51878 ) ;
  assign n51880 = n10794 & ~n51879 ;
  assign n51881 = n38651 ^ n26179 ^ n2874 ;
  assign n51882 = n51881 ^ n30723 ^ 1'b0 ;
  assign n51883 = n4906 | n19747 ;
  assign n51884 = ( n15047 & n32921 ) | ( n15047 & n51883 ) | ( n32921 & n51883 ) ;
  assign n51885 = n51884 ^ n19161 ^ 1'b0 ;
  assign n51886 = n11000 | n51885 ;
  assign n51887 = n42093 ^ n23513 ^ 1'b0 ;
  assign n51888 = n9959 ^ n9773 ^ n135 ;
  assign n51889 = ( n4580 & n8351 ) | ( n4580 & ~n21202 ) | ( n8351 & ~n21202 ) ;
  assign n51890 = n25385 ^ n11052 ^ 1'b0 ;
  assign n51891 = n4039 & n48735 ;
  assign n51892 = ~n26584 & n51891 ;
  assign n51895 = n30406 ^ n6282 ^ 1'b0 ;
  assign n51893 = ( n867 & n5882 ) | ( n867 & ~n43436 ) | ( n5882 & ~n43436 ) ;
  assign n51894 = n5089 & ~n51893 ;
  assign n51896 = n51895 ^ n51894 ^ 1'b0 ;
  assign n51897 = n4275 & n11033 ;
  assign n51898 = n51897 ^ n39742 ^ 1'b0 ;
  assign n51899 = n46699 ^ n694 ^ 1'b0 ;
  assign n51900 = n26773 & n51899 ;
  assign n51901 = n927 | n15314 ;
  assign n51902 = ( n15009 & ~n34377 ) | ( n15009 & n40390 ) | ( ~n34377 & n40390 ) ;
  assign n51903 = n51901 | n51902 ;
  assign n51904 = n4047 & n20446 ;
  assign n51905 = n51904 ^ n43757 ^ n14593 ;
  assign n51906 = n1412 | n15403 ;
  assign n51907 = n42161 ^ n34772 ^ 1'b0 ;
  assign n51908 = n5915 & n11596 ;
  assign n51909 = ~n2928 & n10769 ;
  assign n51910 = n2983 | n51909 ;
  assign n51911 = n51908 | n51910 ;
  assign n51912 = n1818 | n6027 ;
  assign n51913 = n6965 & ~n51912 ;
  assign n51914 = n51913 ^ n1180 ^ 1'b0 ;
  assign n51915 = ~n39443 & n51914 ;
  assign n51916 = n51915 ^ n33979 ^ 1'b0 ;
  assign n51917 = n51911 & n51916 ;
  assign n51918 = ~n8211 & n18782 ;
  assign n51919 = n1871 | n25203 ;
  assign n51920 = n51918 & ~n51919 ;
  assign n51921 = n16430 & ~n22493 ;
  assign n51922 = n21190 | n42717 ;
  assign n51923 = ( ~n28810 & n51921 ) | ( ~n28810 & n51922 ) | ( n51921 & n51922 ) ;
  assign n51924 = n28199 & n51923 ;
  assign n51926 = n41588 ^ n4703 ^ 1'b0 ;
  assign n51925 = ~n10886 & n18904 ;
  assign n51927 = n51926 ^ n51925 ^ 1'b0 ;
  assign n51928 = n44751 ^ n10111 ^ n4743 ;
  assign n51929 = n19800 & n51928 ;
  assign n51930 = n30283 & n51929 ;
  assign n51931 = n21754 | n27000 ;
  assign n51932 = n51931 ^ n36386 ^ 1'b0 ;
  assign n51933 = n23156 ^ n2974 ^ 1'b0 ;
  assign n51934 = n1443 & ~n51933 ;
  assign n51935 = ~n1986 & n51934 ;
  assign n51936 = ~n51932 & n51935 ;
  assign n51937 = n14651 | n51936 ;
  assign n51938 = n29240 | n37554 ;
  assign n51939 = n51938 ^ n28607 ^ 1'b0 ;
  assign n51940 = n51939 ^ n24968 ^ 1'b0 ;
  assign n51941 = ~n11266 & n51940 ;
  assign n51944 = n45163 ^ n33501 ^ n12037 ;
  assign n51945 = n51944 ^ n4838 ^ 1'b0 ;
  assign n51946 = n1932 & n51945 ;
  assign n51942 = n7240 ^ n2671 ^ 1'b0 ;
  assign n51943 = n51942 ^ n32581 ^ n31644 ;
  assign n51947 = n51946 ^ n51943 ^ n1425 ;
  assign n51948 = ~n28430 & n51947 ;
  assign n51949 = n45333 ^ n1762 ^ 1'b0 ;
  assign n51950 = n36738 & n51949 ;
  assign n51951 = ( n11854 & ~n25452 ) | ( n11854 & n39594 ) | ( ~n25452 & n39594 ) ;
  assign n51952 = ~n9033 & n32831 ;
  assign n51953 = n4231 & ~n28796 ;
  assign n51954 = ~n8625 & n51953 ;
  assign n51955 = n44326 ^ n7525 ^ 1'b0 ;
  assign n51956 = n31249 & ~n51955 ;
  assign n51957 = n20605 ^ n8338 ^ 1'b0 ;
  assign n51958 = n5055 & n51957 ;
  assign n51959 = n4430 & ~n25045 ;
  assign n51963 = n44047 ^ n16506 ^ 1'b0 ;
  assign n51960 = ~n11888 & n14416 ;
  assign n51961 = n21075 & n51960 ;
  assign n51962 = n51392 | n51961 ;
  assign n51964 = n51963 ^ n51962 ^ 1'b0 ;
  assign n51965 = n48199 ^ n23716 ^ 1'b0 ;
  assign n51966 = n241 & n27379 ;
  assign n51967 = n51966 ^ n12317 ^ 1'b0 ;
  assign n51968 = ~n14493 & n40632 ;
  assign n51969 = n51968 ^ n31505 ^ 1'b0 ;
  assign n51970 = n51969 ^ n9563 ^ n475 ;
  assign n51971 = n19608 & n21385 ;
  assign n51972 = n51971 ^ n13060 ^ 1'b0 ;
  assign n51973 = n51970 & ~n51972 ;
  assign n51974 = n12051 | n20589 ;
  assign n51975 = n49053 | n51974 ;
  assign n51976 = n18577 ^ n18575 ^ 1'b0 ;
  assign n51977 = n29776 & ~n51976 ;
  assign n51978 = n1155 & n4053 ;
  assign n51979 = ~n51977 & n51978 ;
  assign n51980 = n39049 & n39654 ;
  assign n51981 = n51980 ^ n45221 ^ 1'b0 ;
  assign n51982 = ~n8504 & n51981 ;
  assign n51983 = n45930 & n51982 ;
  assign n51984 = ~n14180 & n36838 ;
  assign n51985 = ~n1770 & n51984 ;
  assign n51986 = n8991 ^ n7751 ^ 1'b0 ;
  assign n51987 = n14719 ^ n1991 ^ 1'b0 ;
  assign n51988 = ~n51986 & n51987 ;
  assign n51989 = n29632 ^ n401 ^ 1'b0 ;
  assign n51990 = n3843 & n51989 ;
  assign n51991 = n2758 & n13307 ;
  assign n51992 = n20955 ^ n9649 ^ n6566 ;
  assign n51993 = ( ~n33504 & n33530 ) | ( ~n33504 & n45916 ) | ( n33530 & n45916 ) ;
  assign n51994 = n26235 ^ n299 ^ 1'b0 ;
  assign n51995 = n40192 ^ n25041 ^ n10452 ;
  assign n51996 = n51995 ^ n27385 ^ 1'b0 ;
  assign n51997 = n15800 & n43918 ;
  assign n51998 = n6700 & n51997 ;
  assign n52002 = n28841 & n44502 ;
  assign n52003 = n16378 & n52002 ;
  assign n51999 = n12042 & n41695 ;
  assign n52000 = n51999 ^ n9179 ^ 1'b0 ;
  assign n52001 = n52000 ^ n30555 ^ n2958 ;
  assign n52004 = n52003 ^ n52001 ^ n5203 ;
  assign n52006 = n21745 & ~n23143 ;
  assign n52005 = n34314 & n45005 ;
  assign n52007 = n52006 ^ n52005 ^ n18380 ;
  assign n52008 = n16173 & n45916 ;
  assign n52009 = n49765 ^ n1712 ^ 1'b0 ;
  assign n52010 = n9226 | n52009 ;
  assign n52011 = n6890 & n20056 ;
  assign n52012 = n15940 & n52011 ;
  assign n52013 = n52012 ^ n46726 ^ 1'b0 ;
  assign n52017 = n16546 | n30101 ;
  assign n52014 = n41965 ^ n14609 ^ 1'b0 ;
  assign n52015 = n52014 ^ n33432 ^ 1'b0 ;
  assign n52016 = ( ~n23 & n1800 ) | ( ~n23 & n52015 ) | ( n1800 & n52015 ) ;
  assign n52018 = n52017 ^ n52016 ^ 1'b0 ;
  assign n52019 = n28680 ^ n26165 ^ 1'b0 ;
  assign n52020 = ( n18715 & ~n27064 ) | ( n18715 & n37370 ) | ( ~n27064 & n37370 ) ;
  assign n52021 = n35982 ^ n33137 ^ 1'b0 ;
  assign n52022 = n52021 ^ n49982 ^ n18403 ;
  assign n52023 = n16710 & n29022 ;
  assign n52024 = n19904 | n52023 ;
  assign n52025 = n41750 & ~n52024 ;
  assign n52026 = n35376 & n52023 ;
  assign n52027 = n42166 ^ n30080 ^ 1'b0 ;
  assign n52028 = n12163 & ~n52027 ;
  assign n52029 = ~n2747 & n35438 ;
  assign n52030 = n10438 & n52029 ;
  assign n52031 = ~n3367 & n29857 ;
  assign n52032 = n28257 ^ n24938 ^ n3426 ;
  assign n52033 = n30188 ^ n17590 ^ 1'b0 ;
  assign n52043 = n9929 | n32303 ;
  assign n52034 = n7655 | n15984 ;
  assign n52035 = n8576 | n52034 ;
  assign n52036 = ~n5311 & n12639 ;
  assign n52037 = n52036 ^ n24601 ^ 1'b0 ;
  assign n52038 = n52037 ^ n28939 ^ n7398 ;
  assign n52039 = ~n29699 & n52038 ;
  assign n52040 = n52039 ^ n12677 ^ 1'b0 ;
  assign n52041 = ( ~n13876 & n52035 ) | ( ~n13876 & n52040 ) | ( n52035 & n52040 ) ;
  assign n52042 = n2067 | n52041 ;
  assign n52044 = n52043 ^ n52042 ^ 1'b0 ;
  assign n52045 = n26451 ^ n22588 ^ 1'b0 ;
  assign n52046 = n38915 & n52045 ;
  assign n52047 = n342 | n46122 ;
  assign n52048 = n19392 & ~n52047 ;
  assign n52049 = n21139 ^ n8962 ^ 1'b0 ;
  assign n52050 = ~n18306 & n52049 ;
  assign n52051 = n19190 | n28511 ;
  assign n52052 = n52050 | n52051 ;
  assign n52053 = n10586 & n52052 ;
  assign n52054 = n52053 ^ n6271 ^ 1'b0 ;
  assign n52055 = n469 & ~n23308 ;
  assign n52056 = n21174 | n52055 ;
  assign n52057 = n52056 ^ n44783 ^ 1'b0 ;
  assign n52058 = n37760 | n47069 ;
  assign n52059 = n52058 ^ n5469 ^ 1'b0 ;
  assign n52060 = n21355 ^ n8667 ^ n1289 ;
  assign n52061 = ( n7031 & n12503 ) | ( n7031 & n17836 ) | ( n12503 & n17836 ) ;
  assign n52062 = ( ~n3056 & n38454 ) | ( ~n3056 & n52061 ) | ( n38454 & n52061 ) ;
  assign n52063 = n134 | n10457 ;
  assign n52064 = n41522 & ~n52063 ;
  assign n52065 = n2347 & ~n25436 ;
  assign n52066 = n52065 ^ n48874 ^ 1'b0 ;
  assign n52067 = n7993 & ~n22909 ;
  assign n52068 = n52067 ^ n19170 ^ 1'b0 ;
  assign n52069 = n6625 ^ n4318 ^ n4215 ;
  assign n52070 = ( n2776 & ~n12077 ) | ( n2776 & n48717 ) | ( ~n12077 & n48717 ) ;
  assign n52071 = n9640 | n26720 ;
  assign n52072 = n19731 | n52071 ;
  assign n52073 = ~n17129 & n22925 ;
  assign n52074 = n10875 & n27863 ;
  assign n52075 = n46006 ^ n35162 ^ 1'b0 ;
  assign n52076 = n4239 & ~n20582 ;
  assign n52077 = n52075 & n52076 ;
  assign n52078 = n14775 & n46269 ;
  assign n52079 = n6085 | n18093 ;
  assign n52080 = n22879 & n31696 ;
  assign n52081 = n2094 & ~n24030 ;
  assign n52082 = n40914 & n52081 ;
  assign n52083 = n52082 ^ n47338 ^ 1'b0 ;
  assign n52084 = n12551 & n19685 ;
  assign n52085 = ~n20059 & n52084 ;
  assign n52086 = n29895 ^ n4657 ^ 1'b0 ;
  assign n52087 = n27314 & ~n30608 ;
  assign n52088 = n52087 ^ n14772 ^ 1'b0 ;
  assign n52089 = ~n9549 & n15075 ;
  assign n52090 = ~n8451 & n20845 ;
  assign n52091 = n29691 & ~n52090 ;
  assign n52092 = n15982 ^ n3698 ^ 1'b0 ;
  assign n52093 = n52091 & ~n52092 ;
  assign n52094 = n9199 & n18984 ;
  assign n52095 = n17308 & ~n22749 ;
  assign n52096 = ~n59 & n52095 ;
  assign n52097 = n3898 | n52096 ;
  assign n52098 = n52097 ^ n10321 ^ 1'b0 ;
  assign n52099 = n11862 & ~n14827 ;
  assign n52100 = n52099 ^ n1129 ^ 1'b0 ;
  assign n52101 = n52100 ^ n35329 ^ 1'b0 ;
  assign n52102 = n3027 & n16672 ;
  assign n52103 = n52102 ^ n30107 ^ 1'b0 ;
  assign n52105 = n9601 ^ x3 ^ 1'b0 ;
  assign n52106 = n17888 | n52105 ;
  assign n52107 = n46652 ^ n38422 ^ 1'b0 ;
  assign n52108 = ~n52106 & n52107 ;
  assign n52104 = ~n243 & n23801 ;
  assign n52109 = n52108 ^ n52104 ^ 1'b0 ;
  assign n52110 = ~n19527 & n23149 ;
  assign n52111 = ~n29710 & n52110 ;
  assign n52112 = n39957 ^ n14821 ^ 1'b0 ;
  assign n52113 = n40020 ^ n12722 ^ 1'b0 ;
  assign n52114 = n12604 & ~n38170 ;
  assign n52115 = ~n47541 & n52114 ;
  assign n52116 = n52113 & n52115 ;
  assign n52117 = n21361 ^ n12756 ^ 1'b0 ;
  assign n52118 = n8775 & n52117 ;
  assign n52119 = n52118 ^ n24804 ^ 1'b0 ;
  assign n52120 = n49753 & ~n52119 ;
  assign n52121 = n23042 & n38311 ;
  assign n52122 = ( n16259 & ~n23928 ) | ( n16259 & n52121 ) | ( ~n23928 & n52121 ) ;
  assign n52123 = n49315 ^ n38405 ^ n3554 ;
  assign n52124 = n41099 ^ n37348 ^ 1'b0 ;
  assign n52125 = ( n29819 & ~n30400 ) | ( n29819 & n52124 ) | ( ~n30400 & n52124 ) ;
  assign n52126 = ~n12638 & n12822 ;
  assign n52127 = n52126 ^ n9564 ^ 1'b0 ;
  assign n52128 = n52127 ^ n46643 ^ 1'b0 ;
  assign n52129 = n49696 ^ n2519 ^ 1'b0 ;
  assign n52130 = n12593 & n22562 ;
  assign n52131 = n24130 & n52130 ;
  assign n52132 = n47827 & ~n52131 ;
  assign n52133 = n517 ^ n101 ^ 1'b0 ;
  assign n52134 = ~n4232 & n20128 ;
  assign n52135 = n52133 & n52134 ;
  assign n52136 = n14251 & ~n52135 ;
  assign n52137 = n4432 & n20111 ;
  assign n52138 = ~n1320 & n9233 ;
  assign n52139 = n6793 ^ n129 ^ 1'b0 ;
  assign n52140 = n44927 ^ n31944 ^ 1'b0 ;
  assign n52141 = n52139 | n52140 ;
  assign n52142 = n52141 ^ n52023 ^ 1'b0 ;
  assign n52143 = n23471 ^ n527 ^ 1'b0 ;
  assign n52144 = ~n13011 & n52143 ;
  assign n52145 = ~n46294 & n52144 ;
  assign n52146 = n12816 & n52145 ;
  assign n52147 = n13011 | n14671 ;
  assign n52148 = n32795 & ~n52147 ;
  assign n52149 = n4810 & n16636 ;
  assign n52150 = n17997 | n28699 ;
  assign n52151 = n29000 | n52150 ;
  assign n52152 = n13903 | n14783 ;
  assign n52153 = n24754 & ~n52152 ;
  assign n52154 = n51677 ^ n16550 ^ n5656 ;
  assign n52155 = n6490 ^ n2434 ^ 1'b0 ;
  assign n52156 = n1040 & ~n3817 ;
  assign n52157 = n52156 ^ n7190 ^ 1'b0 ;
  assign n52158 = ~n5339 & n50578 ;
  assign n52159 = ~n8220 & n52158 ;
  assign n52160 = n46854 ^ n29384 ^ 1'b0 ;
  assign n52161 = ~n3920 & n28395 ;
  assign n52162 = ~n52160 & n52161 ;
  assign n52163 = n27829 ^ n6193 ^ 1'b0 ;
  assign n52164 = n25194 & n52163 ;
  assign n52165 = n7452 | n13274 ;
  assign n52166 = n1105 | n52165 ;
  assign n52167 = n52166 ^ n11682 ^ 1'b0 ;
  assign n52168 = ( ~n20071 & n47102 ) | ( ~n20071 & n52167 ) | ( n47102 & n52167 ) ;
  assign n52169 = n29821 | n52168 ;
  assign n52170 = n13123 | n17149 ;
  assign n52171 = n45576 ^ n31676 ^ 1'b0 ;
  assign n52172 = n12442 & n52171 ;
  assign n52173 = ( n1367 & n4156 ) | ( n1367 & ~n21519 ) | ( n4156 & ~n21519 ) ;
  assign n52174 = n41190 ^ n40434 ^ n1932 ;
  assign n52175 = n52174 ^ n39071 ^ n5781 ;
  assign n52176 = n4569 & ~n13991 ;
  assign n52177 = n2650 & n52176 ;
  assign n52178 = n36101 & ~n52177 ;
  assign n52179 = ( ~n4947 & n10832 ) | ( ~n4947 & n52178 ) | ( n10832 & n52178 ) ;
  assign n52180 = ~n22686 & n45696 ;
  assign n52181 = n4074 | n16394 ;
  assign n52182 = n8833 & ~n21674 ;
  assign n52183 = n52182 ^ n16343 ^ 1'b0 ;
  assign n52184 = ( n24234 & n24996 ) | ( n24234 & ~n52183 ) | ( n24996 & ~n52183 ) ;
  assign n52185 = ~n11930 & n22915 ;
  assign n52186 = n52185 ^ n44582 ^ 1'b0 ;
  assign n52187 = n18349 | n20177 ;
  assign n52188 = n18654 & n27541 ;
  assign n52189 = n52188 ^ n645 ^ 1'b0 ;
  assign n52190 = n8777 ^ n356 ^ 1'b0 ;
  assign n52191 = n8207 & ~n52190 ;
  assign n52192 = ~n23172 & n41636 ;
  assign n52193 = n9169 & ~n52192 ;
  assign n52194 = n52193 ^ n12198 ^ 1'b0 ;
  assign n52195 = ~n3408 & n30789 ;
  assign n52196 = n52194 & n52195 ;
  assign n52197 = n8581 ^ n3655 ^ 1'b0 ;
  assign n52198 = n16652 | n52197 ;
  assign n52199 = n52198 ^ n1079 ^ 1'b0 ;
  assign n52200 = n846 & ~n13555 ;
  assign n52201 = ~n6513 & n52200 ;
  assign n52202 = n4280 | n52201 ;
  assign n52203 = ~n1950 & n43392 ;
  assign n52204 = n52203 ^ n33849 ^ x7 ;
  assign n52205 = ~n8907 & n32096 ;
  assign n52206 = n19299 & n52205 ;
  assign n52207 = n12163 & ~n52206 ;
  assign n52208 = ~n2939 & n18245 ;
  assign n52209 = n52208 ^ n2889 ^ 1'b0 ;
  assign n52210 = n7915 & ~n23669 ;
  assign n52211 = n52210 ^ n45594 ^ 1'b0 ;
  assign n52212 = n46286 ^ n3190 ^ 1'b0 ;
  assign n52213 = n22345 & ~n52212 ;
  assign n52214 = ~n22110 & n52213 ;
  assign n52215 = ~n18893 & n38216 ;
  assign n52216 = n52214 & n52215 ;
  assign n52217 = n827 | n31622 ;
  assign n52218 = n281 & ~n52217 ;
  assign n52219 = n31109 & n41526 ;
  assign n52220 = ( n2196 & n8648 ) | ( n2196 & n52219 ) | ( n8648 & n52219 ) ;
  assign n52221 = ~n31661 & n52220 ;
  assign n52223 = n3608 & n13713 ;
  assign n52224 = ~n13713 & n52223 ;
  assign n52225 = ~n3330 & n52224 ;
  assign n52226 = n18363 & n52225 ;
  assign n52227 = n44578 | n52226 ;
  assign n52222 = n6551 ^ n5725 ^ n730 ;
  assign n52228 = n52227 ^ n52222 ^ 1'b0 ;
  assign n52229 = n24579 ^ n16858 ^ 1'b0 ;
  assign n52230 = n37388 & n52229 ;
  assign n52231 = n10229 | n21751 ;
  assign n52232 = n52231 ^ n29580 ^ 1'b0 ;
  assign n52233 = n16162 | n45749 ;
  assign n52234 = n42507 & ~n52233 ;
  assign n52235 = n47164 ^ n44923 ^ 1'b0 ;
  assign n52236 = n22840 | n52235 ;
  assign n52237 = n2640 | n14849 ;
  assign n52238 = n52237 ^ n6153 ^ 1'b0 ;
  assign n52239 = n6889 & ~n51429 ;
  assign n52240 = n52239 ^ n50963 ^ 1'b0 ;
  assign n52241 = ~n9337 & n39219 ;
  assign n52242 = n52241 ^ n12736 ^ 1'b0 ;
  assign n52243 = ~n14450 & n33813 ;
  assign n52244 = n52243 ^ n42827 ^ n4562 ;
  assign n52245 = n37828 ^ n17030 ^ 1'b0 ;
  assign n52246 = n52245 ^ n1039 ^ 1'b0 ;
  assign n52247 = ~n7285 & n25477 ;
  assign n52248 = ~n19223 & n52247 ;
  assign n52249 = n52248 ^ n6965 ^ 1'b0 ;
  assign n52250 = ~n35910 & n52249 ;
  assign n52251 = ( n1374 & n11330 ) | ( n1374 & n23157 ) | ( n11330 & n23157 ) ;
  assign n52252 = n34583 | n52251 ;
  assign n52253 = n52252 ^ n2939 ^ 1'b0 ;
  assign n52255 = n27490 & n29117 ;
  assign n52254 = n2738 & ~n35415 ;
  assign n52256 = n52255 ^ n52254 ^ 1'b0 ;
  assign n52257 = n8382 ^ n7150 ^ 1'b0 ;
  assign n52258 = ~n5985 & n52257 ;
  assign n52259 = n52258 ^ n4956 ^ 1'b0 ;
  assign n52260 = n52259 ^ n19513 ^ 1'b0 ;
  assign n52261 = n52256 & n52260 ;
  assign n52263 = n19778 ^ n12931 ^ n2034 ;
  assign n52262 = n37564 | n47641 ;
  assign n52264 = n52263 ^ n52262 ^ 1'b0 ;
  assign n52265 = n26695 ^ n16728 ^ 1'b0 ;
  assign n52266 = n1320 & ~n52265 ;
  assign n52267 = n39961 ^ n27854 ^ n13960 ;
  assign n52268 = ~n33917 & n52267 ;
  assign n52269 = ( ~n3005 & n21391 ) | ( ~n3005 & n52268 ) | ( n21391 & n52268 ) ;
  assign n52270 = n52269 ^ n19385 ^ 1'b0 ;
  assign n52271 = n9570 & n31720 ;
  assign n52272 = ~n39838 & n52271 ;
  assign n52273 = n39722 ^ n9875 ^ 1'b0 ;
  assign n52274 = n2618 & ~n36171 ;
  assign n52275 = n14076 & n52274 ;
  assign n52276 = n5867 | n7584 ;
  assign n52277 = n8580 & n34473 ;
  assign n52278 = n35132 & n52277 ;
  assign n52279 = n31431 & ~n52278 ;
  assign n52280 = ~n52276 & n52279 ;
  assign n52282 = n14077 ^ n6497 ^ 1'b0 ;
  assign n52281 = n8153 & n47697 ;
  assign n52283 = n52282 ^ n52281 ^ 1'b0 ;
  assign n52284 = n9111 & ~n43659 ;
  assign n52285 = n52284 ^ n6638 ^ 1'b0 ;
  assign n52286 = n25067 ^ n16658 ^ 1'b0 ;
  assign n52287 = ~n37848 & n52286 ;
  assign n52288 = n50716 & ~n52287 ;
  assign n52289 = ( n17235 & ~n24916 ) | ( n17235 & n36822 ) | ( ~n24916 & n36822 ) ;
  assign n52290 = n13546 & n23161 ;
  assign n52291 = n52290 ^ n24987 ^ 1'b0 ;
  assign n52292 = n45078 & n52291 ;
  assign n52293 = n52292 ^ n33022 ^ 1'b0 ;
  assign n52294 = ( n34464 & ~n51911 ) | ( n34464 & n52293 ) | ( ~n51911 & n52293 ) ;
  assign n52295 = n13218 | n41970 ;
  assign n52296 = n44930 ^ n6212 ^ 1'b0 ;
  assign n52297 = n21125 & n52296 ;
  assign n52298 = n33965 ^ n757 ^ 1'b0 ;
  assign n52299 = n4523 ^ n2845 ^ 1'b0 ;
  assign n52300 = n7380 | n52299 ;
  assign n52301 = n17325 & n52300 ;
  assign n52302 = n34240 ^ n18780 ^ n3313 ;
  assign n52303 = n1491 & ~n28816 ;
  assign n52304 = n40671 & ~n52303 ;
  assign n52305 = n1465 | n34357 ;
  assign n52306 = n5595 & n52305 ;
  assign n52307 = n6934 & n52306 ;
  assign n52308 = ~n927 & n3731 ;
  assign n52309 = n52308 ^ n20153 ^ 1'b0 ;
  assign n52311 = n33253 ^ n22705 ^ 1'b0 ;
  assign n52312 = n24252 & n52311 ;
  assign n52310 = ~n45743 & n51580 ;
  assign n52313 = n52312 ^ n52310 ^ 1'b0 ;
  assign n52314 = n24049 ^ n908 ^ 1'b0 ;
  assign n52315 = n2934 & n33268 ;
  assign n52316 = n51 & n52315 ;
  assign n52317 = n13900 & ~n52316 ;
  assign n52318 = n52317 ^ n961 ^ 1'b0 ;
  assign n52319 = ~n27671 & n43861 ;
  assign n52320 = n3442 & n52319 ;
  assign n52321 = n42513 & ~n43702 ;
  assign n52322 = n22514 ^ n3543 ^ 1'b0 ;
  assign n52323 = n52321 & n52322 ;
  assign n52324 = n2667 & n7795 ;
  assign n52325 = n29948 & n31026 ;
  assign n52326 = ( n1666 & n12337 ) | ( n1666 & n41679 ) | ( n12337 & n41679 ) ;
  assign n52327 = n3540 | n39930 ;
  assign n52328 = n52327 ^ n32707 ^ 1'b0 ;
  assign n52329 = n38439 | n52328 ;
  assign n52330 = n31065 ^ n16606 ^ 1'b0 ;
  assign n52331 = n36579 | n52330 ;
  assign n52332 = n14239 ^ n10597 ^ 1'b0 ;
  assign n52333 = ( n14294 & ~n49707 ) | ( n14294 & n52332 ) | ( ~n49707 & n52332 ) ;
  assign n52334 = ~n22734 & n36034 ;
  assign n52335 = n24082 ^ n13455 ^ 1'b0 ;
  assign n52336 = n3195 & n52335 ;
  assign n52337 = n14152 ^ n3313 ^ 1'b0 ;
  assign n52338 = ~n16307 & n52337 ;
  assign n52339 = n2508 & n52338 ;
  assign n52340 = n52339 ^ n18193 ^ 1'b0 ;
  assign n52341 = n10672 ^ n8051 ^ 1'b0 ;
  assign n52342 = n13218 | n18763 ;
  assign n52343 = ( n19646 & n52341 ) | ( n19646 & ~n52342 ) | ( n52341 & ~n52342 ) ;
  assign n52344 = ( n10576 & n18077 ) | ( n10576 & ~n27339 ) | ( n18077 & ~n27339 ) ;
  assign n52345 = n41588 ^ n23264 ^ 1'b0 ;
  assign n52346 = ~n12211 & n23579 ;
  assign n52347 = n52346 ^ n32746 ^ 1'b0 ;
  assign n52348 = n52102 ^ n23519 ^ 1'b0 ;
  assign n52349 = n16440 | n25358 ;
  assign n52350 = n52349 ^ n8483 ^ 1'b0 ;
  assign n52351 = n40869 & n52350 ;
  assign n52352 = n25910 & n33743 ;
  assign n52353 = ~n19825 & n31478 ;
  assign n52354 = ~n9057 & n52353 ;
  assign n52355 = n8555 & n52354 ;
  assign n52356 = ( n7853 & ~n37595 ) | ( n7853 & n37801 ) | ( ~n37595 & n37801 ) ;
  assign n52357 = ~n3327 & n4939 ;
  assign n52358 = n10654 & n52357 ;
  assign n52359 = n52358 ^ n37348 ^ 1'b0 ;
  assign n52360 = n32 & n52359 ;
  assign n52361 = n52360 ^ n23278 ^ 1'b0 ;
  assign n52362 = n27838 & n52361 ;
  assign n52363 = n52362 ^ n20911 ^ 1'b0 ;
  assign n52364 = ~n3816 & n34112 ;
  assign n52365 = n52364 ^ n23440 ^ 1'b0 ;
  assign n52366 = ( ~n3000 & n13326 ) | ( ~n3000 & n52365 ) | ( n13326 & n52365 ) ;
  assign n52373 = ~n20070 & n35684 ;
  assign n52367 = n17320 & ~n23675 ;
  assign n52368 = n1346 & n52367 ;
  assign n52369 = n4105 & n52368 ;
  assign n52370 = ~n20 & n30760 ;
  assign n52371 = n52370 ^ n47329 ^ 1'b0 ;
  assign n52372 = n52369 & ~n52371 ;
  assign n52374 = n52373 ^ n52372 ^ n8607 ;
  assign n52375 = n6977 & ~n13649 ;
  assign n52376 = n52375 ^ n7890 ^ n5164 ;
  assign n52377 = n23411 & n23534 ;
  assign n52378 = n12129 & n52377 ;
  assign n52379 = n41465 ^ n10897 ^ 1'b0 ;
  assign n52380 = ~n12121 & n52379 ;
  assign n52381 = n10001 & n52380 ;
  assign n52382 = n1196 | n37187 ;
  assign n52383 = n45435 | n52382 ;
  assign n52384 = n6466 ^ n836 ^ 1'b0 ;
  assign n52385 = n17689 ^ n2945 ^ 1'b0 ;
  assign n52386 = ( ~n22826 & n35131 ) | ( ~n22826 & n52385 ) | ( n35131 & n52385 ) ;
  assign n52387 = ~n6042 & n32323 ;
  assign n52388 = n52387 ^ n10589 ^ 1'b0 ;
  assign n52389 = n52388 ^ n25225 ^ 1'b0 ;
  assign n52391 = n7354 ^ n6954 ^ 1'b0 ;
  assign n52392 = n10131 & n52391 ;
  assign n52393 = n52392 ^ n32303 ^ 1'b0 ;
  assign n52390 = n983 | n34241 ;
  assign n52394 = n52393 ^ n52390 ^ n46623 ;
  assign n52395 = n13677 ^ n4459 ^ 1'b0 ;
  assign n52396 = ~n40799 & n52395 ;
  assign n52397 = n52396 ^ n12269 ^ 1'b0 ;
  assign n52398 = n52397 ^ n3514 ^ 1'b0 ;
  assign n52399 = ~n20350 & n21495 ;
  assign n52400 = ~n3343 & n52399 ;
  assign n52401 = n52400 ^ n46537 ^ 1'b0 ;
  assign n52402 = n6713 ^ n3284 ^ 1'b0 ;
  assign n52403 = n13597 & ~n25420 ;
  assign n52404 = n15563 & n52403 ;
  assign n52405 = n36979 & ~n52404 ;
  assign n52406 = n9519 | n39956 ;
  assign n52407 = n52406 ^ n44069 ^ 1'b0 ;
  assign n52408 = n22377 ^ n1293 ^ 1'b0 ;
  assign n52409 = n14331 & n52408 ;
  assign n52410 = n28624 & n52409 ;
  assign n52411 = n41617 & n52410 ;
  assign n52412 = n39337 & n52411 ;
  assign n52413 = ~n923 & n26188 ;
  assign n52414 = n2047 & n52413 ;
  assign n52415 = n3600 & ~n10956 ;
  assign n52416 = n5520 & ~n34488 ;
  assign n52417 = n6076 & n52416 ;
  assign n52418 = n52417 ^ n31869 ^ 1'b0 ;
  assign n52419 = ~n2571 & n5140 ;
  assign n52420 = n24881 ^ n18611 ^ 1'b0 ;
  assign n52421 = n47935 ^ n14022 ^ 1'b0 ;
  assign n52422 = n39329 ^ n3575 ^ 1'b0 ;
  assign n52423 = n27152 ^ n8145 ^ 1'b0 ;
  assign n52424 = n11442 & ~n52423 ;
  assign n52425 = n28850 & ~n52424 ;
  assign n52426 = n15956 ^ n6044 ^ 1'b0 ;
  assign n52427 = n17203 & n52426 ;
  assign n52428 = n3127 | n25164 ;
  assign n52429 = n30043 & ~n52428 ;
  assign n52430 = n32413 ^ n13159 ^ 1'b0 ;
  assign n52431 = n41786 & ~n52430 ;
  assign n52432 = n25388 & n52431 ;
  assign n52433 = n4310 & ~n29668 ;
  assign n52434 = n52433 ^ n39931 ^ 1'b0 ;
  assign n52435 = n5830 | n52434 ;
  assign n52436 = n52435 ^ n19907 ^ 1'b0 ;
  assign n52437 = n13246 & n31688 ;
  assign n52438 = n52437 ^ n12926 ^ 1'b0 ;
  assign n52439 = n14915 ^ n10226 ^ 1'b0 ;
  assign n52440 = n52438 & n52439 ;
  assign n52441 = n11743 | n41589 ;
  assign n52442 = n10263 | n52441 ;
  assign n52443 = n13481 & n17185 ;
  assign n52444 = n32186 ^ n29454 ^ 1'b0 ;
  assign n52445 = n24302 | n52444 ;
  assign n52446 = n21253 & n52445 ;
  assign n52447 = ( n31727 & n43518 ) | ( n31727 & n52446 ) | ( n43518 & n52446 ) ;
  assign n52448 = ~n6638 & n9758 ;
  assign n52449 = n19102 ^ n7468 ^ 1'b0 ;
  assign n52450 = n17963 | n47662 ;
  assign n52451 = n52450 ^ n37354 ^ 1'b0 ;
  assign n52452 = n4092 ^ n1812 ^ 1'b0 ;
  assign n52453 = n33755 & ~n40739 ;
  assign n52454 = n21681 & n52453 ;
  assign n52455 = n7707 | n37997 ;
  assign n52456 = n5093 & ~n41499 ;
  assign n52457 = n48442 & ~n52456 ;
  assign n52458 = ( ~n8950 & n9961 ) | ( ~n8950 & n25652 ) | ( n9961 & n25652 ) ;
  assign n52459 = n3897 | n17030 ;
  assign n52460 = n52459 ^ n6412 ^ 1'b0 ;
  assign n52461 = n43015 & n52460 ;
  assign n52462 = n52461 ^ n12126 ^ 1'b0 ;
  assign n52463 = ~n36308 & n45018 ;
  assign n52464 = n45282 ^ n21643 ^ 1'b0 ;
  assign n52465 = n48293 ^ n4250 ^ 1'b0 ;
  assign n52466 = n52465 ^ n51901 ^ n22018 ;
  assign n52467 = n34317 & ~n49661 ;
  assign n52468 = n5160 & ~n7596 ;
  assign n52469 = n52468 ^ n15396 ^ n2849 ;
  assign n52470 = n52469 ^ n50401 ^ 1'b0 ;
  assign n52471 = n43398 ^ n2302 ^ 1'b0 ;
  assign n52472 = n40925 ^ n21165 ^ n12603 ;
  assign n52473 = n52472 ^ n4006 ^ 1'b0 ;
  assign n52474 = n32407 & ~n52473 ;
  assign n52475 = ~n17395 & n22103 ;
  assign n52476 = n9704 & n52291 ;
  assign n52477 = n49158 | n51939 ;
  assign n52478 = n21868 ^ n18373 ^ 1'b0 ;
  assign n52479 = n7354 & ~n17238 ;
  assign n52480 = n52479 ^ n14246 ^ 1'b0 ;
  assign n52486 = n574 | n3241 ;
  assign n52481 = n838 | n11013 ;
  assign n52482 = n28735 | n52481 ;
  assign n52483 = n24658 | n52482 ;
  assign n52484 = n33927 ^ n5639 ^ 1'b0 ;
  assign n52485 = n52483 & ~n52484 ;
  assign n52487 = n52486 ^ n52485 ^ n230 ;
  assign n52488 = n34596 ^ n22852 ^ n1078 ;
  assign n52489 = n25161 | n46894 ;
  assign n52490 = n52488 | n52489 ;
  assign n52492 = n23569 ^ n16829 ^ 1'b0 ;
  assign n52491 = n11730 & n13642 ;
  assign n52493 = n52492 ^ n52491 ^ 1'b0 ;
  assign n52494 = n5468 | n42301 ;
  assign n52495 = n42109 ^ n27526 ^ 1'b0 ;
  assign n52496 = n1807 | n28939 ;
  assign n52497 = ( n4847 & n35821 ) | ( n4847 & n52496 ) | ( n35821 & n52496 ) ;
  assign n52498 = n14204 & ~n52497 ;
  assign n52499 = n40510 ^ n15577 ^ 1'b0 ;
  assign n52500 = n7248 | n52499 ;
  assign n52501 = n5711 & ~n7870 ;
  assign n52502 = n2631 | n52501 ;
  assign n52503 = n52502 ^ n48229 ^ 1'b0 ;
  assign n52504 = n32717 & ~n52503 ;
  assign n52505 = ~n933 & n32052 ;
  assign n52506 = ~n18048 & n48969 ;
  assign n52507 = n52505 & n52506 ;
  assign n52508 = n3740 & n52507 ;
  assign n52509 = ( n4014 & n10284 ) | ( n4014 & ~n28398 ) | ( n10284 & ~n28398 ) ;
  assign n52510 = n9704 & n18453 ;
  assign n52511 = n6093 ^ n1518 ^ 1'b0 ;
  assign n52512 = n11798 & n15626 ;
  assign n52513 = ~n52511 & n52512 ;
  assign n52514 = n1391 | n5627 ;
  assign n52515 = n7787 & ~n30233 ;
  assign n52516 = n52515 ^ n25343 ^ 1'b0 ;
  assign n52517 = n37788 & n52516 ;
  assign n52518 = n9563 & ~n14590 ;
  assign n52519 = n1290 | n19210 ;
  assign n52520 = n52519 ^ n27319 ^ 1'b0 ;
  assign n52521 = n52518 | n52520 ;
  assign n52522 = n52521 ^ n16517 ^ 1'b0 ;
  assign n52523 = n13881 & ~n52522 ;
  assign n52524 = n31646 ^ n7938 ^ 1'b0 ;
  assign n52525 = n14522 | n41676 ;
  assign n52526 = n8428 & ~n52525 ;
  assign n52527 = n35855 | n52526 ;
  assign n52528 = n1990 & ~n3022 ;
  assign n52529 = n5604 & n7303 ;
  assign n52530 = ~n18332 & n52529 ;
  assign n52537 = n10512 | n25453 ;
  assign n52538 = n28279 & ~n52537 ;
  assign n52534 = n37562 ^ n13208 ^ 1'b0 ;
  assign n52535 = n9727 | n52534 ;
  assign n52536 = n52535 ^ n3214 ^ 1'b0 ;
  assign n52531 = n24394 ^ n8166 ^ n3522 ;
  assign n52532 = n2055 & ~n52531 ;
  assign n52533 = n52532 ^ n10114 ^ 1'b0 ;
  assign n52539 = n52538 ^ n52536 ^ n52533 ;
  assign n52540 = n52539 ^ n24783 ^ n11605 ;
  assign n52541 = ~n36604 & n52540 ;
  assign n52542 = n12801 & n18862 ;
  assign n52543 = n1586 & n13004 ;
  assign n52544 = ~n14889 & n39224 ;
  assign n52545 = n52544 ^ n12286 ^ 1'b0 ;
  assign n52546 = n52545 ^ n29720 ^ 1'b0 ;
  assign n52547 = n52546 ^ n937 ^ n488 ;
  assign n52548 = n848 & n22384 ;
  assign n52549 = n7376 | n12371 ;
  assign n52550 = ~n4957 & n46248 ;
  assign n52551 = n79 & ~n52550 ;
  assign n52552 = n22493 ^ n19002 ^ 1'b0 ;
  assign n52553 = n1311 & ~n18973 ;
  assign n52554 = ~n8443 & n52553 ;
  assign n52555 = ~n20214 & n49630 ;
  assign n52556 = n19000 & n52555 ;
  assign n52557 = ( n9524 & ~n24209 ) | ( n9524 & n44408 ) | ( ~n24209 & n44408 ) ;
  assign n52558 = n52557 ^ n37061 ^ n14709 ;
  assign n52559 = n27339 ^ n20235 ^ n15788 ;
  assign n52560 = n1063 & ~n21705 ;
  assign n52561 = n52560 ^ n4254 ^ 1'b0 ;
  assign n52562 = n52561 ^ n48484 ^ 1'b0 ;
  assign n52565 = n570 & n36930 ;
  assign n52566 = n52565 ^ n15748 ^ 1'b0 ;
  assign n52564 = n27403 | n34943 ;
  assign n52567 = n52566 ^ n52564 ^ 1'b0 ;
  assign n52563 = n27803 & ~n49369 ;
  assign n52568 = n52567 ^ n52563 ^ 1'b0 ;
  assign n52569 = n27107 ^ n16040 ^ n6644 ;
  assign n52570 = n52569 ^ n32956 ^ 1'b0 ;
  assign n52571 = n52570 ^ n33130 ^ n23532 ;
  assign n52572 = n18847 & ~n39176 ;
  assign n52573 = n52572 ^ n37763 ^ n37629 ;
  assign n52574 = n4429 & ~n45798 ;
  assign n52575 = n36938 & n52574 ;
  assign n52576 = n41651 ^ n31106 ^ 1'b0 ;
  assign n52577 = n50997 & n52576 ;
  assign n52578 = n7596 ^ n3240 ^ 1'b0 ;
  assign n52579 = n46812 ^ n37847 ^ 1'b0 ;
  assign n52580 = n52578 & ~n52579 ;
  assign n52581 = n25076 ^ n11103 ^ 1'b0 ;
  assign n52582 = n29172 | n52581 ;
  assign n52583 = n12211 | n52582 ;
  assign n52584 = n52583 ^ n43114 ^ 1'b0 ;
  assign n52585 = n13467 ^ n431 ^ 1'b0 ;
  assign n52586 = n10358 & ~n52585 ;
  assign n52587 = ~n5740 & n52586 ;
  assign n52588 = n30513 & n52587 ;
  assign n52589 = ( ~n16379 & n49907 ) | ( ~n16379 & n52588 ) | ( n49907 & n52588 ) ;
  assign n52590 = ( n310 & n7061 ) | ( n310 & n10586 ) | ( n7061 & n10586 ) ;
  assign n52591 = n52590 ^ n18024 ^ 1'b0 ;
  assign n52592 = n1945 & ~n52591 ;
  assign n52593 = n3188 | n19097 ;
  assign n52594 = n52593 ^ n34361 ^ 1'b0 ;
  assign n52595 = ( n50521 & n52592 ) | ( n50521 & n52594 ) | ( n52592 & n52594 ) ;
  assign n52596 = n2449 & ~n36502 ;
  assign n52598 = n10077 & n32396 ;
  assign n52599 = n52598 ^ n33329 ^ 1'b0 ;
  assign n52597 = n1121 ^ n523 ^ 1'b0 ;
  assign n52600 = n52599 ^ n52597 ^ 1'b0 ;
  assign n52601 = n10478 & ~n52600 ;
  assign n52602 = n52596 & n52601 ;
  assign n52603 = n15095 & ~n52602 ;
  assign n52604 = n52603 ^ n28058 ^ 1'b0 ;
  assign n52605 = n25045 & n25391 ;
  assign n52606 = ~n7842 & n52605 ;
  assign n52607 = ~n11065 & n29511 ;
  assign n52608 = n52606 & n52607 ;
  assign n52609 = n12121 ^ n8806 ^ 1'b0 ;
  assign n52610 = n3634 & n52609 ;
  assign n52611 = ( ~n46486 & n49660 ) | ( ~n46486 & n52610 ) | ( n49660 & n52610 ) ;
  assign n52612 = n27564 | n52611 ;
  assign n52613 = n27906 ^ n4373 ^ 1'b0 ;
  assign n52614 = n34798 | n52613 ;
  assign n52615 = ~n499 & n4317 ;
  assign n52616 = ~n6238 & n52615 ;
  assign n52617 = n42621 ^ n33644 ^ 1'b0 ;
  assign n52618 = n8321 & n26913 ;
  assign n52619 = ( n23095 & n41475 ) | ( n23095 & ~n52618 ) | ( n41475 & ~n52618 ) ;
  assign n52620 = n35322 ^ n25878 ^ 1'b0 ;
  assign n52621 = n7304 | n41121 ;
  assign n52622 = n6118 ^ n361 ^ 1'b0 ;
  assign n52623 = n52622 ^ n14417 ^ n2412 ;
  assign n52624 = n9096 & n35760 ;
  assign n52625 = ~n52623 & n52624 ;
  assign n52628 = ~n11640 & n44713 ;
  assign n52626 = n10473 & ~n45113 ;
  assign n52627 = n13237 & n52626 ;
  assign n52629 = n52628 ^ n52627 ^ 1'b0 ;
  assign n52630 = n46285 ^ n27102 ^ n15566 ;
  assign n52631 = ~n13096 & n52630 ;
  assign n52632 = n477 & ~n1311 ;
  assign n52633 = n52632 ^ n12439 ^ 1'b0 ;
  assign n52634 = ( n22464 & ~n25014 ) | ( n22464 & n47260 ) | ( ~n25014 & n47260 ) ;
  assign n52635 = n43421 ^ n15617 ^ 1'b0 ;
  assign n52636 = n2296 & ~n48788 ;
  assign n52637 = n43416 & n52636 ;
  assign n52638 = n52637 ^ n40414 ^ 1'b0 ;
  assign n52639 = n52635 & n52638 ;
  assign n52640 = n52639 ^ n45379 ^ 1'b0 ;
  assign n52641 = n36001 & ~n48179 ;
  assign n52642 = n52641 ^ n48985 ^ 1'b0 ;
  assign n52645 = ~n1896 & n34226 ;
  assign n52646 = n14219 & n52645 ;
  assign n52643 = n14449 | n29302 ;
  assign n52644 = n52643 ^ n18977 ^ 1'b0 ;
  assign n52647 = n52646 ^ n52644 ^ 1'b0 ;
  assign n52648 = n49982 ^ n9124 ^ 1'b0 ;
  assign n52649 = ~n52647 & n52648 ;
  assign n52650 = n5294 & ~n32955 ;
  assign n52651 = n47383 | n52650 ;
  assign n52652 = n13954 ^ n10147 ^ n5163 ;
  assign n52653 = n7610 & ~n18381 ;
  assign n52654 = n52652 | n52653 ;
  assign n52655 = n52654 ^ n8120 ^ 1'b0 ;
  assign n52656 = n22063 & ~n35636 ;
  assign n52657 = n22078 ^ n19664 ^ n7776 ;
  assign n52658 = n4684 ^ n3581 ^ 1'b0 ;
  assign n52659 = n2816 & ~n52658 ;
  assign n52660 = n30101 | n52659 ;
  assign n52661 = n35369 ^ n35344 ^ 1'b0 ;
  assign n52662 = n52660 & n52661 ;
  assign n52666 = n4915 ^ n2668 ^ n1572 ;
  assign n52663 = n29384 ^ n13747 ^ 1'b0 ;
  assign n52664 = n15660 & ~n52663 ;
  assign n52665 = ~n44006 & n52664 ;
  assign n52667 = n52666 ^ n52665 ^ 1'b0 ;
  assign n52668 = n12409 | n25615 ;
  assign n52669 = n12668 | n23015 ;
  assign n52670 = n52669 ^ n6144 ^ 1'b0 ;
  assign n52671 = n21906 ^ n14741 ^ 1'b0 ;
  assign n52672 = n20246 & n52671 ;
  assign n52673 = n43973 ^ n3807 ^ 1'b0 ;
  assign n52674 = n10154 & n52673 ;
  assign n52675 = n52674 ^ n8052 ^ 1'b0 ;
  assign n52676 = n3749 ^ n3626 ^ n469 ;
  assign n52677 = ( n7818 & ~n42431 ) | ( n7818 & n52676 ) | ( ~n42431 & n52676 ) ;
  assign n52678 = n41972 ^ n4697 ^ 1'b0 ;
  assign n52679 = n52678 ^ n46464 ^ n23072 ;
  assign n52680 = n24936 | n42847 ;
  assign n52681 = n52680 ^ n18053 ^ 1'b0 ;
  assign n52682 = n4275 | n52681 ;
  assign n52683 = n45915 ^ n10667 ^ 1'b0 ;
  assign n52684 = n52682 | n52683 ;
  assign n52685 = n44377 ^ n37200 ^ 1'b0 ;
  assign n52686 = n36848 & ~n52685 ;
  assign n52687 = ~n3850 & n41149 ;
  assign n52688 = ~n5363 & n52687 ;
  assign n52689 = n5673 & ~n41789 ;
  assign n52690 = ~n6902 & n51551 ;
  assign n52691 = n52690 ^ n15203 ^ 1'b0 ;
  assign n52694 = n31677 ^ n24412 ^ 1'b0 ;
  assign n52695 = n19345 & n52694 ;
  assign n52692 = n46592 ^ n21078 ^ 1'b0 ;
  assign n52693 = n25349 | n52692 ;
  assign n52696 = n52695 ^ n52693 ^ 1'b0 ;
  assign n52698 = n52166 ^ n11672 ^ n686 ;
  assign n52697 = ( n3484 & n10220 ) | ( n3484 & ~n41087 ) | ( n10220 & ~n41087 ) ;
  assign n52699 = n52698 ^ n52697 ^ 1'b0 ;
  assign n52700 = n12461 & n24235 ;
  assign n52702 = n12851 | n35243 ;
  assign n52703 = n631 & ~n52702 ;
  assign n52701 = n5212 | n44326 ;
  assign n52704 = n52703 ^ n52701 ^ 1'b0 ;
  assign n52705 = n1134 | n31129 ;
  assign n52706 = n18373 ^ n5892 ^ 1'b0 ;
  assign n52707 = n3151 & ~n52706 ;
  assign n52708 = n52707 ^ n18727 ^ 1'b0 ;
  assign n52709 = n24263 & n52708 ;
  assign n52710 = n6263 & ~n9626 ;
  assign n52711 = n52710 ^ n38326 ^ n34693 ;
  assign n52712 = n14881 ^ n8947 ^ 1'b0 ;
  assign n52713 = n1334 & n6341 ;
  assign n52714 = n3010 | n32580 ;
  assign n52715 = n15461 ^ n13947 ^ 1'b0 ;
  assign n52716 = ~n9688 & n15254 ;
  assign n52717 = n13445 & ~n26107 ;
  assign n52718 = ~n45785 & n52717 ;
  assign n52719 = n9146 & n48494 ;
  assign n52720 = n52719 ^ n16467 ^ 1'b0 ;
  assign n52721 = n34697 ^ n33337 ^ 1'b0 ;
  assign n52722 = n17737 & ~n52721 ;
  assign n52723 = n27416 & n52722 ;
  assign n52724 = n8150 | n15714 ;
  assign n52725 = n2173 | n52724 ;
  assign n52726 = n8101 | n28839 ;
  assign n52727 = n52725 | n52726 ;
  assign n52728 = ( ~n3967 & n13382 ) | ( ~n3967 & n52727 ) | ( n13382 & n52727 ) ;
  assign n52730 = n47876 ^ n30169 ^ 1'b0 ;
  assign n52731 = n31843 & ~n52730 ;
  assign n52729 = n5653 | n49055 ;
  assign n52732 = n52731 ^ n52729 ^ 1'b0 ;
  assign n52733 = ~n11529 & n36516 ;
  assign n52734 = n6514 & n52733 ;
  assign n52735 = n7759 & n10915 ;
  assign n52736 = ~n29026 & n52735 ;
  assign n52737 = n52734 & n52736 ;
  assign n52738 = n20322 ^ n11365 ^ 1'b0 ;
  assign n52739 = n10326 & ~n52738 ;
  assign n52740 = ~n11832 & n52739 ;
  assign n52741 = ( ~n1064 & n4489 ) | ( ~n1064 & n29423 ) | ( n4489 & n29423 ) ;
  assign n52742 = n20885 | n34424 ;
  assign n52743 = n52741 & ~n52742 ;
  assign n52744 = n8195 | n10254 ;
  assign n52745 = n52744 ^ n3408 ^ 1'b0 ;
  assign n52746 = ( n157 & n962 ) | ( n157 & n17096 ) | ( n962 & n17096 ) ;
  assign n52747 = ( n41023 & n50363 ) | ( n41023 & n52746 ) | ( n50363 & n52746 ) ;
  assign n52748 = n38725 ^ n28373 ^ 1'b0 ;
  assign n52749 = n36238 & n52748 ;
  assign n52750 = n20396 & n52749 ;
  assign n52751 = n12030 & n18813 ;
  assign n52752 = n2599 | n52751 ;
  assign n52753 = n52752 ^ n9969 ^ 1'b0 ;
  assign n52754 = n52753 ^ n40893 ^ n15277 ;
  assign n52755 = n7923 & n10739 ;
  assign n52756 = ~n51827 & n52755 ;
  assign n52757 = n3245 & n22271 ;
  assign n52758 = ~n3667 & n7334 ;
  assign n52759 = n52758 ^ n4978 ^ 1'b0 ;
  assign n52760 = n34607 & ~n52759 ;
  assign n52761 = ~n33706 & n43000 ;
  assign n52762 = n5494 & n52761 ;
  assign n52764 = n33239 ^ n9635 ^ 1'b0 ;
  assign n52763 = n10553 & ~n12477 ;
  assign n52765 = n52764 ^ n52763 ^ 1'b0 ;
  assign n52766 = n39722 ^ n31765 ^ n25540 ;
  assign n52767 = n21994 & ~n52766 ;
  assign n52768 = n52767 ^ n46970 ^ 1'b0 ;
  assign n52769 = ~n4335 & n9764 ;
  assign n52770 = n42998 ^ n13689 ^ 1'b0 ;
  assign n52771 = n52770 ^ n29583 ^ n4006 ;
  assign n52772 = n13923 & ~n16313 ;
  assign n52773 = n52772 ^ n823 ^ 1'b0 ;
  assign n52774 = n26551 ^ n17638 ^ 1'b0 ;
  assign n52775 = n23204 | n38634 ;
  assign n52776 = n52775 ^ n51038 ^ 1'b0 ;
  assign n52777 = ( n12695 & n52774 ) | ( n12695 & n52776 ) | ( n52774 & n52776 ) ;
  assign n52778 = ( n6591 & n9868 ) | ( n6591 & ~n14032 ) | ( n9868 & ~n14032 ) ;
  assign n52779 = n41428 ^ n24373 ^ 1'b0 ;
  assign n52780 = ~n1116 & n52779 ;
  assign n52781 = n52780 ^ n25326 ^ 1'b0 ;
  assign n52782 = n15164 & n52781 ;
  assign n52783 = n35653 | n52782 ;
  assign n52784 = n52783 ^ n37291 ^ 1'b0 ;
  assign n52785 = ~n52778 & n52784 ;
  assign n52786 = n19895 | n20931 ;
  assign n52787 = n1587 & ~n52786 ;
  assign n52788 = n52787 ^ n19817 ^ 1'b0 ;
  assign n52789 = n10841 & ~n52788 ;
  assign n52790 = ~n7387 & n37952 ;
  assign n52791 = n48656 ^ n18334 ^ 1'b0 ;
  assign n52792 = n23305 | n28428 ;
  assign n52793 = n19935 ^ n19021 ^ 1'b0 ;
  assign n52794 = n16271 & ~n37318 ;
  assign n52795 = n52794 ^ n2270 ^ 1'b0 ;
  assign n52796 = n37991 ^ n11339 ^ 1'b0 ;
  assign n52797 = n4909 & n52796 ;
  assign n52798 = n2350 | n42296 ;
  assign n52799 = n8174 | n41529 ;
  assign n52801 = ~n1246 & n3655 ;
  assign n52802 = n1066 & n52801 ;
  assign n52803 = n11810 ^ n6695 ^ 1'b0 ;
  assign n52804 = n52802 | n52803 ;
  assign n52800 = ( n3003 & ~n7070 ) | ( n3003 & n30754 ) | ( ~n7070 & n30754 ) ;
  assign n52805 = n52804 ^ n52800 ^ n6114 ;
  assign n52806 = n206 & ~n12969 ;
  assign n52807 = ( n13860 & ~n36796 ) | ( n13860 & n46294 ) | ( ~n36796 & n46294 ) ;
  assign n52808 = n31194 ^ n20501 ^ 1'b0 ;
  assign n52809 = n52807 | n52808 ;
  assign n52810 = n30211 & ~n52430 ;
  assign n52811 = n4497 & ~n37972 ;
  assign n52812 = n52811 ^ n24452 ^ 1'b0 ;
  assign n52813 = n45412 ^ n42671 ^ 1'b0 ;
  assign n52814 = n6355 & n32002 ;
  assign n52815 = ~n46849 & n52814 ;
  assign n52816 = n52815 ^ n4622 ^ 1'b0 ;
  assign n52817 = n21761 & ~n46278 ;
  assign n52818 = n52817 ^ n25658 ^ 1'b0 ;
  assign n52819 = n3256 & n8024 ;
  assign n52820 = n52819 ^ n12890 ^ 1'b0 ;
  assign n52821 = n22704 & ~n26107 ;
  assign n52822 = n52821 ^ n5892 ^ 1'b0 ;
  assign n52826 = n15940 ^ n11213 ^ 1'b0 ;
  assign n52827 = n34782 | n52826 ;
  assign n52823 = ( n5979 & ~n6167 ) | ( n5979 & n18695 ) | ( ~n6167 & n18695 ) ;
  assign n52824 = ( n26975 & ~n50493 ) | ( n26975 & n52823 ) | ( ~n50493 & n52823 ) ;
  assign n52825 = n1004 & ~n52824 ;
  assign n52828 = n52827 ^ n52825 ^ n4410 ;
  assign n52829 = n2165 & n31729 ;
  assign n52830 = ~n5377 & n38018 ;
  assign n52831 = n52830 ^ n42994 ^ 1'b0 ;
  assign n52832 = n52831 ^ n41614 ^ n18816 ;
  assign n52833 = n28511 ^ n8406 ^ 1'b0 ;
  assign n52834 = n50673 & n52833 ;
  assign n52835 = n49822 ^ n7884 ^ 1'b0 ;
  assign n52836 = n34661 | n52835 ;
  assign n52837 = n52836 ^ n25539 ^ 1'b0 ;
  assign n52838 = n29338 & n32768 ;
  assign n52840 = ~n730 & n15624 ;
  assign n52841 = ~n21717 & n52840 ;
  assign n52839 = n8747 ^ n4559 ^ 1'b0 ;
  assign n52842 = n52841 ^ n52839 ^ n26551 ;
  assign n52843 = ( n1091 & n9450 ) | ( n1091 & n14061 ) | ( n9450 & n14061 ) ;
  assign n52844 = n52843 ^ n36924 ^ 1'b0 ;
  assign n52845 = n7787 & n49753 ;
  assign n52846 = n52845 ^ n50409 ^ 1'b0 ;
  assign n52847 = n52846 ^ n381 ^ 1'b0 ;
  assign n52848 = n52847 ^ n4461 ^ 1'b0 ;
  assign n52851 = ( n1126 & n1746 ) | ( n1126 & ~n2027 ) | ( n1746 & ~n2027 ) ;
  assign n52849 = n48050 ^ n20896 ^ 1'b0 ;
  assign n52850 = n49988 & n52849 ;
  assign n52852 = n52851 ^ n52850 ^ n26376 ;
  assign n52853 = n29609 ^ n7610 ^ 1'b0 ;
  assign n52854 = n6563 ^ n4228 ^ 1'b0 ;
  assign n52855 = n50272 ^ n27635 ^ 1'b0 ;
  assign n52856 = n52854 & ~n52855 ;
  assign n52857 = ( n15444 & n52853 ) | ( n15444 & n52856 ) | ( n52853 & n52856 ) ;
  assign n52858 = n41759 ^ n1851 ^ 1'b0 ;
  assign n52859 = n44053 ^ n12033 ^ 1'b0 ;
  assign n52860 = n21506 & ~n52859 ;
  assign n52861 = n27348 ^ n15936 ^ 1'b0 ;
  assign n52862 = n22940 & n52861 ;
  assign n52863 = n2489 & n49827 ;
  assign n52864 = n5436 & n32096 ;
  assign n52865 = n52864 ^ n14775 ^ 1'b0 ;
  assign n52866 = n2631 & ~n24164 ;
  assign n52867 = ~n52865 & n52866 ;
  assign n52869 = n3776 & ~n7118 ;
  assign n52870 = n12873 & n52869 ;
  assign n52868 = n48735 ^ n37715 ^ n7448 ;
  assign n52871 = n52870 ^ n52868 ^ 1'b0 ;
  assign n52872 = ( n35 & n4889 ) | ( n35 & ~n20764 ) | ( n4889 & ~n20764 ) ;
  assign n52873 = ~n7676 & n9226 ;
  assign n52874 = n52873 ^ n44257 ^ 1'b0 ;
  assign n52875 = n11405 ^ n5790 ^ 1'b0 ;
  assign n52876 = n20589 | n24644 ;
  assign n52877 = n52876 ^ n7913 ^ 1'b0 ;
  assign n52878 = n15789 ^ n2445 ^ 1'b0 ;
  assign n52879 = n10296 & ~n52878 ;
  assign n52880 = n3926 & n9169 ;
  assign n52881 = n52880 ^ n455 ^ 1'b0 ;
  assign n52882 = n4635 ^ n763 ^ 1'b0 ;
  assign n52883 = ~n52881 & n52882 ;
  assign n52884 = n10373 & n28130 ;
  assign n52885 = n52751 & n52884 ;
  assign n52886 = n15533 & ~n51019 ;
  assign n52887 = n14425 & n52886 ;
  assign n52888 = n43756 ^ n32453 ^ 1'b0 ;
  assign n52889 = n44284 ^ n21363 ^ n11383 ;
  assign n52890 = n6415 & ~n14156 ;
  assign n52891 = n10985 ^ n10245 ^ 1'b0 ;
  assign n52892 = n1391 & ~n52891 ;
  assign n52893 = ~n2040 & n4712 ;
  assign n52894 = ~n52892 & n52893 ;
  assign n52895 = n7167 & ~n43447 ;
  assign n52896 = ( n9571 & n16556 ) | ( n9571 & ~n25881 ) | ( n16556 & ~n25881 ) ;
  assign n52897 = n5554 | n52896 ;
  assign n52898 = n7654 & ~n29888 ;
  assign n52899 = n3082 & ~n12143 ;
  assign n52900 = n17824 | n52899 ;
  assign n52901 = n52900 ^ n50705 ^ 1'b0 ;
  assign n52902 = ~n52898 & n52901 ;
  assign n52903 = ~n25614 & n48047 ;
  assign n52904 = n2036 ^ n615 ^ n186 ;
  assign n52905 = n16047 ^ n10305 ^ 1'b0 ;
  assign n52906 = ~n52904 & n52905 ;
  assign n52907 = ( ~n412 & n7893 ) | ( ~n412 & n38139 ) | ( n7893 & n38139 ) ;
  assign n52908 = n6925 | n12314 ;
  assign n52909 = n2581 & n29531 ;
  assign n52910 = n52909 ^ n52393 ^ 1'b0 ;
  assign n52911 = n14996 & n43610 ;
  assign n52913 = n6493 | n26810 ;
  assign n52912 = n6245 & n36001 ;
  assign n52914 = n52913 ^ n52912 ^ 1'b0 ;
  assign n52915 = n1120 & ~n17441 ;
  assign n52916 = ~n31539 & n52915 ;
  assign n52917 = n7411 & n13412 ;
  assign n52918 = n34120 ^ n30472 ^ 1'b0 ;
  assign n52919 = n19050 ^ n2597 ^ 1'b0 ;
  assign n52920 = n8182 & n12146 ;
  assign n52921 = n18526 & ~n29845 ;
  assign n52922 = n18162 ^ n4204 ^ 1'b0 ;
  assign n52923 = ~n14960 & n30057 ;
  assign n52924 = n6316 & n52923 ;
  assign n52925 = n9040 ^ n3519 ^ n259 ;
  assign n52926 = n7413 | n52925 ;
  assign n52927 = n29222 | n52926 ;
  assign n52928 = n21863 | n26755 ;
  assign n52929 = ~n12695 & n35909 ;
  assign n52932 = ~n890 & n1389 ;
  assign n52930 = n35678 ^ n12109 ^ 1'b0 ;
  assign n52931 = ~n10491 & n52930 ;
  assign n52933 = n52932 ^ n52931 ^ 1'b0 ;
  assign n52934 = n48130 ^ n24789 ^ 1'b0 ;
  assign n52936 = n14439 | n37670 ;
  assign n52937 = n35605 | n52936 ;
  assign n52935 = n5222 & n20129 ;
  assign n52938 = n52937 ^ n52935 ^ n49186 ;
  assign n52939 = n46469 ^ n12883 ^ n2486 ;
  assign n52940 = n52938 | n52939 ;
  assign n52941 = n8945 | n37918 ;
  assign n52942 = n11177 & ~n52941 ;
  assign n52943 = n47948 ^ n23852 ^ n16155 ;
  assign n52944 = n30460 ^ n16670 ^ 1'b0 ;
  assign n52945 = ~n52943 & n52944 ;
  assign n52946 = n12456 | n40112 ;
  assign n52947 = n18893 ^ n5301 ^ n4578 ;
  assign n52948 = n52946 & ~n52947 ;
  assign n52949 = n5625 & n52948 ;
  assign n52950 = ~n27471 & n52949 ;
  assign n52952 = n36906 ^ n26135 ^ 1'b0 ;
  assign n52951 = n37057 | n48770 ;
  assign n52953 = n52952 ^ n52951 ^ 1'b0 ;
  assign n52954 = ~n7916 & n34844 ;
  assign n52955 = n17080 ^ n9251 ^ 1'b0 ;
  assign n52956 = n36571 ^ n28918 ^ n10764 ;
  assign n52957 = ~n15282 & n52956 ;
  assign n52958 = n52957 ^ n50897 ^ 1'b0 ;
  assign n52959 = n25806 ^ n16242 ^ 1'b0 ;
  assign n52960 = n16169 | n52959 ;
  assign n52961 = n25519 ^ n21007 ^ 1'b0 ;
  assign n52962 = n38968 | n52961 ;
  assign n52963 = n7208 & n40523 ;
  assign n52964 = ~n12877 & n52963 ;
  assign n52965 = n52964 ^ n48832 ^ n1791 ;
  assign n52966 = n4002 & ~n14064 ;
  assign n52967 = n32825 ^ n18280 ^ n8018 ;
  assign n52968 = n39199 & ~n52967 ;
  assign n52969 = n52968 ^ n15504 ^ 1'b0 ;
  assign n52970 = n12391 & n35865 ;
  assign n52973 = n18573 ^ n7400 ^ n1296 ;
  assign n52971 = n51944 ^ n42683 ^ n12061 ;
  assign n52972 = n52971 ^ n28761 ^ n27405 ;
  assign n52974 = n52973 ^ n52972 ^ n2544 ;
  assign n52975 = n28761 ^ n814 ^ 1'b0 ;
  assign n52976 = n52975 ^ n14428 ^ n4770 ;
  assign n52977 = n52976 ^ n40803 ^ 1'b0 ;
  assign n52978 = ~n3741 & n52977 ;
  assign n52979 = ~n52974 & n52978 ;
  assign n52980 = ~n3027 & n6909 ;
  assign n52981 = n52980 ^ n4188 ^ 1'b0 ;
  assign n52982 = n21967 & ~n52981 ;
  assign n52983 = n52982 ^ n19083 ^ 1'b0 ;
  assign n52984 = ~n50897 & n52983 ;
  assign n52985 = n52984 ^ n41978 ^ 1'b0 ;
  assign n52986 = n7993 & n38955 ;
  assign n52987 = ~n20101 & n52986 ;
  assign n52988 = n35198 ^ n19436 ^ 1'b0 ;
  assign n52989 = ~n3192 & n52988 ;
  assign n52990 = n52989 ^ n34665 ^ 1'b0 ;
  assign n52991 = n52990 ^ n3345 ^ 1'b0 ;
  assign n52992 = n52987 | n52991 ;
  assign n52993 = n50570 ^ n8403 ^ 1'b0 ;
  assign n52994 = n52426 ^ n16792 ^ n4118 ;
  assign n52995 = n19158 ^ n13666 ^ 1'b0 ;
  assign n52996 = n52994 & n52995 ;
  assign n52997 = n13230 ^ n13112 ^ 1'b0 ;
  assign n52998 = n7915 & ~n52997 ;
  assign n52999 = n12606 ^ n819 ^ 1'b0 ;
  assign n53000 = n32823 | n52999 ;
  assign n53001 = n19324 & ~n53000 ;
  assign n53002 = n2648 & ~n53001 ;
  assign n53005 = n9511 ^ n1856 ^ 1'b0 ;
  assign n53003 = n22815 ^ n14386 ^ 1'b0 ;
  assign n53004 = ~n10348 & n53003 ;
  assign n53006 = n53005 ^ n53004 ^ 1'b0 ;
  assign n53007 = n5486 | n50914 ;
  assign n53008 = ( n12339 & ~n26025 ) | ( n12339 & n53007 ) | ( ~n26025 & n53007 ) ;
  assign n53009 = ( n15324 & ~n53006 ) | ( n15324 & n53008 ) | ( ~n53006 & n53008 ) ;
  assign n53012 = n2566 & n13949 ;
  assign n53013 = ~n11791 & n53012 ;
  assign n53014 = n1992 | n53013 ;
  assign n53015 = n53014 ^ n7126 ^ 1'b0 ;
  assign n53016 = n39539 | n53015 ;
  assign n53010 = n28368 & n32125 ;
  assign n53011 = n10707 | n53010 ;
  assign n53017 = n53016 ^ n53011 ^ 1'b0 ;
  assign n53018 = n3530 & ~n18742 ;
  assign n53019 = n39612 & n53018 ;
  assign n53020 = n40230 ^ n16444 ^ 1'b0 ;
  assign n53021 = n5760 & n47185 ;
  assign n53022 = ~n8409 & n15569 ;
  assign n53023 = n53022 ^ n21926 ^ 1'b0 ;
  assign n53024 = n23656 ^ n13333 ^ n4690 ;
  assign n53025 = n46909 ^ n6597 ^ 1'b0 ;
  assign n53026 = n1300 & ~n8458 ;
  assign n53027 = n26810 & n53026 ;
  assign n53028 = n26297 & n49089 ;
  assign n53029 = ~n8595 & n53028 ;
  assign n53030 = ( n42789 & n53027 ) | ( n42789 & ~n53029 ) | ( n53027 & ~n53029 ) ;
  assign n53031 = ~n4287 & n16755 ;
  assign n53032 = n11733 & ~n44143 ;
  assign n53033 = n53032 ^ n16124 ^ 1'b0 ;
  assign n53034 = n1493 | n45285 ;
  assign n53035 = n11197 & ~n53034 ;
  assign n53036 = n29931 | n53035 ;
  assign n53037 = n53036 ^ n34042 ^ 1'b0 ;
  assign n53038 = n12915 & n25237 ;
  assign n53039 = n9242 | n53038 ;
  assign n53040 = n19399 ^ n15444 ^ n1022 ;
  assign n53041 = n20781 ^ n17360 ^ 1'b0 ;
  assign n53042 = n34920 | n53041 ;
  assign n53043 = n38248 ^ n26783 ^ n8941 ;
  assign n53044 = ~n53042 & n53043 ;
  assign n53045 = n47543 ^ n14080 ^ 1'b0 ;
  assign n53046 = n1139 & n53045 ;
  assign n53047 = ~n16687 & n51176 ;
  assign n53048 = n53047 ^ n20707 ^ 1'b0 ;
  assign n53049 = n6496 | n42703 ;
  assign n53050 = n53048 | n53049 ;
  assign n53051 = n9778 & ~n37638 ;
  assign n53052 = ~n36273 & n53051 ;
  assign n53053 = n3606 & n53052 ;
  assign n53054 = n43370 ^ n37258 ^ 1'b0 ;
  assign n53055 = n22529 | n53054 ;
  assign n53056 = n2139 & ~n48784 ;
  assign n53057 = n53056 ^ n4635 ^ 1'b0 ;
  assign n53058 = ( n29638 & n34973 ) | ( n29638 & ~n53057 ) | ( n34973 & ~n53057 ) ;
  assign n53059 = n2483 & ~n53058 ;
  assign n53060 = n53059 ^ n16522 ^ 1'b0 ;
  assign n53062 = n33077 ^ n7634 ^ n1267 ;
  assign n53063 = n53062 ^ n23214 ^ 1'b0 ;
  assign n53064 = n24372 | n53063 ;
  assign n53061 = n44080 ^ n25050 ^ n6154 ;
  assign n53065 = n53064 ^ n53061 ^ n4267 ;
  assign n53066 = n20289 ^ n8342 ^ 1'b0 ;
  assign n53067 = n8647 ^ n3843 ^ n3523 ;
  assign n53068 = n13821 ^ n5469 ^ 1'b0 ;
  assign n53069 = n53067 | n53068 ;
  assign n53070 = ~n243 & n9171 ;
  assign n53071 = ( ~n1808 & n7915 ) | ( ~n1808 & n25973 ) | ( n7915 & n25973 ) ;
  assign n53072 = ( n29966 & ~n53070 ) | ( n29966 & n53071 ) | ( ~n53070 & n53071 ) ;
  assign n53073 = n53072 ^ n18123 ^ 1'b0 ;
  assign n53074 = n31411 ^ n2719 ^ 1'b0 ;
  assign n53079 = n6277 & n16630 ;
  assign n53075 = n10185 | n18228 ;
  assign n53076 = n53075 ^ n26729 ^ 1'b0 ;
  assign n53077 = n53076 ^ n8175 ^ n334 ;
  assign n53078 = ~n2577 & n53077 ;
  assign n53080 = n53079 ^ n53078 ^ 1'b0 ;
  assign n53081 = n50668 ^ n16251 ^ 1'b0 ;
  assign n53082 = n21876 & ~n24421 ;
  assign n53083 = ~n47697 & n53082 ;
  assign n53084 = n43095 ^ n11832 ^ 1'b0 ;
  assign n53085 = n12422 | n53084 ;
  assign n53086 = ( n6071 & n12149 ) | ( n6071 & n53085 ) | ( n12149 & n53085 ) ;
  assign n53087 = ~n5389 & n13479 ;
  assign n53088 = n33172 & ~n34207 ;
  assign n53089 = n17149 & ~n40158 ;
  assign n53090 = n53089 ^ n35364 ^ 1'b0 ;
  assign n53091 = n42871 ^ n3751 ^ 1'b0 ;
  assign n53092 = ~n53090 & n53091 ;
  assign n53093 = n14004 | n37628 ;
  assign n53094 = n39568 | n53093 ;
  assign n53095 = n21079 | n44281 ;
  assign n53097 = n28835 ^ n3479 ^ n2538 ;
  assign n53096 = ~n9646 & n51595 ;
  assign n53098 = n53097 ^ n53096 ^ 1'b0 ;
  assign n53099 = n32510 & n53098 ;
  assign n53100 = n53099 ^ n21703 ^ 1'b0 ;
  assign n53101 = n1455 & ~n11891 ;
  assign n53102 = n53101 ^ n7368 ^ 1'b0 ;
  assign n53103 = n18208 & n53102 ;
  assign n53104 = ( ~n5044 & n9227 ) | ( ~n5044 & n12425 ) | ( n9227 & n12425 ) ;
  assign n53105 = n46005 ^ n19549 ^ 1'b0 ;
  assign n53106 = n39588 ^ n6273 ^ 1'b0 ;
  assign n53107 = n33896 | n53106 ;
  assign n53108 = n25160 & ~n53107 ;
  assign n53109 = n53108 ^ n1178 ^ 1'b0 ;
  assign n53110 = n2589 & ~n53006 ;
  assign n53111 = ~n8491 & n53110 ;
  assign n53112 = n12054 & n14331 ;
  assign n53113 = n53112 ^ n1531 ^ 1'b0 ;
  assign n53114 = n2818 & ~n42217 ;
  assign n53115 = n53113 & n53114 ;
  assign n53119 = n32323 ^ n17508 ^ n10721 ;
  assign n53116 = ~n22488 & n26514 ;
  assign n53117 = ~n607 & n53116 ;
  assign n53118 = n6454 | n53117 ;
  assign n53120 = n53119 ^ n53118 ^ 1'b0 ;
  assign n53121 = ~n10868 & n36099 ;
  assign n53122 = n53121 ^ n14981 ^ 1'b0 ;
  assign n53123 = n25889 ^ n12175 ^ 1'b0 ;
  assign n53124 = ( n10065 & ~n13757 ) | ( n10065 & n21870 ) | ( ~n13757 & n21870 ) ;
  assign n53125 = n53124 ^ n43807 ^ 1'b0 ;
  assign n53126 = n42697 ^ n3067 ^ 1'b0 ;
  assign n53127 = ~n16178 & n53126 ;
  assign n53128 = n2341 & n15009 ;
  assign n53129 = n51510 ^ n791 ^ 1'b0 ;
  assign n53130 = n42867 | n53129 ;
  assign n53131 = n14715 | n29685 ;
  assign n53132 = n53131 ^ n5820 ^ 1'b0 ;
  assign n53133 = n29683 ^ n22751 ^ 1'b0 ;
  assign n53134 = n23335 ^ n3779 ^ 1'b0 ;
  assign n53136 = ( n5294 & n7479 ) | ( n5294 & n48136 ) | ( n7479 & n48136 ) ;
  assign n53135 = n2615 & ~n12106 ;
  assign n53137 = n53136 ^ n53135 ^ n34724 ;
  assign n53138 = ~n378 & n53137 ;
  assign n53139 = ~n44857 & n53138 ;
  assign n53140 = ( ~n26800 & n53134 ) | ( ~n26800 & n53139 ) | ( n53134 & n53139 ) ;
  assign n53141 = n53133 | n53140 ;
  assign n53142 = n5870 & ~n18737 ;
  assign n53143 = n26498 ^ n13164 ^ 1'b0 ;
  assign n53144 = ~n53142 & n53143 ;
  assign n53145 = n15781 & ~n47925 ;
  assign n53146 = n25011 | n30046 ;
  assign n53147 = n6381 | n20355 ;
  assign n53148 = n53147 ^ n34362 ^ n23030 ;
  assign n53149 = n826 & n40137 ;
  assign n53150 = n13866 & n53149 ;
  assign n53151 = n777 & n6406 ;
  assign n53152 = n53150 & n53151 ;
  assign n53153 = ( n6353 & ~n27419 ) | ( n6353 & n53152 ) | ( ~n27419 & n53152 ) ;
  assign n53154 = n45384 ^ n26513 ^ 1'b0 ;
  assign n53155 = n7399 & ~n7846 ;
  assign n53156 = n53155 ^ n30558 ^ 1'b0 ;
  assign n53157 = n53156 ^ n52639 ^ n30076 ;
  assign n53158 = n53157 ^ n39675 ^ n18643 ;
  assign n53159 = n17502 ^ n5423 ^ 1'b0 ;
  assign n53160 = n3923 & ~n53159 ;
  assign n53161 = ~n30816 & n39590 ;
  assign n53164 = n51101 ^ n25953 ^ n17491 ;
  assign n53162 = n31305 ^ n12507 ^ 1'b0 ;
  assign n53163 = n29877 & n53162 ;
  assign n53165 = n53164 ^ n53163 ^ 1'b0 ;
  assign n53166 = n36839 | n53165 ;
  assign n53167 = n21373 & ~n33273 ;
  assign n53168 = n53167 ^ n33430 ^ 1'b0 ;
  assign n53169 = n3686 | n53168 ;
  assign n53170 = n26341 | n53169 ;
  assign n53171 = n53170 ^ n26430 ^ 1'b0 ;
  assign n53172 = n4974 & ~n30638 ;
  assign n53173 = n53172 ^ n14441 ^ 1'b0 ;
  assign n53174 = n53173 ^ n19226 ^ 1'b0 ;
  assign n53175 = n31411 | n53174 ;
  assign n53176 = n7657 ^ n1992 ^ 1'b0 ;
  assign n53177 = n53176 ^ n15919 ^ 1'b0 ;
  assign n53178 = n7091 ^ n1029 ^ 1'b0 ;
  assign n53179 = n53178 ^ n26455 ^ 1'b0 ;
  assign n53180 = n53177 | n53179 ;
  assign n53183 = n1996 | n43119 ;
  assign n53184 = n53183 ^ n20822 ^ 1'b0 ;
  assign n53181 = ( n11180 & n16500 ) | ( n11180 & ~n30842 ) | ( n16500 & ~n30842 ) ;
  assign n53182 = n21655 & n53181 ;
  assign n53185 = n53184 ^ n53182 ^ n9242 ;
  assign n53192 = n827 & n5693 ;
  assign n53193 = ~n827 & n53192 ;
  assign n53194 = n53193 ^ n15864 ^ 1'b0 ;
  assign n53186 = ~n3690 & n9659 ;
  assign n53187 = n3690 & n53186 ;
  assign n53188 = n41722 | n53187 ;
  assign n53189 = n53187 & ~n53188 ;
  assign n53190 = n28541 | n53189 ;
  assign n53191 = n27232 & ~n53190 ;
  assign n53195 = n53194 ^ n53191 ^ 1'b0 ;
  assign n53196 = n53195 ^ n28576 ^ n20407 ;
  assign n53197 = n14807 ^ n2086 ^ 1'b0 ;
  assign n53198 = ( n25354 & ~n53196 ) | ( n25354 & n53197 ) | ( ~n53196 & n53197 ) ;
  assign n53199 = ~n538 & n15653 ;
  assign n53200 = n53199 ^ n11078 ^ 1'b0 ;
  assign n53201 = n18312 | n53200 ;
  assign n53202 = n12826 | n53201 ;
  assign n53203 = n18212 & n25392 ;
  assign n53204 = ~n11009 & n53203 ;
  assign n53207 = n14370 & n40076 ;
  assign n53205 = n11853 & n40230 ;
  assign n53206 = n1078 & n53205 ;
  assign n53208 = n53207 ^ n53206 ^ 1'b0 ;
  assign n53209 = n45847 ^ n37353 ^ n29321 ;
  assign n53210 = n53209 ^ n3685 ^ 1'b0 ;
  assign n53211 = n4317 & n5083 ;
  assign n53212 = n9284 & n53211 ;
  assign n53213 = n7526 & ~n32289 ;
  assign n53214 = ~n47488 & n53213 ;
  assign n53215 = n12807 & ~n36005 ;
  assign n53216 = n20347 ^ n11614 ^ 1'b0 ;
  assign n53217 = n20698 & n21218 ;
  assign n53218 = ( n2114 & n16403 ) | ( n2114 & ~n46719 ) | ( n16403 & ~n46719 ) ;
  assign n53219 = n53218 ^ n11460 ^ 1'b0 ;
  assign n53220 = n30962 & ~n53219 ;
  assign n53221 = n53220 ^ n1351 ^ 1'b0 ;
  assign n53222 = n11577 & n16917 ;
  assign n53223 = ~n14551 & n33161 ;
  assign n53224 = ( ~n39138 & n53222 ) | ( ~n39138 & n53223 ) | ( n53222 & n53223 ) ;
  assign n53225 = n11830 | n35365 ;
  assign n53226 = n21902 ^ n2666 ^ 1'b0 ;
  assign n53227 = n48968 ^ n33482 ^ 1'b0 ;
  assign n53228 = n30929 ^ n2211 ^ 1'b0 ;
  assign n53229 = n25645 ^ n13157 ^ 1'b0 ;
  assign n53230 = n42677 | n53229 ;
  assign n53231 = n53230 ^ n3606 ^ 1'b0 ;
  assign n53232 = n6593 & n47080 ;
  assign n53233 = n53232 ^ n23890 ^ 1'b0 ;
  assign n53234 = n2815 & ~n53233 ;
  assign n53235 = n53081 ^ n15730 ^ 1'b0 ;
  assign n53236 = n53234 & ~n53235 ;
  assign n53237 = n39325 ^ n27044 ^ n26926 ;
  assign n53238 = ~n2123 & n18339 ;
  assign n53239 = n18330 & ~n45755 ;
  assign n53240 = n37673 | n47041 ;
  assign n53241 = n11196 & ~n53240 ;
  assign n53242 = n3514 | n12855 ;
  assign n53243 = n33018 ^ n9919 ^ 1'b0 ;
  assign n53244 = n7535 ^ n854 ^ 1'b0 ;
  assign n53245 = n28378 | n53244 ;
  assign n53246 = ~n15736 & n53245 ;
  assign n53247 = ~n12847 & n16319 ;
  assign n53248 = n18675 | n38580 ;
  assign n53250 = n33706 ^ n16499 ^ 1'b0 ;
  assign n53251 = ~n7522 & n53250 ;
  assign n53249 = n7506 ^ n3455 ^ 1'b0 ;
  assign n53252 = n53251 ^ n53249 ^ n6394 ;
  assign n53253 = ~n170 & n32395 ;
  assign n53254 = ~n7101 & n16316 ;
  assign n53255 = n38216 & n53254 ;
  assign n53256 = n38218 ^ n20955 ^ 1'b0 ;
  assign n53257 = ~n53255 & n53256 ;
  assign n53258 = ~n3011 & n53257 ;
  assign n53259 = ~n41296 & n53258 ;
  assign n53260 = n15338 & ~n21191 ;
  assign n53261 = n53260 ^ n38060 ^ 1'b0 ;
  assign n53262 = n8443 & ~n26139 ;
  assign n53263 = n53262 ^ n48726 ^ 1'b0 ;
  assign n53264 = n6524 & ~n39962 ;
  assign n53265 = n53264 ^ n7291 ^ 1'b0 ;
  assign n53266 = n25927 ^ n16402 ^ n517 ;
  assign n53267 = ( n4503 & n8345 ) | ( n4503 & ~n37716 ) | ( n8345 & ~n37716 ) ;
  assign n53268 = n11495 ^ n4745 ^ 1'b0 ;
  assign n53269 = n7739 | n53268 ;
  assign n53270 = n53269 ^ n47126 ^ 1'b0 ;
  assign n53271 = n5346 & n50409 ;
  assign n53272 = ~n4004 & n53271 ;
  assign n53273 = n53272 ^ n33947 ^ 1'b0 ;
  assign n53274 = ( ~n39168 & n53270 ) | ( ~n39168 & n53273 ) | ( n53270 & n53273 ) ;
  assign n53275 = n28573 & ~n29071 ;
  assign n53276 = n15173 & n24909 ;
  assign n53277 = n34996 & ~n53276 ;
  assign n53282 = ~n24580 & n52676 ;
  assign n53283 = n53282 ^ n3656 ^ 1'b0 ;
  assign n53284 = ~n3920 & n53283 ;
  assign n53279 = n37013 ^ n22869 ^ 1'b0 ;
  assign n53280 = n8676 & n53279 ;
  assign n53278 = ~n1500 & n50448 ;
  assign n53281 = n53280 ^ n53278 ^ 1'b0 ;
  assign n53285 = n53284 ^ n53281 ^ 1'b0 ;
  assign n53286 = n26184 | n29312 ;
  assign n53287 = n53286 ^ n46349 ^ 1'b0 ;
  assign n53288 = n28096 ^ n15077 ^ n7025 ;
  assign n53289 = n53288 ^ n28604 ^ 1'b0 ;
  assign n53291 = n27729 ^ n580 ^ 1'b0 ;
  assign n53290 = n11173 & n43141 ;
  assign n53292 = n53291 ^ n53290 ^ n17334 ;
  assign n53293 = n34810 ^ n10711 ^ 1'b0 ;
  assign n53294 = n35794 ^ n21679 ^ 1'b0 ;
  assign n53295 = ~n22814 & n53294 ;
  assign n53296 = n53295 ^ n19948 ^ 1'b0 ;
  assign n53297 = n53293 & n53296 ;
  assign n53298 = n8362 ^ n5823 ^ 1'b0 ;
  assign n53299 = n10948 | n53298 ;
  assign n53300 = n51154 & n53299 ;
  assign n53301 = n53300 ^ n15076 ^ 1'b0 ;
  assign n53302 = n1586 & n18200 ;
  assign n53303 = n53301 & n53302 ;
  assign n53304 = n12637 & ~n21331 ;
  assign n53305 = ~n3256 & n53304 ;
  assign n53306 = ~n42701 & n52765 ;
  assign n53307 = n7627 | n20727 ;
  assign n53308 = n53307 ^ n16176 ^ 1'b0 ;
  assign n53309 = n13332 & n53308 ;
  assign n53311 = n25596 ^ n22987 ^ 1'b0 ;
  assign n53310 = n32770 ^ n3506 ^ 1'b0 ;
  assign n53312 = n53311 ^ n53310 ^ n9020 ;
  assign n53315 = n26845 ^ n7322 ^ 1'b0 ;
  assign n53313 = n6375 | n16445 ;
  assign n53314 = n53313 ^ n39417 ^ 1'b0 ;
  assign n53316 = n53315 ^ n53314 ^ n23379 ;
  assign n53317 = n36640 & n52725 ;
  assign n53318 = n53316 & n53317 ;
  assign n53319 = n20086 ^ n3638 ^ 1'b0 ;
  assign n53320 = ~n35963 & n53319 ;
  assign n53321 = n53320 ^ n49745 ^ 1'b0 ;
  assign n53323 = ( n14608 & n24348 ) | ( n14608 & ~n48209 ) | ( n24348 & ~n48209 ) ;
  assign n53322 = ~n1367 & n4239 ;
  assign n53324 = n53323 ^ n53322 ^ 1'b0 ;
  assign n53325 = ~n5423 & n10391 ;
  assign n53326 = n53325 ^ n15765 ^ 1'b0 ;
  assign n53327 = ~n53324 & n53326 ;
  assign n53328 = n9967 & ~n52616 ;
  assign n53329 = n1492 & n53328 ;
  assign n53330 = n18585 & n53329 ;
  assign n53331 = n50950 ^ n31288 ^ n1933 ;
  assign n53332 = n53330 & ~n53331 ;
  assign n53333 = n47800 ^ n34887 ^ 1'b0 ;
  assign n53334 = n8305 & ~n26571 ;
  assign n53335 = n10288 & ~n29454 ;
  assign n53336 = n6402 & n53335 ;
  assign n53337 = n6060 & n10269 ;
  assign n53338 = ( n6551 & n9706 ) | ( n6551 & n53337 ) | ( n9706 & n53337 ) ;
  assign n53339 = ~n9162 & n25276 ;
  assign n53340 = ~n20859 & n53339 ;
  assign n53341 = ( n51252 & n53338 ) | ( n51252 & n53340 ) | ( n53338 & n53340 ) ;
  assign n53342 = n12683 & n36541 ;
  assign n53343 = ( n15520 & n16440 ) | ( n15520 & ~n38713 ) | ( n16440 & ~n38713 ) ;
  assign n53344 = n46852 & n53343 ;
  assign n53345 = n53342 & n53344 ;
  assign n53346 = n12439 & ~n36791 ;
  assign n53347 = n53346 ^ n1351 ^ 1'b0 ;
  assign n53350 = n30416 | n33713 ;
  assign n53348 = n2904 | n34746 ;
  assign n53349 = ~n9145 & n53348 ;
  assign n53351 = n53350 ^ n53349 ^ 1'b0 ;
  assign n53352 = n32995 & ~n35434 ;
  assign n53353 = n53352 ^ n1936 ^ 1'b0 ;
  assign n53354 = n6324 & n53353 ;
  assign n53355 = n3441 & n10213 ;
  assign n53356 = ~n4745 & n53355 ;
  assign n53357 = n52507 & ~n53356 ;
  assign n53358 = n41621 ^ n20057 ^ 1'b0 ;
  assign n53359 = ( ~n18210 & n19646 ) | ( ~n18210 & n30227 ) | ( n19646 & n30227 ) ;
  assign n53360 = n42522 | n53359 ;
  assign n53361 = n976 & ~n7888 ;
  assign n53362 = n53361 ^ n1276 ^ 1'b0 ;
  assign n53363 = n39657 ^ n28906 ^ 1'b0 ;
  assign n53364 = n53362 | n53363 ;
  assign n53365 = n10163 & n14875 ;
  assign n53366 = ~n5380 & n39671 ;
  assign n53367 = n53366 ^ n4356 ^ 1'b0 ;
  assign n53368 = ~n3216 & n21411 ;
  assign n53369 = n2327 & n53368 ;
  assign n53370 = n46376 ^ n41519 ^ n16806 ;
  assign n53371 = n13486 & n39946 ;
  assign n53372 = ~n1444 & n53371 ;
  assign n53373 = n3441 & ~n48738 ;
  assign n53374 = n53373 ^ n5706 ^ 1'b0 ;
  assign n53375 = n49827 & ~n53374 ;
  assign n53376 = n49754 & n53375 ;
  assign n53377 = n32619 | n41563 ;
  assign n53378 = n24185 ^ n1290 ^ 1'b0 ;
  assign n53379 = n53377 & n53378 ;
  assign n53380 = n14429 & n39488 ;
  assign n53381 = n31348 & n53380 ;
  assign n53382 = n31174 & ~n53381 ;
  assign n53383 = n16402 | n42322 ;
  assign n53384 = n53382 | n53383 ;
  assign n53385 = n20781 & ~n51153 ;
  assign n53386 = n53385 ^ n28008 ^ 1'b0 ;
  assign n53387 = n33372 ^ n12860 ^ 1'b0 ;
  assign n53388 = ( n12789 & n19256 ) | ( n12789 & ~n26289 ) | ( n19256 & ~n26289 ) ;
  assign n53389 = n7812 & n16925 ;
  assign n53390 = n17876 ^ n12289 ^ 1'b0 ;
  assign n53391 = n39764 ^ n9226 ^ 1'b0 ;
  assign n53392 = ~n15704 & n51915 ;
  assign n53393 = n11533 & n43904 ;
  assign n53394 = n24761 | n34712 ;
  assign n53395 = n53394 ^ n9838 ^ 1'b0 ;
  assign n53396 = n4096 & ~n4834 ;
  assign n53397 = n1684 | n3245 ;
  assign n53398 = n18828 | n53397 ;
  assign n53399 = n36113 & n53398 ;
  assign n53401 = ~n7536 & n20008 ;
  assign n53400 = n27668 ^ n15737 ^ n12328 ;
  assign n53402 = n53401 ^ n53400 ^ n1319 ;
  assign n53403 = n115 & ~n1105 ;
  assign n53404 = ~n115 & n53403 ;
  assign n53405 = n2471 | n53404 ;
  assign n53406 = n53405 ^ n37004 ^ n4654 ;
  assign n53407 = n13842 & ~n53406 ;
  assign n53408 = n53406 & n53407 ;
  assign n53409 = ( n17136 & n26799 ) | ( n17136 & ~n53408 ) | ( n26799 & ~n53408 ) ;
  assign n53410 = n17712 | n22472 ;
  assign n53411 = n45829 ^ n852 ^ 1'b0 ;
  assign n53412 = n15154 & ~n53411 ;
  assign n53413 = n4953 ^ n63 ^ 1'b0 ;
  assign n53414 = n36346 ^ n25728 ^ 1'b0 ;
  assign n53415 = n13813 & ~n41292 ;
  assign n53416 = n53415 ^ n53313 ^ 1'b0 ;
  assign n53417 = n2239 | n8912 ;
  assign n53418 = n53417 ^ n13097 ^ 1'b0 ;
  assign n53419 = n28534 & ~n35342 ;
  assign n53420 = n11753 & ~n48851 ;
  assign n53421 = n34232 ^ n24518 ^ n20724 ;
  assign n53422 = n21867 ^ n13546 ^ 1'b0 ;
  assign n53423 = n19246 ^ n9899 ^ n4787 ;
  assign n53424 = ~n9782 & n23795 ;
  assign n53425 = n7900 & n53424 ;
  assign n53426 = n11729 & ~n13633 ;
  assign n53427 = n1312 & n53426 ;
  assign n53428 = n35035 ^ n2696 ^ 1'b0 ;
  assign n53429 = n53428 ^ n48417 ^ 1'b0 ;
  assign n53430 = ~n951 & n8427 ;
  assign n53431 = n53430 ^ n28827 ^ 1'b0 ;
  assign n53432 = n24662 | n31011 ;
  assign n53433 = n14009 | n53432 ;
  assign n53434 = ( n1310 & n14370 ) | ( n1310 & ~n33881 ) | ( n14370 & ~n33881 ) ;
  assign n53435 = n53434 ^ n48801 ^ n5645 ;
  assign n53436 = n24115 ^ x1 ^ 1'b0 ;
  assign n53437 = n16130 & n53436 ;
  assign n53438 = n20710 & ~n53437 ;
  assign n53439 = n18875 ^ n16099 ^ 1'b0 ;
  assign n53440 = n53439 ^ n25627 ^ n23423 ;
  assign n53441 = ~n2855 & n34891 ;
  assign n53442 = ~n17979 & n53441 ;
  assign n53443 = n12366 ^ n8428 ^ n1289 ;
  assign n53444 = n50127 & n53443 ;
  assign n53445 = n53444 ^ n17147 ^ 1'b0 ;
  assign n53446 = n15256 & ~n47911 ;
  assign n53447 = n53446 ^ n8858 ^ 1'b0 ;
  assign n53448 = n13067 | n14057 ;
  assign n53449 = n15672 & ~n53448 ;
  assign n53450 = n53449 ^ n8254 ^ 1'b0 ;
  assign n53451 = n53447 & ~n53450 ;
  assign n53454 = n8330 | n49938 ;
  assign n53455 = n2705 | n53454 ;
  assign n53452 = n254 & ~n1409 ;
  assign n53453 = n21267 & n53452 ;
  assign n53456 = n53455 ^ n53453 ^ n27935 ;
  assign n53457 = n9819 & n21775 ;
  assign n53459 = n12894 & ~n35909 ;
  assign n53460 = ~n14682 & n53459 ;
  assign n53461 = n34931 | n53460 ;
  assign n53458 = ( n620 & ~n7260 ) | ( n620 & n53455 ) | ( ~n7260 & n53455 ) ;
  assign n53462 = n53461 ^ n53458 ^ n2140 ;
  assign n53463 = ( ~n25088 & n25283 ) | ( ~n25088 & n37351 ) | ( n25283 & n37351 ) ;
  assign n53464 = n5509 & ~n53463 ;
  assign n53465 = ~n26783 & n53464 ;
  assign n53466 = n8008 | n49780 ;
  assign n53467 = n53466 ^ n18654 ^ 1'b0 ;
  assign n53468 = n19529 ^ n154 ^ 1'b0 ;
  assign n53469 = n39702 ^ n22612 ^ 1'b0 ;
  assign n53470 = n53468 & ~n53469 ;
  assign n53471 = ~n6740 & n10263 ;
  assign n53472 = n2408 & n53471 ;
  assign n53473 = ~n3473 & n18003 ;
  assign n53474 = n8929 & n53473 ;
  assign n53475 = ~n53472 & n53474 ;
  assign n53476 = n17738 ^ n16261 ^ 1'b0 ;
  assign n53477 = n23 & ~n53476 ;
  assign n53478 = n52335 ^ n1411 ^ 1'b0 ;
  assign n53479 = ~n12451 & n24038 ;
  assign n53480 = n48944 | n53479 ;
  assign n53481 = n53480 ^ n7055 ^ 1'b0 ;
  assign n53482 = n17558 & ~n53481 ;
  assign n53483 = ~n5781 & n8647 ;
  assign n53484 = n53483 ^ n15009 ^ 1'b0 ;
  assign n53485 = ( ~n3863 & n37553 ) | ( ~n3863 & n53484 ) | ( n37553 & n53484 ) ;
  assign n53486 = n53485 ^ n52271 ^ n37011 ;
  assign n53487 = ~n6368 & n19431 ;
  assign n53488 = ~n6105 & n53487 ;
  assign n53489 = n53488 ^ n82 ^ 1'b0 ;
  assign n53490 = n53489 ^ n37224 ^ 1'b0 ;
  assign n53491 = n53490 ^ n42915 ^ 1'b0 ;
  assign n53492 = n19450 & n23411 ;
  assign n53493 = n53492 ^ n45627 ^ 1'b0 ;
  assign n53495 = n42322 ^ n19614 ^ 1'b0 ;
  assign n53494 = n209 & n37068 ;
  assign n53496 = n53495 ^ n53494 ^ 1'b0 ;
  assign n53497 = n43404 | n44790 ;
  assign n53498 = ( n2648 & n6795 ) | ( n2648 & n13522 ) | ( n6795 & n13522 ) ;
  assign n53499 = n29113 & ~n29207 ;
  assign n53500 = n53499 ^ n48455 ^ 1'b0 ;
  assign n53501 = n30776 ^ n18909 ^ n6497 ;
  assign n53502 = n2050 & n53501 ;
  assign n53503 = n53502 ^ n10154 ^ 1'b0 ;
  assign n53504 = n40328 ^ n33253 ^ 1'b0 ;
  assign n53505 = n49030 ^ n22419 ^ n10002 ;
  assign n53506 = n30138 ^ n982 ^ 1'b0 ;
  assign n53507 = n53506 ^ n23569 ^ 1'b0 ;
  assign n53508 = n36367 | n53507 ;
  assign n53509 = n19195 & ~n38948 ;
  assign n53510 = n46625 & n53509 ;
  assign n53511 = n6481 & n14978 ;
  assign n53512 = n53511 ^ n26109 ^ 1'b0 ;
  assign n53513 = ~n44358 & n53512 ;
  assign n53514 = n17338 ^ n3593 ^ 1'b0 ;
  assign n53515 = n53513 & ~n53514 ;
  assign n53516 = n53479 ^ n13903 ^ 1'b0 ;
  assign n53517 = n32358 ^ n12707 ^ n5186 ;
  assign n53518 = n53517 ^ n3731 ^ 1'b0 ;
  assign n53519 = n50942 ^ n33099 ^ 1'b0 ;
  assign n53520 = n453 | n29196 ;
  assign n53521 = n7374 | n53520 ;
  assign n53522 = n53521 ^ n20638 ^ 1'b0 ;
  assign n53523 = n53522 ^ n20292 ^ 1'b0 ;
  assign n53524 = n1311 | n1962 ;
  assign n53525 = n5131 & ~n53524 ;
  assign n53526 = n11570 & n53525 ;
  assign n53527 = n37565 | n53526 ;
  assign n53528 = n13722 ^ n3614 ^ 1'b0 ;
  assign n53531 = n4670 & ~n5562 ;
  assign n53529 = ~n3773 & n7649 ;
  assign n53530 = ~n2425 & n53529 ;
  assign n53532 = n53531 ^ n53530 ^ 1'b0 ;
  assign n53533 = n29643 & n53532 ;
  assign n53534 = n52804 ^ n9601 ^ 1'b0 ;
  assign n53535 = n5570 & ~n14702 ;
  assign n53536 = n9586 ^ n4572 ^ 1'b0 ;
  assign n53537 = n53535 & n53536 ;
  assign n53538 = n43624 ^ n16313 ^ n10511 ;
  assign n53539 = n53136 ^ n25199 ^ 1'b0 ;
  assign n53540 = n41518 & n53539 ;
  assign n53541 = ~n53538 & n53540 ;
  assign n53542 = n41550 & ~n53541 ;
  assign n53543 = ( ~n21996 & n45207 ) | ( ~n21996 & n51947 ) | ( n45207 & n51947 ) ;
  assign n53544 = n53543 ^ n20316 ^ n11759 ;
  assign n53545 = ~n7858 & n8337 ;
  assign n53546 = ~n28120 & n53545 ;
  assign n53547 = n3581 & ~n53546 ;
  assign n53548 = ~n38289 & n53547 ;
  assign n53549 = n46102 ^ n35162 ^ 1'b0 ;
  assign n53550 = ( n47256 & n53548 ) | ( n47256 & n53549 ) | ( n53548 & n53549 ) ;
  assign n53551 = n10993 & n26035 ;
  assign n53552 = n53551 ^ n37013 ^ n6073 ;
  assign n53553 = ~n4888 & n29532 ;
  assign n53554 = ~n10042 & n26391 ;
  assign n53555 = ~n47166 & n53554 ;
  assign n53559 = n37591 ^ n8536 ^ n2677 ;
  assign n53556 = n25625 & ~n41759 ;
  assign n53557 = ~n13180 & n53556 ;
  assign n53558 = n9734 & ~n53557 ;
  assign n53560 = n53559 ^ n53558 ^ 1'b0 ;
  assign n53561 = n13496 ^ n1865 ^ 1'b0 ;
  assign n53562 = n30021 ^ n22090 ^ 1'b0 ;
  assign n53563 = n49731 & n53562 ;
  assign n53564 = n53561 | n53563 ;
  assign n53565 = n8641 & ~n36708 ;
  assign n53566 = n21005 | n38917 ;
  assign n53567 = n19041 ^ n12375 ^ n686 ;
  assign n53568 = ( n14979 & ~n17608 ) | ( n14979 & n53567 ) | ( ~n17608 & n53567 ) ;
  assign n53569 = n5715 ^ n332 ^ 1'b0 ;
  assign n53570 = n14456 ^ n7790 ^ 1'b0 ;
  assign n53571 = n53570 ^ n41856 ^ 1'b0 ;
  assign n53572 = ~n53569 & n53571 ;
  assign n53573 = n5506 & n37788 ;
  assign n53574 = n53573 ^ n19743 ^ 1'b0 ;
  assign n53575 = ( n42157 & n53572 ) | ( n42157 & n53574 ) | ( n53572 & n53574 ) ;
  assign n53576 = n5722 | n17927 ;
  assign n53577 = n18804 ^ n9049 ^ 1'b0 ;
  assign n53578 = n4088 | n53577 ;
  assign n53579 = n43610 ^ n43227 ^ 1'b0 ;
  assign n53580 = n98 | n37674 ;
  assign n53581 = n16284 | n53580 ;
  assign n53582 = n18664 & ~n53581 ;
  assign n53583 = n53579 & n53582 ;
  assign n53584 = n2317 | n4859 ;
  assign n53586 = ~n24408 & n40579 ;
  assign n53585 = n14116 & n14296 ;
  assign n53587 = n53586 ^ n53585 ^ 1'b0 ;
  assign n53588 = n23923 & n43436 ;
  assign n53589 = n16374 | n16542 ;
  assign n53590 = n53589 ^ n24647 ^ 1'b0 ;
  assign n53591 = n3389 ^ n375 ^ 1'b0 ;
  assign n53592 = ~n10312 & n53591 ;
  assign n53593 = n53592 ^ n2873 ^ 1'b0 ;
  assign n53594 = n18680 ^ n14335 ^ 1'b0 ;
  assign n53595 = n18164 ^ n10436 ^ 1'b0 ;
  assign n53596 = n53595 ^ n35561 ^ 1'b0 ;
  assign n53597 = n19957 & ~n35335 ;
  assign n53598 = n53597 ^ n17068 ^ 1'b0 ;
  assign n53599 = n2766 | n6758 ;
  assign n53600 = n53599 ^ n24300 ^ 1'b0 ;
  assign n53601 = ~n11811 & n13296 ;
  assign n53602 = n31717 ^ n10406 ^ 1'b0 ;
  assign n53603 = n53601 & ~n53602 ;
  assign n53604 = n30164 ^ n27117 ^ n25761 ;
  assign n53605 = n53603 & n53604 ;
  assign n53606 = ( n19856 & n41287 ) | ( n19856 & n42891 ) | ( n41287 & n42891 ) ;
  assign n53607 = n18692 & n35762 ;
  assign n53608 = n53607 ^ n28786 ^ n22720 ;
  assign n53609 = n24473 ^ n11746 ^ 1'b0 ;
  assign n53610 = n1918 & ~n53609 ;
  assign n53611 = n43531 & ~n46393 ;
  assign n53612 = n26336 & n28380 ;
  assign n53613 = n18322 | n20954 ;
  assign n53614 = n16935 & ~n53613 ;
  assign n53615 = n21807 ^ n2934 ^ 1'b0 ;
  assign n53616 = ~n30317 & n53615 ;
  assign n53617 = n6150 & n6771 ;
  assign n53618 = n18387 & ~n53617 ;
  assign n53619 = n34424 ^ n33501 ^ n5022 ;
  assign n53620 = n4658 & ~n42715 ;
  assign n53621 = n53620 ^ n41837 ^ 1'b0 ;
  assign n53622 = n25812 ^ n5604 ^ 1'b0 ;
  assign n53623 = ~n22556 & n53622 ;
  assign n53624 = n16260 & ~n34828 ;
  assign n53625 = n53624 ^ n15203 ^ 1'b0 ;
  assign n53626 = n8056 & n33725 ;
  assign n53627 = n13986 & n53626 ;
  assign n53628 = ( n12529 & ~n28375 ) | ( n12529 & n46694 ) | ( ~n28375 & n46694 ) ;
  assign n53629 = n53628 ^ n2747 ^ 1'b0 ;
  assign n53630 = n14711 | n53629 ;
  assign n53631 = n49492 | n53630 ;
  assign n53632 = n11531 ^ n5537 ^ 1'b0 ;
  assign n53633 = n43810 | n53632 ;
  assign n53634 = n11753 | n23070 ;
  assign n53635 = ( n5010 & n41885 ) | ( n5010 & n53634 ) | ( n41885 & n53634 ) ;
  assign n53636 = ~n21781 & n25131 ;
  assign n53639 = n27645 ^ n18726 ^ n14675 ;
  assign n53638 = n38614 ^ n36333 ^ 1'b0 ;
  assign n53637 = n31224 ^ n919 ^ 1'b0 ;
  assign n53640 = n53639 ^ n53638 ^ n53637 ;
  assign n53641 = n28402 ^ n11295 ^ 1'b0 ;
  assign n53642 = ~n15593 & n53641 ;
  assign n53643 = n53642 ^ n3248 ^ 1'b0 ;
  assign n53644 = ~n4305 & n7354 ;
  assign n53645 = n4221 & n13680 ;
  assign n53646 = n53645 ^ n25968 ^ 1'b0 ;
  assign n53647 = n53646 ^ n25253 ^ n12789 ;
  assign n53648 = n53647 ^ n39182 ^ 1'b0 ;
  assign n53649 = ~n3471 & n11379 ;
  assign n53650 = n53648 & n53649 ;
  assign n53651 = n5372 & n8902 ;
  assign n53652 = n5850 | n53651 ;
  assign n53653 = n53652 ^ n47283 ^ n10329 ;
  assign n53655 = ( n659 & n1509 ) | ( n659 & n50378 ) | ( n1509 & n50378 ) ;
  assign n53656 = n18977 & ~n53655 ;
  assign n53657 = n53656 ^ n21078 ^ 1'b0 ;
  assign n53654 = n53452 ^ n42837 ^ 1'b0 ;
  assign n53658 = n53657 ^ n53654 ^ 1'b0 ;
  assign n53659 = ~n14873 & n19780 ;
  assign n53660 = ~n115 & n53659 ;
  assign n53661 = n2568 & ~n53660 ;
  assign n53662 = n53661 ^ n39832 ^ n960 ;
  assign n53663 = n4512 ^ n44 ^ 1'b0 ;
  assign n53664 = n3478 | n53663 ;
  assign n53665 = n20357 & n53664 ;
  assign n53666 = n12063 & ~n12071 ;
  assign n53667 = n43590 & n53666 ;
  assign n53668 = n2330 & ~n4553 ;
  assign n53669 = n50115 & n53668 ;
  assign n53670 = n34828 ^ n29970 ^ 1'b0 ;
  assign n53671 = n20968 ^ n3987 ^ 1'b0 ;
  assign n53672 = n49899 ^ n16635 ^ 1'b0 ;
  assign n53673 = n2901 & ~n53672 ;
  assign n53674 = n1772 & ~n14736 ;
  assign n53675 = n44457 & ~n53674 ;
  assign n53676 = ( n1728 & n17979 ) | ( n1728 & ~n18136 ) | ( n17979 & ~n18136 ) ;
  assign n53677 = n16828 | n45433 ;
  assign n53678 = n23299 & n53677 ;
  assign n53679 = ~n11914 & n36651 ;
  assign n53684 = n37746 ^ n30356 ^ n2977 ;
  assign n53680 = n19703 ^ n15687 ^ n2216 ;
  assign n53681 = n35433 ^ n15408 ^ 1'b0 ;
  assign n53682 = ( n18531 & n53680 ) | ( n18531 & ~n53681 ) | ( n53680 & ~n53681 ) ;
  assign n53683 = n19997 & n53682 ;
  assign n53685 = n53684 ^ n53683 ^ 1'b0 ;
  assign n53686 = ~n6441 & n10819 ;
  assign n53687 = n53686 ^ n17712 ^ 1'b0 ;
  assign n53688 = n514 & ~n53687 ;
  assign n53689 = ~n4949 & n12286 ;
  assign n53690 = ~n1095 & n53689 ;
  assign n53691 = n33168 ^ n11740 ^ 1'b0 ;
  assign n53692 = n16452 | n51769 ;
  assign n53693 = ( n22645 & n50329 ) | ( n22645 & n53692 ) | ( n50329 & n53692 ) ;
  assign n53694 = n16540 & n17162 ;
  assign n53695 = n32848 ^ n17226 ^ 1'b0 ;
  assign n53696 = n10701 & ~n53695 ;
  assign n53697 = n10501 & n25903 ;
  assign n53698 = n53697 ^ n42511 ^ 1'b0 ;
  assign n53699 = n585 | n53698 ;
  assign n53700 = n10962 | n31846 ;
  assign n53701 = n53700 ^ n4977 ^ 1'b0 ;
  assign n53702 = n5722 & n40570 ;
  assign n53703 = n49689 & n53702 ;
  assign n53704 = n48547 ^ n15013 ^ 1'b0 ;
  assign n53705 = n12576 ^ n6954 ^ 1'b0 ;
  assign n53706 = n6820 & ~n53705 ;
  assign n53707 = n11810 & ~n42844 ;
  assign n53708 = n17077 & n53707 ;
  assign n53709 = ( ~n27489 & n53706 ) | ( ~n27489 & n53708 ) | ( n53706 & n53708 ) ;
  assign n53710 = ( ~n2218 & n13228 ) | ( ~n2218 & n30608 ) | ( n13228 & n30608 ) ;
  assign n53711 = n9548 | n23837 ;
  assign n53712 = ~n523 & n24443 ;
  assign n53713 = n53712 ^ n601 ^ 1'b0 ;
  assign n53714 = n16409 | n53713 ;
  assign n53715 = n4265 & n22907 ;
  assign n53716 = ~n10971 & n27472 ;
  assign n53717 = n3737 & n53716 ;
  assign n53718 = n53717 ^ n17401 ^ 1'b0 ;
  assign n53719 = ~n13391 & n53718 ;
  assign n53720 = n14996 & n40096 ;
  assign n53721 = n11593 & n22515 ;
  assign n53722 = n53721 ^ n37776 ^ 1'b0 ;
  assign n53723 = n33833 | n34398 ;
  assign n53724 = n53723 ^ n4957 ^ 1'b0 ;
  assign n53725 = ~n14145 & n53724 ;
  assign n53726 = ( n6287 & n7119 ) | ( n6287 & ~n19869 ) | ( n7119 & ~n19869 ) ;
  assign n53727 = n53726 ^ n28749 ^ n8073 ;
  assign n53728 = n21336 ^ n11902 ^ n293 ;
  assign n53729 = n47533 ^ n32567 ^ 1'b0 ;
  assign n53730 = n51385 & ~n53729 ;
  assign n53731 = ~n16089 & n36529 ;
  assign n53732 = n18672 ^ n14231 ^ 1'b0 ;
  assign n53733 = n49782 | n53732 ;
  assign n53734 = n11492 ^ n7099 ^ n3738 ;
  assign n53735 = n4173 | n14731 ;
  assign n53736 = n18626 & n19450 ;
  assign n53737 = n53736 ^ n50343 ^ 1'b0 ;
  assign n53738 = ~n5450 & n14492 ;
  assign n53739 = n49540 & n53738 ;
  assign n53740 = n53737 & n53739 ;
  assign n53741 = n27602 ^ n10212 ^ 1'b0 ;
  assign n53742 = n21679 | n53741 ;
  assign n53743 = ~n5356 & n23290 ;
  assign n53744 = ~n7104 & n53743 ;
  assign n53745 = n5353 & n9293 ;
  assign n53746 = n53744 & n53745 ;
  assign n53747 = n16915 & ~n17308 ;
  assign n53748 = n34969 ^ n20086 ^ 1'b0 ;
  assign n53749 = n21775 | n53748 ;
  assign n53750 = n6191 | n53749 ;
  assign n53751 = n53750 ^ n9470 ^ 1'b0 ;
  assign n53752 = ( n11718 & n35198 ) | ( n11718 & n52040 ) | ( n35198 & n52040 ) ;
  assign n53753 = n11503 & ~n53752 ;
  assign n53754 = ~n10999 & n53753 ;
  assign n53755 = ~n5696 & n13533 ;
  assign n53756 = n53755 ^ n5078 ^ 1'b0 ;
  assign n53757 = n53756 ^ n28737 ^ 1'b0 ;
  assign n53758 = n26012 & n44475 ;
  assign n53759 = n6888 & ~n53758 ;
  assign n53760 = n4168 & n53759 ;
  assign n53761 = n3964 & n40800 ;
  assign n53762 = n53761 ^ n41816 ^ n2661 ;
  assign n53763 = n10974 ^ n6674 ^ 1'b0 ;
  assign n53764 = ~n23733 & n53763 ;
  assign n53765 = ( n4966 & n19418 ) | ( n4966 & ~n36621 ) | ( n19418 & ~n36621 ) ;
  assign n53766 = ~n3161 & n22653 ;
  assign n53767 = n2256 | n5414 ;
  assign n53768 = n53766 & ~n53767 ;
  assign n53769 = n52899 ^ n21741 ^ 1'b0 ;
  assign n53770 = n40779 ^ n14857 ^ 1'b0 ;
  assign n53772 = n26410 ^ n6676 ^ 1'b0 ;
  assign n53773 = n22068 & ~n53772 ;
  assign n53771 = ~n18171 & n31173 ;
  assign n53774 = n53773 ^ n53771 ^ 1'b0 ;
  assign n53775 = n41141 ^ n22584 ^ 1'b0 ;
  assign n53776 = n12139 & n53775 ;
  assign n53777 = n4231 & n31870 ;
  assign n53778 = ~n53776 & n53777 ;
  assign n53782 = n36519 ^ n31132 ^ n15618 ;
  assign n53779 = ~n4590 & n13110 ;
  assign n53780 = n2807 & n53779 ;
  assign n53781 = n21202 | n53780 ;
  assign n53783 = n53782 ^ n53781 ^ 1'b0 ;
  assign n53784 = n29593 | n32468 ;
  assign n53785 = n8103 & ~n13028 ;
  assign n53786 = n53785 ^ n21184 ^ n1138 ;
  assign n53788 = n28290 | n33896 ;
  assign n53789 = n12290 | n53788 ;
  assign n53790 = n10333 & ~n53789 ;
  assign n53791 = n16797 ^ n272 ^ 1'b0 ;
  assign n53792 = ~n53790 & n53791 ;
  assign n53787 = n19080 | n19807 ;
  assign n53793 = n53792 ^ n53787 ^ 1'b0 ;
  assign n53794 = n53793 ^ n38287 ^ 1'b0 ;
  assign n53795 = n53794 ^ n3142 ^ 1'b0 ;
  assign n53796 = n53795 ^ n16661 ^ 1'b0 ;
  assign n53797 = n33001 ^ n29955 ^ 1'b0 ;
  assign n53798 = ~n18444 & n53797 ;
  assign n53799 = n8241 & n50832 ;
  assign n53800 = n38916 & ~n45530 ;
  assign n53801 = n53800 ^ n40604 ^ 1'b0 ;
  assign n53802 = n53801 ^ n7235 ^ 1'b0 ;
  assign n53803 = n53799 & n53802 ;
  assign n53804 = n21532 ^ n5239 ^ 1'b0 ;
  assign n53805 = ~n42317 & n53804 ;
  assign n53806 = ~n37292 & n53805 ;
  assign n53807 = n14183 ^ n8130 ^ 1'b0 ;
  assign n53808 = n10878 & n53807 ;
  assign n53809 = n27671 & n53808 ;
  assign n53810 = n7631 ^ n3606 ^ 1'b0 ;
  assign n53811 = n12551 & ~n53810 ;
  assign n53812 = n8630 ^ n2108 ^ 1'b0 ;
  assign n53813 = n48736 | n53812 ;
  assign n53814 = n11717 & n17278 ;
  assign n53815 = ~n26941 & n53814 ;
  assign n53816 = n37877 ^ n5903 ^ 1'b0 ;
  assign n53817 = n10444 ^ n8780 ^ n8026 ;
  assign n53818 = n20509 | n33938 ;
  assign n53819 = n53818 ^ n36744 ^ 1'b0 ;
  assign n53820 = n17980 & n53819 ;
  assign n53821 = ~n46088 & n53820 ;
  assign n53822 = ~n13009 & n13818 ;
  assign n53823 = n53822 ^ n29068 ^ 1'b0 ;
  assign n53824 = n14204 & ~n20151 ;
  assign n53825 = ~n50240 & n53824 ;
  assign n53826 = n24465 ^ n4258 ^ 1'b0 ;
  assign n53827 = n29710 & ~n53826 ;
  assign n53830 = n42403 ^ n17407 ^ n10755 ;
  assign n53828 = n11418 & ~n28917 ;
  assign n53829 = n53828 ^ n4058 ^ 1'b0 ;
  assign n53831 = n53830 ^ n53829 ^ 1'b0 ;
  assign n53832 = n53831 ^ n12239 ^ 1'b0 ;
  assign n53833 = n16083 ^ n9146 ^ n7345 ;
  assign n53834 = ( n17604 & n26717 ) | ( n17604 & ~n46975 ) | ( n26717 & ~n46975 ) ;
  assign n53835 = n13284 & ~n50313 ;
  assign n53836 = ( n5261 & n25368 ) | ( n5261 & n53835 ) | ( n25368 & n53835 ) ;
  assign n53837 = ( n4700 & n38524 ) | ( n4700 & n53313 ) | ( n38524 & n53313 ) ;
  assign n53838 = n9332 & ~n33903 ;
  assign n53839 = n53838 ^ n24718 ^ 1'b0 ;
  assign n53840 = n14500 & ~n45095 ;
  assign n53841 = ( ~n12263 & n38172 ) | ( ~n12263 & n51139 ) | ( n38172 & n51139 ) ;
  assign n53842 = n50444 ^ n23404 ^ 1'b0 ;
  assign n53843 = ~n53841 & n53842 ;
  assign n53844 = n24779 ^ n1311 ^ 1'b0 ;
  assign n53845 = n34443 ^ n3345 ^ 1'b0 ;
  assign n53846 = n53845 ^ n42216 ^ n4368 ;
  assign n53847 = n45710 ^ n3982 ^ 1'b0 ;
  assign n53848 = n6362 | n53847 ;
  assign n53849 = n82 | n521 ;
  assign n53850 = n53849 ^ n27525 ^ n884 ;
  assign n53851 = n8190 & n13037 ;
  assign n53852 = n28374 & n53851 ;
  assign n53853 = n53852 ^ n19389 ^ 1'b0 ;
  assign n53854 = n52004 ^ n46114 ^ 1'b0 ;
  assign n53855 = n15083 & ~n30983 ;
  assign n53856 = n40492 ^ n10451 ^ n3837 ;
  assign n53857 = n25760 ^ n16383 ^ 1'b0 ;
  assign n53858 = ~n17003 & n27295 ;
  assign n53859 = n53858 ^ n4743 ^ 1'b0 ;
  assign n53860 = n20061 ^ n7295 ^ 1'b0 ;
  assign n53861 = ~n37623 & n53860 ;
  assign n53863 = n17683 ^ n6974 ^ n5455 ;
  assign n53862 = n4875 & ~n13543 ;
  assign n53864 = n53863 ^ n53862 ^ 1'b0 ;
  assign n53865 = ~n7376 & n8607 ;
  assign n53866 = n53865 ^ n35521 ^ n6584 ;
  assign n53867 = n53866 ^ n14097 ^ 1'b0 ;
  assign n53868 = n7614 | n53867 ;
  assign n53869 = n13250 & n44780 ;
  assign n53870 = n11023 ^ n5236 ^ 1'b0 ;
  assign n53871 = n12618 & ~n26873 ;
  assign n53872 = n53871 ^ n22391 ^ 1'b0 ;
  assign n53873 = n22776 ^ n11438 ^ 1'b0 ;
  assign n53874 = n5456 | n53873 ;
  assign n53875 = ~n3741 & n29423 ;
  assign n53876 = n35659 ^ n8119 ^ 1'b0 ;
  assign n53877 = ( n20512 & n53875 ) | ( n20512 & n53876 ) | ( n53875 & n53876 ) ;
  assign n53878 = n14808 & n37173 ;
  assign n53879 = n34516 & n43148 ;
  assign n53880 = ~n3455 & n14114 ;
  assign n53881 = n25436 & n53880 ;
  assign n53882 = n12107 | n43259 ;
  assign n53883 = n16918 | n34998 ;
  assign n53884 = n47105 & ~n53883 ;
  assign n53885 = n21671 & ~n51211 ;
  assign n53886 = n4662 | n50125 ;
  assign n53887 = n5160 & ~n53886 ;
  assign n53888 = n11781 ^ n1072 ^ 1'b0 ;
  assign n53889 = n53888 ^ n41209 ^ n30967 ;
  assign n53891 = n23 | n7796 ;
  assign n53892 = n16706 | n53891 ;
  assign n53890 = n1167 & ~n13943 ;
  assign n53893 = n53892 ^ n53890 ^ 1'b0 ;
  assign n53894 = n11458 & n16853 ;
  assign n53896 = n1843 & n15316 ;
  assign n53897 = ( ~n17170 & n25326 ) | ( ~n17170 & n53896 ) | ( n25326 & n53896 ) ;
  assign n53895 = n3866 | n7234 ;
  assign n53898 = n53897 ^ n53895 ^ 1'b0 ;
  assign n53899 = n3708 ^ n3384 ^ n2873 ;
  assign n53900 = n53899 ^ n32119 ^ 1'b0 ;
  assign n53901 = ~n22552 & n53900 ;
  assign n53902 = ~n23554 & n23781 ;
  assign n53903 = ~n39722 & n53902 ;
  assign n53904 = n25576 & ~n45958 ;
  assign n53905 = n53904 ^ n3051 ^ 1'b0 ;
  assign n53907 = n471 | n10040 ;
  assign n53906 = ~n11932 & n15186 ;
  assign n53908 = n53907 ^ n53906 ^ 1'b0 ;
  assign n53909 = n49812 ^ n13139 ^ n5806 ;
  assign n53910 = ( n30966 & n43798 ) | ( n30966 & n47301 ) | ( n43798 & n47301 ) ;
  assign n53911 = n53910 ^ n27979 ^ n15912 ;
  assign n53912 = n11126 & ~n19931 ;
  assign n53913 = n20444 & n53912 ;
  assign n53915 = ~n744 & n24873 ;
  assign n53914 = n5333 & n38233 ;
  assign n53916 = n53915 ^ n53914 ^ 1'b0 ;
  assign n53917 = n29857 ^ n13547 ^ n9029 ;
  assign n53918 = n40314 | n47881 ;
  assign n53919 = n53918 ^ n52430 ^ n5578 ;
  assign n53920 = n25979 ^ n16828 ^ 1'b0 ;
  assign n53924 = n12461 ^ n971 ^ 1'b0 ;
  assign n53922 = n4331 & n22149 ;
  assign n53923 = n53922 ^ n9331 ^ 1'b0 ;
  assign n53925 = n53924 ^ n53923 ^ 1'b0 ;
  assign n53926 = n16554 | n53925 ;
  assign n53921 = n22155 & ~n34918 ;
  assign n53927 = n53926 ^ n53921 ^ 1'b0 ;
  assign n53928 = n4974 & ~n12916 ;
  assign n53929 = n11169 ^ n7092 ^ 1'b0 ;
  assign n53930 = n3348 | n53929 ;
  assign n53931 = n5716 & n53930 ;
  assign n53932 = ~n53928 & n53931 ;
  assign n53933 = ~n7433 & n25010 ;
  assign n53934 = n53933 ^ n40166 ^ 1'b0 ;
  assign n53935 = n18686 ^ n4892 ^ 1'b0 ;
  assign n53936 = n11341 & n53935 ;
  assign n53937 = n24110 ^ n8088 ^ 1'b0 ;
  assign n53938 = n22261 | n53937 ;
  assign n53939 = n53938 ^ n10852 ^ 1'b0 ;
  assign n53940 = n14373 | n52783 ;
  assign n53941 = n18813 ^ n13783 ^ 1'b0 ;
  assign n53942 = n46100 & ~n53941 ;
  assign n53943 = n17501 & n32135 ;
  assign n53944 = n1717 & n53943 ;
  assign n53945 = n36861 & n53944 ;
  assign n53946 = ( ~n20083 & n53942 ) | ( ~n20083 & n53945 ) | ( n53942 & n53945 ) ;
  assign n53947 = ~n2114 & n4733 ;
  assign n53948 = n4545 & n36634 ;
  assign n53949 = n53948 ^ n33764 ^ 1'b0 ;
  assign n53950 = ~n53947 & n53949 ;
  assign n53951 = n20370 ^ n8313 ^ 1'b0 ;
  assign n53952 = ~n22990 & n53951 ;
  assign n53953 = n18745 & n53952 ;
  assign n53954 = ~n33488 & n53953 ;
  assign n53955 = n4719 | n19210 ;
  assign n53956 = n25442 & n31445 ;
  assign n53957 = n21973 & n52753 ;
  assign n53958 = n8509 ^ n1305 ^ 1'b0 ;
  assign n53959 = n53957 & n53958 ;
  assign n53960 = n13379 | n37907 ;
  assign n53961 = n53960 ^ n32888 ^ 1'b0 ;
  assign n53962 = n17166 ^ n6398 ^ 1'b0 ;
  assign n53963 = n11867 & n53962 ;
  assign n53964 = n19140 ^ n8528 ^ 1'b0 ;
  assign n53965 = n1441 & ~n53964 ;
  assign n53966 = n53963 & n53965 ;
  assign n53967 = n53966 ^ n25973 ^ 1'b0 ;
  assign n53968 = n9358 & ~n9683 ;
  assign n53969 = n4167 & ~n15796 ;
  assign n53970 = ( n29560 & n53968 ) | ( n29560 & ~n53969 ) | ( n53968 & ~n53969 ) ;
  assign n53971 = ~n36418 & n47329 ;
  assign n53972 = n53971 ^ n15754 ^ 1'b0 ;
  assign n53973 = n3333 & n53972 ;
  assign n53974 = n53973 ^ n19598 ^ 1'b0 ;
  assign n53975 = n19435 & n33617 ;
  assign n53976 = n20163 ^ n16507 ^ 1'b0 ;
  assign n53978 = n2720 | n47820 ;
  assign n53979 = n32023 | n53978 ;
  assign n53977 = n10149 & n11717 ;
  assign n53980 = n53979 ^ n53977 ^ 1'b0 ;
  assign n53981 = n51580 ^ n6890 ^ 1'b0 ;
  assign n53982 = n11233 & n53981 ;
  assign n53983 = ~n14052 & n29417 ;
  assign n53984 = ( n8715 & ~n16471 ) | ( n8715 & n18612 ) | ( ~n16471 & n18612 ) ;
  assign n53985 = n42077 | n53984 ;
  assign n53987 = n16419 ^ n14518 ^ 1'b0 ;
  assign n53988 = ~n22196 & n53987 ;
  assign n53986 = n35188 & ~n40731 ;
  assign n53989 = n53988 ^ n53986 ^ n23359 ;
  assign n53990 = n12789 & n53989 ;
  assign n53991 = ~n3156 & n42987 ;
  assign n53992 = n299 | n15627 ;
  assign n53993 = ~n52910 & n53992 ;
  assign n53994 = n14439 ^ n10821 ^ 1'b0 ;
  assign n53995 = n19019 ^ n9452 ^ n2919 ;
  assign n53999 = n1702 | n28609 ;
  assign n53996 = n11796 ^ n2873 ^ 1'b0 ;
  assign n53997 = n22161 & n53996 ;
  assign n53998 = n26091 | n53997 ;
  assign n54000 = n53999 ^ n53998 ^ 1'b0 ;
  assign n54001 = ~n53995 & n54000 ;
  assign n54003 = n29140 ^ n14928 ^ 1'b0 ;
  assign n54004 = n2569 | n54003 ;
  assign n54002 = n3778 & ~n4160 ;
  assign n54005 = n54004 ^ n54002 ^ n3375 ;
  assign n54006 = n45306 ^ n1346 ^ 1'b0 ;
  assign n54007 = n2732 & n54006 ;
  assign n54008 = n54007 ^ n36102 ^ 1'b0 ;
  assign n54009 = ~n45379 & n54008 ;
  assign n54010 = ~n20748 & n28721 ;
  assign n54011 = n13738 ^ n2225 ^ 1'b0 ;
  assign n54012 = n17652 ^ n13300 ^ 1'b0 ;
  assign n54013 = n49938 | n54012 ;
  assign n54014 = n18 & n13019 ;
  assign n54015 = n10072 & ~n15338 ;
  assign n54016 = n54015 ^ n5625 ^ 1'b0 ;
  assign n54017 = n11882 ^ n7583 ^ n5793 ;
  assign n54018 = n13644 ^ n6998 ^ 1'b0 ;
  assign n54019 = ( ~n10569 & n21024 ) | ( ~n10569 & n54018 ) | ( n21024 & n54018 ) ;
  assign n54021 = n14045 ^ n217 ^ 1'b0 ;
  assign n54022 = n43793 & ~n54021 ;
  assign n54020 = n1563 & ~n8181 ;
  assign n54023 = n54022 ^ n54020 ^ 1'b0 ;
  assign n54024 = n16393 & n18709 ;
  assign n54025 = ~n13558 & n54024 ;
  assign n54026 = n54025 ^ n39931 ^ 1'b0 ;
  assign n54027 = n2039 & n54026 ;
  assign n54029 = ~n874 & n9239 ;
  assign n54028 = ~n4296 & n19026 ;
  assign n54030 = n54029 ^ n54028 ^ 1'b0 ;
  assign n54031 = n104 | n13489 ;
  assign n54032 = n41186 & ~n52320 ;
  assign n54033 = n54032 ^ n51489 ^ 1'b0 ;
  assign n54034 = n6939 & ~n42043 ;
  assign n54035 = n8143 ^ n3648 ^ 1'b0 ;
  assign n54036 = n11801 & n54035 ;
  assign n54037 = n23841 & ~n54036 ;
  assign n54038 = n47108 ^ n2384 ^ 1'b0 ;
  assign n54039 = n916 & n5852 ;
  assign n54040 = ~n5852 & n54039 ;
  assign n54041 = n54040 ^ n9428 ^ 1'b0 ;
  assign n54042 = n54041 ^ n3321 ^ 1'b0 ;
  assign n54043 = ~n34372 & n54042 ;
  assign n54044 = n20340 ^ n813 ^ 1'b0 ;
  assign n54045 = n5392 | n16660 ;
  assign n54046 = n54045 ^ n40943 ^ 1'b0 ;
  assign n54047 = n54046 ^ n47252 ^ 1'b0 ;
  assign n54048 = n11717 | n44103 ;
  assign n54053 = n29068 ^ n15912 ^ n15622 ;
  assign n54051 = n10292 | n49628 ;
  assign n54052 = n30856 | n54051 ;
  assign n54049 = ~n20335 & n38026 ;
  assign n54050 = n54049 ^ n15437 ^ 1'b0 ;
  assign n54054 = n54053 ^ n54052 ^ n54050 ;
  assign n54055 = n53015 ^ n28706 ^ 1'b0 ;
  assign n54056 = n16874 & n54055 ;
  assign n54057 = n38199 ^ n24910 ^ 1'b0 ;
  assign n54058 = n54056 & ~n54057 ;
  assign n54059 = n15341 & n54058 ;
  assign n54060 = n13140 ^ n3912 ^ n134 ;
  assign n54061 = n1142 & ~n27117 ;
  assign n54062 = n5838 | n10050 ;
  assign n54063 = n54062 ^ n10354 ^ 1'b0 ;
  assign n54064 = ~n32602 & n54063 ;
  assign n54065 = n320 | n54064 ;
  assign n54066 = n1647 | n20525 ;
  assign n54067 = n32903 ^ n19596 ^ n8655 ;
  assign n54068 = ( n7400 & ~n10883 ) | ( n7400 & n54067 ) | ( ~n10883 & n54067 ) ;
  assign n54069 = n1961 | n15590 ;
  assign n54070 = ( ~n2108 & n29548 ) | ( ~n2108 & n54069 ) | ( n29548 & n54069 ) ;
  assign n54071 = n19825 ^ n8557 ^ 1'b0 ;
  assign n54072 = n37567 & n54071 ;
  assign n54073 = ~n5912 & n23605 ;
  assign n54074 = n25275 ^ n11482 ^ 1'b0 ;
  assign n54075 = ~n28029 & n54074 ;
  assign n54076 = n48374 ^ n31402 ^ 1'b0 ;
  assign n54077 = ~n5757 & n13769 ;
  assign n54078 = ~n7019 & n54077 ;
  assign n54079 = ( ~n24553 & n31772 ) | ( ~n24553 & n34647 ) | ( n31772 & n34647 ) ;
  assign n54080 = n8750 ^ n7962 ^ n3634 ;
  assign n54081 = ( n7323 & ~n34181 ) | ( n7323 & n54080 ) | ( ~n34181 & n54080 ) ;
  assign n54082 = n37450 ^ n18595 ^ 1'b0 ;
  assign n54083 = n10147 & n26170 ;
  assign n54084 = n53506 ^ n22299 ^ n15070 ;
  assign n54085 = ~n54083 & n54084 ;
  assign n54086 = n54085 ^ n23804 ^ 1'b0 ;
  assign n54087 = n25358 ^ n23839 ^ 1'b0 ;
  assign n54088 = ~n43959 & n54087 ;
  assign n54089 = n4062 & ~n17514 ;
  assign n54090 = n23622 ^ n6126 ^ 1'b0 ;
  assign n54091 = n33899 & n54090 ;
  assign n54092 = ~n25562 & n36837 ;
  assign n54093 = n41217 & n54092 ;
  assign n54094 = n9818 ^ n4574 ^ 1'b0 ;
  assign n54095 = n54093 | n54094 ;
  assign n54096 = n16256 | n54095 ;
  assign n54097 = n8240 & ~n12233 ;
  assign n54098 = n54097 ^ n29645 ^ 1'b0 ;
  assign n54099 = n43564 & ~n54098 ;
  assign n54107 = ~n1166 & n1907 ;
  assign n54108 = ~n1907 & n54107 ;
  assign n54109 = n567 & n54108 ;
  assign n54110 = n54109 ^ n23941 ^ 1'b0 ;
  assign n54100 = n28355 ^ n15552 ^ 1'b0 ;
  assign n54101 = ~n21679 & n54100 ;
  assign n54102 = n54101 ^ n29774 ^ 1'b0 ;
  assign n54103 = ( ~n1845 & n26114 ) | ( ~n1845 & n54102 ) | ( n26114 & n54102 ) ;
  assign n54104 = n10885 | n20324 ;
  assign n54105 = n54104 ^ n26289 ^ 1'b0 ;
  assign n54106 = n54103 & n54105 ;
  assign n54111 = n54110 ^ n54106 ^ 1'b0 ;
  assign n54112 = n3901 | n29060 ;
  assign n54113 = ~n4463 & n14423 ;
  assign n54114 = n18213 ^ n829 ^ 1'b0 ;
  assign n54115 = ( n2967 & ~n22662 ) | ( n2967 & n44362 ) | ( ~n22662 & n44362 ) ;
  assign n54116 = n27940 ^ n21945 ^ 1'b0 ;
  assign n54117 = n2474 & n54116 ;
  assign n54119 = n28476 ^ n4239 ^ n3124 ;
  assign n54120 = n54119 ^ n19942 ^ 1'b0 ;
  assign n54118 = ~n16005 & n18630 ;
  assign n54121 = n54120 ^ n54118 ^ 1'b0 ;
  assign n54124 = n4801 | n12992 ;
  assign n54122 = n31030 ^ n1822 ^ 1'b0 ;
  assign n54123 = n20285 | n54122 ;
  assign n54125 = n54124 ^ n54123 ^ n16043 ;
  assign n54126 = n51549 ^ n11409 ^ 1'b0 ;
  assign n54127 = n11508 ^ n1676 ^ 1'b0 ;
  assign n54128 = ( n28398 & ~n54126 ) | ( n28398 & n54127 ) | ( ~n54126 & n54127 ) ;
  assign n54129 = n22525 | n28758 ;
  assign n54130 = n24674 | n54129 ;
  assign n54131 = n44373 ^ n16238 ^ 1'b0 ;
  assign n54132 = n54130 & n54131 ;
  assign n54133 = n12985 | n28403 ;
  assign n54134 = n3811 & ~n54133 ;
  assign n54135 = n12547 ^ n716 ^ 1'b0 ;
  assign n54136 = n50173 ^ n2866 ^ 1'b0 ;
  assign n54137 = n54135 & n54136 ;
  assign n54138 = n14545 | n18143 ;
  assign n54139 = n54138 ^ n44584 ^ 1'b0 ;
  assign n54140 = ( n4538 & n20426 ) | ( n4538 & ~n24036 ) | ( n20426 & ~n24036 ) ;
  assign n54141 = n47456 | n54140 ;
  assign n54143 = n20314 ^ n6877 ^ n5012 ;
  assign n54142 = n49479 ^ n47231 ^ n4803 ;
  assign n54144 = n54143 ^ n54142 ^ n7413 ;
  assign n54145 = n12425 ^ n2825 ^ 1'b0 ;
  assign n54146 = n9101 & ~n54145 ;
  assign n54147 = ( ~n10240 & n38307 ) | ( ~n10240 & n54146 ) | ( n38307 & n54146 ) ;
  assign n54148 = n9935 & ~n43188 ;
  assign n54149 = ~n13253 & n54148 ;
  assign n54151 = n6134 | n12143 ;
  assign n54150 = ~n13256 & n38497 ;
  assign n54152 = n54151 ^ n54150 ^ 1'b0 ;
  assign n54153 = n9175 & n54152 ;
  assign n54154 = n54153 ^ n22530 ^ 1'b0 ;
  assign n54155 = n49167 ^ n38660 ^ n15083 ;
  assign n54157 = n19335 | n24864 ;
  assign n54158 = n54157 ^ n32465 ^ 1'b0 ;
  assign n54156 = n40433 ^ n41 ^ 1'b0 ;
  assign n54159 = n54158 ^ n54156 ^ n11154 ;
  assign n54160 = ( n33289 & ~n46327 ) | ( n33289 & n47939 ) | ( ~n46327 & n47939 ) ;
  assign n54161 = n9357 & n47002 ;
  assign n54162 = n17226 & n25477 ;
  assign n54163 = n31884 ^ n11987 ^ 1'b0 ;
  assign n54164 = n7151 | n54163 ;
  assign n54165 = ~n2933 & n10424 ;
  assign n54166 = n54165 ^ n20248 ^ 1'b0 ;
  assign n54167 = n1026 & ~n31908 ;
  assign n54168 = n54167 ^ n17285 ^ 1'b0 ;
  assign n54169 = n40451 ^ n19164 ^ 1'b0 ;
  assign n54170 = ~n12371 & n54169 ;
  assign n54171 = n7428 & n10734 ;
  assign n54172 = n54171 ^ n23333 ^ 1'b0 ;
  assign n54173 = n50942 ^ n15330 ^ 1'b0 ;
  assign n54174 = ( n622 & ~n54172 ) | ( n622 & n54173 ) | ( ~n54172 & n54173 ) ;
  assign n54175 = n2100 | n5968 ;
  assign n54176 = n54175 ^ n51196 ^ 1'b0 ;
  assign n54177 = n9902 & ~n54176 ;
  assign n54178 = n40578 & n45306 ;
  assign n54179 = n9288 & ~n16726 ;
  assign n54180 = n54178 & n54179 ;
  assign n54181 = ( n1886 & n15226 ) | ( n1886 & ~n41178 ) | ( n15226 & ~n41178 ) ;
  assign n54182 = n54181 ^ n17520 ^ 1'b0 ;
  assign n54183 = n17567 & ~n54182 ;
  assign n54184 = n16917 | n29968 ;
  assign n54185 = n22664 & ~n54184 ;
  assign n54186 = n39674 | n54185 ;
  assign n54187 = n17687 ^ n15260 ^ 1'b0 ;
  assign n54188 = n34219 ^ n18424 ^ 1'b0 ;
  assign n54189 = n54187 & n54188 ;
  assign n54190 = n5068 ^ n3936 ^ 1'b0 ;
  assign n54191 = n54189 & n54190 ;
  assign n54192 = n40875 ^ n11706 ^ 1'b0 ;
  assign n54193 = ~n15328 & n46244 ;
  assign n54194 = n54192 & n54193 ;
  assign n54195 = n22104 ^ n19418 ^ 1'b0 ;
  assign n54196 = n51572 & n52097 ;
  assign n54197 = n16450 ^ n4515 ^ 1'b0 ;
  assign n54198 = n4475 & ~n14141 ;
  assign n54199 = n54198 ^ n48167 ^ n19007 ;
  assign n54200 = n10149 & ~n46571 ;
  assign n54201 = n8950 & n54200 ;
  assign n54202 = n17008 | n18264 ;
  assign n54203 = n24519 & ~n54202 ;
  assign n54204 = n3060 & ~n8991 ;
  assign n54205 = n11247 & n54204 ;
  assign n54206 = n6045 | n15982 ;
  assign n54207 = n4845 ^ n1650 ^ 1'b0 ;
  assign n54208 = n18675 | n54207 ;
  assign n54209 = n10791 & n25724 ;
  assign n54210 = n54209 ^ n40436 ^ 1'b0 ;
  assign n54211 = n54208 & ~n54210 ;
  assign n54212 = ~n1209 & n41772 ;
  assign n54213 = n9313 | n23996 ;
  assign n54214 = n54213 ^ n46423 ^ n16532 ;
  assign n54215 = n35773 ^ n23174 ^ 1'b0 ;
  assign n54216 = n37847 & n54215 ;
  assign n54217 = n13708 | n46022 ;
  assign n54218 = n54217 ^ n36128 ^ 1'b0 ;
  assign n54219 = ( ~n5870 & n6664 ) | ( ~n5870 & n19304 ) | ( n6664 & n19304 ) ;
  assign n54220 = n14939 & ~n54219 ;
  assign n54221 = n54220 ^ n19803 ^ 1'b0 ;
  assign n54222 = n42461 & n54221 ;
  assign n54223 = n26782 ^ n9095 ^ 1'b0 ;
  assign n54224 = n4105 & ~n54223 ;
  assign n54225 = n28529 ^ n12589 ^ 1'b0 ;
  assign n54226 = n47320 ^ n21887 ^ 1'b0 ;
  assign n54227 = n5436 | n47469 ;
  assign n54228 = ( n18799 & n46107 ) | ( n18799 & ~n54227 ) | ( n46107 & ~n54227 ) ;
  assign n54230 = ~n15507 & n40729 ;
  assign n54231 = ~n3075 & n54230 ;
  assign n54229 = n30516 ^ n17197 ^ 1'b0 ;
  assign n54232 = n54231 ^ n54229 ^ n23842 ;
  assign n54233 = n12107 | n14154 ;
  assign n54234 = n21913 & ~n54233 ;
  assign n54235 = n12208 | n12438 ;
  assign n54236 = n54235 ^ n13550 ^ 1'b0 ;
  assign n54237 = n14252 | n26278 ;
  assign n54238 = n2070 | n54237 ;
  assign n54239 = n6504 & n53670 ;
  assign n54240 = n54239 ^ n12408 ^ 1'b0 ;
  assign n54241 = n38191 ^ n1499 ^ n823 ;
  assign n54242 = ~n4994 & n54241 ;
  assign n54243 = n34839 ^ n27875 ^ 1'b0 ;
  assign n54246 = n17200 & ~n42327 ;
  assign n54247 = n54246 ^ n23302 ^ 1'b0 ;
  assign n54244 = ~n10506 & n10844 ;
  assign n54245 = ( n8853 & n23258 ) | ( n8853 & ~n54244 ) | ( n23258 & ~n54244 ) ;
  assign n54248 = n54247 ^ n54245 ^ 1'b0 ;
  assign n54249 = n17138 & ~n32961 ;
  assign n54250 = n7046 & n54249 ;
  assign n54251 = n34320 ^ n4694 ^ 1'b0 ;
  assign n54252 = ~n54250 & n54251 ;
  assign n54253 = ~n498 & n34421 ;
  assign n54254 = n54253 ^ n1444 ^ 1'b0 ;
  assign n54255 = n10807 | n11219 ;
  assign n54256 = n54255 ^ n3923 ^ 1'b0 ;
  assign n54257 = n7427 & n15975 ;
  assign n54258 = ( n2040 & n3452 ) | ( n2040 & n4807 ) | ( n3452 & n4807 ) ;
  assign n54259 = n7124 & ~n8122 ;
  assign n54260 = ~n54258 & n54259 ;
  assign n54261 = n4408 | n54260 ;
  assign n54262 = n38141 ^ n25802 ^ 1'b0 ;
  assign n54263 = ( ~n10263 & n15610 ) | ( ~n10263 & n21398 ) | ( n15610 & n21398 ) ;
  assign n54264 = n46484 ^ n42700 ^ 1'b0 ;
  assign n54265 = n6238 & n8404 ;
  assign n54266 = n54265 ^ n48915 ^ n29809 ;
  assign n54267 = n20056 ^ n10279 ^ n3295 ;
  assign n54268 = ~n35242 & n54267 ;
  assign n54269 = n30516 | n33514 ;
  assign n54270 = n21587 ^ n10307 ^ n2769 ;
  assign n54271 = n8925 & n54270 ;
  assign n54272 = n70 & ~n2640 ;
  assign n54273 = ~n19146 & n54272 ;
  assign n54274 = n54273 ^ n15452 ^ 1'b0 ;
  assign n54275 = n28325 & ~n53811 ;
  assign n54276 = n11423 ^ n2323 ^ 1'b0 ;
  assign n54277 = n7575 & ~n11676 ;
  assign n54278 = n12830 & n54277 ;
  assign n54279 = n54278 ^ n37323 ^ 1'b0 ;
  assign n54280 = n54276 & n54279 ;
  assign n54281 = n577 & ~n51614 ;
  assign n54282 = n7808 & n54281 ;
  assign n54283 = ~n7268 & n23901 ;
  assign n54284 = n54283 ^ n8232 ^ 1'b0 ;
  assign n54285 = n35369 ^ n637 ^ 1'b0 ;
  assign n54286 = ~n285 & n15402 ;
  assign n54287 = ~n1903 & n31854 ;
  assign n54288 = n24114 & n54287 ;
  assign n54289 = n16736 | n54288 ;
  assign n54290 = n6322 | n25898 ;
  assign n54291 = n13829 ^ n11676 ^ 1'b0 ;
  assign n54292 = n15923 | n54291 ;
  assign n54293 = n54292 ^ n19487 ^ 1'b0 ;
  assign n54294 = n8374 | n54293 ;
  assign n54295 = ~n54290 & n54294 ;
  assign n54296 = n9127 ^ n1859 ^ 1'b0 ;
  assign n54297 = ( ~n4825 & n22745 ) | ( ~n4825 & n54296 ) | ( n22745 & n54296 ) ;
  assign n54298 = n54297 ^ n36656 ^ 1'b0 ;
  assign n54299 = n33642 ^ n7434 ^ 1'b0 ;
  assign n54300 = n36523 & ~n45927 ;
  assign n54301 = ~n24220 & n39359 ;
  assign n54302 = n29578 ^ n4271 ^ 1'b0 ;
  assign n54303 = n54301 & ~n54302 ;
  assign n54304 = n54303 ^ n33566 ^ 1'b0 ;
  assign n54305 = ~n40551 & n45746 ;
  assign n54306 = n28084 ^ n5444 ^ 1'b0 ;
  assign n54307 = ( n3614 & ~n5137 ) | ( n3614 & n25184 ) | ( ~n5137 & n25184 ) ;
  assign n54308 = n43678 ^ n26162 ^ n13534 ;
  assign n54309 = ( ~n10517 & n30474 ) | ( ~n10517 & n54308 ) | ( n30474 & n54308 ) ;
  assign n54310 = n8783 ^ n7340 ^ 1'b0 ;
  assign n54311 = n14023 & n54310 ;
  assign n54312 = n15306 & ~n54311 ;
  assign n54313 = n16383 & n35048 ;
  assign n54314 = n54313 ^ n5606 ^ 1'b0 ;
  assign n54315 = n621 | n43624 ;
  assign n54316 = n17513 ^ n15999 ^ 1'b0 ;
  assign n54317 = n7219 | n54316 ;
  assign n54318 = n11532 ^ n1091 ^ 1'b0 ;
  assign n54319 = ~n54317 & n54318 ;
  assign n54320 = ( n6081 & n28600 ) | ( n6081 & n33312 ) | ( n28600 & n33312 ) ;
  assign n54321 = n908 | n54320 ;
  assign n54322 = n17049 & ~n33703 ;
  assign n54324 = n38199 ^ n15324 ^ 1'b0 ;
  assign n54325 = n30453 | n54324 ;
  assign n54326 = n54325 ^ n21736 ^ n2344 ;
  assign n54323 = n7267 & n23205 ;
  assign n54327 = n54326 ^ n54323 ^ 1'b0 ;
  assign n54328 = ( n23443 & ~n54322 ) | ( n23443 & n54327 ) | ( ~n54322 & n54327 ) ;
  assign n54329 = n46395 ^ n11998 ^ 1'b0 ;
  assign n54330 = n23239 ^ n14273 ^ n6191 ;
  assign n54331 = ~n13181 & n16415 ;
  assign n54332 = n54331 ^ n52481 ^ 1'b0 ;
  assign n54334 = n8463 ^ n2986 ^ 1'b0 ;
  assign n54333 = n788 & ~n12504 ;
  assign n54335 = n54334 ^ n54333 ^ 1'b0 ;
  assign n54336 = n42444 ^ n31984 ^ n23903 ;
  assign n54337 = n42120 ^ n39962 ^ 1'b0 ;
  assign n54338 = n20153 ^ n18773 ^ 1'b0 ;
  assign n54339 = n11949 & n54338 ;
  assign n54340 = n54339 ^ n49091 ^ n30071 ;
  assign n54341 = n24189 ^ n9934 ^ 1'b0 ;
  assign n54342 = n2117 | n54341 ;
  assign n54343 = n19153 & n27391 ;
  assign n54344 = n11321 & n23089 ;
  assign n54345 = ~n960 & n54344 ;
  assign n54346 = n22916 | n54345 ;
  assign n54347 = n9029 ^ n1400 ^ 1'b0 ;
  assign n54348 = n6948 | n54347 ;
  assign n54349 = n54346 | n54348 ;
  assign n54350 = n48887 & ~n54349 ;
  assign n54351 = ~n18164 & n54350 ;
  assign n54352 = ~n9633 & n20301 ;
  assign n54353 = n32864 & n54352 ;
  assign n54354 = n53206 ^ n49885 ^ 1'b0 ;
  assign n54355 = n50218 & n50361 ;
  assign n54356 = ~n1885 & n4894 ;
  assign n54357 = ~n10428 & n54356 ;
  assign n54358 = n54357 ^ n45139 ^ 1'b0 ;
  assign n54359 = n9671 & n54358 ;
  assign n54360 = n2222 | n9087 ;
  assign n54361 = n25238 ^ n21040 ^ n3016 ;
  assign n54362 = n47929 ^ n38352 ^ n10374 ;
  assign n54363 = ~n762 & n3883 ;
  assign n54364 = n14866 ^ n9284 ^ 1'b0 ;
  assign n54365 = n19193 & n20750 ;
  assign n54366 = n54364 & n54365 ;
  assign n54367 = ~n5802 & n6348 ;
  assign n54368 = ~n27508 & n33571 ;
  assign n54369 = n1400 & n20099 ;
  assign n54370 = n13969 & n39539 ;
  assign n54371 = ( ~n54368 & n54369 ) | ( ~n54368 & n54370 ) | ( n54369 & n54370 ) ;
  assign n54372 = n26926 ^ n10743 ^ n1319 ;
  assign n54373 = n2048 & ~n33972 ;
  assign n54374 = n54373 ^ n45094 ^ 1'b0 ;
  assign n54375 = n33925 ^ n27100 ^ 1'b0 ;
  assign n54376 = n22247 | n54375 ;
  assign n54377 = n38524 & n43287 ;
  assign n54378 = n8351 & ~n54377 ;
  assign n54379 = n22992 | n54378 ;
  assign n54380 = ( n1376 & n9110 ) | ( n1376 & n21499 ) | ( n9110 & n21499 ) ;
  assign n54381 = n52369 ^ n2602 ^ 1'b0 ;
  assign n54382 = n54380 & n54381 ;
  assign n54383 = n28090 ^ n25194 ^ 1'b0 ;
  assign n54384 = n15600 & ~n54383 ;
  assign n54385 = n51112 ^ n16475 ^ 1'b0 ;
  assign n54386 = n8057 | n29115 ;
  assign n54387 = n31439 | n35093 ;
  assign n54388 = ~n3768 & n35364 ;
  assign n54389 = ~n10254 & n54388 ;
  assign n54390 = n2614 | n12770 ;
  assign n54391 = n8229 | n54390 ;
  assign n54392 = n2135 & n20353 ;
  assign n54393 = n53557 & n54392 ;
  assign n54394 = ( n12089 & n16115 ) | ( n12089 & n27810 ) | ( n16115 & n27810 ) ;
  assign n54395 = n8199 & ~n48291 ;
  assign n54396 = n10154 ^ n8906 ^ 1'b0 ;
  assign n54397 = ~n35129 & n54396 ;
  assign n54398 = n7544 ^ n5569 ^ 1'b0 ;
  assign n54399 = n30470 | n54398 ;
  assign n54400 = n31087 | n54399 ;
  assign n54401 = n44877 ^ n22642 ^ 1'b0 ;
  assign n54402 = n54400 & ~n54401 ;
  assign n54404 = n18038 ^ n15987 ^ 1'b0 ;
  assign n54405 = n469 & n54404 ;
  assign n54403 = ~n16920 & n29910 ;
  assign n54406 = n54405 ^ n54403 ^ 1'b0 ;
  assign n54407 = n32861 & n52603 ;
  assign n54408 = ( n8170 & n13889 ) | ( n8170 & ~n39350 ) | ( n13889 & ~n39350 ) ;
  assign n54409 = n29816 & n54408 ;
  assign n54410 = n54409 ^ n29403 ^ 1'b0 ;
  assign n54411 = n13517 & n31306 ;
  assign n54412 = n11692 & n33732 ;
  assign n54413 = n46911 ^ n27092 ^ 1'b0 ;
  assign n54414 = ~n21809 & n54083 ;
  assign n54415 = n23124 | n33638 ;
  assign n54416 = n46469 ^ n4233 ^ 1'b0 ;
  assign n54417 = n1039 | n20831 ;
  assign n54418 = n38320 | n54417 ;
  assign n54419 = ~n2225 & n45594 ;
  assign n54420 = n9020 & n54419 ;
  assign n54421 = n22375 | n49429 ;
  assign n54426 = ~n21448 & n31483 ;
  assign n54422 = ~n18466 & n23283 ;
  assign n54423 = n9863 | n28359 ;
  assign n54424 = n54423 ^ n63 ^ 1'b0 ;
  assign n54425 = n54422 | n54424 ;
  assign n54427 = n54426 ^ n54425 ^ 1'b0 ;
  assign n54428 = n16 | n11701 ;
  assign n54429 = n865 & n2177 ;
  assign n54430 = n54429 ^ n29845 ^ 1'b0 ;
  assign n54431 = n13598 ^ n1932 ^ 1'b0 ;
  assign n54432 = ~n23351 & n54431 ;
  assign n54433 = n16200 ^ n6164 ^ 1'b0 ;
  assign n54434 = ( n299 & n8738 ) | ( n299 & ~n12935 ) | ( n8738 & ~n12935 ) ;
  assign n54435 = n54434 ^ n15671 ^ 1'b0 ;
  assign n54436 = n558 | n22673 ;
  assign n54437 = n9995 | n30586 ;
  assign n54438 = n46457 ^ n29634 ^ 1'b0 ;
  assign n54439 = n5941 | n11256 ;
  assign n54440 = n46588 & ~n54439 ;
  assign n54441 = n54440 ^ n30943 ^ 1'b0 ;
  assign n54443 = n15021 | n17542 ;
  assign n54444 = n32634 ^ n5312 ^ 1'b0 ;
  assign n54445 = n54443 | n54444 ;
  assign n54442 = n37358 & ~n40272 ;
  assign n54446 = n54445 ^ n54442 ^ 1'b0 ;
  assign n54447 = n54446 ^ n34871 ^ 1'b0 ;
  assign n54448 = n31726 ^ n7588 ^ 1'b0 ;
  assign n54449 = n30267 | n54448 ;
  assign n54450 = n29842 | n40642 ;
  assign n54451 = n54450 ^ n39138 ^ 1'b0 ;
  assign n54452 = n30196 ^ n26271 ^ n6548 ;
  assign n54453 = n16603 ^ n15323 ^ 1'b0 ;
  assign n54454 = n5582 & ~n8301 ;
  assign n54455 = n54454 ^ n2818 ^ 1'b0 ;
  assign n54456 = n54455 ^ n415 ^ 1'b0 ;
  assign n54457 = n54453 & ~n54456 ;
  assign n54458 = n54457 ^ n52943 ^ 1'b0 ;
  assign n54459 = n3742 ^ n1018 ^ 1'b0 ;
  assign n54460 = ~n16836 & n39001 ;
  assign n54461 = n54460 ^ n27156 ^ 1'b0 ;
  assign n54462 = n29889 & n54461 ;
  assign n54463 = ~n14827 & n38393 ;
  assign n54464 = ~n54462 & n54463 ;
  assign n54465 = n25368 & ~n54464 ;
  assign n54466 = n54465 ^ n10707 ^ 1'b0 ;
  assign n54467 = n35572 ^ n25714 ^ 1'b0 ;
  assign n54468 = ~n838 & n7033 ;
  assign n54469 = ( n5974 & n9094 ) | ( n5974 & n9116 ) | ( n9094 & n9116 ) ;
  assign n54470 = ~n22515 & n54469 ;
  assign n54471 = n52888 ^ n888 ^ 1'b0 ;
  assign n54472 = n41792 & ~n48684 ;
  assign n54473 = n38738 ^ n10222 ^ 1'b0 ;
  assign n54474 = n19407 & n26937 ;
  assign n54475 = ~n54473 & n54474 ;
  assign n54476 = n32408 | n36043 ;
  assign n54477 = n12707 | n15886 ;
  assign n54478 = n31426 ^ n6460 ^ 1'b0 ;
  assign n54479 = n54478 ^ n38279 ^ n35571 ;
  assign n54480 = n8019 & n43978 ;
  assign n54481 = n54480 ^ n8853 ^ 1'b0 ;
  assign n54482 = n7767 & ~n54481 ;
  assign n54483 = n12155 & n54482 ;
  assign n54484 = n17062 ^ n16979 ^ 1'b0 ;
  assign n54486 = n2977 & n4785 ;
  assign n54485 = n8878 | n40301 ;
  assign n54487 = n54486 ^ n54485 ^ 1'b0 ;
  assign n54488 = n16783 ^ n1952 ^ 1'b0 ;
  assign n54489 = n24660 & ~n54488 ;
  assign n54490 = n20679 ^ n9809 ^ 1'b0 ;
  assign n54491 = n37471 | n54490 ;
  assign n54492 = n23814 & n34542 ;
  assign n54493 = n17614 ^ n13180 ^ 1'b0 ;
  assign n54494 = n54493 ^ n42431 ^ n4560 ;
  assign n54495 = n39303 ^ n10507 ^ 1'b0 ;
  assign n54496 = n12708 & n38171 ;
  assign n54497 = n54496 ^ n30304 ^ 1'b0 ;
  assign n54498 = n1882 & n10676 ;
  assign n54499 = n42243 & n54498 ;
  assign n54500 = n8298 & ~n40345 ;
  assign n54501 = n2350 | n41714 ;
  assign n54502 = ( n31206 & ~n37866 ) | ( n31206 & n41703 ) | ( ~n37866 & n41703 ) ;
  assign n54503 = n54502 ^ n39045 ^ n27553 ;
  assign n54504 = n19529 ^ n14459 ^ 1'b0 ;
  assign n54505 = n25312 & ~n54504 ;
  assign n54506 = n10635 ^ n8526 ^ 1'b0 ;
  assign n54507 = ~n918 & n54506 ;
  assign n54508 = n52800 ^ n3926 ^ 1'b0 ;
  assign n54509 = n12095 | n16268 ;
  assign n54510 = n29817 ^ n5072 ^ 1'b0 ;
  assign n54515 = n12005 | n17820 ;
  assign n54516 = n54515 ^ n16415 ^ 1'b0 ;
  assign n54517 = n41068 ^ n33677 ^ 1'b0 ;
  assign n54518 = ~n24100 & n54517 ;
  assign n54519 = ~n54516 & n54518 ;
  assign n54520 = ~n1764 & n1891 ;
  assign n54521 = ( n11859 & n54519 ) | ( n11859 & ~n54520 ) | ( n54519 & ~n54520 ) ;
  assign n54522 = n54521 ^ n50848 ^ 1'b0 ;
  assign n54512 = n13400 ^ n1586 ^ 1'b0 ;
  assign n54513 = n6581 & ~n54512 ;
  assign n54511 = n42399 | n54185 ;
  assign n54514 = n54513 ^ n54511 ^ 1'b0 ;
  assign n54523 = n54522 ^ n54514 ^ 1'b0 ;
  assign n54524 = ( ~n27104 & n29561 ) | ( ~n27104 & n37285 ) | ( n29561 & n37285 ) ;
  assign n54525 = n33337 ^ n31694 ^ 1'b0 ;
  assign n54526 = n37 & ~n3784 ;
  assign n54527 = ~n54525 & n54526 ;
  assign n54528 = n54527 ^ n9026 ^ 1'b0 ;
  assign n54529 = n3998 | n22387 ;
  assign n54530 = n54529 ^ n40171 ^ 1'b0 ;
  assign n54531 = n10911 | n10993 ;
  assign n54532 = n18796 ^ n11272 ^ 1'b0 ;
  assign n54533 = n577 & ~n54532 ;
  assign n54534 = ( n16873 & n20967 ) | ( n16873 & ~n23666 ) | ( n20967 & ~n23666 ) ;
  assign n54535 = n2044 & ~n54534 ;
  assign n54536 = n16546 ^ n10467 ^ 1'b0 ;
  assign n54537 = ~n20355 & n29242 ;
  assign n54538 = n4944 & ~n54537 ;
  assign n54539 = ~n28877 & n54538 ;
  assign n54540 = n31335 | n54539 ;
  assign n54541 = n2412 & ~n18247 ;
  assign n54542 = n50225 ^ n12111 ^ 1'b0 ;
  assign n54543 = n14791 & n44605 ;
  assign n54545 = ( ~n18511 & n31953 ) | ( ~n18511 & n34982 ) | ( n31953 & n34982 ) ;
  assign n54544 = ~n16402 & n52189 ;
  assign n54546 = n54545 ^ n54544 ^ 1'b0 ;
  assign n54547 = n47963 ^ n34527 ^ n15382 ;
  assign n54548 = n2674 ^ n1248 ^ 1'b0 ;
  assign n54549 = n43856 | n54548 ;
  assign n54550 = n54549 ^ n30993 ^ 1'b0 ;
  assign n54551 = n17239 & n34343 ;
  assign n54552 = n29368 | n37150 ;
  assign n54553 = n13522 & ~n26217 ;
  assign n54554 = n27556 | n37727 ;
  assign n54555 = n17712 | n24447 ;
  assign n54556 = n54555 ^ n20353 ^ 1'b0 ;
  assign n54557 = ( n10118 & n33423 ) | ( n10118 & n54556 ) | ( n33423 & n54556 ) ;
  assign n54558 = ( n4316 & n13497 ) | ( n4316 & n14867 ) | ( n13497 & n14867 ) ;
  assign n54559 = ( n168 & n362 ) | ( n168 & n54558 ) | ( n362 & n54558 ) ;
  assign n54560 = ~n13453 & n15383 ;
  assign n54561 = n54560 ^ n15024 ^ 1'b0 ;
  assign n54562 = n478 & n830 ;
  assign n54563 = ~n1328 & n43233 ;
  assign n54564 = n44125 ^ n13795 ^ 1'b0 ;
  assign n54565 = n54563 | n54564 ;
  assign n54566 = n10313 ^ n4694 ^ 1'b0 ;
  assign n54567 = n35410 | n54566 ;
  assign n54568 = n30873 | n54567 ;
  assign n54569 = n54565 & ~n54568 ;
  assign n54570 = n25672 ^ n7423 ^ 1'b0 ;
  assign n54571 = ~n19679 & n37156 ;
  assign n54572 = n54571 ^ n34647 ^ 1'b0 ;
  assign n54573 = n19463 & ~n20269 ;
  assign n54574 = n29752 ^ n16540 ^ 1'b0 ;
  assign n54575 = n53865 ^ n12849 ^ n10333 ;
  assign n54576 = n36622 ^ n33304 ^ n14603 ;
  assign n54577 = n2666 & ~n3791 ;
  assign n54578 = n54577 ^ n20277 ^ 1'b0 ;
  assign n54579 = ~n4006 & n54578 ;
  assign n54580 = n30394 | n47070 ;
  assign n54581 = n54580 ^ n738 ^ 1'b0 ;
  assign n54582 = n54581 ^ n15505 ^ 1'b0 ;
  assign n54583 = ~n1882 & n54582 ;
  assign n54584 = n36304 ^ n21090 ^ 1'b0 ;
  assign n54585 = n8967 & ~n22835 ;
  assign n54586 = n35215 & n39951 ;
  assign n54587 = n54586 ^ n10948 ^ 1'b0 ;
  assign n54588 = ~n54585 & n54587 ;
  assign n54590 = n41983 ^ n21605 ^ 1'b0 ;
  assign n54591 = n3193 & ~n54590 ;
  assign n54589 = ~n16735 & n23526 ;
  assign n54592 = n54591 ^ n54589 ^ 1'b0 ;
  assign n54593 = n47121 ^ n44375 ^ n8542 ;
  assign n54594 = ( n10007 & n19716 ) | ( n10007 & n54593 ) | ( n19716 & n54593 ) ;
  assign n54598 = n1311 ^ x3 ^ 1'b0 ;
  assign n54595 = n8139 & ~n20843 ;
  assign n54596 = n4028 & n54595 ;
  assign n54597 = n29335 & n54596 ;
  assign n54599 = n54598 ^ n54597 ^ 1'b0 ;
  assign n54600 = ~n779 & n24891 ;
  assign n54601 = n54600 ^ n911 ^ 1'b0 ;
  assign n54603 = n15290 & n16594 ;
  assign n54602 = n22686 & n32986 ;
  assign n54604 = n54603 ^ n54602 ^ 1'b0 ;
  assign n54605 = n4794 & n11430 ;
  assign n54606 = n7896 & n46852 ;
  assign n54607 = ~n38789 & n54606 ;
  assign n54608 = n40183 & n54607 ;
  assign n54611 = n34484 ^ n13077 ^ 1'b0 ;
  assign n54612 = ~n9813 & n54611 ;
  assign n54609 = n30898 & ~n53209 ;
  assign n54610 = n54609 ^ n48438 ^ 1'b0 ;
  assign n54613 = n54612 ^ n54610 ^ n50251 ;
  assign n54614 = n28125 & n31078 ;
  assign n54615 = n54614 ^ n27984 ^ 1'b0 ;
  assign n54616 = n13211 & ~n49512 ;
  assign n54617 = n5722 & n54616 ;
  assign n54618 = n18786 ^ n2721 ^ 1'b0 ;
  assign n54619 = n15258 ^ n11949 ^ 1'b0 ;
  assign n54620 = ~n49618 & n54619 ;
  assign n54621 = n33119 ^ n4830 ^ 1'b0 ;
  assign n54622 = n54620 & n54621 ;
  assign n54623 = n26389 & ~n49430 ;
  assign n54624 = n4545 ^ n4141 ^ 1'b0 ;
  assign n54625 = n3692 & ~n54624 ;
  assign n54626 = n54625 ^ n22361 ^ 1'b0 ;
  assign n54627 = ( n5732 & n12720 ) | ( n5732 & ~n14175 ) | ( n12720 & ~n14175 ) ;
  assign n54628 = n18196 | n54627 ;
  assign n54629 = n11147 | n54628 ;
  assign n54630 = n44435 & n54629 ;
  assign n54631 = ~n2830 & n54630 ;
  assign n54632 = n15660 & ~n54631 ;
  assign n54633 = n9303 & n54632 ;
  assign n54634 = n28843 ^ n4580 ^ 1'b0 ;
  assign n54635 = n3642 & n54634 ;
  assign n54636 = n10140 | n22912 ;
  assign n54637 = n54635 | n54636 ;
  assign n54638 = n25338 ^ n22682 ^ 1'b0 ;
  assign n54639 = ~n12522 & n54638 ;
  assign n54640 = n53576 ^ n48822 ^ 1'b0 ;
  assign n54641 = n13326 & ~n54640 ;
  assign n54642 = n21433 ^ n3469 ^ 1'b0 ;
  assign n54643 = n24676 | n47155 ;
  assign n54644 = n54643 ^ n23225 ^ 1'b0 ;
  assign n54645 = n35491 ^ n401 ^ 1'b0 ;
  assign n54647 = n48070 ^ n16103 ^ n6620 ;
  assign n54646 = n35410 & ~n39745 ;
  assign n54648 = n54647 ^ n54646 ^ 1'b0 ;
  assign n54649 = n18843 ^ n2597 ^ 1'b0 ;
  assign n54650 = n13234 & ~n54649 ;
  assign n54651 = n11706 & ~n19429 ;
  assign n54652 = n30716 & n54651 ;
  assign n54653 = n16049 ^ n5987 ^ 1'b0 ;
  assign n54654 = n7795 & ~n54653 ;
  assign n54655 = n54654 ^ n35958 ^ 1'b0 ;
  assign n54656 = n5183 & ~n19014 ;
  assign n54657 = ( ~n6153 & n6862 ) | ( ~n6153 & n9634 ) | ( n6862 & n9634 ) ;
  assign n54658 = n15566 ^ n2551 ^ 1'b0 ;
  assign n54659 = n10049 | n54658 ;
  assign n54660 = ~n5844 & n54659 ;
  assign n54661 = n47476 & ~n54660 ;
  assign n54662 = n54661 ^ n29849 ^ 1'b0 ;
  assign n54663 = ~n9103 & n44317 ;
  assign n54664 = ( n3248 & n38875 ) | ( n3248 & ~n45967 ) | ( n38875 & ~n45967 ) ;
  assign n54665 = n30873 ^ n9224 ^ 1'b0 ;
  assign n54666 = ~n54664 & n54665 ;
  assign n54667 = n32004 & ~n44582 ;
  assign n54668 = n53201 ^ n10634 ^ 1'b0 ;
  assign n54669 = n15254 ^ x3 ^ 1'b0 ;
  assign n54670 = n18629 & ~n54669 ;
  assign n54671 = n22702 & ~n54670 ;
  assign n54672 = n1401 & n52839 ;
  assign n54673 = n31306 | n44660 ;
  assign n54674 = n44600 & ~n54673 ;
  assign n54675 = ~n17507 & n36508 ;
  assign n54676 = n54675 ^ n46419 ^ 1'b0 ;
  assign n54677 = n7993 & n29040 ;
  assign n54678 = n54677 ^ n9577 ^ 1'b0 ;
  assign n54679 = n19839 ^ n13428 ^ 1'b0 ;
  assign n54680 = n54678 & ~n54679 ;
  assign n54681 = ~n4923 & n54680 ;
  assign n54682 = n54681 ^ n31259 ^ 1'b0 ;
  assign n54683 = n50788 ^ n9109 ^ 1'b0 ;
  assign n54684 = n18904 ^ n10820 ^ n1124 ;
  assign n54685 = ( ~n11177 & n30132 ) | ( ~n11177 & n54684 ) | ( n30132 & n54684 ) ;
  assign n54686 = n5864 | n12456 ;
  assign n54687 = n54686 ^ n47244 ^ n5585 ;
  assign n54688 = n38835 & n54687 ;
  assign n54689 = n6639 ^ n6545 ^ 1'b0 ;
  assign n54690 = n28285 & ~n54689 ;
  assign n54691 = n22453 & ~n45218 ;
  assign n54692 = ~n28649 & n48890 ;
  assign n54693 = ~n36072 & n48881 ;
  assign n54694 = ~n54692 & n54693 ;
  assign n54695 = n51764 ^ n21185 ^ n151 ;
  assign n54696 = ( ~n2432 & n7915 ) | ( ~n2432 & n21787 ) | ( n7915 & n21787 ) ;
  assign n54697 = ( n12854 & n43619 ) | ( n12854 & n51032 ) | ( n43619 & n51032 ) ;
  assign n54698 = n41494 ^ n8856 ^ 1'b0 ;
  assign n54699 = n5427 | n54698 ;
  assign n54700 = n41186 ^ n32834 ^ 1'b0 ;
  assign n54701 = n6733 & ~n23558 ;
  assign n54702 = n7377 | n23590 ;
  assign n54703 = n54701 | n54702 ;
  assign n54704 = n14069 ^ n11535 ^ 1'b0 ;
  assign n54705 = n23433 | n54704 ;
  assign n54706 = ~n7908 & n23004 ;
  assign n54707 = n9509 & n54706 ;
  assign n54708 = n3879 | n4367 ;
  assign n54709 = n54707 & ~n54708 ;
  assign n54710 = n4906 & ~n54709 ;
  assign n54711 = n54710 ^ n13034 ^ 1'b0 ;
  assign n54712 = n54711 ^ n1167 ^ 1'b0 ;
  assign n54713 = n691 & n22307 ;
  assign n54714 = n18723 ^ n16828 ^ 1'b0 ;
  assign n54715 = ~n40862 & n54714 ;
  assign n54716 = n29471 ^ n15192 ^ 1'b0 ;
  assign n54717 = ( n2526 & ~n9905 ) | ( n2526 & n9909 ) | ( ~n9905 & n9909 ) ;
  assign n54718 = ( n24976 & ~n54716 ) | ( n24976 & n54717 ) | ( ~n54716 & n54717 ) ;
  assign n54719 = n28407 | n32470 ;
  assign n54720 = n35419 | n38163 ;
  assign n54721 = n54720 ^ n15328 ^ 1'b0 ;
  assign n54722 = n1085 | n16829 ;
  assign n54723 = ~n54721 & n54722 ;
  assign n54724 = ~n6686 & n17280 ;
  assign n54725 = n4992 & ~n9006 ;
  assign n54726 = n2377 & ~n5008 ;
  assign n54727 = n5008 & n54726 ;
  assign n54728 = n12093 & ~n54727 ;
  assign n54729 = ~n12093 & n54728 ;
  assign n54730 = n1400 | n54729 ;
  assign n54731 = n1699 & n54730 ;
  assign n54732 = ~n54730 & n54731 ;
  assign n54733 = n54732 ^ n31539 ^ n18268 ;
  assign n54734 = n54733 ^ n2278 ^ 1'b0 ;
  assign n54735 = n54725 & ~n54734 ;
  assign n54736 = n17761 ^ n10774 ^ 1'b0 ;
  assign n54737 = n54736 ^ n28984 ^ n28325 ;
  assign n54738 = n54737 ^ n6589 ^ 1'b0 ;
  assign n54739 = n948 | n28184 ;
  assign n54740 = n54739 ^ n29604 ^ n16347 ;
  assign n54741 = ( n14715 & ~n44667 ) | ( n14715 & n54740 ) | ( ~n44667 & n54740 ) ;
  assign n54745 = n18648 ^ n1412 ^ 1'b0 ;
  assign n54746 = n3762 | n54745 ;
  assign n54743 = n21022 ^ n3094 ^ 1'b0 ;
  assign n54744 = n3898 & ~n54743 ;
  assign n54742 = n43423 ^ n33905 ^ n18598 ;
  assign n54747 = n54746 ^ n54744 ^ n54742 ;
  assign n54748 = n6254 & ~n36742 ;
  assign n54749 = n4914 & n54748 ;
  assign n54750 = n15849 ^ n6554 ^ 1'b0 ;
  assign n54751 = ~n131 & n2541 ;
  assign n54752 = n54751 ^ n37208 ^ 1'b0 ;
  assign n54753 = n16120 & n42911 ;
  assign n54754 = ~n16060 & n54753 ;
  assign n54755 = n54754 ^ n14146 ^ n5066 ;
  assign n54756 = n45331 ^ n19317 ^ n4469 ;
  assign n54757 = n7496 & ~n54756 ;
  assign n54758 = n10868 ^ n9191 ^ 1'b0 ;
  assign n54759 = n4539 & ~n36979 ;
  assign n54760 = n35818 ^ n34026 ^ 1'b0 ;
  assign n54761 = ~n32863 & n54760 ;
  assign n54762 = n21394 | n30704 ;
  assign n54763 = n966 & ~n54762 ;
  assign n54764 = ( n3891 & n5427 ) | ( n3891 & ~n16419 ) | ( n5427 & ~n16419 ) ;
  assign n54765 = n54764 ^ n21827 ^ 1'b0 ;
  assign n54766 = n12008 | n43122 ;
  assign n54767 = n45610 | n54766 ;
  assign n54768 = ~n6570 & n8004 ;
  assign n54769 = n20238 ^ n2098 ^ 1'b0 ;
  assign n54770 = n35178 ^ n19144 ^ 1'b0 ;
  assign n54771 = n4541 & ~n54770 ;
  assign n54772 = ( n10382 & ~n30979 ) | ( n10382 & n52335 ) | ( ~n30979 & n52335 ) ;
  assign n54773 = n54771 & n54772 ;
  assign n54774 = n9498 ^ n4394 ^ 1'b0 ;
  assign n54775 = n54774 ^ n21833 ^ n6638 ;
  assign n54777 = n19222 ^ n18793 ^ 1'b0 ;
  assign n54776 = n3876 & ~n37018 ;
  assign n54778 = n54777 ^ n54776 ^ 1'b0 ;
  assign n54779 = n1037 & ~n8542 ;
  assign n54780 = n2157 & n54779 ;
  assign n54781 = ~n38646 & n54780 ;
  assign n54782 = n3455 & ~n54781 ;
  assign n54783 = ~n30078 & n54782 ;
  assign n54784 = n4920 & n8260 ;
  assign n54785 = n37141 ^ n28545 ^ 1'b0 ;
  assign n54786 = n39522 ^ n24169 ^ n1082 ;
  assign n54787 = n35240 & ~n44531 ;
  assign n54788 = n54787 ^ n4105 ^ 1'b0 ;
  assign n54789 = n54788 ^ n53132 ^ 1'b0 ;
  assign n54790 = n14597 & n54789 ;
  assign n54791 = n30816 ^ n11508 ^ 1'b0 ;
  assign n54792 = n5163 | n16822 ;
  assign n54793 = n54792 ^ n2667 ^ 1'b0 ;
  assign n54794 = ( n14980 & n15702 ) | ( n14980 & n54793 ) | ( n15702 & n54793 ) ;
  assign n54795 = ( n7927 & n24131 ) | ( n7927 & ~n54794 ) | ( n24131 & ~n54794 ) ;
  assign n54796 = n7067 | n54795 ;
  assign n54797 = n53257 | n54796 ;
  assign n54798 = n31327 ^ n4269 ^ 1'b0 ;
  assign n54799 = n11773 & ~n54798 ;
  assign n54800 = n54799 ^ n5795 ^ 1'b0 ;
  assign n54801 = ~n15341 & n16776 ;
  assign n54802 = ( n5102 & n25058 ) | ( n5102 & n54801 ) | ( n25058 & n54801 ) ;
  assign n54803 = ~n30699 & n54802 ;
  assign n54804 = n54803 ^ n27477 ^ 1'b0 ;
  assign n54805 = n2840 | n51943 ;
  assign n54806 = n54804 | n54805 ;
  assign n54807 = n54806 ^ n32697 ^ 1'b0 ;
  assign n54808 = n12457 ^ n7280 ^ 1'b0 ;
  assign n54809 = n26300 ^ n7707 ^ n2869 ;
  assign n54810 = n37353 & ~n54809 ;
  assign n54811 = n1603 ^ n87 ^ 1'b0 ;
  assign n54812 = n8008 & n54811 ;
  assign n54813 = n27479 & n36788 ;
  assign n54814 = ~n54812 & n54813 ;
  assign n54815 = n22947 & ~n36664 ;
  assign n54816 = n45667 & n54815 ;
  assign n54817 = n27514 | n41542 ;
  assign n54818 = n54816 & ~n54817 ;
  assign n54819 = n577 & ~n6332 ;
  assign n54820 = n54819 ^ n34371 ^ 1'b0 ;
  assign n54821 = n54007 ^ n22202 ^ 1'b0 ;
  assign n54822 = ( n10261 & n26857 ) | ( n10261 & n45710 ) | ( n26857 & n45710 ) ;
  assign n54823 = n54822 ^ n47596 ^ 1'b0 ;
  assign n54824 = n44804 & n54823 ;
  assign n54825 = ( n157 & n2680 ) | ( n157 & n54824 ) | ( n2680 & n54824 ) ;
  assign n54826 = n54825 ^ n2251 ^ 1'b0 ;
  assign n54827 = n54821 | n54826 ;
  assign n54828 = n20689 & ~n41496 ;
  assign n54829 = n11851 & n28216 ;
  assign n54830 = ~n44000 & n54829 ;
  assign n54831 = n26230 ^ n25244 ^ 1'b0 ;
  assign n54832 = ~n54830 & n54831 ;
  assign n54833 = n2932 & ~n13747 ;
  assign n54834 = n54833 ^ n34905 ^ 1'b0 ;
  assign n54835 = n38163 & n54834 ;
  assign n54836 = n32548 ^ n20734 ^ n11614 ;
  assign n54837 = n54836 ^ n40267 ^ n21469 ;
  assign n54838 = n7352 ^ n4604 ^ 1'b0 ;
  assign n54839 = n54838 ^ n38509 ^ 1'b0 ;
  assign n54840 = n52166 ^ n42270 ^ n906 ;
  assign n54841 = n54840 ^ n3413 ^ 1'b0 ;
  assign n54842 = n12107 | n34569 ;
  assign n54843 = n9160 ^ n7330 ^ 1'b0 ;
  assign n54844 = n20350 & n54843 ;
  assign n54846 = ~n33953 & n36663 ;
  assign n54845 = n29601 & n39985 ;
  assign n54847 = n54846 ^ n54845 ^ 1'b0 ;
  assign n54848 = n25409 ^ n14071 ^ 1'b0 ;
  assign n54850 = n9987 ^ n3560 ^ 1'b0 ;
  assign n54851 = n15 & n54850 ;
  assign n54849 = ~n10969 & n47994 ;
  assign n54852 = n54851 ^ n54849 ^ 1'b0 ;
  assign n54854 = n16103 & n19681 ;
  assign n54853 = ~n670 & n42762 ;
  assign n54855 = n54854 ^ n54853 ^ 1'b0 ;
  assign n54856 = n54855 ^ n23065 ^ n15159 ;
  assign n54857 = n14757 & n22253 ;
  assign n54858 = ( n50900 & n53134 ) | ( n50900 & n54857 ) | ( n53134 & n54857 ) ;
  assign n54859 = n47100 ^ n6935 ^ 1'b0 ;
  assign n54860 = n31932 & n47427 ;
  assign n54861 = n50877 ^ n20548 ^ 1'b0 ;
  assign n54862 = ~n54860 & n54861 ;
  assign n54863 = n9258 ^ n997 ^ n695 ;
  assign n54864 = n54863 ^ n47572 ^ n29799 ;
  assign n54865 = n19805 | n43752 ;
  assign n54866 = n35821 | n54865 ;
  assign n54867 = n54864 & ~n54866 ;
  assign n54868 = n16850 & ~n20876 ;
  assign n54869 = ~n26736 & n54868 ;
  assign n54870 = ~n29406 & n54869 ;
  assign n54871 = n4684 | n38380 ;
  assign n54872 = n54871 ^ n4252 ^ n4134 ;
  assign n54873 = ~n2933 & n25627 ;
  assign n54874 = ( n1022 & ~n28940 ) | ( n1022 & n54873 ) | ( ~n28940 & n54873 ) ;
  assign n54876 = n22611 & ~n37309 ;
  assign n54875 = ( n908 & ~n15080 ) | ( n908 & n16810 ) | ( ~n15080 & n16810 ) ;
  assign n54877 = n54876 ^ n54875 ^ 1'b0 ;
  assign n54879 = n13343 & n22253 ;
  assign n54880 = n54879 ^ n27078 ^ 1'b0 ;
  assign n54881 = n53472 | n54880 ;
  assign n54882 = n54881 ^ n3075 ^ 1'b0 ;
  assign n54878 = ~n22681 & n45126 ;
  assign n54883 = n54882 ^ n54878 ^ 1'b0 ;
  assign n54884 = n40984 ^ n15405 ^ 1'b0 ;
  assign n54885 = n17299 ^ x11 ^ 1'b0 ;
  assign n54886 = ~n2358 & n38816 ;
  assign n54887 = ~n54885 & n54886 ;
  assign n54888 = n7213 & ~n54887 ;
  assign n54889 = ~n23697 & n54888 ;
  assign n54890 = n12892 & ~n54889 ;
  assign n54891 = ~n5982 & n32580 ;
  assign n54892 = n54891 ^ n13374 ^ 1'b0 ;
  assign n54893 = ~n16846 & n54892 ;
  assign n54894 = n21339 & n54893 ;
  assign n54895 = n50933 ^ n7428 ^ 1'b0 ;
  assign n54896 = n8074 & ~n32214 ;
  assign n54897 = n38345 & ~n54896 ;
  assign n54898 = n41679 ^ n35683 ^ 1'b0 ;
  assign n54899 = n23854 | n47059 ;
  assign n54900 = n18454 & ~n54899 ;
  assign n54901 = n34252 & ~n54900 ;
  assign n54902 = n28978 & ~n39480 ;
  assign n54903 = n9143 & ~n12548 ;
  assign n54904 = n36543 ^ n256 ^ 1'b0 ;
  assign n54905 = n8813 & ~n26308 ;
  assign n54906 = n54905 ^ n822 ^ 1'b0 ;
  assign n54907 = n8943 & ~n9283 ;
  assign n54908 = n54907 ^ n4417 ^ 1'b0 ;
  assign n54909 = n8872 & ~n35450 ;
  assign n54910 = n54909 ^ n48733 ^ n839 ;
  assign n54911 = ~n15452 & n21200 ;
  assign n54912 = n35635 ^ n32007 ^ 1'b0 ;
  assign n54913 = n5704 & n54912 ;
  assign n54914 = n6309 & n54913 ;
  assign n54915 = n33285 ^ n21271 ^ 1'b0 ;
  assign n54916 = n24691 & ~n54915 ;
  assign n54917 = n21017 ^ n1037 ^ 1'b0 ;
  assign n54918 = n43596 & n54917 ;
  assign n54919 = n54918 ^ n34191 ^ 1'b0 ;
  assign n54920 = n36019 | n54919 ;
  assign n54921 = n40561 & ~n52245 ;
  assign n54922 = n54921 ^ n53674 ^ 1'b0 ;
  assign n54923 = n46294 & n54922 ;
  assign n54924 = n2135 & n5914 ;
  assign n54925 = ~n13737 & n54924 ;
  assign n54926 = n3286 & ~n54925 ;
  assign n54927 = n4903 & ~n54926 ;
  assign n54928 = n1525 & n54927 ;
  assign n54929 = n11707 & ~n13222 ;
  assign n54930 = n11983 ^ n4552 ^ 1'b0 ;
  assign n54931 = n54930 ^ n53897 ^ n40159 ;
  assign n54932 = n42222 ^ n17751 ^ 1'b0 ;
  assign n54933 = ~n54931 & n54932 ;
  assign n54934 = n32352 & n44540 ;
  assign n54935 = n47125 & n54934 ;
  assign n54936 = n54935 ^ n41383 ^ 1'b0 ;
  assign n54937 = n43027 ^ n30513 ^ 1'b0 ;
  assign n54938 = n34770 ^ n31858 ^ n2427 ;
  assign n54939 = n13094 ^ n10093 ^ n1019 ;
  assign n54940 = n10712 ^ n4097 ^ 1'b0 ;
  assign n54941 = n54939 & ~n54940 ;
  assign n54942 = n41623 ^ n21716 ^ 1'b0 ;
  assign n54943 = ~n21148 & n54942 ;
  assign n54944 = n36776 ^ n5736 ^ 1'b0 ;
  assign n54945 = n54943 & n54944 ;
  assign n54946 = n8655 ^ n4146 ^ 1'b0 ;
  assign n54947 = n491 & ~n54946 ;
  assign n54948 = n7354 & n54947 ;
  assign n54949 = n52535 ^ n44363 ^ n20371 ;
  assign n54950 = ( n11934 & ~n12298 ) | ( n11934 & n54949 ) | ( ~n12298 & n54949 ) ;
  assign n54951 = ~n2551 & n22751 ;
  assign n54952 = n41153 & ~n54951 ;
  assign n54953 = n23099 ^ n2719 ^ 1'b0 ;
  assign n54954 = n34401 ^ n31530 ^ 1'b0 ;
  assign n54955 = n25900 | n54954 ;
  assign n54956 = n54955 ^ n51283 ^ 1'b0 ;
  assign n54957 = ~n27029 & n54956 ;
  assign n54958 = n4685 & ~n12375 ;
  assign n54959 = n36322 ^ n33843 ^ 1'b0 ;
  assign n54960 = n2660 & ~n54959 ;
  assign n54961 = n10108 ^ n8937 ^ n607 ;
  assign n54962 = ~n34239 & n54961 ;
  assign n54963 = ~n9774 & n54962 ;
  assign n54964 = n45867 ^ n35057 ^ 1'b0 ;
  assign n54965 = n5944 & ~n54964 ;
  assign n54966 = n4830 | n53140 ;
  assign n54967 = n4247 ^ n3997 ^ n1046 ;
  assign n54968 = n54967 ^ n37957 ^ 1'b0 ;
  assign n54969 = n46903 ^ n37214 ^ n2177 ;
  assign n54970 = n37897 ^ n29154 ^ 1'b0 ;
  assign n54971 = n4772 & n48956 ;
  assign n54972 = ~n25499 & n54971 ;
  assign n54973 = ~n942 & n38747 ;
  assign n54974 = n20430 & n42041 ;
  assign n54975 = n54974 ^ n20641 ^ 1'b0 ;
  assign n54977 = n17658 ^ n14893 ^ 1'b0 ;
  assign n54978 = ~n31306 & n54977 ;
  assign n54976 = n16459 & n52397 ;
  assign n54979 = n54978 ^ n54976 ^ 1'b0 ;
  assign n54980 = n20019 ^ n7307 ^ 1'b0 ;
  assign n54981 = ~n15058 & n54980 ;
  assign n54982 = n19370 ^ n9538 ^ 1'b0 ;
  assign n54983 = n43430 | n54982 ;
  assign n54984 = ~n21723 & n30542 ;
  assign n54985 = n54984 ^ n52360 ^ 1'b0 ;
  assign n54986 = n6477 | n11079 ;
  assign n54987 = n7751 & n9228 ;
  assign n54988 = ( n14719 & n46747 ) | ( n14719 & ~n54987 ) | ( n46747 & ~n54987 ) ;
  assign n54989 = n593 | n4083 ;
  assign n54990 = n33619 & ~n54989 ;
  assign n54995 = n13208 ^ n119 ^ 1'b0 ;
  assign n54991 = ( ~n686 & n22157 ) | ( ~n686 & n23876 ) | ( n22157 & n23876 ) ;
  assign n54992 = n4542 & n54991 ;
  assign n54993 = n54992 ^ n26950 ^ 1'b0 ;
  assign n54994 = ~n11231 & n54993 ;
  assign n54996 = n54995 ^ n54994 ^ 1'b0 ;
  assign n54997 = n34001 ^ n1410 ^ 1'b0 ;
  assign n54998 = n6000 & ~n54997 ;
  assign n55000 = ~n8266 & n38497 ;
  assign n55001 = n55000 ^ n23743 ^ 1'b0 ;
  assign n54999 = ( n28827 & n36626 ) | ( n28827 & n39608 ) | ( n36626 & n39608 ) ;
  assign n55002 = n55001 ^ n54999 ^ 1'b0 ;
  assign n55003 = n10071 & ~n52378 ;
  assign n55004 = ~n1272 & n55003 ;
  assign n55005 = ~n29231 & n47890 ;
  assign n55006 = ~n30373 & n55005 ;
  assign n55007 = n2602 | n13620 ;
  assign n55008 = n55007 ^ n52622 ^ 1'b0 ;
  assign n55009 = ( n11782 & n33648 ) | ( n11782 & ~n55008 ) | ( n33648 & ~n55008 ) ;
  assign n55010 = n8142 & n16390 ;
  assign n55011 = n55010 ^ n24268 ^ 1'b0 ;
  assign n55012 = n12885 | n18416 ;
  assign n55013 = n55011 | n55012 ;
  assign n55014 = n7110 | n55013 ;
  assign n55015 = n2105 ^ n1826 ^ 1'b0 ;
  assign n55016 = n2271 & ~n55015 ;
  assign n55017 = n3342 & ~n15173 ;
  assign n55018 = n55017 ^ n7971 ^ 1'b0 ;
  assign n55019 = n10415 ^ n278 ^ 1'b0 ;
  assign n55020 = n17293 ^ n11138 ^ 1'b0 ;
  assign n55021 = n55019 & ~n55020 ;
  assign n55022 = n22611 ^ n20831 ^ 1'b0 ;
  assign n55023 = n8909 & n13081 ;
  assign n55024 = n48709 & n55023 ;
  assign n55025 = ~n10127 & n18268 ;
  assign n55026 = n55025 ^ n37161 ^ 1'b0 ;
  assign n55027 = n55026 ^ n49782 ^ 1'b0 ;
  assign n55028 = n48518 & n55027 ;
  assign n55029 = n15364 & ~n25984 ;
  assign n55030 = n55029 ^ n2449 ^ 1'b0 ;
  assign n55031 = n23852 ^ n4275 ^ n458 ;
  assign n55032 = n47681 ^ n30975 ^ 1'b0 ;
  assign n55033 = n55031 | n55032 ;
  assign n55034 = n17700 | n26850 ;
  assign n55035 = ( n40973 & ~n48021 ) | ( n40973 & n55034 ) | ( ~n48021 & n55034 ) ;
  assign n55036 = ( n24601 & n32486 ) | ( n24601 & n38230 ) | ( n32486 & n38230 ) ;
  assign n55037 = n55036 ^ n4922 ^ 1'b0 ;
  assign n55038 = n38713 | n55037 ;
  assign n55039 = n55035 & ~n55038 ;
  assign n55040 = n8242 & ~n51713 ;
  assign n55042 = n25371 | n37653 ;
  assign n55043 = n47852 | n55042 ;
  assign n55041 = n7868 | n13992 ;
  assign n55044 = n55043 ^ n55041 ^ 1'b0 ;
  assign n55045 = n3848 | n18399 ;
  assign n55046 = n8615 | n55045 ;
  assign n55047 = n55046 ^ n18651 ^ 1'b0 ;
  assign n55048 = n48789 ^ n28728 ^ n19350 ;
  assign n55049 = n55048 ^ n2120 ^ 1'b0 ;
  assign n55050 = n36490 | n38352 ;
  assign n55051 = n16398 & ~n28600 ;
  assign n55052 = ~n5037 & n18419 ;
  assign n55053 = ~n863 & n55052 ;
  assign n55054 = n55051 | n55053 ;
  assign n55055 = n15972 & n26382 ;
  assign n55056 = ~n39867 & n55055 ;
  assign n55057 = n35419 | n41231 ;
  assign n55058 = n34337 & ~n55057 ;
  assign n55059 = n6846 & ~n16557 ;
  assign n55060 = ~n14207 & n55059 ;
  assign n55061 = ~n11727 & n49387 ;
  assign n55062 = n24155 ^ n9724 ^ 1'b0 ;
  assign n55063 = n8281 & ~n55062 ;
  assign n55064 = n26426 ^ n4168 ^ 1'b0 ;
  assign n55065 = ~n6498 & n55064 ;
  assign n55066 = ~n55063 & n55065 ;
  assign n55067 = n6607 & ~n32432 ;
  assign n55068 = n18634 & n37396 ;
  assign n55069 = n6691 ^ n2230 ^ x3 ;
  assign n55070 = n55069 ^ n6343 ^ 1'b0 ;
  assign n55071 = n55070 ^ n46605 ^ 1'b0 ;
  assign n55072 = n3112 & ~n55071 ;
  assign n55073 = n6128 & n55072 ;
  assign n55074 = ( n10218 & n38825 ) | ( n10218 & ~n40679 ) | ( n38825 & ~n40679 ) ;
  assign n55075 = ( n12442 & ~n32908 ) | ( n12442 & n55074 ) | ( ~n32908 & n55074 ) ;
  assign n55076 = n17898 ^ n16189 ^ 1'b0 ;
  assign n55077 = ~n13885 & n55076 ;
  assign n55078 = n22979 & n49186 ;
  assign n55079 = n9184 & n15472 ;
  assign n55080 = n3773 | n34428 ;
  assign n55081 = n55079 | n55080 ;
  assign n55082 = n41474 ^ n40697 ^ 1'b0 ;
  assign n55083 = ( ~n4877 & n34839 ) | ( ~n4877 & n37064 ) | ( n34839 & n37064 ) ;
  assign n55084 = n53603 ^ n1364 ^ 1'b0 ;
  assign n55085 = n19021 ^ n15179 ^ 1'b0 ;
  assign n55086 = n7295 | n55085 ;
  assign n55087 = n23035 | n49425 ;
  assign n55088 = n13207 | n55087 ;
  assign n55089 = n40248 ^ n38809 ^ n28435 ;
  assign n55090 = n44580 & n55089 ;
  assign n55091 = n44661 ^ n35884 ^ 1'b0 ;
  assign n55092 = n8968 | n55091 ;
  assign n55093 = n5552 & ~n55092 ;
  assign n55094 = ~n33153 & n55093 ;
  assign n55095 = n22913 ^ n18247 ^ n1723 ;
  assign n55096 = n55095 ^ n39195 ^ 1'b0 ;
  assign n55097 = ( n3257 & n12964 ) | ( n3257 & n22327 ) | ( n12964 & n22327 ) ;
  assign n55098 = n25253 ^ n8163 ^ 1'b0 ;
  assign n55099 = n53859 ^ n11720 ^ 1'b0 ;
  assign n55100 = ~n15109 & n55099 ;
  assign n55101 = n23910 ^ n7493 ^ 1'b0 ;
  assign n55102 = n37318 ^ n26829 ^ 1'b0 ;
  assign n55103 = n4806 ^ n117 ^ 1'b0 ;
  assign n55104 = n37581 ^ n30509 ^ 1'b0 ;
  assign n55105 = n8086 & ~n52358 ;
  assign n55106 = ~n25312 & n55105 ;
  assign n55107 = n55106 ^ n28188 ^ n434 ;
  assign n55108 = n27570 | n30313 ;
  assign n55109 = n25494 | n43562 ;
  assign n55110 = n55109 ^ n20347 ^ 1'b0 ;
  assign n55111 = n777 & ~n55110 ;
  assign n55112 = n55108 & n55111 ;
  assign n55113 = n35455 ^ n23652 ^ 1'b0 ;
  assign n55114 = n4789 | n55113 ;
  assign n55115 = n732 & ~n7534 ;
  assign n55116 = n55115 ^ n5780 ^ 1'b0 ;
  assign n55117 = n1083 & n2147 ;
  assign n55118 = n55117 ^ n14479 ^ n9781 ;
  assign n55119 = n24705 | n55118 ;
  assign n55120 = n46327 ^ n31678 ^ n13078 ;
  assign n55121 = n55120 ^ n38317 ^ 1'b0 ;
  assign n55122 = n30998 & ~n55121 ;
  assign n55123 = n55119 & n55122 ;
  assign n55124 = n8421 & ~n55123 ;
  assign n55125 = n55124 ^ n7298 ^ 1'b0 ;
  assign n55126 = n17861 | n38278 ;
  assign n55127 = ( n45586 & n54244 ) | ( n45586 & ~n55126 ) | ( n54244 & ~n55126 ) ;
  assign n55128 = n39096 ^ n35682 ^ n17039 ;
  assign n55129 = n55128 ^ n18045 ^ n5573 ;
  assign n55130 = n38504 ^ n12868 ^ 1'b0 ;
  assign n55131 = n39168 ^ n21744 ^ 1'b0 ;
  assign n55132 = ~n43501 & n55131 ;
  assign n55133 = n6581 & n30472 ;
  assign n55134 = n6866 & n55133 ;
  assign n55135 = n28712 | n55134 ;
  assign n55136 = n39462 & ~n55135 ;
  assign n55137 = n4599 | n30839 ;
  assign n55138 = n30552 ^ n14135 ^ 1'b0 ;
  assign n55139 = n42636 ^ n13559 ^ 1'b0 ;
  assign n55140 = n55138 & n55139 ;
  assign n55141 = n21550 | n43308 ;
  assign n55142 = n18643 & n37697 ;
  assign n55143 = n55142 ^ n7668 ^ 1'b0 ;
  assign n55144 = n26214 & n53511 ;
  assign n55145 = ~n55143 & n55144 ;
  assign n55146 = n3515 & n54891 ;
  assign n55147 = n55146 ^ n3336 ^ 1'b0 ;
  assign n55148 = n20706 ^ n17247 ^ 1'b0 ;
  assign n55149 = n14479 ^ n1060 ^ 1'b0 ;
  assign n55150 = n49163 & ~n55149 ;
  assign n55151 = ~n5402 & n32585 ;
  assign n55152 = n19695 & n55151 ;
  assign n55153 = n2570 & n20855 ;
  assign n55154 = n55153 ^ n16398 ^ 1'b0 ;
  assign n55155 = n29406 | n38688 ;
  assign n55156 = n21476 | n44713 ;
  assign n55157 = n43528 | n55156 ;
  assign n55158 = n46271 ^ n43131 ^ 1'b0 ;
  assign n55159 = n3698 & ~n21968 ;
  assign n55160 = n55159 ^ n15383 ^ 1'b0 ;
  assign n55161 = ~n8150 & n29194 ;
  assign n55162 = ~n6171 & n18648 ;
  assign n55163 = n32125 | n46534 ;
  assign n55164 = n53947 | n55163 ;
  assign n55165 = n10517 | n11969 ;
  assign n55166 = n17001 & n55165 ;
  assign n55167 = n36535 ^ n21573 ^ n3608 ;
  assign n55168 = n37691 ^ n14460 ^ n12890 ;
  assign n55169 = n27978 ^ n17110 ^ n2080 ;
  assign n55170 = n39976 ^ n10528 ^ 1'b0 ;
  assign n55171 = ( ~n1463 & n25612 ) | ( ~n1463 & n55170 ) | ( n25612 & n55170 ) ;
  assign n55172 = n45517 ^ n30189 ^ 1'b0 ;
  assign n55173 = n24116 & n55172 ;
  assign n55174 = n15083 & ~n22128 ;
  assign n55175 = ~n7017 & n55174 ;
  assign n55176 = n55175 ^ n494 ^ 1'b0 ;
  assign n55177 = n7273 | n28204 ;
  assign n55178 = n37778 & ~n55177 ;
  assign n55179 = ( n5506 & ~n12284 ) | ( n5506 & n49857 ) | ( ~n12284 & n49857 ) ;
  assign n55180 = n55179 ^ n49179 ^ n777 ;
  assign n55181 = ~n2733 & n55180 ;
  assign n55183 = n848 & n24897 ;
  assign n55184 = ~n9273 & n55183 ;
  assign n55182 = n523 & ~n31279 ;
  assign n55185 = n55184 ^ n55182 ^ 1'b0 ;
  assign n55186 = n19852 ^ n17199 ^ n9321 ;
  assign n55187 = n33299 | n49086 ;
  assign n55188 = n8864 ^ n5625 ^ 1'b0 ;
  assign n55189 = n51853 & ~n55188 ;
  assign n55190 = ( n16567 & n55187 ) | ( n16567 & n55189 ) | ( n55187 & n55189 ) ;
  assign n55191 = n8455 ^ n4055 ^ 1'b0 ;
  assign n55192 = n11535 | n55191 ;
  assign n55193 = n3624 | n53531 ;
  assign n55194 = n48235 ^ n6844 ^ 1'b0 ;
  assign n55195 = n33587 ^ n33349 ^ 1'b0 ;
  assign n55196 = n7142 & ~n55195 ;
  assign n55197 = n55196 ^ n1794 ^ 1'b0 ;
  assign n55198 = n11486 ^ n8265 ^ n6343 ;
  assign n55199 = ~n3632 & n9773 ;
  assign n55200 = n10769 & n49877 ;
  assign n55201 = n51679 ^ n44 ^ 1'b0 ;
  assign n55202 = n37067 | n55201 ;
  assign n55203 = n7316 ^ n2905 ^ 1'b0 ;
  assign n55204 = n51342 & n55203 ;
  assign n55205 = n2001 & ~n3475 ;
  assign n55206 = n5316 & n55205 ;
  assign n55207 = n3240 | n10485 ;
  assign n55208 = ( n35046 & n35552 ) | ( n35046 & ~n55207 ) | ( n35552 & ~n55207 ) ;
  assign n55209 = n55206 & n55208 ;
  assign n55210 = n2960 | n9006 ;
  assign n55211 = n55210 ^ n35945 ^ n8919 ;
  assign n55212 = n55211 ^ n13684 ^ 1'b0 ;
  assign n55220 = n4317 & ~n10163 ;
  assign n55221 = n33913 & n55220 ;
  assign n55213 = n12259 ^ n12145 ^ n8945 ;
  assign n55214 = n33137 & ~n55213 ;
  assign n55215 = n13591 & n55214 ;
  assign n55216 = n4333 ^ n617 ^ 1'b0 ;
  assign n55217 = ~n25080 & n55216 ;
  assign n55218 = ~n17664 & n55217 ;
  assign n55219 = ( ~n1138 & n55215 ) | ( ~n1138 & n55218 ) | ( n55215 & n55218 ) ;
  assign n55222 = n55221 ^ n55219 ^ 1'b0 ;
  assign n55223 = n3392 & n24783 ;
  assign n55224 = n24844 ^ n2435 ^ 1'b0 ;
  assign n55225 = n27417 & n32207 ;
  assign n55226 = n7014 & ~n55225 ;
  assign n55227 = ~n55224 & n55226 ;
  assign n55228 = ~n30707 & n46941 ;
  assign n55229 = n55228 ^ n6153 ^ 1'b0 ;
  assign n55230 = ~n38 & n33553 ;
  assign n55231 = ~n25260 & n55230 ;
  assign n55232 = n39387 ^ n16896 ^ 1'b0 ;
  assign n55233 = n9165 & n36091 ;
  assign n55234 = ~n55232 & n55233 ;
  assign n55235 = n2375 | n7087 ;
  assign n55236 = n17727 | n55235 ;
  assign n55237 = n28892 ^ n1186 ^ 1'b0 ;
  assign n55238 = n24558 ^ n8227 ^ n6426 ;
  assign n55239 = n7676 ^ n5924 ^ 1'b0 ;
  assign n55240 = n11802 | n55239 ;
  assign n55241 = n5094 | n55240 ;
  assign n55242 = n1035 & n6326 ;
  assign n55243 = n31343 ^ n11472 ^ 1'b0 ;
  assign n55244 = n25159 ^ n9528 ^ 1'b0 ;
  assign n55245 = n21290 | n55244 ;
  assign n55246 = n27307 | n43462 ;
  assign n55247 = ( n648 & ~n37024 ) | ( n648 & n53965 ) | ( ~n37024 & n53965 ) ;
  assign n55248 = n22612 | n43383 ;
  assign n55249 = ~n27258 & n55248 ;
  assign n55250 = n55249 ^ n34283 ^ 1'b0 ;
  assign n55251 = n55250 ^ n11009 ^ n3671 ;
  assign n55252 = n5898 & ~n37866 ;
  assign n55253 = n15552 & ~n50186 ;
  assign n55254 = ( n5010 & n55252 ) | ( n5010 & n55253 ) | ( n55252 & n55253 ) ;
  assign n55255 = n1562 | n35489 ;
  assign n55256 = n55255 ^ n6729 ^ 1'b0 ;
  assign n55257 = n4245 & n44359 ;
  assign n55258 = n33534 ^ n23666 ^ n5259 ;
  assign n55259 = n27560 ^ n1292 ^ 1'b0 ;
  assign n55260 = n40788 ^ n9292 ^ 1'b0 ;
  assign n55261 = n48576 ^ n32200 ^ n4192 ;
  assign n55262 = n55261 ^ n39458 ^ 1'b0 ;
  assign n55263 = n53866 ^ n5519 ^ n4183 ;
  assign n55266 = n21823 ^ n19696 ^ n709 ;
  assign n55267 = n13717 & ~n22064 ;
  assign n55268 = n55266 & n55267 ;
  assign n55264 = n4231 ^ n2689 ^ 1'b0 ;
  assign n55265 = n14757 | n55264 ;
  assign n55269 = n55268 ^ n55265 ^ n39899 ;
  assign n55270 = ( n47427 & n55263 ) | ( n47427 & ~n55269 ) | ( n55263 & ~n55269 ) ;
  assign n55271 = ( n55260 & n55262 ) | ( n55260 & ~n55270 ) | ( n55262 & ~n55270 ) ;
  assign n55272 = ~n15978 & n19182 ;
  assign n55273 = n55272 ^ n24108 ^ 1'b0 ;
  assign n55275 = n2370 & n15362 ;
  assign n55276 = n55275 ^ n15294 ^ 1'b0 ;
  assign n55277 = n20945 & n55276 ;
  assign n55278 = ~n38632 & n55277 ;
  assign n55274 = n28883 & ~n29608 ;
  assign n55279 = n55278 ^ n55274 ^ 1'b0 ;
  assign n55280 = n55279 ^ n20795 ^ 1'b0 ;
  assign n55281 = n12906 & n18447 ;
  assign n55282 = n8143 & n55281 ;
  assign n55283 = n55282 ^ n41159 ^ 1'b0 ;
  assign n55284 = n427 & n34966 ;
  assign n55285 = n55284 ^ n36023 ^ 1'b0 ;
  assign n55286 = ~n34989 & n55285 ;
  assign n55287 = ( n7917 & n16246 ) | ( n7917 & n46991 ) | ( n16246 & n46991 ) ;
  assign n55288 = n42878 ^ n5749 ^ 1'b0 ;
  assign n55289 = n2523 | n14969 ;
  assign n55290 = n55289 ^ n9322 ^ n5592 ;
  assign n55291 = n7996 | n11215 ;
  assign n55292 = n35908 ^ n5782 ^ 1'b0 ;
  assign n55293 = ~n55291 & n55292 ;
  assign n55294 = n7282 | n38907 ;
  assign n55295 = n29366 ^ n3648 ^ 1'b0 ;
  assign n55296 = n553 | n16391 ;
  assign n55297 = n55296 ^ n10396 ^ 1'b0 ;
  assign n55298 = n55297 ^ n34450 ^ 1'b0 ;
  assign n55299 = n34576 ^ n33195 ^ n20729 ;
  assign n55300 = n888 | n55299 ;
  assign n55301 = ~n718 & n21985 ;
  assign n55302 = n55301 ^ n4696 ^ 1'b0 ;
  assign n55303 = n37870 ^ n11867 ^ n4505 ;
  assign n55304 = n55302 | n55303 ;
  assign n55305 = n7728 & ~n28511 ;
  assign n55306 = n55305 ^ n41703 ^ 1'b0 ;
  assign n55308 = n5053 & n38218 ;
  assign n55307 = n17605 & ~n17700 ;
  assign n55309 = n55308 ^ n55307 ^ 1'b0 ;
  assign n55310 = n43688 ^ n35719 ^ n892 ;
  assign n55311 = n50044 ^ n29769 ^ 1'b0 ;
  assign n55312 = n3128 & ~n55311 ;
  assign n55313 = n55312 ^ n33690 ^ n5569 ;
  assign n55314 = n6804 | n48475 ;
  assign n55315 = n53338 | n55314 ;
  assign n55316 = n1436 & ~n11633 ;
  assign n55317 = n8950 & n55316 ;
  assign n55318 = n55317 ^ n4953 ^ 1'b0 ;
  assign n55319 = ~n685 & n50900 ;
  assign n55320 = n43124 ^ n31423 ^ 1'b0 ;
  assign n55321 = n4056 & n11919 ;
  assign n55322 = n13576 & n55321 ;
  assign n55323 = n54400 | n55322 ;
  assign n55324 = n12867 & n55323 ;
  assign n55325 = n40699 ^ n33270 ^ n28883 ;
  assign n55326 = n47983 ^ n44600 ^ 1'b0 ;
  assign n55327 = ( n15767 & ~n28100 ) | ( n15767 & n55326 ) | ( ~n28100 & n55326 ) ;
  assign n55328 = ( n4004 & n7141 ) | ( n4004 & n15580 ) | ( n7141 & n15580 ) ;
  assign n55329 = n55328 ^ n10046 ^ n2257 ;
  assign n55330 = n24531 ^ n20513 ^ 1'b0 ;
  assign n55331 = n17339 & n55330 ;
  assign n55332 = n16388 & ~n31675 ;
  assign n55333 = ~n14712 & n55332 ;
  assign n55334 = n55331 | n55333 ;
  assign n55335 = n532 & ~n38522 ;
  assign n55336 = n6217 | n15189 ;
  assign n55337 = n6217 & ~n55336 ;
  assign n55338 = n55337 ^ n32553 ^ n11874 ;
  assign n55339 = n22783 ^ n7419 ^ 1'b0 ;
  assign n55340 = n20436 & n55339 ;
  assign n55341 = n13393 & n55340 ;
  assign n55342 = ~n55338 & n55341 ;
  assign n55343 = n39595 ^ n6361 ^ 1'b0 ;
  assign n55344 = ~n18454 & n55343 ;
  assign n55345 = ( ~n36746 & n41908 ) | ( ~n36746 & n46626 ) | ( n41908 & n46626 ) ;
  assign n55346 = ~n23901 & n55345 ;
  assign n55347 = n55346 ^ n19216 ^ 1'b0 ;
  assign n55348 = n4502 & ~n9704 ;
  assign n55349 = n54331 & n55348 ;
  assign n55350 = n37201 ^ n13088 ^ n5740 ;
  assign n55351 = n3730 & ~n36886 ;
  assign n55352 = n4497 & ~n34249 ;
  assign n55353 = n3358 & ~n52778 ;
  assign n55354 = n55353 ^ n43817 ^ 1'b0 ;
  assign n55355 = n38593 ^ n17130 ^ n3312 ;
  assign n55356 = n55355 ^ n48577 ^ n492 ;
  assign n55357 = ~n20545 & n25515 ;
  assign n55358 = ~n55356 & n55357 ;
  assign n55359 = n19527 ^ n4385 ^ n835 ;
  assign n55360 = n55359 ^ n16171 ^ n8709 ;
  assign n55361 = n15741 ^ n4140 ^ 1'b0 ;
  assign n55362 = n55360 | n55361 ;
  assign n55363 = n9081 | n33756 ;
  assign n55366 = n13736 & n48396 ;
  assign n55364 = n15748 ^ n11778 ^ 1'b0 ;
  assign n55365 = n55364 ^ n51172 ^ n18969 ;
  assign n55367 = n55366 ^ n55365 ^ 1'b0 ;
  assign n55368 = n48144 ^ n6524 ^ 1'b0 ;
  assign n55369 = ( ~n6504 & n43645 ) | ( ~n6504 & n55368 ) | ( n43645 & n55368 ) ;
  assign n55370 = n10845 ^ n3187 ^ 1'b0 ;
  assign n55371 = ( n19294 & n39595 ) | ( n19294 & ~n55370 ) | ( n39595 & ~n55370 ) ;
  assign n55372 = ~n1031 & n54141 ;
  assign n55373 = n55372 ^ n26673 ^ 1'b0 ;
  assign n55374 = n20607 & ~n51660 ;
  assign n55375 = n49436 ^ n23798 ^ 1'b0 ;
  assign n55376 = ~n55374 & n55375 ;
  assign n55377 = n11573 & n30574 ;
  assign n55378 = n30989 | n54309 ;
  assign n55379 = n27767 & ~n55378 ;
  assign n55380 = n3355 | n50059 ;
  assign n55381 = ( n12106 & ~n17851 ) | ( n12106 & n51599 ) | ( ~n17851 & n51599 ) ;
  assign n55382 = n7514 ^ n1817 ^ 1'b0 ;
  assign n55383 = ~n37119 & n55382 ;
  assign n55384 = ( n1679 & n27178 ) | ( n1679 & ~n55383 ) | ( n27178 & ~n55383 ) ;
  assign n55385 = ~n5175 & n16629 ;
  assign n55386 = ~n21521 & n30926 ;
  assign n55387 = ~n30919 & n55386 ;
  assign n55388 = n15646 & n31328 ;
  assign n55389 = n55388 ^ n14071 ^ 1'b0 ;
  assign n55390 = n55389 ^ n53981 ^ 1'b0 ;
  assign n55391 = ~n7479 & n55390 ;
  assign n55392 = n31011 | n55391 ;
  assign n55393 = n4185 & n12502 ;
  assign n55394 = n1926 & n55393 ;
  assign n55395 = ~n17354 & n20105 ;
  assign n55396 = ~n37406 & n55395 ;
  assign n55397 = n55396 ^ n21163 ^ 1'b0 ;
  assign n55398 = ( n45593 & n49883 ) | ( n45593 & n51002 ) | ( n49883 & n51002 ) ;
  assign n55399 = n36865 | n55398 ;
  assign n55400 = n5069 & n14067 ;
  assign n55401 = n53534 ^ n22639 ^ 1'b0 ;
  assign n55402 = n55400 & ~n55401 ;
  assign n55403 = n37214 & n39489 ;
  assign n55404 = ( ~n523 & n2304 ) | ( ~n523 & n29314 ) | ( n2304 & n29314 ) ;
  assign n55405 = n27474 ^ n1614 ^ 1'b0 ;
  assign n55406 = n6076 | n17778 ;
  assign n55407 = n2333 | n55406 ;
  assign n55408 = ( n252 & n18548 ) | ( n252 & n55407 ) | ( n18548 & n55407 ) ;
  assign n55409 = n31330 & ~n55408 ;
  assign n55410 = n44288 | n55409 ;
  assign n55411 = n55410 ^ n4631 ^ 1'b0 ;
  assign n55412 = n55411 ^ n17961 ^ 1'b0 ;
  assign n55413 = n10312 | n55412 ;
  assign n55414 = n3898 & ~n26879 ;
  assign n55415 = n55414 ^ n16823 ^ 1'b0 ;
  assign n55416 = n1546 | n6710 ;
  assign n55417 = n55415 | n55416 ;
  assign n55418 = n23726 ^ n22658 ^ 1'b0 ;
  assign n55419 = n13768 | n55418 ;
  assign n55420 = n55419 ^ n46442 ^ 1'b0 ;
  assign n55421 = n2808 & ~n19379 ;
  assign n55422 = ~n36194 & n55421 ;
  assign n55423 = n15861 & ~n28409 ;
  assign n55424 = n55423 ^ n49924 ^ 1'b0 ;
  assign n55425 = n37914 ^ n7358 ^ 1'b0 ;
  assign n55426 = n8485 & ~n36730 ;
  assign n55427 = n5661 & ~n13614 ;
  assign n55428 = n39581 & n55427 ;
  assign n55429 = n16589 & ~n46668 ;
  assign n55430 = n49289 & n55429 ;
  assign n55431 = n11915 ^ n11062 ^ n4275 ;
  assign n55432 = n55431 ^ n55328 ^ 1'b0 ;
  assign n55433 = n20753 | n55432 ;
  assign n55434 = ~n16006 & n22788 ;
  assign n55435 = ~n43443 & n55434 ;
  assign n55436 = n20206 | n34547 ;
  assign n55437 = n55436 ^ n45905 ^ 1'b0 ;
  assign n55438 = n3175 & ~n26250 ;
  assign n55439 = n26944 & ~n45251 ;
  assign n55440 = n54273 ^ n25126 ^ n3901 ;
  assign n55441 = n32703 & n32825 ;
  assign n55442 = ~n34049 & n39940 ;
  assign n55443 = ( n55440 & ~n55441 ) | ( n55440 & n55442 ) | ( ~n55441 & n55442 ) ;
  assign n55444 = n19909 ^ n11369 ^ 1'b0 ;
  assign n55445 = n6078 & n6640 ;
  assign n55446 = ~n14258 & n55445 ;
  assign n55447 = n25903 | n55446 ;
  assign n55448 = n55447 ^ n14905 ^ 1'b0 ;
  assign n55449 = n26004 | n55448 ;
  assign n55450 = n2531 & n54722 ;
  assign n55451 = ~n15403 & n55450 ;
  assign n55452 = n34542 | n43481 ;
  assign n55453 = n55452 ^ n40931 ^ 1'b0 ;
  assign n55454 = n2504 & ~n55453 ;
  assign n55455 = n26288 ^ n11021 ^ n3950 ;
  assign n55456 = n44390 & ~n45541 ;
  assign n55457 = n55456 ^ n845 ^ 1'b0 ;
  assign n55458 = n55455 | n55457 ;
  assign n55459 = n55458 ^ n3294 ^ 1'b0 ;
  assign n55460 = n10085 & ~n31588 ;
  assign n55461 = n33128 ^ n8775 ^ 1'b0 ;
  assign n55462 = n31901 ^ n3339 ^ 1'b0 ;
  assign n55463 = n14282 ^ n2201 ^ 1'b0 ;
  assign n55464 = n37313 ^ n416 ^ 1'b0 ;
  assign n55465 = n28191 | n55464 ;
  assign n55466 = n14962 ^ n2232 ^ n345 ;
  assign n55467 = n39235 & n55466 ;
  assign n55468 = n38265 & n55467 ;
  assign n55469 = n44163 ^ n38437 ^ 1'b0 ;
  assign n55470 = n52888 ^ n15376 ^ 1'b0 ;
  assign n55471 = n15395 & ~n55470 ;
  assign n55472 = n19191 ^ n2211 ^ 1'b0 ;
  assign n55473 = n3358 & n55472 ;
  assign n55474 = n24140 ^ n21832 ^ n10326 ;
  assign n55475 = ( n10091 & n55473 ) | ( n10091 & ~n55474 ) | ( n55473 & ~n55474 ) ;
  assign n55476 = x7 & n1698 ;
  assign n55477 = ~x7 & n55476 ;
  assign n55478 = ~n2328 & n55477 ;
  assign n55479 = n5195 & ~n55478 ;
  assign n55480 = ~n345 & n9623 ;
  assign n55481 = ~n9623 & n55480 ;
  assign n55482 = n829 & ~n55481 ;
  assign n55483 = n55479 | n55482 ;
  assign n55484 = n12413 & n55483 ;
  assign n55485 = n35342 ^ n15043 ^ 1'b0 ;
  assign n55486 = n108 & n415 ;
  assign n55487 = n41259 & n55486 ;
  assign n55488 = n30315 | n48958 ;
  assign n55489 = n26470 ^ n10134 ^ 1'b0 ;
  assign n55490 = ~n55488 & n55489 ;
  assign n55491 = ( n2504 & n22847 ) | ( n2504 & n24661 ) | ( n22847 & n24661 ) ;
  assign n55492 = n24674 | n55491 ;
  assign n55493 = n40622 ^ n13164 ^ 1'b0 ;
  assign n55494 = n41776 ^ n21242 ^ 1'b0 ;
  assign n55496 = n37588 | n38054 ;
  assign n55495 = n6709 & n23580 ;
  assign n55497 = n55496 ^ n55495 ^ 1'b0 ;
  assign n55498 = n14843 ^ n10374 ^ n8511 ;
  assign n55499 = ~n736 & n55498 ;
  assign n55500 = ~n7168 & n55499 ;
  assign n55501 = n36599 ^ n33819 ^ 1'b0 ;
  assign n55502 = n16973 & ~n39572 ;
  assign n55503 = n55502 ^ n25578 ^ 1'b0 ;
  assign n55504 = n43959 ^ n25601 ^ 1'b0 ;
  assign n55505 = n3180 & n55504 ;
  assign n55506 = n55503 | n55505 ;
  assign n55507 = ( ~n10519 & n46604 ) | ( ~n10519 & n55506 ) | ( n46604 & n55506 ) ;
  assign n55508 = n24809 | n25766 ;
  assign n55509 = n6004 | n55508 ;
  assign n55510 = n23550 & n55509 ;
  assign n55511 = n55510 ^ n36604 ^ n2432 ;
  assign n55512 = n11804 & ~n45121 ;
  assign n55513 = ~n17230 & n55512 ;
  assign n55514 = n55513 ^ n13011 ^ 1'b0 ;
  assign n55515 = ~n53717 & n55514 ;
  assign n55517 = n22004 ^ n8281 ^ 1'b0 ;
  assign n55518 = ~n35213 & n55517 ;
  assign n55516 = n15111 & ~n17204 ;
  assign n55519 = n55518 ^ n55516 ^ 1'b0 ;
  assign n55520 = n21037 ^ n13013 ^ 1'b0 ;
  assign n55523 = n55210 ^ n8919 ^ 1'b0 ;
  assign n55522 = n655 & ~n22261 ;
  assign n55524 = n55523 ^ n55522 ^ 1'b0 ;
  assign n55521 = n22907 ^ n3464 ^ 1'b0 ;
  assign n55525 = n55524 ^ n55521 ^ n7391 ;
  assign n55526 = n55525 ^ n33089 ^ n8756 ;
  assign n55527 = n55526 ^ n48397 ^ 1'b0 ;
  assign n55528 = n42677 ^ n39698 ^ n38985 ;
  assign n55529 = n8657 & ~n12770 ;
  assign n55530 = n55529 ^ n41125 ^ 1'b0 ;
  assign n55531 = n24707 | n52418 ;
  assign n55532 = n11097 & n16321 ;
  assign n55533 = n46 & ~n55532 ;
  assign n55534 = n55533 ^ n41931 ^ 1'b0 ;
  assign n55535 = ~n9072 & n39913 ;
  assign n55536 = ( n18184 & n25184 ) | ( n18184 & ~n32150 ) | ( n25184 & ~n32150 ) ;
  assign n55537 = n36940 | n55536 ;
  assign n55538 = n55535 & ~n55537 ;
  assign n55539 = n13947 ^ n5713 ^ 1'b0 ;
  assign n55540 = n6131 | n20475 ;
  assign n55541 = n55540 ^ n17236 ^ 1'b0 ;
  assign n55542 = n24681 | n40327 ;
  assign n55543 = n26165 | n55542 ;
  assign n55544 = n14127 ^ n3591 ^ 1'b0 ;
  assign n55545 = n14917 & n16642 ;
  assign n55546 = ~n46509 & n49885 ;
  assign n55547 = n49152 ^ n42232 ^ n28250 ;
  assign n55548 = n19383 & ~n55547 ;
  assign n55549 = n55548 ^ n18248 ^ 1'b0 ;
  assign n55550 = ( n32199 & n36983 ) | ( n32199 & ~n55549 ) | ( n36983 & ~n55549 ) ;
  assign n55551 = n2405 & ~n46584 ;
  assign n55552 = ~n9918 & n55551 ;
  assign n55553 = n55552 ^ n50889 ^ n12668 ;
  assign n55554 = n3560 & n38447 ;
  assign n55555 = n51739 ^ n46716 ^ n20268 ;
  assign n55556 = n19038 | n55555 ;
  assign n55557 = n24912 ^ n2873 ^ 1'b0 ;
  assign n55558 = n27000 ^ n22403 ^ 1'b0 ;
  assign n55559 = n5747 & n55558 ;
  assign n55560 = n21878 & n55559 ;
  assign n55561 = n55557 & n55560 ;
  assign n55562 = n11275 | n55561 ;
  assign n55563 = n55562 ^ n9339 ^ 1'b0 ;
  assign n55565 = n7796 ^ n7028 ^ 1'b0 ;
  assign n55566 = n3266 & n55565 ;
  assign n55564 = n8097 & ~n29720 ;
  assign n55567 = n55566 ^ n55564 ^ 1'b0 ;
  assign n55568 = ( n434 & ~n38683 ) | ( n434 & n44601 ) | ( ~n38683 & n44601 ) ;
  assign n55569 = n39642 ^ n29652 ^ n82 ;
  assign n55570 = n55569 ^ n18299 ^ 1'b0 ;
  assign n55571 = n40795 | n55570 ;
  assign n55572 = n55571 ^ n23208 ^ 1'b0 ;
  assign n55573 = n55568 | n55572 ;
  assign n55574 = n9415 & n15005 ;
  assign n55575 = n55574 ^ n25455 ^ 1'b0 ;
  assign n55576 = n45565 ^ n3054 ^ 1'b0 ;
  assign n55577 = n20425 ^ n7033 ^ 1'b0 ;
  assign n55578 = n26977 | n55577 ;
  assign n55579 = n10224 & n26847 ;
  assign n55580 = n10345 & n13523 ;
  assign n55581 = n17542 ^ n10288 ^ 1'b0 ;
  assign n55582 = n15638 | n22546 ;
  assign n55583 = n3973 & n36985 ;
  assign n55584 = n39357 ^ n10975 ^ 1'b0 ;
  assign n55585 = n20209 & n55584 ;
  assign n55586 = ( ~n44646 & n55583 ) | ( ~n44646 & n55585 ) | ( n55583 & n55585 ) ;
  assign n55587 = n18836 | n22929 ;
  assign n55588 = ( n7534 & ~n10320 ) | ( n7534 & n17692 ) | ( ~n10320 & n17692 ) ;
  assign n55589 = n16070 & ~n19324 ;
  assign n55590 = n28378 ^ n8278 ^ 1'b0 ;
  assign n55591 = n50349 & ~n55590 ;
  assign n55593 = n12037 & ~n16138 ;
  assign n55592 = ~n25164 & n32554 ;
  assign n55594 = n55593 ^ n55592 ^ 1'b0 ;
  assign n55596 = n7038 | n25988 ;
  assign n55597 = n1006 & ~n55596 ;
  assign n55595 = n2174 & n48232 ;
  assign n55598 = n55597 ^ n55595 ^ 1'b0 ;
  assign n55599 = n15370 ^ n1527 ^ n1231 ;
  assign n55600 = ~n48440 & n55599 ;
  assign n55601 = n38134 ^ n5732 ^ 1'b0 ;
  assign n55602 = n1069 & ~n55601 ;
  assign n55603 = n34777 ^ n26997 ^ 1'b0 ;
  assign n55604 = n35036 ^ n22524 ^ 1'b0 ;
  assign n55605 = n2569 & ~n55604 ;
  assign n55606 = n4405 & n12191 ;
  assign n55607 = n40596 ^ n9924 ^ 1'b0 ;
  assign n55608 = ~n55606 & n55607 ;
  assign n55609 = ~n4840 & n46928 ;
  assign n55610 = n7293 & ~n49697 ;
  assign n55611 = n55610 ^ n31999 ^ 1'b0 ;
  assign n55612 = n29593 ^ n8557 ^ 1'b0 ;
  assign n55613 = n37212 ^ n10528 ^ 1'b0 ;
  assign n55614 = n55612 & n55613 ;
  assign n55615 = n46908 & n55614 ;
  assign n55616 = n55615 ^ n25045 ^ 1'b0 ;
  assign n55617 = n6168 | n55616 ;
  assign n55618 = n55617 ^ n54848 ^ 1'b0 ;
  assign n55619 = n45145 ^ n4240 ^ 1'b0 ;
  assign n55620 = n18819 & n39299 ;
  assign n55622 = n13688 & ~n17891 ;
  assign n55621 = n4363 | n28872 ;
  assign n55623 = n55622 ^ n55621 ^ 1'b0 ;
  assign n55624 = ( n13143 & n20612 ) | ( n13143 & ~n55623 ) | ( n20612 & ~n55623 ) ;
  assign n55625 = n10975 & ~n31744 ;
  assign n55626 = n29586 ^ n2258 ^ 1'b0 ;
  assign n55627 = n9392 & ~n55626 ;
  assign n55628 = n55627 ^ n16670 ^ n9146 ;
  assign n55629 = n25325 & n42829 ;
  assign n55630 = n41975 ^ n9678 ^ 1'b0 ;
  assign n55631 = n53398 & n55630 ;
  assign n55632 = n21301 ^ n20720 ^ n12161 ;
  assign n55633 = n33599 | n55632 ;
  assign n55634 = n34965 & n53158 ;
  assign n55635 = n1367 | n14014 ;
  assign n55636 = n55635 ^ n26561 ^ 1'b0 ;
  assign n55637 = n19897 & n30798 ;
  assign n55641 = ( n4207 & n12728 ) | ( n4207 & ~n16523 ) | ( n12728 & ~n16523 ) ;
  assign n55638 = n8874 & ~n15034 ;
  assign n55639 = n4077 & n55638 ;
  assign n55640 = n2449 | n55639 ;
  assign n55642 = n55641 ^ n55640 ^ 1'b0 ;
  assign n55643 = n55642 ^ n25881 ^ n676 ;
  assign n55644 = n574 & n43528 ;
  assign n55645 = n55644 ^ n29910 ^ 1'b0 ;
  assign n55646 = n4126 & n36033 ;
  assign n55647 = n25706 & n30816 ;
  assign n55648 = n16205 & ~n54739 ;
  assign n55649 = n55648 ^ n5419 ^ 1'b0 ;
  assign n55650 = n24905 ^ n3667 ^ 1'b0 ;
  assign n55651 = ~n22161 & n22173 ;
  assign n55652 = n55616 ^ n35882 ^ n17693 ;
  assign n55653 = ( n11164 & ~n39682 ) | ( n11164 & n55652 ) | ( ~n39682 & n55652 ) ;
  assign n55654 = n55651 | n55653 ;
  assign n55655 = n31132 ^ n9598 ^ 1'b0 ;
  assign n55656 = n2728 & n55655 ;
  assign n55657 = ( n3056 & ~n15772 ) | ( n3056 & n43816 ) | ( ~n15772 & n43816 ) ;
  assign n55658 = n23672 ^ n19559 ^ 1'b0 ;
  assign n55659 = n55657 & ~n55658 ;
  assign n55660 = n5741 & ~n26091 ;
  assign n55661 = ~n6166 & n55660 ;
  assign n55662 = n20496 ^ n10375 ^ 1'b0 ;
  assign n55663 = n55661 | n55662 ;
  assign n55664 = n10938 ^ n8603 ^ 1'b0 ;
  assign n55665 = ~n46271 & n55664 ;
  assign n55666 = n54972 ^ n4997 ^ 1'b0 ;
  assign n55667 = n31794 | n55666 ;
  assign n55668 = ( n32 & ~n13396 ) | ( n32 & n49470 ) | ( ~n13396 & n49470 ) ;
  assign n55669 = ~n4014 & n29162 ;
  assign n55670 = n953 & ~n5550 ;
  assign n55671 = n3428 & n55670 ;
  assign n55672 = n659 & n17531 ;
  assign n55673 = ~n30201 & n55672 ;
  assign n55674 = ( n49750 & n55671 ) | ( n49750 & n55673 ) | ( n55671 & n55673 ) ;
  assign n55675 = ~n38922 & n49050 ;
  assign n55676 = n55675 ^ n32266 ^ 1'b0 ;
  assign n55677 = ~n3199 & n9760 ;
  assign n55678 = n1186 | n17459 ;
  assign n55679 = n11555 | n55678 ;
  assign n55680 = n19982 & ~n55679 ;
  assign n55681 = n32873 ^ n18465 ^ 1'b0 ;
  assign n55682 = n38743 | n55681 ;
  assign n55683 = n6305 & n55682 ;
  assign n55684 = n36832 | n51329 ;
  assign n55685 = n5997 & n10950 ;
  assign n55686 = n55685 ^ n22706 ^ 1'b0 ;
  assign n55687 = n18812 ^ n8858 ^ 1'b0 ;
  assign n55688 = ( n28031 & n44831 ) | ( n28031 & n47550 ) | ( n44831 & n47550 ) ;
  assign n55689 = n14388 | n33091 ;
  assign n55690 = n31249 & ~n55689 ;
  assign n55691 = n1918 & n6282 ;
  assign n55692 = n37321 & n55691 ;
  assign n55693 = n954 & ~n1594 ;
  assign n55694 = n108 & n19931 ;
  assign n55695 = n48627 ^ n33782 ^ 1'b0 ;
  assign n55696 = n27759 & n55695 ;
  assign n55697 = n4810 & n46589 ;
  assign n55698 = ~n982 & n55697 ;
  assign n55699 = n1871 | n52494 ;
  assign n55700 = n55699 ^ n23941 ^ 1'b0 ;
  assign n55701 = ( ~n15328 & n19226 ) | ( ~n15328 & n33573 ) | ( n19226 & n33573 ) ;
  assign n55702 = n29650 | n55701 ;
  assign n55703 = ~n11788 & n53807 ;
  assign n55704 = n55703 ^ n32861 ^ 1'b0 ;
  assign n55705 = n21403 ^ n14048 ^ 1'b0 ;
  assign n55706 = ~n14202 & n25766 ;
  assign n55707 = ~n9055 & n15350 ;
  assign n55708 = n55707 ^ n20626 ^ 1'b0 ;
  assign n55709 = n4048 | n18351 ;
  assign n55710 = n9193 & ~n41344 ;
  assign n55711 = ~n55709 & n55710 ;
  assign n55712 = n55711 ^ n31195 ^ 1'b0 ;
  assign n55713 = ~n55708 & n55712 ;
  assign n55714 = n7818 | n17814 ;
  assign n55715 = n14895 & n55714 ;
  assign n55716 = n55715 ^ n24172 ^ 1'b0 ;
  assign n55717 = ~n6351 & n55716 ;
  assign n55718 = n32643 & n55717 ;
  assign n55719 = n34846 | n54158 ;
  assign n55720 = n27256 & n55719 ;
  assign n55721 = n6549 | n21195 ;
  assign n55722 = n26988 & ~n48533 ;
  assign n55723 = n55721 & n55722 ;
  assign n55724 = n15991 | n34251 ;
  assign n55725 = n8114 & ~n55724 ;
  assign n55726 = n55164 ^ n23390 ^ 1'b0 ;
  assign n55727 = n13433 & n35433 ;
  assign n55728 = n8996 ^ n4717 ^ 1'b0 ;
  assign n55729 = n18424 & n55728 ;
  assign n55730 = n55729 ^ n15953 ^ n5800 ;
  assign n55731 = n46655 ^ n7035 ^ 1'b0 ;
  assign n55732 = n55671 ^ n21980 ^ n12089 ;
  assign n55733 = n51067 ^ n24018 ^ 1'b0 ;
  assign n55734 = n2145 | n43405 ;
  assign n55735 = n9709 | n55734 ;
  assign n55736 = n953 | n10924 ;
  assign n55737 = n396 & ~n55736 ;
  assign n55738 = n2114 & ~n21350 ;
  assign n55739 = n7776 | n23893 ;
  assign n55740 = n55739 ^ n35306 ^ 1'b0 ;
  assign n55741 = n55740 ^ n29668 ^ n9778 ;
  assign n55742 = n12077 & ~n32485 ;
  assign n55743 = ~n7641 & n55742 ;
  assign n55744 = n55743 ^ n2597 ^ 1'b0 ;
  assign n55745 = ( ~n25791 & n52375 ) | ( ~n25791 & n55744 ) | ( n52375 & n55744 ) ;
  assign n55746 = n39870 ^ n12259 ^ n10349 ;
  assign n55747 = n11264 | n54672 ;
  assign n55748 = ~n10276 & n45243 ;
  assign n55749 = n19240 ^ n18292 ^ 1'b0 ;
  assign n55750 = ~n7335 & n55749 ;
  assign n55751 = n3060 | n42077 ;
  assign n55752 = n31139 & n55751 ;
  assign n55753 = n11531 ^ n6722 ^ 1'b0 ;
  assign n55754 = n42820 ^ n723 ^ 1'b0 ;
  assign n55755 = n46107 ^ n22859 ^ 1'b0 ;
  assign n55756 = n26206 ^ n7796 ^ 1'b0 ;
  assign n55757 = ( n31929 & ~n35558 ) | ( n31929 & n37113 ) | ( ~n35558 & n37113 ) ;
  assign n55758 = n44362 ^ n34371 ^ 1'b0 ;
  assign n55759 = ~n30356 & n55758 ;
  assign n55760 = n20733 ^ n13258 ^ 1'b0 ;
  assign n55761 = n12155 | n55760 ;
  assign n55762 = n7551 & ~n44306 ;
  assign n55763 = n5923 & n32576 ;
  assign n55764 = ~n3478 & n55763 ;
  assign n55765 = ~n49981 & n55764 ;
  assign n55766 = n41885 ^ n15863 ^ 1'b0 ;
  assign n55767 = n5433 | n55766 ;
  assign n55768 = n55767 ^ n6265 ^ 1'b0 ;
  assign n55772 = ~n5866 & n29631 ;
  assign n55773 = n55772 ^ n29294 ^ 1'b0 ;
  assign n55769 = n12998 | n49315 ;
  assign n55770 = n55769 ^ n3901 ^ 1'b0 ;
  assign n55771 = n11059 & n55770 ;
  assign n55774 = n55773 ^ n55771 ^ 1'b0 ;
  assign n55775 = n29790 & n55774 ;
  assign n55776 = ~n40776 & n55775 ;
  assign n55777 = n19411 & n36652 ;
  assign n55778 = n55776 & n55777 ;
  assign n55779 = n37574 | n55778 ;
  assign n55780 = ( ~n797 & n36675 ) | ( ~n797 & n42114 ) | ( n36675 & n42114 ) ;
  assign n55781 = n1357 & n35836 ;
  assign n55782 = n55781 ^ n28749 ^ 1'b0 ;
  assign n55783 = n55782 ^ n23311 ^ n5725 ;
  assign n55784 = n32547 ^ n4847 ^ 1'b0 ;
  assign n55785 = n48901 & n55784 ;
  assign n55786 = n55785 ^ n3710 ^ 1'b0 ;
  assign n55787 = n34851 & n55786 ;
  assign n55788 = n27897 ^ n24523 ^ n15725 ;
  assign n55789 = ( n5442 & ~n28279 ) | ( n5442 & n55788 ) | ( ~n28279 & n55788 ) ;
  assign n55790 = n55789 ^ n5140 ^ 1'b0 ;
  assign n55791 = ~n1138 & n55790 ;
  assign n55792 = n33938 ^ n21802 ^ 1'b0 ;
  assign n55793 = n10349 & ~n55792 ;
  assign n55794 = n55793 ^ n34886 ^ 1'b0 ;
  assign n55795 = ~n3703 & n55794 ;
  assign n55796 = ( n14978 & n18688 ) | ( n14978 & ~n29703 ) | ( n18688 & ~n29703 ) ;
  assign n55797 = n14214 & ~n41451 ;
  assign n55798 = n55797 ^ n51328 ^ n16622 ;
  assign n55799 = n46114 ^ n17731 ^ n3805 ;
  assign n55800 = ( n11826 & n12325 ) | ( n11826 & ~n55799 ) | ( n12325 & ~n55799 ) ;
  assign n55801 = n8551 ^ n5762 ^ 1'b0 ;
  assign n55802 = n7218 & ~n55801 ;
  assign n55803 = n24914 & n55802 ;
  assign n55804 = n37778 ^ n4507 ^ 1'b0 ;
  assign n55805 = n55803 | n55804 ;
  assign n55806 = ~n18369 & n26172 ;
  assign n55807 = n45374 ^ n16573 ^ 1'b0 ;
  assign n55808 = n33148 & ~n55807 ;
  assign n55809 = ~n9433 & n55808 ;
  assign n55810 = n4008 & ~n24288 ;
  assign n55811 = n24985 | n43220 ;
  assign n55812 = n55810 | n55811 ;
  assign n55813 = n654 & n28255 ;
  assign n55814 = ~n16260 & n55813 ;
  assign n55815 = n6840 & ~n22029 ;
  assign n55816 = n55814 & n55815 ;
  assign n55817 = n18531 & ~n23332 ;
  assign n55818 = n50155 ^ n9914 ^ n177 ;
  assign n55819 = ( n19373 & ~n42288 ) | ( n19373 & n55818 ) | ( ~n42288 & n55818 ) ;
  assign n55820 = n50523 ^ n16695 ^ 1'b0 ;
  assign n55821 = n99 & n20262 ;
  assign n55822 = ~n13749 & n55821 ;
  assign n55823 = n7197 & ~n7214 ;
  assign n55824 = n11244 | n16948 ;
  assign n55825 = ( n4971 & n11011 ) | ( n4971 & ~n55824 ) | ( n11011 & ~n55824 ) ;
  assign n55826 = n37426 ^ n7867 ^ 1'b0 ;
  assign n55827 = ~n55825 & n55826 ;
  assign n55828 = ~n11065 & n35601 ;
  assign n55829 = ( n6350 & n45433 ) | ( n6350 & ~n55828 ) | ( n45433 & ~n55828 ) ;
  assign n55836 = n29267 ^ n23539 ^ n20819 ;
  assign n55830 = n39741 ^ n32008 ^ 1'b0 ;
  assign n55831 = n19606 & n43064 ;
  assign n55832 = ~n55830 & n55831 ;
  assign n55833 = ~n1957 & n22774 ;
  assign n55834 = ~n2217 & n55833 ;
  assign n55835 = ( n28306 & ~n55832 ) | ( n28306 & n55834 ) | ( ~n55832 & n55834 ) ;
  assign n55837 = n55836 ^ n55835 ^ n25658 ;
  assign n55838 = n45266 ^ n43529 ^ n13222 ;
  assign n55839 = n4697 ^ n1596 ^ 1'b0 ;
  assign n55840 = n40832 & n55839 ;
  assign n55841 = n15638 & n27483 ;
  assign n55842 = ~n17820 & n55841 ;
  assign n55843 = ~n25488 & n55842 ;
  assign n55844 = n30373 & ~n55843 ;
  assign n55845 = ~n55840 & n55844 ;
  assign n55846 = n10035 | n36315 ;
  assign n55847 = n55845 & ~n55846 ;
  assign n55848 = n3255 ^ n1312 ^ 1'b0 ;
  assign n55849 = n18123 & ~n20282 ;
  assign n55850 = n55849 ^ n2083 ^ 1'b0 ;
  assign n55851 = n51161 ^ n6000 ^ 1'b0 ;
  assign n55852 = ~n6001 & n48842 ;
  assign n55853 = n43592 ^ n38168 ^ n31547 ;
  assign n55854 = n17399 ^ n3760 ^ 1'b0 ;
  assign n55855 = n15886 | n51524 ;
  assign n55856 = n1818 & ~n44657 ;
  assign n55857 = n34733 ^ n30997 ^ 1'b0 ;
  assign n55858 = n11329 | n55857 ;
  assign n55859 = n55858 ^ n12263 ^ n4222 ;
  assign n55860 = n18316 & ~n55859 ;
  assign n55861 = ~n43735 & n48669 ;
  assign n55862 = n5713 & n27945 ;
  assign n55863 = n46986 ^ n6707 ^ 1'b0 ;
  assign n55864 = n55862 | n55863 ;
  assign n55865 = ( n7144 & n11961 ) | ( n7144 & ~n30702 ) | ( n11961 & ~n30702 ) ;
  assign n55866 = n45932 & n55843 ;
  assign n55867 = n30557 ^ n18283 ^ n5599 ;
  assign n55868 = ( ~n44118 & n51773 ) | ( ~n44118 & n55867 ) | ( n51773 & n55867 ) ;
  assign n55870 = ( n2160 & ~n4009 ) | ( n2160 & n34087 ) | ( ~n4009 & n34087 ) ;
  assign n55869 = ~n11603 & n17162 ;
  assign n55871 = n55870 ^ n55869 ^ 1'b0 ;
  assign n55872 = n9233 & n11864 ;
  assign n55873 = n33343 & n55872 ;
  assign n55874 = n13522 | n55873 ;
  assign n55875 = ~n18368 & n42142 ;
  assign n55876 = n55875 ^ n11908 ^ 1'b0 ;
  assign n55877 = ~n43494 & n55876 ;
  assign n55878 = n9022 & ~n48093 ;
  assign n55879 = n43219 & n55878 ;
  assign n55880 = n47696 ^ n29471 ^ 1'b0 ;
  assign n55881 = n47155 & ~n55880 ;
  assign n55882 = n3607 & ~n4227 ;
  assign n55883 = n14587 & n55882 ;
  assign n55884 = n38666 ^ n31076 ^ 1'b0 ;
  assign n55885 = n41145 ^ n16984 ^ 1'b0 ;
  assign n55886 = n55885 ^ n36251 ^ 1'b0 ;
  assign n55887 = ~n6183 & n12156 ;
  assign n55888 = n36041 ^ n25970 ^ n8414 ;
  assign n55889 = ~n55887 & n55888 ;
  assign n55890 = n19823 & ~n22376 ;
  assign n55891 = n55890 ^ n15622 ^ 1'b0 ;
  assign n55892 = n11969 ^ n6003 ^ 1'b0 ;
  assign n55893 = n55891 & n55892 ;
  assign n55894 = n16614 & ~n48311 ;
  assign n55895 = ~n1105 & n23008 ;
  assign n55896 = n9919 & ~n55895 ;
  assign n55897 = n2949 & n55896 ;
  assign n55898 = n32347 & n33580 ;
  assign n55899 = n55897 & n55898 ;
  assign n55900 = n31285 & n44874 ;
  assign n55901 = n55900 ^ n10212 ^ 1'b0 ;
  assign n55902 = n37141 ^ n228 ^ 1'b0 ;
  assign n55903 = n19894 & ~n22852 ;
  assign n55904 = ~n3830 & n8323 ;
  assign n55905 = ~n6144 & n55904 ;
  assign n55906 = ~n17360 & n55905 ;
  assign n55907 = n7468 | n10408 ;
  assign n55908 = n572 & ~n55907 ;
  assign n55909 = n25576 ^ n17254 ^ 1'b0 ;
  assign n55910 = n29148 & n55909 ;
  assign n55911 = ~n29208 & n55910 ;
  assign n55912 = n43671 ^ n13007 ^ 1'b0 ;
  assign n55913 = n20879 & ~n21975 ;
  assign n55914 = ~n55912 & n55913 ;
  assign n55915 = n3077 & ~n7949 ;
  assign n55916 = n55915 ^ n24985 ^ 1'b0 ;
  assign n55917 = ( n19551 & ~n26041 ) | ( n19551 & n27163 ) | ( ~n26041 & n27163 ) ;
  assign n55918 = n15501 | n55917 ;
  assign n55919 = n5302 | n55918 ;
  assign n55920 = n38559 & n39166 ;
  assign n55921 = ( n39922 & ~n55919 ) | ( n39922 & n55920 ) | ( ~n55919 & n55920 ) ;
  assign n55922 = n6341 & ~n26152 ;
  assign n55923 = n55922 ^ n321 ^ 1'b0 ;
  assign n55924 = ~n22805 & n55923 ;
  assign n55925 = ~n16341 & n55924 ;
  assign n55926 = ~n55921 & n55925 ;
  assign n55927 = n54003 ^ n45281 ^ 1'b0 ;
  assign n55928 = n19657 ^ n3593 ^ 1'b0 ;
  assign n55929 = n32125 & n55928 ;
  assign n55930 = ( n5428 & n11025 ) | ( n5428 & ~n55929 ) | ( n11025 & ~n55929 ) ;
  assign n55931 = ( ~n9093 & n11330 ) | ( ~n9093 & n13210 ) | ( n11330 & n13210 ) ;
  assign n55932 = ~n14307 & n49897 ;
  assign n55933 = n55932 ^ n18234 ^ 1'b0 ;
  assign n55934 = n48709 ^ n22042 ^ 1'b0 ;
  assign n55935 = n5310 & n17401 ;
  assign n55936 = n36841 ^ n11847 ^ 1'b0 ;
  assign n55937 = ~n28365 & n55936 ;
  assign n55938 = n4584 | n16785 ;
  assign n55939 = n29847 | n55938 ;
  assign n55940 = n23084 ^ n15504 ^ n11902 ;
  assign n55941 = n9781 & n53988 ;
  assign n55942 = n15958 & ~n23756 ;
  assign n55944 = n35836 & ~n37817 ;
  assign n55943 = n11323 & n46167 ;
  assign n55945 = n55944 ^ n55943 ^ 1'b0 ;
  assign n55946 = n20922 ^ n777 ^ n508 ;
  assign n55947 = n55946 ^ n16008 ^ 1'b0 ;
  assign n55948 = n24894 & ~n55947 ;
  assign n55950 = n23560 & n43148 ;
  assign n55951 = ~n43191 & n55950 ;
  assign n55949 = n4901 & ~n40511 ;
  assign n55952 = n55951 ^ n55949 ^ 1'b0 ;
  assign n55953 = n22114 ^ n8190 ^ n940 ;
  assign n55954 = n10679 & n42650 ;
  assign n55955 = n55269 | n55954 ;
  assign n55956 = n15254 ^ n3135 ^ n1853 ;
  assign n55957 = n12771 & ~n30772 ;
  assign n55958 = n5324 & ~n14409 ;
  assign n55959 = n55958 ^ n4201 ^ 1'b0 ;
  assign n55960 = n32073 ^ n26434 ^ 1'b0 ;
  assign n55961 = n33347 ^ n10875 ^ n8432 ;
  assign n55962 = n55961 ^ n30342 ^ 1'b0 ;
  assign n55963 = ~n8103 & n52235 ;
  assign n55964 = n42441 ^ n12296 ^ n11712 ;
  assign n55965 = n55964 ^ n22826 ^ 1'b0 ;
  assign n55966 = ~n245 & n9181 ;
  assign n55967 = n23900 | n50043 ;
  assign n55968 = n55966 & ~n55967 ;
  assign n55969 = ~n11406 & n12188 ;
  assign n55970 = n55969 ^ n5952 ^ 1'b0 ;
  assign n55971 = n49736 ^ n27649 ^ n12373 ;
  assign n55972 = n55971 ^ n5822 ^ 1'b0 ;
  assign n55973 = n55972 ^ n51178 ^ 1'b0 ;
  assign n55974 = ( ~n3802 & n13663 ) | ( ~n3802 & n33652 ) | ( n13663 & n33652 ) ;
  assign n55975 = n2825 & ~n23109 ;
  assign n55976 = ( n840 & n32583 ) | ( n840 & n55975 ) | ( n32583 & n55975 ) ;
  assign n55977 = n41097 ^ n31244 ^ n9974 ;
  assign n55978 = n55977 ^ n16810 ^ 1'b0 ;
  assign n55979 = n7358 & n55978 ;
  assign n55980 = ~n2684 & n55979 ;
  assign n55981 = n36168 & ~n40595 ;
  assign n55982 = ~n55980 & n55981 ;
  assign n55983 = n9701 | n38024 ;
  assign n55984 = n3997 & n17452 ;
  assign n55985 = n55984 ^ n1435 ^ 1'b0 ;
  assign n55986 = n55985 ^ n30913 ^ 1'b0 ;
  assign n55987 = n6653 | n20453 ;
  assign n55988 = n51928 | n55987 ;
  assign n55989 = ~n10245 & n33647 ;
  assign n55990 = ~n46585 & n55989 ;
  assign n55991 = ~n954 & n5797 ;
  assign n55992 = n55991 ^ n3810 ^ 1'b0 ;
  assign n55993 = n55992 ^ n2352 ^ 1'b0 ;
  assign n55994 = ( n8413 & ~n13900 ) | ( n8413 & n16288 ) | ( ~n13900 & n16288 ) ;
  assign n55995 = n33098 | n55994 ;
  assign n55996 = n55993 | n55995 ;
  assign n55997 = n9707 | n12961 ;
  assign n55998 = n14786 & n55997 ;
  assign n55999 = n19364 & n55998 ;
  assign n56000 = n55999 ^ n14169 ^ 1'b0 ;
  assign n56001 = ~n30233 & n56000 ;
  assign n56002 = n56001 ^ n36243 ^ 1'b0 ;
  assign n56003 = ~n41808 & n56002 ;
  assign n56004 = n31529 ^ n4577 ^ 1'b0 ;
  assign n56005 = n24061 | n56004 ;
  assign n56006 = n56005 ^ n36502 ^ n19703 ;
  assign n56007 = n37122 ^ n35210 ^ n5197 ;
  assign n56008 = n26936 ^ n19592 ^ 1'b0 ;
  assign n56009 = n6771 & ~n12075 ;
  assign n56010 = n30700 & n56009 ;
  assign n56011 = n56008 & n56010 ;
  assign n56012 = n47373 | n56011 ;
  assign n56013 = n24801 & ~n55342 ;
  assign n56016 = n8672 & ~n14188 ;
  assign n56014 = n30127 & n40718 ;
  assign n56015 = n56014 ^ n2282 ^ 1'b0 ;
  assign n56017 = n56016 ^ n56015 ^ 1'b0 ;
  assign n56018 = n3890 & n20747 ;
  assign n56019 = n5740 & n56018 ;
  assign n56020 = n41026 | n56019 ;
  assign n56021 = n620 & ~n56020 ;
  assign n56022 = n2044 & n47769 ;
  assign n56023 = n27100 & n56022 ;
  assign n56024 = ( n1929 & n31591 ) | ( n1929 & ~n52399 ) | ( n31591 & ~n52399 ) ;
  assign n56025 = ~n13964 & n30122 ;
  assign n56026 = n2841 & ~n21029 ;
  assign n56027 = n56026 ^ n46950 ^ 1'b0 ;
  assign n56028 = n2528 & ~n56027 ;
  assign n56029 = ( ~n18443 & n56025 ) | ( ~n18443 & n56028 ) | ( n56025 & n56028 ) ;
  assign n56030 = n18955 ^ n15744 ^ n12631 ;
  assign n56031 = ~n10813 & n56030 ;
  assign n56032 = n28440 | n42752 ;
  assign n56033 = n960 | n52582 ;
  assign n56034 = n8239 ^ n6937 ^ 1'b0 ;
  assign n56035 = n47880 & n56034 ;
  assign n56036 = n15779 & ~n39606 ;
  assign n56037 = n24462 ^ n5744 ^ 1'b0 ;
  assign n56038 = n20836 & n35611 ;
  assign n56039 = n23203 ^ n9194 ^ n5500 ;
  assign n56040 = n3122 | n7916 ;
  assign n56041 = n17487 | n56040 ;
  assign n56042 = n15136 & ~n56041 ;
  assign n56043 = n27094 | n44177 ;
  assign n56044 = n56042 & ~n56043 ;
  assign n56045 = ( n8504 & n15780 ) | ( n8504 & ~n56044 ) | ( n15780 & ~n56044 ) ;
  assign n56046 = n5563 & ~n12863 ;
  assign n56047 = n52854 ^ n40887 ^ 1'b0 ;
  assign n56048 = ~n15091 & n56047 ;
  assign n56049 = n1574 & n35349 ;
  assign n56050 = n56049 ^ n21038 ^ 1'b0 ;
  assign n56051 = n32306 ^ n20237 ^ n5130 ;
  assign n56052 = ( n14766 & n33247 ) | ( n14766 & ~n42023 ) | ( n33247 & ~n42023 ) ;
  assign n56053 = n9764 & n56052 ;
  assign n56054 = ( ~n29317 & n33472 ) | ( ~n29317 & n44523 ) | ( n33472 & n44523 ) ;
  assign n56055 = n42064 ^ n38999 ^ 1'b0 ;
  assign n56056 = n50281 | n56055 ;
  assign n56057 = n12475 | n45537 ;
  assign n56058 = n56057 ^ n22674 ^ 1'b0 ;
  assign n56059 = n23578 ^ n18619 ^ 1'b0 ;
  assign n56062 = n10868 | n15477 ;
  assign n56063 = n56062 ^ n48123 ^ 1'b0 ;
  assign n56060 = ~n7273 & n35612 ;
  assign n56061 = n56060 ^ n23401 ^ 1'b0 ;
  assign n56064 = n56063 ^ n56061 ^ n1017 ;
  assign n56065 = ~n25169 & n28427 ;
  assign n56066 = n15083 ^ n11934 ^ n2571 ;
  assign n56067 = n34783 ^ n23761 ^ n11925 ;
  assign n56068 = ( ~n19645 & n43436 ) | ( ~n19645 & n56067 ) | ( n43436 & n56067 ) ;
  assign n56069 = ( n56065 & ~n56066 ) | ( n56065 & n56068 ) | ( ~n56066 & n56068 ) ;
  assign n56070 = n4201 & ~n46684 ;
  assign n56071 = ( ~n2268 & n7864 ) | ( ~n2268 & n41534 ) | ( n7864 & n41534 ) ;
  assign n56072 = n56070 & ~n56071 ;
  assign n56073 = n28594 & ~n51140 ;
  assign n56074 = n1378 & n56073 ;
  assign n56075 = n11015 ^ n6230 ^ 1'b0 ;
  assign n56076 = n11873 & ~n27972 ;
  assign n56077 = n56076 ^ n21132 ^ 1'b0 ;
  assign n56078 = n22622 | n25542 ;
  assign n56079 = n56078 ^ n19319 ^ 1'b0 ;
  assign n56080 = ~n34735 & n43730 ;
  assign n56081 = ~n56079 & n56080 ;
  assign n56082 = n21264 ^ n1896 ^ 1'b0 ;
  assign n56084 = n25983 & n34371 ;
  assign n56083 = n26257 | n39083 ;
  assign n56085 = n56084 ^ n56083 ^ 1'b0 ;
  assign n56086 = n56085 ^ n40788 ^ 1'b0 ;
  assign n56087 = n18720 & ~n50933 ;
  assign n56088 = ~n8827 & n48193 ;
  assign n56089 = n8850 | n31650 ;
  assign n56090 = n299 & n23720 ;
  assign n56091 = n43416 & ~n56090 ;
  assign n56092 = n34387 ^ n25766 ^ 1'b0 ;
  assign n56093 = n4638 & n56092 ;
  assign n56094 = ~n8893 & n56093 ;
  assign n56095 = n56094 ^ n40247 ^ 1'b0 ;
  assign n56096 = n40729 ^ n19774 ^ 1'b0 ;
  assign n56097 = n7773 & ~n56096 ;
  assign n56098 = n56097 ^ n35609 ^ 1'b0 ;
  assign n56099 = ~n4848 & n56098 ;
  assign n56100 = ( n11241 & n30113 ) | ( n11241 & ~n48066 ) | ( n30113 & ~n48066 ) ;
  assign n56101 = n9103 ^ n3214 ^ 1'b0 ;
  assign n56102 = ~n18712 & n56101 ;
  assign n56103 = n56102 ^ n6374 ^ n2511 ;
  assign n56104 = n52543 ^ n47948 ^ 1'b0 ;
  assign y0 = x6 ;
  assign y1 = n13 ;
  assign y2 = n15 ;
  assign y3 = ~1'b0 ;
  assign y4 = ~1'b0 ;
  assign y5 = ~1'b0 ;
  assign y6 = n22 ;
  assign y7 = x3 ;
  assign y8 = n23 ;
  assign y9 = ~1'b0 ;
  assign y10 = ~n33 ;
  assign y11 = ~n38 ;
  assign y12 = ~n39 ;
  assign y13 = ~n42 ;
  assign y14 = ~1'b0 ;
  assign y15 = ~n44 ;
  assign y16 = n46 ;
  assign y17 = ~n48 ;
  assign y18 = ~n51 ;
  assign y19 = n53 ;
  assign y20 = n54 ;
  assign y21 = x10 ;
  assign y22 = ~n55 ;
  assign y23 = ~n61 ;
  assign y24 = ~n62 ;
  assign y25 = ~n63 ;
  assign y26 = n68 ;
  assign y27 = ~1'b0 ;
  assign y28 = ~n74 ;
  assign y29 = ~n75 ;
  assign y30 = ~n78 ;
  assign y31 = n79 ;
  assign y32 = n41 ;
  assign y33 = ~1'b0 ;
  assign y34 = n82 ;
  assign y35 = 1'b0 ;
  assign y36 = ~n63 ;
  assign y37 = x3 ;
  assign y38 = n85 ;
  assign y39 = n89 ;
  assign y40 = n91 ;
  assign y41 = ~n97 ;
  assign y42 = ~n102 ;
  assign y43 = ~1'b0 ;
  assign y44 = n41 ;
  assign y45 = n105 ;
  assign y46 = n37 ;
  assign y47 = n108 ;
  assign y48 = ~1'b0 ;
  assign y49 = n109 ;
  assign y50 = ~n112 ;
  assign y51 = ~1'b0 ;
  assign y52 = ~n117 ;
  assign y53 = n118 ;
  assign y54 = n119 ;
  assign y55 = ~1'b0 ;
  assign y56 = ~n125 ;
  assign y57 = n130 ;
  assign y58 = ~1'b0 ;
  assign y59 = ~1'b0 ;
  assign y60 = n132 ;
  assign y61 = ~n135 ;
  assign y62 = 1'b0 ;
  assign y63 = ~n98 ;
  assign y64 = n136 ;
  assign y65 = ~n139 ;
  assign y66 = ~n142 ;
  assign y67 = ~n147 ;
  assign y68 = ~1'b0 ;
  assign y69 = ~n151 ;
  assign y70 = ~1'b0 ;
  assign y71 = n152 ;
  assign y72 = ~1'b0 ;
  assign y73 = ~n153 ;
  assign y74 = ~1'b0 ;
  assign y75 = ~1'b0 ;
  assign y76 = ~n156 ;
  assign y77 = ~n159 ;
  assign y78 = n165 ;
  assign y79 = n172 ;
  assign y80 = n174 ;
  assign y81 = ~n176 ;
  assign y82 = n177 ;
  assign y83 = ~n40 ;
  assign y84 = ~n179 ;
  assign y85 = ~n183 ;
  assign y86 = ~n185 ;
  assign y87 = ~n190 ;
  assign y88 = ~1'b0 ;
  assign y89 = n192 ;
  assign y90 = 1'b0 ;
  assign y91 = n197 ;
  assign y92 = ~n139 ;
  assign y93 = ~n205 ;
  assign y94 = ~n208 ;
  assign y95 = ~n210 ;
  assign y96 = ~1'b0 ;
  assign y97 = n213 ;
  assign y98 = ~1'b0 ;
  assign y99 = ~1'b0 ;
  assign y100 = ~n214 ;
  assign y101 = ~n141 ;
  assign y102 = ~n217 ;
  assign y103 = ~n218 ;
  assign y104 = ~n220 ;
  assign y105 = ~n222 ;
  assign y106 = ~1'b0 ;
  assign y107 = ~n205 ;
  assign y108 = n224 ;
  assign y109 = ~n225 ;
  assign y110 = n230 ;
  assign y111 = ~n238 ;
  assign y112 = n241 ;
  assign y113 = ~n242 ;
  assign y114 = ~n243 ;
  assign y115 = n250 ;
  assign y116 = ~n252 ;
  assign y117 = ~1'b0 ;
  assign y118 = n254 ;
  assign y119 = ~n255 ;
  assign y120 = n259 ;
  assign y121 = ~n260 ;
  assign y122 = ~n265 ;
  assign y123 = ~1'b0 ;
  assign y124 = ~n269 ;
  assign y125 = ~n272 ;
  assign y126 = ~1'b0 ;
  assign y127 = ~1'b0 ;
  assign y128 = n281 ;
  assign y129 = n283 ;
  assign y130 = n289 ;
  assign y131 = ~1'b0 ;
  assign y132 = n291 ;
  assign y133 = ~n293 ;
  assign y134 = n305 ;
  assign y135 = 1'b0 ;
  assign y136 = n283 ;
  assign y137 = n306 ;
  assign y138 = ~1'b0 ;
  assign y139 = n309 ;
  assign y140 = n312 ;
  assign y141 = n317 ;
  assign y142 = ~n319 ;
  assign y143 = ~1'b0 ;
  assign y144 = ~1'b0 ;
  assign y145 = ~n321 ;
  assign y146 = ~n322 ;
  assign y147 = ~1'b0 ;
  assign y148 = ~1'b0 ;
  assign y149 = x10 ;
  assign y150 = n329 ;
  assign y151 = ~1'b0 ;
  assign y152 = ~n332 ;
  assign y153 = n338 ;
  assign y154 = n341 ;
  assign y155 = ~n345 ;
  assign y156 = n353 ;
  assign y157 = ~1'b0 ;
  assign y158 = ~1'b0 ;
  assign y159 = ~n355 ;
  assign y160 = n358 ;
  assign y161 = ~n373 ;
  assign y162 = ~n374 ;
  assign y163 = ~n379 ;
  assign y164 = ~1'b0 ;
  assign y165 = n386 ;
  assign y166 = n388 ;
  assign y167 = n390 ;
  assign y168 = ~n392 ;
  assign y169 = n394 ;
  assign y170 = ~1'b0 ;
  assign y171 = ~n401 ;
  assign y172 = n403 ;
  assign y173 = ~1'b0 ;
  assign y174 = n406 ;
  assign y175 = n409 ;
  assign y176 = n415 ;
  assign y177 = ~n416 ;
  assign y178 = n417 ;
  assign y179 = ~n421 ;
  assign y180 = ~n423 ;
  assign y181 = n424 ;
  assign y182 = n428 ;
  assign y183 = n37 ;
  assign y184 = n431 ;
  assign y185 = n435 ;
  assign y186 = n436 ;
  assign y187 = 1'b0 ;
  assign y188 = ~n437 ;
  assign y189 = n438 ;
  assign y190 = ~n439 ;
  assign y191 = ~n446 ;
  assign y192 = n447 ;
  assign y193 = ~1'b0 ;
  assign y194 = n452 ;
  assign y195 = ~n453 ;
  assign y196 = n459 ;
  assign y197 = ~1'b0 ;
  assign y198 = n463 ;
  assign y199 = 1'b0 ;
  assign y200 = ~1'b0 ;
  assign y201 = ~1'b0 ;
  assign y202 = n464 ;
  assign y203 = ~n466 ;
  assign y204 = n467 ;
  assign y205 = n469 ;
  assign y206 = ~1'b0 ;
  assign y207 = n477 ;
  assign y208 = ~n478 ;
  assign y209 = ~n481 ;
  assign y210 = ~1'b0 ;
  assign y211 = ~1'b0 ;
  assign y212 = ~n484 ;
  assign y213 = ~n485 ;
  assign y214 = ~n494 ;
  assign y215 = n498 ;
  assign y216 = ~n499 ;
  assign y217 = ~1'b0 ;
  assign y218 = ~n500 ;
  assign y219 = ~n502 ;
  assign y220 = ~1'b0 ;
  assign y221 = ~n513 ;
  assign y222 = ~1'b0 ;
  assign y223 = ~1'b0 ;
  assign y224 = ~n515 ;
  assign y225 = n519 ;
  assign y226 = ~n44 ;
  assign y227 = ~1'b0 ;
  assign y228 = ~n523 ;
  assign y229 = ~1'b0 ;
  assign y230 = ~n529 ;
  assign y231 = n530 ;
  assign y232 = ~n221 ;
  assign y233 = n532 ;
  assign y234 = ~1'b0 ;
  assign y235 = 1'b0 ;
  assign y236 = n533 ;
  assign y237 = ~1'b0 ;
  assign y238 = ~n538 ;
  assign y239 = ~1'b0 ;
  assign y240 = ~n542 ;
  assign y241 = n544 ;
  assign y242 = n545 ;
  assign y243 = ~n547 ;
  assign y244 = ~n553 ;
  assign y245 = n554 ;
  assign y246 = ~n556 ;
  assign y247 = ~1'b0 ;
  assign y248 = ~1'b0 ;
  assign y249 = ~n557 ;
  assign y250 = ~1'b0 ;
  assign y251 = n560 ;
  assign y252 = ~n561 ;
  assign y253 = n563 ;
  assign y254 = ~n569 ;
  assign y255 = n574 ;
  assign y256 = ~1'b0 ;
  assign y257 = n578 ;
  assign y258 = ~1'b0 ;
  assign y259 = n580 ;
  assign y260 = ~n587 ;
  assign y261 = ~n588 ;
  assign y262 = n590 ;
  assign y263 = ~n593 ;
  assign y264 = ~1'b0 ;
  assign y265 = n594 ;
  assign y266 = ~n597 ;
  assign y267 = ~n601 ;
  assign y268 = ~1'b0 ;
  assign y269 = ~1'b0 ;
  assign y270 = ~n604 ;
  assign y271 = ~1'b0 ;
  assign y272 = n605 ;
  assign y273 = ~n608 ;
  assign y274 = ~n611 ;
  assign y275 = ~1'b0 ;
  assign y276 = n612 ;
  assign y277 = ~n617 ;
  assign y278 = ~n627 ;
  assign y279 = ~n628 ;
  assign y280 = n629 ;
  assign y281 = n633 ;
  assign y282 = ~n636 ;
  assign y283 = ~n640 ;
  assign y284 = ~n401 ;
  assign y285 = ~n641 ;
  assign y286 = ~n645 ;
  assign y287 = n647 ;
  assign y288 = n650 ;
  assign y289 = n656 ;
  assign y290 = n661 ;
  assign y291 = n666 ;
  assign y292 = ~1'b0 ;
  assign y293 = ~1'b0 ;
  assign y294 = ~1'b0 ;
  assign y295 = ~n668 ;
  assign y296 = ~1'b0 ;
  assign y297 = ~n670 ;
  assign y298 = ~n685 ;
  assign y299 = n688 ;
  assign y300 = ~1'b0 ;
  assign y301 = n690 ;
  assign y302 = ~n691 ;
  assign y303 = ~1'b0 ;
  assign y304 = ~n692 ;
  assign y305 = n697 ;
  assign y306 = ~n698 ;
  assign y307 = n702 ;
  assign y308 = ~1'b0 ;
  assign y309 = ~n706 ;
  assign y310 = n708 ;
  assign y311 = ~n710 ;
  assign y312 = ~1'b0 ;
  assign y313 = ~1'b0 ;
  assign y314 = 1'b0 ;
  assign y315 = ~1'b0 ;
  assign y316 = ~n714 ;
  assign y317 = ~1'b0 ;
  assign y318 = ~n719 ;
  assign y319 = ~n720 ;
  assign y320 = ~1'b0 ;
  assign y321 = ~n726 ;
  assign y322 = n729 ;
  assign y323 = ~n730 ;
  assign y324 = ~n733 ;
  assign y325 = n735 ;
  assign y326 = ~n736 ;
  assign y327 = ~n739 ;
  assign y328 = ~n740 ;
  assign y329 = ~1'b0 ;
  assign y330 = n742 ;
  assign y331 = ~1'b0 ;
  assign y332 = ~1'b0 ;
  assign y333 = ~n749 ;
  assign y334 = n750 ;
  assign y335 = ~1'b0 ;
  assign y336 = ~1'b0 ;
  assign y337 = ~n752 ;
  assign y338 = ~n755 ;
  assign y339 = ~n756 ;
  assign y340 = ~1'b0 ;
  assign y341 = n761 ;
  assign y342 = n766 ;
  assign y343 = ~n769 ;
  assign y344 = n771 ;
  assign y345 = ~1'b0 ;
  assign y346 = ~n776 ;
  assign y347 = n777 ;
  assign y348 = ~1'b0 ;
  assign y349 = n780 ;
  assign y350 = ~n787 ;
  assign y351 = n794 ;
  assign y352 = n800 ;
  assign y353 = ~1'b0 ;
  assign y354 = ~1'b0 ;
  assign y355 = ~n802 ;
  assign y356 = n803 ;
  assign y357 = ~n804 ;
  assign y358 = n808 ;
  assign y359 = ~1'b0 ;
  assign y360 = ~n811 ;
  assign y361 = ~1'b0 ;
  assign y362 = n814 ;
  assign y363 = ~n817 ;
  assign y364 = ~n819 ;
  assign y365 = ~1'b0 ;
  assign y366 = ~n824 ;
  assign y367 = n836 ;
  assign y368 = ~1'b0 ;
  assign y369 = ~n837 ;
  assign y370 = ~n841 ;
  assign y371 = ~n844 ;
  assign y372 = n845 ;
  assign y373 = n846 ;
  assign y374 = ~n852 ;
  assign y375 = n854 ;
  assign y376 = n860 ;
  assign y377 = n861 ;
  assign y378 = n863 ;
  assign y379 = ~n866 ;
  assign y380 = ~n868 ;
  assign y381 = ~n871 ;
  assign y382 = ~n875 ;
  assign y383 = n563 ;
  assign y384 = ~1'b0 ;
  assign y385 = n877 ;
  assign y386 = ~n879 ;
  assign y387 = n881 ;
  assign y388 = ~1'b0 ;
  assign y389 = ~n884 ;
  assign y390 = n889 ;
  assign y391 = ~1'b0 ;
  assign y392 = ~n890 ;
  assign y393 = n891 ;
  assign y394 = ~n900 ;
  assign y395 = ~1'b0 ;
  assign y396 = ~n902 ;
  assign y397 = n903 ;
  assign y398 = ~n905 ;
  assign y399 = ~n906 ;
  assign y400 = n909 ;
  assign y401 = ~n915 ;
  assign y402 = ~n921 ;
  assign y403 = ~n744 ;
  assign y404 = n922 ;
  assign y405 = ~1'b0 ;
  assign y406 = n925 ;
  assign y407 = ~1'b0 ;
  assign y408 = ~n926 ;
  assign y409 = n929 ;
  assign y410 = n931 ;
  assign y411 = ~n934 ;
  assign y412 = ~n938 ;
  assign y413 = ~1'b0 ;
  assign y414 = ~1'b0 ;
  assign y415 = ~1'b0 ;
  assign y416 = ~n944 ;
  assign y417 = n945 ;
  assign y418 = ~n946 ;
  assign y419 = n947 ;
  assign y420 = ~1'b0 ;
  assign y421 = ~n949 ;
  assign y422 = ~n957 ;
  assign y423 = n958 ;
  assign y424 = n959 ;
  assign y425 = ~1'b0 ;
  assign y426 = n963 ;
  assign y427 = n966 ;
  assign y428 = ~1'b0 ;
  assign y429 = ~1'b0 ;
  assign y430 = ~1'b0 ;
  assign y431 = ~n968 ;
  assign y432 = ~1'b0 ;
  assign y433 = ~n969 ;
  assign y434 = ~1'b0 ;
  assign y435 = n973 ;
  assign y436 = n974 ;
  assign y437 = n975 ;
  assign y438 = ~1'b0 ;
  assign y439 = ~n976 ;
  assign y440 = ~n230 ;
  assign y441 = n985 ;
  assign y442 = ~n990 ;
  assign y443 = n991 ;
  assign y444 = n993 ;
  assign y445 = ~1'b0 ;
  assign y446 = n994 ;
  assign y447 = ~n996 ;
  assign y448 = n997 ;
  assign y449 = n998 ;
  assign y450 = n1003 ;
  assign y451 = n1004 ;
  assign y452 = ~n1009 ;
  assign y453 = n1015 ;
  assign y454 = ~n1018 ;
  assign y455 = ~n1023 ;
  assign y456 = ~n1024 ;
  assign y457 = n1025 ;
  assign y458 = n1028 ;
  assign y459 = n1029 ;
  assign y460 = n1030 ;
  assign y461 = ~1'b0 ;
  assign y462 = n1032 ;
  assign y463 = ~n1033 ;
  assign y464 = n1037 ;
  assign y465 = n1046 ;
  assign y466 = ~n1048 ;
  assign y467 = ~n1049 ;
  assign y468 = ~n1050 ;
  assign y469 = n1051 ;
  assign y470 = ~1'b0 ;
  assign y471 = ~n1052 ;
  assign y472 = ~1'b0 ;
  assign y473 = ~n1060 ;
  assign y474 = n1062 ;
  assign y475 = ~n1064 ;
  assign y476 = ~1'b0 ;
  assign y477 = ~n1068 ;
  assign y478 = n1071 ;
  assign y479 = ~n101 ;
  assign y480 = n1072 ;
  assign y481 = 1'b0 ;
  assign y482 = ~n1079 ;
  assign y483 = n1083 ;
  assign y484 = ~n1084 ;
  assign y485 = n1087 ;
  assign y486 = ~1'b0 ;
  assign y487 = n1089 ;
  assign y488 = ~n1090 ;
  assign y489 = ~n1093 ;
  assign y490 = ~1'b0 ;
  assign y491 = n1097 ;
  assign y492 = ~n1104 ;
  assign y493 = ~n1105 ;
  assign y494 = n1107 ;
  assign y495 = n1108 ;
  assign y496 = ~n1115 ;
  assign y497 = ~1'b0 ;
  assign y498 = ~n1116 ;
  assign y499 = n1120 ;
  assign y500 = ~n1122 ;
  assign y501 = ~n1127 ;
  assign y502 = n1131 ;
  assign y503 = ~n809 ;
  assign y504 = ~n1135 ;
  assign y505 = ~n1138 ;
  assign y506 = ~n1142 ;
  assign y507 = ~1'b0 ;
  assign y508 = n1145 ;
  assign y509 = n1147 ;
  assign y510 = n1149 ;
  assign y511 = ~n1150 ;
  assign y512 = ~1'b0 ;
  assign y513 = n1153 ;
  assign y514 = n1156 ;
  assign y515 = n1153 ;
  assign y516 = ~n1162 ;
  assign y517 = ~n1164 ;
  assign y518 = ~1'b0 ;
  assign y519 = n1170 ;
  assign y520 = ~n1171 ;
  assign y521 = ~n1173 ;
  assign y522 = 1'b0 ;
  assign y523 = ~n1181 ;
  assign y524 = ~1'b0 ;
  assign y525 = ~1'b0 ;
  assign y526 = ~1'b0 ;
  assign y527 = n1182 ;
  assign y528 = ~n1183 ;
  assign y529 = n1186 ;
  assign y530 = ~1'b0 ;
  assign y531 = n1188 ;
  assign y532 = ~n1193 ;
  assign y533 = ~n1198 ;
  assign y534 = n1202 ;
  assign y535 = n866 ;
  assign y536 = 1'b0 ;
  assign y537 = n1204 ;
  assign y538 = n1209 ;
  assign y539 = n1210 ;
  assign y540 = ~n957 ;
  assign y541 = ~n1223 ;
  assign y542 = 1'b0 ;
  assign y543 = ~1'b0 ;
  assign y544 = n711 ;
  assign y545 = n1226 ;
  assign y546 = n1230 ;
  assign y547 = ~1'b0 ;
  assign y548 = ~n1232 ;
  assign y549 = ~n1233 ;
  assign y550 = ~n1235 ;
  assign y551 = ~n1238 ;
  assign y552 = n1244 ;
  assign y553 = n1245 ;
  assign y554 = ~n1251 ;
  assign y555 = ~1'b0 ;
  assign y556 = ~n1255 ;
  assign y557 = n1258 ;
  assign y558 = n1261 ;
  assign y559 = n1262 ;
  assign y560 = n1270 ;
  assign y561 = n1277 ;
  assign y562 = ~n1279 ;
  assign y563 = ~n1285 ;
  assign y564 = ~1'b0 ;
  assign y565 = n1293 ;
  assign y566 = n1302 ;
  assign y567 = n1307 ;
  assign y568 = n1308 ;
  assign y569 = n1309 ;
  assign y570 = ~1'b0 ;
  assign y571 = ~n1314 ;
  assign y572 = n1316 ;
  assign y573 = ~n1317 ;
  assign y574 = ~n1322 ;
  assign y575 = ~n1327 ;
  assign y576 = ~n1328 ;
  assign y577 = ~1'b0 ;
  assign y578 = ~n1330 ;
  assign y579 = ~n1332 ;
  assign y580 = n1336 ;
  assign y581 = ~n1337 ;
  assign y582 = ~n1339 ;
  assign y583 = n1341 ;
  assign y584 = n1343 ;
  assign y585 = n1346 ;
  assign y586 = n115 ;
  assign y587 = ~1'b0 ;
  assign y588 = ~1'b0 ;
  assign y589 = n1355 ;
  assign y590 = ~n1363 ;
  assign y591 = ~n1365 ;
  assign y592 = n1368 ;
  assign y593 = ~1'b0 ;
  assign y594 = ~n1371 ;
  assign y595 = n1382 ;
  assign y596 = n1383 ;
  assign y597 = ~n1391 ;
  assign y598 = ~1'b0 ;
  assign y599 = ~n1397 ;
  assign y600 = ~1'b0 ;
  assign y601 = n1400 ;
  assign y602 = n1401 ;
  assign y603 = ~n1402 ;
  assign y604 = ~n1403 ;
  assign y605 = n1175 ;
  assign y606 = n1406 ;
  assign y607 = ~1'b0 ;
  assign y608 = ~1'b0 ;
  assign y609 = 1'b0 ;
  assign y610 = ~n1414 ;
  assign y611 = ~n1416 ;
  assign y612 = n1418 ;
  assign y613 = ~1'b0 ;
  assign y614 = ~1'b0 ;
  assign y615 = n963 ;
  assign y616 = ~n1421 ;
  assign y617 = ~1'b0 ;
  assign y618 = n523 ;
  assign y619 = n1210 ;
  assign y620 = ~n884 ;
  assign y621 = 1'b0 ;
  assign y622 = ~n1423 ;
  assign y623 = ~n1425 ;
  assign y624 = n1426 ;
  assign y625 = n1431 ;
  assign y626 = ~n1435 ;
  assign y627 = ~n1437 ;
  assign y628 = ~1'b0 ;
  assign y629 = ~1'b0 ;
  assign y630 = n1443 ;
  assign y631 = n1455 ;
  assign y632 = ~1'b0 ;
  assign y633 = ~1'b0 ;
  assign y634 = n1456 ;
  assign y635 = n1457 ;
  assign y636 = ~n1462 ;
  assign y637 = ~1'b0 ;
  assign y638 = n1471 ;
  assign y639 = ~n1478 ;
  assign y640 = ~n1481 ;
  assign y641 = n1483 ;
  assign y642 = n1484 ;
  assign y643 = ~n1485 ;
  assign y644 = ~1'b0 ;
  assign y645 = ~1'b0 ;
  assign y646 = n1488 ;
  assign y647 = ~1'b0 ;
  assign y648 = ~1'b0 ;
  assign y649 = ~1'b0 ;
  assign y650 = ~1'b0 ;
  assign y651 = ~n191 ;
  assign y652 = n1489 ;
  assign y653 = n1490 ;
  assign y654 = n1496 ;
  assign y655 = ~n1503 ;
  assign y656 = ~n1505 ;
  assign y657 = n1506 ;
  assign y658 = ~n1511 ;
  assign y659 = ~n1512 ;
  assign y660 = ~n1515 ;
  assign y661 = ~n1518 ;
  assign y662 = n1520 ;
  assign y663 = n1523 ;
  assign y664 = n1167 ;
  assign y665 = ~1'b0 ;
  assign y666 = ~n1532 ;
  assign y667 = ~n1533 ;
  assign y668 = ~n1537 ;
  assign y669 = n1538 ;
  assign y670 = n1539 ;
  assign y671 = n556 ;
  assign y672 = ~n1540 ;
  assign y673 = ~1'b0 ;
  assign y674 = 1'b0 ;
  assign y675 = n1543 ;
  assign y676 = ~n1545 ;
  assign y677 = ~n1546 ;
  assign y678 = n1549 ;
  assign y679 = n1550 ;
  assign y680 = ~1'b0 ;
  assign y681 = 1'b0 ;
  assign y682 = 1'b0 ;
  assign y683 = ~1'b0 ;
  assign y684 = ~1'b0 ;
  assign y685 = n1552 ;
  assign y686 = ~n1553 ;
  assign y687 = ~n1556 ;
  assign y688 = ~n1563 ;
  assign y689 = ~1'b0 ;
  assign y690 = n1565 ;
  assign y691 = ~1'b0 ;
  assign y692 = ~1'b0 ;
  assign y693 = ~n1568 ;
  assign y694 = ~n1573 ;
  assign y695 = ~n368 ;
  assign y696 = n1574 ;
  assign y697 = n1577 ;
  assign y698 = n1578 ;
  assign y699 = ~n1581 ;
  assign y700 = ~n1583 ;
  assign y701 = ~n1585 ;
  assign y702 = ~1'b0 ;
  assign y703 = ~1'b0 ;
  assign y704 = n1586 ;
  assign y705 = ~n1589 ;
  assign y706 = ~1'b0 ;
  assign y707 = ~n1592 ;
  assign y708 = ~n1594 ;
  assign y709 = n1596 ;
  assign y710 = ~n1602 ;
  assign y711 = n32 ;
  assign y712 = ~1'b0 ;
  assign y713 = n1606 ;
  assign y714 = ~1'b0 ;
  assign y715 = ~1'b0 ;
  assign y716 = ~n1609 ;
  assign y717 = ~n1613 ;
  assign y718 = n1623 ;
  assign y719 = ~n1625 ;
  assign y720 = ~n1628 ;
  assign y721 = ~n1630 ;
  assign y722 = ~1'b0 ;
  assign y723 = ~n1634 ;
  assign y724 = n1635 ;
  assign y725 = ~n1638 ;
  assign y726 = n1641 ;
  assign y727 = ~1'b0 ;
  assign y728 = n1642 ;
  assign y729 = ~n1643 ;
  assign y730 = ~n73 ;
  assign y731 = n1645 ;
  assign y732 = n1650 ;
  assign y733 = n944 ;
  assign y734 = ~1'b0 ;
  assign y735 = ~1'b0 ;
  assign y736 = ~n1652 ;
  assign y737 = ~n1653 ;
  assign y738 = ~n1654 ;
  assign y739 = ~n1658 ;
  assign y740 = ~n1660 ;
  assign y741 = ~n1665 ;
  assign y742 = ~n1668 ;
  assign y743 = ~n1670 ;
  assign y744 = ~n1690 ;
  assign y745 = ~1'b0 ;
  assign y746 = ~n1691 ;
  assign y747 = n1694 ;
  assign y748 = ~1'b0 ;
  assign y749 = ~n78 ;
  assign y750 = n619 ;
  assign y751 = n1699 ;
  assign y752 = n1710 ;
  assign y753 = ~n1712 ;
  assign y754 = ~1'b0 ;
  assign y755 = ~n496 ;
  assign y756 = ~1'b0 ;
  assign y757 = 1'b0 ;
  assign y758 = ~1'b0 ;
  assign y759 = ~1'b0 ;
  assign y760 = ~n1716 ;
  assign y761 = ~1'b0 ;
  assign y762 = n1721 ;
  assign y763 = n1722 ;
  assign y764 = ~1'b0 ;
  assign y765 = ~1'b0 ;
  assign y766 = 1'b0 ;
  assign y767 = ~1'b0 ;
  assign y768 = ~n1105 ;
  assign y769 = n1724 ;
  assign y770 = ~1'b0 ;
  assign y771 = n1726 ;
  assign y772 = n1727 ;
  assign y773 = ~1'b0 ;
  assign y774 = n1731 ;
  assign y775 = n1734 ;
  assign y776 = ~1'b0 ;
  assign y777 = n1736 ;
  assign y778 = n1737 ;
  assign y779 = n1745 ;
  assign y780 = ~1'b0 ;
  assign y781 = n1746 ;
  assign y782 = ~n1751 ;
  assign y783 = ~1'b0 ;
  assign y784 = n1758 ;
  assign y785 = n1760 ;
  assign y786 = n1761 ;
  assign y787 = ~n1766 ;
  assign y788 = ~1'b0 ;
  assign y789 = ~n1768 ;
  assign y790 = ~n1771 ;
  assign y791 = ~n1786 ;
  assign y792 = ~1'b0 ;
  assign y793 = ~1'b0 ;
  assign y794 = ~n1787 ;
  assign y795 = n1793 ;
  assign y796 = n1803 ;
  assign y797 = n1807 ;
  assign y798 = n1808 ;
  assign y799 = n1809 ;
  assign y800 = n1810 ;
  assign y801 = n1811 ;
  assign y802 = n1812 ;
  assign y803 = ~n1818 ;
  assign y804 = n1822 ;
  assign y805 = ~n1823 ;
  assign y806 = n1824 ;
  assign y807 = n1825 ;
  assign y808 = n1826 ;
  assign y809 = ~1'b0 ;
  assign y810 = ~1'b0 ;
  assign y811 = ~1'b0 ;
  assign y812 = ~1'b0 ;
  assign y813 = ~1'b0 ;
  assign y814 = n1828 ;
  assign y815 = ~n1830 ;
  assign y816 = ~1'b0 ;
  assign y817 = ~n1838 ;
  assign y818 = ~n1840 ;
  assign y819 = ~1'b0 ;
  assign y820 = n757 ;
  assign y821 = ~n1841 ;
  assign y822 = ~1'b0 ;
  assign y823 = n1843 ;
  assign y824 = n1846 ;
  assign y825 = ~n1851 ;
  assign y826 = ~1'b0 ;
  assign y827 = n1852 ;
  assign y828 = ~1'b0 ;
  assign y829 = ~n1864 ;
  assign y830 = ~1'b0 ;
  assign y831 = ~n1866 ;
  assign y832 = ~n1868 ;
  assign y833 = n1878 ;
  assign y834 = n1881 ;
  assign y835 = n1882 ;
  assign y836 = ~1'b0 ;
  assign y837 = n1883 ;
  assign y838 = n1888 ;
  assign y839 = n1890 ;
  assign y840 = 1'b0 ;
  assign y841 = ~n1891 ;
  assign y842 = ~n1893 ;
  assign y843 = ~1'b0 ;
  assign y844 = ~n1894 ;
  assign y845 = ~1'b0 ;
  assign y846 = n1900 ;
  assign y847 = n1904 ;
  assign y848 = ~1'b0 ;
  assign y849 = ~n1905 ;
  assign y850 = ~n1913 ;
  assign y851 = n220 ;
  assign y852 = ~n1921 ;
  assign y853 = ~1'b0 ;
  assign y854 = ~n1927 ;
  assign y855 = ~n1928 ;
  assign y856 = n1201 ;
  assign y857 = ~1'b0 ;
  assign y858 = n1931 ;
  assign y859 = ~n1933 ;
  assign y860 = ~n1934 ;
  assign y861 = n1940 ;
  assign y862 = n1943 ;
  assign y863 = ~n1945 ;
  assign y864 = n1948 ;
  assign y865 = ~n1952 ;
  assign y866 = ~n1957 ;
  assign y867 = ~1'b0 ;
  assign y868 = ~1'b0 ;
  assign y869 = ~n1958 ;
  assign y870 = ~n1960 ;
  assign y871 = ~1'b0 ;
  assign y872 = n1962 ;
  assign y873 = n1967 ;
  assign y874 = ~1'b0 ;
  assign y875 = ~n1972 ;
  assign y876 = ~n1976 ;
  assign y877 = 1'b0 ;
  assign y878 = ~n1982 ;
  assign y879 = n1984 ;
  assign y880 = ~n1986 ;
  assign y881 = ~n1988 ;
  assign y882 = n1995 ;
  assign y883 = ~n1997 ;
  assign y884 = ~1'b0 ;
  assign y885 = ~1'b0 ;
  assign y886 = ~1'b0 ;
  assign y887 = ~1'b0 ;
  assign y888 = ~1'b0 ;
  assign y889 = ~n1999 ;
  assign y890 = ~n2002 ;
  assign y891 = ~n2006 ;
  assign y892 = ~n2011 ;
  assign y893 = n2015 ;
  assign y894 = ~1'b0 ;
  assign y895 = ~n2017 ;
  assign y896 = n2022 ;
  assign y897 = ~n2027 ;
  assign y898 = ~n2028 ;
  assign y899 = ~n247 ;
  assign y900 = n2029 ;
  assign y901 = n2030 ;
  assign y902 = ~1'b0 ;
  assign y903 = n2037 ;
  assign y904 = n2039 ;
  assign y905 = n2049 ;
  assign y906 = n2053 ;
  assign y907 = ~1'b0 ;
  assign y908 = n2059 ;
  assign y909 = ~1'b0 ;
  assign y910 = n2062 ;
  assign y911 = ~n2067 ;
  assign y912 = ~n2068 ;
  assign y913 = ~n2071 ;
  assign y914 = ~n2072 ;
  assign y915 = n2076 ;
  assign y916 = n2092 ;
  assign y917 = n2097 ;
  assign y918 = ~1'b0 ;
  assign y919 = ~n2100 ;
  assign y920 = ~n2102 ;
  assign y921 = ~n2111 ;
  assign y922 = n2113 ;
  assign y923 = ~1'b0 ;
  assign y924 = n2115 ;
  assign y925 = ~n2119 ;
  assign y926 = n2122 ;
  assign y927 = ~1'b0 ;
  assign y928 = ~1'b0 ;
  assign y929 = n2125 ;
  assign y930 = n2129 ;
  assign y931 = n2130 ;
  assign y932 = ~1'b0 ;
  assign y933 = ~1'b0 ;
  assign y934 = n2132 ;
  assign y935 = ~n2134 ;
  assign y936 = ~n2139 ;
  assign y937 = ~n2142 ;
  assign y938 = ~n2145 ;
  assign y939 = n2147 ;
  assign y940 = n2150 ;
  assign y941 = ~1'b0 ;
  assign y942 = ~1'b0 ;
  assign y943 = ~1'b0 ;
  assign y944 = ~1'b0 ;
  assign y945 = ~1'b0 ;
  assign y946 = n2154 ;
  assign y947 = n2158 ;
  assign y948 = ~n2161 ;
  assign y949 = n2169 ;
  assign y950 = ~n2172 ;
  assign y951 = n2174 ;
  assign y952 = ~n2177 ;
  assign y953 = ~n2178 ;
  assign y954 = n2180 ;
  assign y955 = ~n2181 ;
  assign y956 = ~n2187 ;
  assign y957 = n2188 ;
  assign y958 = ~n2194 ;
  assign y959 = n2199 ;
  assign y960 = ~n2202 ;
  assign y961 = ~1'b0 ;
  assign y962 = ~n2205 ;
  assign y963 = ~1'b0 ;
  assign y964 = n2206 ;
  assign y965 = ~n2208 ;
  assign y966 = n2211 ;
  assign y967 = ~1'b0 ;
  assign y968 = ~1'b0 ;
  assign y969 = n2213 ;
  assign y970 = ~n2223 ;
  assign y971 = ~n2225 ;
  assign y972 = n2226 ;
  assign y973 = ~n2236 ;
  assign y974 = n2241 ;
  assign y975 = ~1'b0 ;
  assign y976 = ~1'b0 ;
  assign y977 = n2247 ;
  assign y978 = ~1'b0 ;
  assign y979 = n2249 ;
  assign y980 = n2251 ;
  assign y981 = ~n2253 ;
  assign y982 = ~n2256 ;
  assign y983 = n2258 ;
  assign y984 = ~n2264 ;
  assign y985 = ~n2148 ;
  assign y986 = ~n2268 ;
  assign y987 = n2270 ;
  assign y988 = n2277 ;
  assign y989 = ~1'b0 ;
  assign y990 = ~1'b0 ;
  assign y991 = ~n2278 ;
  assign y992 = n2281 ;
  assign y993 = n451 ;
  assign y994 = ~1'b0 ;
  assign y995 = ~n2283 ;
  assign y996 = ~n2286 ;
  assign y997 = n2289 ;
  assign y998 = n2294 ;
  assign y999 = ~n2298 ;
  assign y1000 = ~1'b0 ;
  assign y1001 = ~n2300 ;
  assign y1002 = ~n2309 ;
  assign y1003 = ~n2311 ;
  assign y1004 = ~n2312 ;
  assign y1005 = ~n2317 ;
  assign y1006 = ~1'b0 ;
  assign y1007 = n2319 ;
  assign y1008 = ~1'b0 ;
  assign y1009 = ~n176 ;
  assign y1010 = ~n2322 ;
  assign y1011 = n2324 ;
  assign y1012 = n2326 ;
  assign y1013 = ~n2330 ;
  assign y1014 = n2334 ;
  assign y1015 = n2335 ;
  assign y1016 = ~1'b0 ;
  assign y1017 = ~1'b0 ;
  assign y1018 = ~1'b0 ;
  assign y1019 = n2338 ;
  assign y1020 = ~n2341 ;
  assign y1021 = ~1'b0 ;
  assign y1022 = n2346 ;
  assign y1023 = ~n1201 ;
  assign y1024 = ~1'b0 ;
  assign y1025 = n2347 ;
  assign y1026 = ~n2350 ;
  assign y1027 = n2352 ;
  assign y1028 = ~1'b0 ;
  assign y1029 = ~n2356 ;
  assign y1030 = n2357 ;
  assign y1031 = ~n1518 ;
  assign y1032 = n2360 ;
  assign y1033 = ~n2367 ;
  assign y1034 = n2370 ;
  assign y1035 = ~n2281 ;
  assign y1036 = ~1'b0 ;
  assign y1037 = ~n2372 ;
  assign y1038 = ~n2375 ;
  assign y1039 = n2377 ;
  assign y1040 = ~n2389 ;
  assign y1041 = ~1'b0 ;
  assign y1042 = ~n2390 ;
  assign y1043 = ~n2393 ;
  assign y1044 = ~n2399 ;
  assign y1045 = ~1'b0 ;
  assign y1046 = ~n2403 ;
  assign y1047 = ~1'b0 ;
  assign y1048 = n2405 ;
  assign y1049 = ~1'b0 ;
  assign y1050 = ~n2409 ;
  assign y1051 = n2411 ;
  assign y1052 = n2413 ;
  assign y1053 = n2414 ;
  assign y1054 = n2421 ;
  assign y1055 = ~1'b0 ;
  assign y1056 = ~1'b0 ;
  assign y1057 = ~n2422 ;
  assign y1058 = ~1'b0 ;
  assign y1059 = ~1'b0 ;
  assign y1060 = ~1'b0 ;
  assign y1061 = ~1'b0 ;
  assign y1062 = n2428 ;
  assign y1063 = ~n2429 ;
  assign y1064 = n2374 ;
  assign y1065 = n2433 ;
  assign y1066 = ~n2445 ;
  assign y1067 = ~n2451 ;
  assign y1068 = ~n2452 ;
  assign y1069 = ~1'b0 ;
  assign y1070 = ~n2453 ;
  assign y1071 = ~n2454 ;
  assign y1072 = n2457 ;
  assign y1073 = n2460 ;
  assign y1074 = ~n2466 ;
  assign y1075 = n2470 ;
  assign y1076 = ~n2472 ;
  assign y1077 = ~n2476 ;
  assign y1078 = n2479 ;
  assign y1079 = ~1'b0 ;
  assign y1080 = ~1'b0 ;
  assign y1081 = n2482 ;
  assign y1082 = n2483 ;
  assign y1083 = n2485 ;
  assign y1084 = ~1'b0 ;
  assign y1085 = ~1'b0 ;
  assign y1086 = n2488 ;
  assign y1087 = ~n2489 ;
  assign y1088 = n2490 ;
  assign y1089 = ~n2494 ;
  assign y1090 = ~1'b0 ;
  assign y1091 = ~n2495 ;
  assign y1092 = ~1'b0 ;
  assign y1093 = ~n1389 ;
  assign y1094 = n2497 ;
  assign y1095 = n2500 ;
  assign y1096 = ~n2503 ;
  assign y1097 = ~1'b0 ;
  assign y1098 = n2505 ;
  assign y1099 = n2508 ;
  assign y1100 = n2514 ;
  assign y1101 = ~1'b0 ;
  assign y1102 = n2516 ;
  assign y1103 = n2517 ;
  assign y1104 = ~1'b0 ;
  assign y1105 = ~n2519 ;
  assign y1106 = ~n2521 ;
  assign y1107 = n2523 ;
  assign y1108 = n2531 ;
  assign y1109 = ~n2537 ;
  assign y1110 = ~1'b0 ;
  assign y1111 = n2539 ;
  assign y1112 = n2545 ;
  assign y1113 = n2546 ;
  assign y1114 = n2552 ;
  assign y1115 = n2555 ;
  assign y1116 = ~1'b0 ;
  assign y1117 = ~n2557 ;
  assign y1118 = ~1'b0 ;
  assign y1119 = ~n2558 ;
  assign y1120 = n2560 ;
  assign y1121 = ~1'b0 ;
  assign y1122 = ~1'b0 ;
  assign y1123 = ~n2561 ;
  assign y1124 = ~n2563 ;
  assign y1125 = ~1'b0 ;
  assign y1126 = ~n2568 ;
  assign y1127 = n2575 ;
  assign y1128 = ~n2577 ;
  assign y1129 = ~n2580 ;
  assign y1130 = n2582 ;
  assign y1131 = ~1'b0 ;
  assign y1132 = ~1'b0 ;
  assign y1133 = n2586 ;
  assign y1134 = ~n2587 ;
  assign y1135 = n2589 ;
  assign y1136 = ~1'b0 ;
  assign y1137 = ~n2599 ;
  assign y1138 = ~n2602 ;
  assign y1139 = ~n2607 ;
  assign y1140 = ~n2610 ;
  assign y1141 = ~n2614 ;
  assign y1142 = ~n2616 ;
  assign y1143 = ~1'b0 ;
  assign y1144 = n2620 ;
  assign y1145 = ~n2622 ;
  assign y1146 = ~1'b0 ;
  assign y1147 = n2623 ;
  assign y1148 = n1822 ;
  assign y1149 = n2625 ;
  assign y1150 = ~1'b0 ;
  assign y1151 = ~n2627 ;
  assign y1152 = ~n2630 ;
  assign y1153 = ~1'b0 ;
  assign y1154 = ~n2646 ;
  assign y1155 = ~1'b0 ;
  assign y1156 = n2649 ;
  assign y1157 = ~n2650 ;
  assign y1158 = ~n2653 ;
  assign y1159 = ~n2657 ;
  assign y1160 = n2660 ;
  assign y1161 = n2662 ;
  assign y1162 = ~1'b0 ;
  assign y1163 = ~n2664 ;
  assign y1164 = ~1'b0 ;
  assign y1165 = n2667 ;
  assign y1166 = ~n2668 ;
  assign y1167 = ~n2672 ;
  assign y1168 = ~1'b0 ;
  assign y1169 = n2673 ;
  assign y1170 = n2678 ;
  assign y1171 = n2679 ;
  assign y1172 = n2684 ;
  assign y1173 = n2686 ;
  assign y1174 = n2689 ;
  assign y1175 = ~n2692 ;
  assign y1176 = n2702 ;
  assign y1177 = ~1'b0 ;
  assign y1178 = n2705 ;
  assign y1179 = ~n2706 ;
  assign y1180 = ~n2712 ;
  assign y1181 = n2713 ;
  assign y1182 = ~1'b0 ;
  assign y1183 = ~n2718 ;
  assign y1184 = ~n2720 ;
  assign y1185 = n2723 ;
  assign y1186 = ~1'b0 ;
  assign y1187 = ~1'b0 ;
  assign y1188 = ~n2725 ;
  assign y1189 = n2727 ;
  assign y1190 = ~1'b0 ;
  assign y1191 = ~1'b0 ;
  assign y1192 = ~1'b0 ;
  assign y1193 = n2729 ;
  assign y1194 = n2733 ;
  assign y1195 = ~1'b0 ;
  assign y1196 = ~n2735 ;
  assign y1197 = ~1'b0 ;
  assign y1198 = n2736 ;
  assign y1199 = n2738 ;
  assign y1200 = ~n2740 ;
  assign y1201 = ~1'b0 ;
  assign y1202 = ~1'b0 ;
  assign y1203 = n2741 ;
  assign y1204 = ~1'b0 ;
  assign y1205 = 1'b0 ;
  assign y1206 = ~n1545 ;
  assign y1207 = n2743 ;
  assign y1208 = ~1'b0 ;
  assign y1209 = n2746 ;
  assign y1210 = ~n2747 ;
  assign y1211 = ~1'b0 ;
  assign y1212 = ~1'b0 ;
  assign y1213 = ~1'b0 ;
  assign y1214 = n2749 ;
  assign y1215 = n526 ;
  assign y1216 = ~n33 ;
  assign y1217 = n2751 ;
  assign y1218 = ~1'b0 ;
  assign y1219 = ~x3 ;
  assign y1220 = n2757 ;
  assign y1221 = ~1'b0 ;
  assign y1222 = ~1'b0 ;
  assign y1223 = ~n2761 ;
  assign y1224 = n2763 ;
  assign y1225 = n2764 ;
  assign y1226 = n2765 ;
  assign y1227 = n1001 ;
  assign y1228 = ~n2766 ;
  assign y1229 = ~n2768 ;
  assign y1230 = ~n13 ;
  assign y1231 = ~1'b0 ;
  assign y1232 = n2772 ;
  assign y1233 = n2781 ;
  assign y1234 = ~n2783 ;
  assign y1235 = ~1'b0 ;
  assign y1236 = n2794 ;
  assign y1237 = ~n2802 ;
  assign y1238 = ~n2805 ;
  assign y1239 = ~n2807 ;
  assign y1240 = n2815 ;
  assign y1241 = n2671 ;
  assign y1242 = n2816 ;
  assign y1243 = ~1'b0 ;
  assign y1244 = ~n2817 ;
  assign y1245 = n2819 ;
  assign y1246 = n2820 ;
  assign y1247 = n2825 ;
  assign y1248 = ~1'b0 ;
  assign y1249 = n2831 ;
  assign y1250 = ~1'b0 ;
  assign y1251 = n2833 ;
  assign y1252 = ~n2836 ;
  assign y1253 = n2839 ;
  assign y1254 = ~n2840 ;
  assign y1255 = ~1'b0 ;
  assign y1256 = ~1'b0 ;
  assign y1257 = ~n2843 ;
  assign y1258 = ~1'b0 ;
  assign y1259 = ~1'b0 ;
  assign y1260 = n2845 ;
  assign y1261 = ~n2848 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = ~n2853 ;
  assign y1265 = ~1'b0 ;
  assign y1266 = ~n2855 ;
  assign y1267 = ~n2859 ;
  assign y1268 = ~n2863 ;
  assign y1269 = ~n2866 ;
  assign y1270 = ~1'b0 ;
  assign y1271 = ~1'b0 ;
  assign y1272 = n2867 ;
  assign y1273 = n903 ;
  assign y1274 = n2868 ;
  assign y1275 = ~1'b0 ;
  assign y1276 = ~1'b0 ;
  assign y1277 = ~1'b0 ;
  assign y1278 = ~n2871 ;
  assign y1279 = ~n1889 ;
  assign y1280 = ~1'b0 ;
  assign y1281 = ~n2872 ;
  assign y1282 = ~1'b0 ;
  assign y1283 = n2877 ;
  assign y1284 = ~n2879 ;
  assign y1285 = ~1'b0 ;
  assign y1286 = ~n2882 ;
  assign y1287 = ~1'b0 ;
  assign y1288 = ~1'b0 ;
  assign y1289 = ~n2885 ;
  assign y1290 = n2886 ;
  assign y1291 = n2888 ;
  assign y1292 = ~n2556 ;
  assign y1293 = ~n2892 ;
  assign y1294 = ~n2893 ;
  assign y1295 = n2895 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = n2904 ;
  assign y1298 = ~n2905 ;
  assign y1299 = n2907 ;
  assign y1300 = n2909 ;
  assign y1301 = n2911 ;
  assign y1302 = n2916 ;
  assign y1303 = n2917 ;
  assign y1304 = n2918 ;
  assign y1305 = ~n2923 ;
  assign y1306 = n2925 ;
  assign y1307 = ~1'b0 ;
  assign y1308 = ~1'b0 ;
  assign y1309 = 1'b0 ;
  assign y1310 = ~n2926 ;
  assign y1311 = ~n1322 ;
  assign y1312 = n2932 ;
  assign y1313 = ~1'b0 ;
  assign y1314 = ~n2933 ;
  assign y1315 = ~1'b0 ;
  assign y1316 = n2934 ;
  assign y1317 = ~n2935 ;
  assign y1318 = ~1'b0 ;
  assign y1319 = n2937 ;
  assign y1320 = n2939 ;
  assign y1321 = ~n2943 ;
  assign y1322 = n2952 ;
  assign y1323 = ~1'b0 ;
  assign y1324 = n2954 ;
  assign y1325 = ~1'b0 ;
  assign y1326 = ~n2955 ;
  assign y1327 = ~1'b0 ;
  assign y1328 = ~1'b0 ;
  assign y1329 = n2958 ;
  assign y1330 = n2961 ;
  assign y1331 = ~n2967 ;
  assign y1332 = n2969 ;
  assign y1333 = n2972 ;
  assign y1334 = ~n2974 ;
  assign y1335 = 1'b0 ;
  assign y1336 = n2980 ;
  assign y1337 = n260 ;
  assign y1338 = ~n2982 ;
  assign y1339 = ~1'b0 ;
  assign y1340 = n2985 ;
  assign y1341 = n2989 ;
  assign y1342 = ~n691 ;
  assign y1343 = n2990 ;
  assign y1344 = ~1'b0 ;
  assign y1345 = ~n2992 ;
  assign y1346 = ~n2994 ;
  assign y1347 = ~n2997 ;
  assign y1348 = n2999 ;
  assign y1349 = ~n3001 ;
  assign y1350 = ~1'b0 ;
  assign y1351 = n3006 ;
  assign y1352 = ~n3007 ;
  assign y1353 = ~1'b0 ;
  assign y1354 = n3008 ;
  assign y1355 = n3009 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = n962 ;
  assign y1358 = ~n3010 ;
  assign y1359 = ~1'b0 ;
  assign y1360 = ~1'b0 ;
  assign y1361 = ~n3011 ;
  assign y1362 = n682 ;
  assign y1363 = n3018 ;
  assign y1364 = n3030 ;
  assign y1365 = n3033 ;
  assign y1366 = n3035 ;
  assign y1367 = ~1'b0 ;
  assign y1368 = n3038 ;
  assign y1369 = n3039 ;
  assign y1370 = 1'b0 ;
  assign y1371 = ~1'b0 ;
  assign y1372 = n3064 ;
  assign y1373 = ~1'b0 ;
  assign y1374 = ~n3071 ;
  assign y1375 = ~n3076 ;
  assign y1376 = ~1'b0 ;
  assign y1377 = n3077 ;
  assign y1378 = n3079 ;
  assign y1379 = ~1'b0 ;
  assign y1380 = n3080 ;
  assign y1381 = ~n3087 ;
  assign y1382 = ~1'b0 ;
  assign y1383 = n3089 ;
  assign y1384 = n3096 ;
  assign y1385 = ~1'b0 ;
  assign y1386 = ~n3097 ;
  assign y1387 = ~1'b0 ;
  assign y1388 = ~n3102 ;
  assign y1389 = ~n3104 ;
  assign y1390 = n68 ;
  assign y1391 = n3106 ;
  assign y1392 = ~n3107 ;
  assign y1393 = ~1'b0 ;
  assign y1394 = ~n3109 ;
  assign y1395 = n3111 ;
  assign y1396 = n3113 ;
  assign y1397 = n3114 ;
  assign y1398 = 1'b0 ;
  assign y1399 = ~n3116 ;
  assign y1400 = n3120 ;
  assign y1401 = n3121 ;
  assign y1402 = n3122 ;
  assign y1403 = n3124 ;
  assign y1404 = n3128 ;
  assign y1405 = ~n3138 ;
  assign y1406 = ~1'b0 ;
  assign y1407 = ~1'b0 ;
  assign y1408 = ~1'b0 ;
  assign y1409 = ~n3141 ;
  assign y1410 = ~1'b0 ;
  assign y1411 = n3153 ;
  assign y1412 = ~1'b0 ;
  assign y1413 = ~n3154 ;
  assign y1414 = ~1'b0 ;
  assign y1415 = ~1'b0 ;
  assign y1416 = ~1'b0 ;
  assign y1417 = ~n2667 ;
  assign y1418 = n3155 ;
  assign y1419 = n3156 ;
  assign y1420 = n3158 ;
  assign y1421 = ~1'b0 ;
  assign y1422 = ~n3159 ;
  assign y1423 = n3163 ;
  assign y1424 = ~n3167 ;
  assign y1425 = n3174 ;
  assign y1426 = ~1'b0 ;
  assign y1427 = ~n3176 ;
  assign y1428 = ~n3179 ;
  assign y1429 = ~1'b0 ;
  assign y1430 = n3183 ;
  assign y1431 = n3185 ;
  assign y1432 = n3191 ;
  assign y1433 = n3196 ;
  assign y1434 = n3205 ;
  assign y1435 = ~n3214 ;
  assign y1436 = ~n3085 ;
  assign y1437 = n2791 ;
  assign y1438 = ~n3224 ;
  assign y1439 = ~n3235 ;
  assign y1440 = ~n3236 ;
  assign y1441 = n3237 ;
  assign y1442 = ~1'b0 ;
  assign y1443 = ~1'b0 ;
  assign y1444 = ~n3242 ;
  assign y1445 = ~1'b0 ;
  assign y1446 = n3243 ;
  assign y1447 = ~1'b0 ;
  assign y1448 = n3246 ;
  assign y1449 = ~1'b0 ;
  assign y1450 = n3248 ;
  assign y1451 = ~n3252 ;
  assign y1452 = n3254 ;
  assign y1453 = ~n3259 ;
  assign y1454 = n3268 ;
  assign y1455 = ~n3270 ;
  assign y1456 = n3275 ;
  assign y1457 = n3276 ;
  assign y1458 = n352 ;
  assign y1459 = n3279 ;
  assign y1460 = ~1'b0 ;
  assign y1461 = ~n3282 ;
  assign y1462 = ~n3284 ;
  assign y1463 = ~1'b0 ;
  assign y1464 = ~n3286 ;
  assign y1465 = ~n3292 ;
  assign y1466 = ~n3298 ;
  assign y1467 = ~n3304 ;
  assign y1468 = n3309 ;
  assign y1469 = ~n3314 ;
  assign y1470 = n3321 ;
  assign y1471 = ~n3327 ;
  assign y1472 = n3332 ;
  assign y1473 = n3333 ;
  assign y1474 = n3336 ;
  assign y1475 = ~1'b0 ;
  assign y1476 = ~n3341 ;
  assign y1477 = n3342 ;
  assign y1478 = ~n3346 ;
  assign y1479 = ~n3350 ;
  assign y1480 = n3354 ;
  assign y1481 = n1312 ;
  assign y1482 = n3355 ;
  assign y1483 = ~1'b0 ;
  assign y1484 = n3358 ;
  assign y1485 = ~n3363 ;
  assign y1486 = ~n3365 ;
  assign y1487 = n3368 ;
  assign y1488 = ~1'b0 ;
  assign y1489 = ~1'b0 ;
  assign y1490 = n3370 ;
  assign y1491 = n3376 ;
  assign y1492 = ~1'b0 ;
  assign y1493 = n709 ;
  assign y1494 = n3377 ;
  assign y1495 = n3382 ;
  assign y1496 = ~1'b0 ;
  assign y1497 = ~n3384 ;
  assign y1498 = n3385 ;
  assign y1499 = ~n3386 ;
  assign y1500 = ~n3389 ;
  assign y1501 = n3395 ;
  assign y1502 = ~n3406 ;
  assign y1503 = n3410 ;
  assign y1504 = ~n3412 ;
  assign y1505 = n3416 ;
  assign y1506 = n3418 ;
  assign y1507 = ~n3421 ;
  assign y1508 = ~1'b0 ;
  assign y1509 = ~1'b0 ;
  assign y1510 = n3423 ;
  assign y1511 = ~n3425 ;
  assign y1512 = n3433 ;
  assign y1513 = ~1'b0 ;
  assign y1514 = ~1'b0 ;
  assign y1515 = ~n3435 ;
  assign y1516 = ~1'b0 ;
  assign y1517 = ~n1201 ;
  assign y1518 = ~n3443 ;
  assign y1519 = ~n3450 ;
  assign y1520 = n3452 ;
  assign y1521 = n3454 ;
  assign y1522 = ~n3455 ;
  assign y1523 = ~n3460 ;
  assign y1524 = n3464 ;
  assign y1525 = n3467 ;
  assign y1526 = ~n3473 ;
  assign y1527 = ~n3478 ;
  assign y1528 = ~n3482 ;
  assign y1529 = ~n3483 ;
  assign y1530 = ~n3484 ;
  assign y1531 = ~n3493 ;
  assign y1532 = ~1'b0 ;
  assign y1533 = ~1'b0 ;
  assign y1534 = n2541 ;
  assign y1535 = ~n3498 ;
  assign y1536 = ~n3503 ;
  assign y1537 = n3505 ;
  assign y1538 = n3506 ;
  assign y1539 = n3514 ;
  assign y1540 = n3515 ;
  assign y1541 = ~n2449 ;
  assign y1542 = ~n3517 ;
  assign y1543 = ~1'b0 ;
  assign y1544 = ~1'b0 ;
  assign y1545 = ~1'b0 ;
  assign y1546 = ~1'b0 ;
  assign y1547 = n3518 ;
  assign y1548 = ~1'b0 ;
  assign y1549 = ~1'b0 ;
  assign y1550 = ~n3519 ;
  assign y1551 = n3530 ;
  assign y1552 = ~n411 ;
  assign y1553 = ~n3540 ;
  assign y1554 = ~n3546 ;
  assign y1555 = ~n3550 ;
  assign y1556 = n3555 ;
  assign y1557 = n3558 ;
  assign y1558 = ~n3574 ;
  assign y1559 = ~n3578 ;
  assign y1560 = ~n3581 ;
  assign y1561 = n3585 ;
  assign y1562 = ~n3588 ;
  assign y1563 = ~n3597 ;
  assign y1564 = ~n3599 ;
  assign y1565 = ~1'b0 ;
  assign y1566 = ~n3600 ;
  assign y1567 = x11 ;
  assign y1568 = n3607 ;
  assign y1569 = ~n3477 ;
  assign y1570 = ~n3608 ;
  assign y1571 = n3610 ;
  assign y1572 = n3620 ;
  assign y1573 = n3622 ;
  assign y1574 = ~1'b0 ;
  assign y1575 = n3626 ;
  assign y1576 = ~n3630 ;
  assign y1577 = n3634 ;
  assign y1578 = ~1'b0 ;
  assign y1579 = ~1'b0 ;
  assign y1580 = ~1'b0 ;
  assign y1581 = n3635 ;
  assign y1582 = ~1'b0 ;
  assign y1583 = ~1'b0 ;
  assign y1584 = ~n3636 ;
  assign y1585 = ~1'b0 ;
  assign y1586 = n3637 ;
  assign y1587 = n3639 ;
  assign y1588 = ~n3640 ;
  assign y1589 = ~n3641 ;
  assign y1590 = n3644 ;
  assign y1591 = ~1'b0 ;
  assign y1592 = n3655 ;
  assign y1593 = n3656 ;
  assign y1594 = ~1'b0 ;
  assign y1595 = ~n3662 ;
  assign y1596 = ~1'b0 ;
  assign y1597 = ~n3663 ;
  assign y1598 = ~n3669 ;
  assign y1599 = n3677 ;
  assign y1600 = ~1'b0 ;
  assign y1601 = ~1'b0 ;
  assign y1602 = ~1'b0 ;
  assign y1603 = n3680 ;
  assign y1604 = n3692 ;
  assign y1605 = ~1'b0 ;
  assign y1606 = n3693 ;
  assign y1607 = ~n3694 ;
  assign y1608 = ~n3696 ;
  assign y1609 = ~n3706 ;
  assign y1610 = ~n3707 ;
  assign y1611 = ~n3712 ;
  assign y1612 = ~n3714 ;
  assign y1613 = n3719 ;
  assign y1614 = ~n3722 ;
  assign y1615 = ~1'b0 ;
  assign y1616 = n3725 ;
  assign y1617 = ~n3727 ;
  assign y1618 = n3731 ;
  assign y1619 = ~n3736 ;
  assign y1620 = ~n3741 ;
  assign y1621 = ~n3747 ;
  assign y1622 = ~1'b0 ;
  assign y1623 = ~1'b0 ;
  assign y1624 = ~1'b0 ;
  assign y1625 = n3754 ;
  assign y1626 = ~n3760 ;
  assign y1627 = ~n3768 ;
  assign y1628 = ~n3769 ;
  assign y1629 = n777 ;
  assign y1630 = ~n3770 ;
  assign y1631 = ~1'b0 ;
  assign y1632 = n3777 ;
  assign y1633 = 1'b0 ;
  assign y1634 = n3778 ;
  assign y1635 = ~n3784 ;
  assign y1636 = n3789 ;
  assign y1637 = n3792 ;
  assign y1638 = n3795 ;
  assign y1639 = ~n3798 ;
  assign y1640 = n1694 ;
  assign y1641 = n3804 ;
  assign y1642 = n3805 ;
  assign y1643 = n3812 ;
  assign y1644 = ~n3814 ;
  assign y1645 = ~n3816 ;
  assign y1646 = ~n3817 ;
  assign y1647 = ~1'b0 ;
  assign y1648 = ~1'b0 ;
  assign y1649 = 1'b0 ;
  assign y1650 = n3819 ;
  assign y1651 = ~n3830 ;
  assign y1652 = ~n3832 ;
  assign y1653 = n3835 ;
  assign y1654 = n3846 ;
  assign y1655 = ~n3847 ;
  assign y1656 = ~n3848 ;
  assign y1657 = ~1'b0 ;
  assign y1658 = ~1'b0 ;
  assign y1659 = ~n3850 ;
  assign y1660 = ~n3851 ;
  assign y1661 = ~n3855 ;
  assign y1662 = n3860 ;
  assign y1663 = n3864 ;
  assign y1664 = ~1'b0 ;
  assign y1665 = ~1'b0 ;
  assign y1666 = ~1'b0 ;
  assign y1667 = ~1'b0 ;
  assign y1668 = ~n3866 ;
  assign y1669 = n3867 ;
  assign y1670 = ~n3871 ;
  assign y1671 = n3874 ;
  assign y1672 = n3876 ;
  assign y1673 = ~n3877 ;
  assign y1674 = n3878 ;
  assign y1675 = ~1'b0 ;
  assign y1676 = ~1'b0 ;
  assign y1677 = ~1'b0 ;
  assign y1678 = n3880 ;
  assign y1679 = ~n3881 ;
  assign y1680 = n3883 ;
  assign y1681 = ~n3885 ;
  assign y1682 = ~1'b0 ;
  assign y1683 = ~1'b0 ;
  assign y1684 = ~n3891 ;
  assign y1685 = n3893 ;
  assign y1686 = ~n3894 ;
  assign y1687 = n63 ;
  assign y1688 = ~1'b0 ;
  assign y1689 = n3901 ;
  assign y1690 = ~n3902 ;
  assign y1691 = n3905 ;
  assign y1692 = ~n3906 ;
  assign y1693 = ~1'b0 ;
  assign y1694 = n3908 ;
  assign y1695 = ~n3914 ;
  assign y1696 = n3916 ;
  assign y1697 = ~1'b0 ;
  assign y1698 = ~1'b0 ;
  assign y1699 = ~1'b0 ;
  assign y1700 = ~n3920 ;
  assign y1701 = ~n3922 ;
  assign y1702 = n3930 ;
  assign y1703 = n3931 ;
  assign y1704 = n3934 ;
  assign y1705 = ~n3936 ;
  assign y1706 = ~1'b0 ;
  assign y1707 = ~n3940 ;
  assign y1708 = n3941 ;
  assign y1709 = ~n3945 ;
  assign y1710 = ~n3948 ;
  assign y1711 = ~n3949 ;
  assign y1712 = ~1'b0 ;
  assign y1713 = n3950 ;
  assign y1714 = ~n3951 ;
  assign y1715 = ~n3953 ;
  assign y1716 = n2925 ;
  assign y1717 = ~n2070 ;
  assign y1718 = ~1'b0 ;
  assign y1719 = n3957 ;
  assign y1720 = n3961 ;
  assign y1721 = 1'b0 ;
  assign y1722 = n3964 ;
  assign y1723 = ~n3971 ;
  assign y1724 = ~n3982 ;
  assign y1725 = ~n3984 ;
  assign y1726 = n3987 ;
  assign y1727 = ~n3993 ;
  assign y1728 = n3994 ;
  assign y1729 = n3997 ;
  assign y1730 = n2004 ;
  assign y1731 = n4000 ;
  assign y1732 = n4002 ;
  assign y1733 = n4004 ;
  assign y1734 = n4006 ;
  assign y1735 = n4011 ;
  assign y1736 = ~n4021 ;
  assign y1737 = ~1'b0 ;
  assign y1738 = ~n4024 ;
  assign y1739 = ~n4027 ;
  assign y1740 = n2747 ;
  assign y1741 = ~n4032 ;
  assign y1742 = ~n4036 ;
  assign y1743 = ~n3027 ;
  assign y1744 = n4039 ;
  assign y1745 = n4043 ;
  assign y1746 = ~1'b0 ;
  assign y1747 = ~1'b0 ;
  assign y1748 = ~n4045 ;
  assign y1749 = n4047 ;
  assign y1750 = ~1'b0 ;
  assign y1751 = ~1'b0 ;
  assign y1752 = n4050 ;
  assign y1753 = ~1'b0 ;
  assign y1754 = n4053 ;
  assign y1755 = ~1'b0 ;
  assign y1756 = n4056 ;
  assign y1757 = n4057 ;
  assign y1758 = ~n4065 ;
  assign y1759 = ~n4070 ;
  assign y1760 = ~n4071 ;
  assign y1761 = ~n4074 ;
  assign y1762 = ~n4078 ;
  assign y1763 = ~n4079 ;
  assign y1764 = n4083 ;
  assign y1765 = ~1'b0 ;
  assign y1766 = n4084 ;
  assign y1767 = n4092 ;
  assign y1768 = ~n4095 ;
  assign y1769 = n4097 ;
  assign y1770 = ~n4099 ;
  assign y1771 = n4104 ;
  assign y1772 = ~n2254 ;
  assign y1773 = n4113 ;
  assign y1774 = ~1'b0 ;
  assign y1775 = n4114 ;
  assign y1776 = ~1'b0 ;
  assign y1777 = n4115 ;
  assign y1778 = n4121 ;
  assign y1779 = ~1'b0 ;
  assign y1780 = ~1'b0 ;
  assign y1781 = ~1'b0 ;
  assign y1782 = ~n4123 ;
  assign y1783 = ~1'b0 ;
  assign y1784 = ~n4124 ;
  assign y1785 = ~1'b0 ;
  assign y1786 = ~1'b0 ;
  assign y1787 = ~n4128 ;
  assign y1788 = n4135 ;
  assign y1789 = ~n4141 ;
  assign y1790 = n4142 ;
  assign y1791 = n1367 ;
  assign y1792 = n4150 ;
  assign y1793 = ~n4151 ;
  assign y1794 = ~n4154 ;
  assign y1795 = ~n4160 ;
  assign y1796 = ~n4165 ;
  assign y1797 = ~n68 ;
  assign y1798 = n4171 ;
  assign y1799 = ~n4175 ;
  assign y1800 = n4177 ;
  assign y1801 = n4179 ;
  assign y1802 = n4181 ;
  assign y1803 = n4185 ;
  assign y1804 = ~n4186 ;
  assign y1805 = ~n4187 ;
  assign y1806 = ~n4191 ;
  assign y1807 = n4195 ;
  assign y1808 = n4196 ;
  assign y1809 = n4197 ;
  assign y1810 = ~1'b0 ;
  assign y1811 = ~1'b0 ;
  assign y1812 = ~n4200 ;
  assign y1813 = ~1'b0 ;
  assign y1814 = ~n350 ;
  assign y1815 = 1'b0 ;
  assign y1816 = ~n4207 ;
  assign y1817 = ~n4210 ;
  assign y1818 = ~1'b0 ;
  assign y1819 = ~1'b0 ;
  assign y1820 = ~n4211 ;
  assign y1821 = n4215 ;
  assign y1822 = n4217 ;
  assign y1823 = n4218 ;
  assign y1824 = n4219 ;
  assign y1825 = ~n4223 ;
  assign y1826 = n4225 ;
  assign y1827 = n4228 ;
  assign y1828 = ~n4230 ;
  assign y1829 = n4233 ;
  assign y1830 = n4234 ;
  assign y1831 = ~1'b0 ;
  assign y1832 = ~1'b0 ;
  assign y1833 = ~n4237 ;
  assign y1834 = ~n4239 ;
  assign y1835 = ~n4241 ;
  assign y1836 = n4242 ;
  assign y1837 = n4249 ;
  assign y1838 = n4251 ;
  assign y1839 = ~1'b0 ;
  assign y1840 = ~n4252 ;
  assign y1841 = ~n4253 ;
  assign y1842 = ~n4256 ;
  assign y1843 = n471 ;
  assign y1844 = n4257 ;
  assign y1845 = ~1'b0 ;
  assign y1846 = 1'b0 ;
  assign y1847 = ~1'b0 ;
  assign y1848 = n4259 ;
  assign y1849 = ~n4263 ;
  assign y1850 = ~n4264 ;
  assign y1851 = n4265 ;
  assign y1852 = ~1'b0 ;
  assign y1853 = ~1'b0 ;
  assign y1854 = ~n4271 ;
  assign y1855 = ~n4274 ;
  assign y1856 = ~1'b0 ;
  assign y1857 = n4278 ;
  assign y1858 = ~n4280 ;
  assign y1859 = n4285 ;
  assign y1860 = ~n4286 ;
  assign y1861 = ~1'b0 ;
  assign y1862 = ~1'b0 ;
  assign y1863 = 1'b0 ;
  assign y1864 = ~1'b0 ;
  assign y1865 = n4287 ;
  assign y1866 = ~n4294 ;
  assign y1867 = n4297 ;
  assign y1868 = ~1'b0 ;
  assign y1869 = n4303 ;
  assign y1870 = n4304 ;
  assign y1871 = 1'b0 ;
  assign y1872 = ~1'b0 ;
  assign y1873 = ~1'b0 ;
  assign y1874 = ~1'b0 ;
  assign y1875 = ~1'b0 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = ~n4305 ;
  assign y1878 = ~n4308 ;
  assign y1879 = n4311 ;
  assign y1880 = ~n4313 ;
  assign y1881 = ~1'b0 ;
  assign y1882 = ~n4315 ;
  assign y1883 = ~n4318 ;
  assign y1884 = ~1'b0 ;
  assign y1885 = ~n4320 ;
  assign y1886 = n4324 ;
  assign y1887 = ~n4325 ;
  assign y1888 = ~n4326 ;
  assign y1889 = ~n4328 ;
  assign y1890 = ~1'b0 ;
  assign y1891 = n4331 ;
  assign y1892 = ~n799 ;
  assign y1893 = ~n4334 ;
  assign y1894 = ~1'b0 ;
  assign y1895 = n4336 ;
  assign y1896 = ~n4337 ;
  assign y1897 = ~1'b0 ;
  assign y1898 = ~n4338 ;
  assign y1899 = ~n1875 ;
  assign y1900 = ~n4341 ;
  assign y1901 = n4342 ;
  assign y1902 = ~n4105 ;
  assign y1903 = n4347 ;
  assign y1904 = ~n4348 ;
  assign y1905 = n4350 ;
  assign y1906 = n4354 ;
  assign y1907 = n4355 ;
  assign y1908 = n4356 ;
  assign y1909 = ~n4359 ;
  assign y1910 = ~1'b0 ;
  assign y1911 = ~n4363 ;
  assign y1912 = n4364 ;
  assign y1913 = ~1'b0 ;
  assign y1914 = ~1'b0 ;
  assign y1915 = ~1'b0 ;
  assign y1916 = ~n4365 ;
  assign y1917 = ~n4367 ;
  assign y1918 = 1'b0 ;
  assign y1919 = ~n3469 ;
  assign y1920 = n4369 ;
  assign y1921 = ~n4371 ;
  assign y1922 = n4372 ;
  assign y1923 = n1459 ;
  assign y1924 = ~n4373 ;
  assign y1925 = n4380 ;
  assign y1926 = ~n4381 ;
  assign y1927 = ~n4382 ;
  assign y1928 = ~n4383 ;
  assign y1929 = n4388 ;
  assign y1930 = n4390 ;
  assign y1931 = ~1'b0 ;
  assign y1932 = n4394 ;
  assign y1933 = ~1'b0 ;
  assign y1934 = ~1'b0 ;
  assign y1935 = ~n4397 ;
  assign y1936 = ~n4403 ;
  assign y1937 = ~1'b0 ;
  assign y1938 = ~1'b0 ;
  assign y1939 = ~1'b0 ;
  assign y1940 = ~n4406 ;
  assign y1941 = ~n4408 ;
  assign y1942 = ~n4411 ;
  assign y1943 = n2421 ;
  assign y1944 = ~n4412 ;
  assign y1945 = ~n4419 ;
  assign y1946 = n4421 ;
  assign y1947 = ~1'b0 ;
  assign y1948 = n4422 ;
  assign y1949 = ~1'b0 ;
  assign y1950 = n4425 ;
  assign y1951 = ~n4426 ;
  assign y1952 = ~1'b0 ;
  assign y1953 = 1'b0 ;
  assign y1954 = n4429 ;
  assign y1955 = n4439 ;
  assign y1956 = ~n4442 ;
  assign y1957 = ~n4447 ;
  assign y1958 = n4455 ;
  assign y1959 = n4460 ;
  assign y1960 = n4465 ;
  assign y1961 = n4473 ;
  assign y1962 = ~n4479 ;
  assign y1963 = ~1'b0 ;
  assign y1964 = n4480 ;
  assign y1965 = ~n4483 ;
  assign y1966 = n4487 ;
  assign y1967 = n4497 ;
  assign y1968 = ~n4505 ;
  assign y1969 = ~n4506 ;
  assign y1970 = n4507 ;
  assign y1971 = ~1'b0 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = ~1'b0 ;
  assign y1974 = n4510 ;
  assign y1975 = ~1'b0 ;
  assign y1976 = n4512 ;
  assign y1977 = ~n4516 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = ~n4523 ;
  assign y1980 = n4528 ;
  assign y1981 = n4529 ;
  assign y1982 = n4530 ;
  assign y1983 = ~n4531 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = ~1'b0 ;
  assign y1986 = ~1'b0 ;
  assign y1987 = n4534 ;
  assign y1988 = n4536 ;
  assign y1989 = n4537 ;
  assign y1990 = n4542 ;
  assign y1991 = n4545 ;
  assign y1992 = n4548 ;
  assign y1993 = ~n4553 ;
  assign y1994 = ~n4555 ;
  assign y1995 = ~n4557 ;
  assign y1996 = ~n4558 ;
  assign y1997 = ~n4560 ;
  assign y1998 = n4562 ;
  assign y1999 = n4569 ;
  assign y2000 = ~1'b0 ;
  assign y2001 = ~1'b0 ;
  assign y2002 = n4571 ;
  assign y2003 = ~1'b0 ;
  assign y2004 = n4572 ;
  assign y2005 = ~n4578 ;
  assign y2006 = ~1'b0 ;
  assign y2007 = ~n4579 ;
  assign y2008 = n4587 ;
  assign y2009 = n3288 ;
  assign y2010 = ~1'b0 ;
  assign y2011 = ~n4590 ;
  assign y2012 = ~n216 ;
  assign y2013 = ~1'b0 ;
  assign y2014 = n601 ;
  assign y2015 = ~1'b0 ;
  assign y2016 = n4596 ;
  assign y2017 = ~1'b0 ;
  assign y2018 = n4599 ;
  assign y2019 = ~n4605 ;
  assign y2020 = ~n4610 ;
  assign y2021 = n4612 ;
  assign y2022 = ~n4615 ;
  assign y2023 = ~1'b0 ;
  assign y2024 = n4618 ;
  assign y2025 = n3508 ;
  assign y2026 = n4620 ;
  assign y2027 = n4629 ;
  assign y2028 = ~n4631 ;
  assign y2029 = 1'b0 ;
  assign y2030 = ~n4635 ;
  assign y2031 = n4639 ;
  assign y2032 = n4640 ;
  assign y2033 = n4642 ;
  assign y2034 = ~n2677 ;
  assign y2035 = ~1'b0 ;
  assign y2036 = ~n4644 ;
  assign y2037 = n4647 ;
  assign y2038 = ~n4648 ;
  assign y2039 = ~n3199 ;
  assign y2040 = n3004 ;
  assign y2041 = ~1'b0 ;
  assign y2042 = n4650 ;
  assign y2043 = n4654 ;
  assign y2044 = ~n4657 ;
  assign y2045 = ~n1773 ;
  assign y2046 = n4658 ;
  assign y2047 = ~n4662 ;
  assign y2048 = ~1'b0 ;
  assign y2049 = ~1'b0 ;
  assign y2050 = ~1'b0 ;
  assign y2051 = n4663 ;
  assign y2052 = ~n4667 ;
  assign y2053 = ~n4668 ;
  assign y2054 = n4670 ;
  assign y2055 = ~n4674 ;
  assign y2056 = n4677 ;
  assign y2057 = ~1'b0 ;
  assign y2058 = n4685 ;
  assign y2059 = ~n4689 ;
  assign y2060 = 1'b0 ;
  assign y2061 = ~1'b0 ;
  assign y2062 = ~n2815 ;
  assign y2063 = n4691 ;
  assign y2064 = ~n3466 ;
  assign y2065 = ~1'b0 ;
  assign y2066 = ~n4698 ;
  assign y2067 = n4701 ;
  assign y2068 = n4702 ;
  assign y2069 = n4711 ;
  assign y2070 = n4712 ;
  assign y2071 = ~n4713 ;
  assign y2072 = ~1'b0 ;
  assign y2073 = n4715 ;
  assign y2074 = n4717 ;
  assign y2075 = n4207 ;
  assign y2076 = 1'b0 ;
  assign y2077 = n4721 ;
  assign y2078 = ~1'b0 ;
  assign y2079 = ~n4742 ;
  assign y2080 = n4745 ;
  assign y2081 = n4747 ;
  assign y2082 = ~n4749 ;
  assign y2083 = ~1'b0 ;
  assign y2084 = n4752 ;
  assign y2085 = ~n4758 ;
  assign y2086 = ~1'b0 ;
  assign y2087 = n4769 ;
  assign y2088 = n4770 ;
  assign y2089 = n4772 ;
  assign y2090 = n4779 ;
  assign y2091 = ~1'b0 ;
  assign y2092 = ~n4780 ;
  assign y2093 = ~n4781 ;
  assign y2094 = n1545 ;
  assign y2095 = ~n4786 ;
  assign y2096 = ~n4792 ;
  assign y2097 = n4804 ;
  assign y2098 = ~1'b0 ;
  assign y2099 = n4807 ;
  assign y2100 = n4810 ;
  assign y2101 = ~1'b0 ;
  assign y2102 = ~n4817 ;
  assign y2103 = ~1'b0 ;
  assign y2104 = n4819 ;
  assign y2105 = n4826 ;
  assign y2106 = ~n4827 ;
  assign y2107 = ~n4832 ;
  assign y2108 = ~n4834 ;
  assign y2109 = ~n4838 ;
  assign y2110 = ~1'b0 ;
  assign y2111 = n4842 ;
  assign y2112 = n4845 ;
  assign y2113 = ~n4851 ;
  assign y2114 = n4854 ;
  assign y2115 = n4856 ;
  assign y2116 = n4857 ;
  assign y2117 = ~1'b0 ;
  assign y2118 = ~x3 ;
  assign y2119 = n4860 ;
  assign y2120 = ~n4863 ;
  assign y2121 = ~1'b0 ;
  assign y2122 = ~n4864 ;
  assign y2123 = n4875 ;
  assign y2124 = ~n4878 ;
  assign y2125 = ~n4886 ;
  assign y2126 = n4894 ;
  assign y2127 = n4899 ;
  assign y2128 = n4900 ;
  assign y2129 = n4903 ;
  assign y2130 = ~1'b0 ;
  assign y2131 = ~1'b0 ;
  assign y2132 = ~n4904 ;
  assign y2133 = n4906 ;
  assign y2134 = ~n4908 ;
  assign y2135 = n4911 ;
  assign y2136 = n4916 ;
  assign y2137 = ~n4918 ;
  assign y2138 = ~n4923 ;
  assign y2139 = n4925 ;
  assign y2140 = n4928 ;
  assign y2141 = ~1'b0 ;
  assign y2142 = n4931 ;
  assign y2143 = n1623 ;
  assign y2144 = ~1'b0 ;
  assign y2145 = n4933 ;
  assign y2146 = n601 ;
  assign y2147 = ~n4937 ;
  assign y2148 = n4939 ;
  assign y2149 = ~n4941 ;
  assign y2150 = ~n4944 ;
  assign y2151 = n4945 ;
  assign y2152 = ~n4949 ;
  assign y2153 = ~1'b0 ;
  assign y2154 = ~1'b0 ;
  assign y2155 = ~1'b0 ;
  assign y2156 = n4953 ;
  assign y2157 = ~n4961 ;
  assign y2158 = ~n4964 ;
  assign y2159 = n4965 ;
  assign y2160 = n4967 ;
  assign y2161 = n4968 ;
  assign y2162 = n4969 ;
  assign y2163 = n4970 ;
  assign y2164 = n4976 ;
  assign y2165 = n4977 ;
  assign y2166 = ~n4978 ;
  assign y2167 = ~n4980 ;
  assign y2168 = n4981 ;
  assign y2169 = n1812 ;
  assign y2170 = n4983 ;
  assign y2171 = ~1'b0 ;
  assign y2172 = ~1'b0 ;
  assign y2173 = ~1'b0 ;
  assign y2174 = ~n4990 ;
  assign y2175 = n4992 ;
  assign y2176 = ~n4993 ;
  assign y2177 = n4998 ;
  assign y2178 = n4999 ;
  assign y2179 = n5004 ;
  assign y2180 = ~n5007 ;
  assign y2181 = ~n5009 ;
  assign y2182 = n5011 ;
  assign y2183 = ~1'b0 ;
  assign y2184 = n5013 ;
  assign y2185 = ~n5014 ;
  assign y2186 = n5016 ;
  assign y2187 = ~n5018 ;
  assign y2188 = ~n5029 ;
  assign y2189 = n5040 ;
  assign y2190 = ~n5042 ;
  assign y2191 = ~n5043 ;
  assign y2192 = ~n5045 ;
  assign y2193 = ~n5048 ;
  assign y2194 = ~1'b0 ;
  assign y2195 = ~n5051 ;
  assign y2196 = ~n5057 ;
  assign y2197 = n5058 ;
  assign y2198 = n5073 ;
  assign y2199 = n5082 ;
  assign y2200 = ~n5084 ;
  assign y2201 = n5089 ;
  assign y2202 = ~n5091 ;
  assign y2203 = 1'b0 ;
  assign y2204 = ~n5097 ;
  assign y2205 = ~n5101 ;
  assign y2206 = n5108 ;
  assign y2207 = n5109 ;
  assign y2208 = ~1'b0 ;
  assign y2209 = ~n5110 ;
  assign y2210 = ~n5112 ;
  assign y2211 = ~1'b0 ;
  assign y2212 = ~1'b0 ;
  assign y2213 = ~n5113 ;
  assign y2214 = ~n5119 ;
  assign y2215 = ~n5120 ;
  assign y2216 = n5122 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = ~1'b0 ;
  assign y2219 = ~1'b0 ;
  assign y2220 = ~n5124 ;
  assign y2221 = ~1'b0 ;
  assign y2222 = ~n5127 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = ~1'b0 ;
  assign y2225 = ~n5131 ;
  assign y2226 = n5135 ;
  assign y2227 = n5136 ;
  assign y2228 = n5140 ;
  assign y2229 = n5144 ;
  assign y2230 = ~n5147 ;
  assign y2231 = n2327 ;
  assign y2232 = ~n5153 ;
  assign y2233 = ~n5157 ;
  assign y2234 = ~1'b0 ;
  assign y2235 = ~1'b0 ;
  assign y2236 = ~1'b0 ;
  assign y2237 = ~n5161 ;
  assign y2238 = ~1'b0 ;
  assign y2239 = ~1'b0 ;
  assign y2240 = ~n5165 ;
  assign y2241 = n5166 ;
  assign y2242 = ~n5175 ;
  assign y2243 = ~n5176 ;
  assign y2244 = ~n5178 ;
  assign y2245 = ~n5180 ;
  assign y2246 = n5182 ;
  assign y2247 = ~n5186 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = ~1'b0 ;
  assign y2250 = ~n5188 ;
  assign y2251 = n1295 ;
  assign y2252 = ~1'b0 ;
  assign y2253 = ~n2602 ;
  assign y2254 = n5189 ;
  assign y2255 = ~1'b0 ;
  assign y2256 = ~n5199 ;
  assign y2257 = ~1'b0 ;
  assign y2258 = ~1'b0 ;
  assign y2259 = ~1'b0 ;
  assign y2260 = n310 ;
  assign y2261 = n5200 ;
  assign y2262 = n5204 ;
  assign y2263 = n5206 ;
  assign y2264 = ~n5207 ;
  assign y2265 = n4381 ;
  assign y2266 = ~1'b0 ;
  assign y2267 = ~n5214 ;
  assign y2268 = n5220 ;
  assign y2269 = n5224 ;
  assign y2270 = 1'b0 ;
  assign y2271 = ~1'b0 ;
  assign y2272 = n5225 ;
  assign y2273 = ~1'b0 ;
  assign y2274 = ~n5228 ;
  assign y2275 = n5237 ;
  assign y2276 = n5240 ;
  assign y2277 = n5242 ;
  assign y2278 = 1'b0 ;
  assign y2279 = ~1'b0 ;
  assign y2280 = n5244 ;
  assign y2281 = ~n1668 ;
  assign y2282 = ~n5247 ;
  assign y2283 = ~n5250 ;
  assign y2284 = n5252 ;
  assign y2285 = n5253 ;
  assign y2286 = ~1'b0 ;
  assign y2287 = ~n5254 ;
  assign y2288 = ~n5255 ;
  assign y2289 = ~n5258 ;
  assign y2290 = n3898 ;
  assign y2291 = n5262 ;
  assign y2292 = n5270 ;
  assign y2293 = ~1'b0 ;
  assign y2294 = ~1'b0 ;
  assign y2295 = n5272 ;
  assign y2296 = 1'b0 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = ~n5274 ;
  assign y2299 = ~n5277 ;
  assign y2300 = n5279 ;
  assign y2301 = n5280 ;
  assign y2302 = ~n5286 ;
  assign y2303 = ~n5287 ;
  assign y2304 = ~1'b0 ;
  assign y2305 = ~n5298 ;
  assign y2306 = n5304 ;
  assign y2307 = ~1'b0 ;
  assign y2308 = n5307 ;
  assign y2309 = ~1'b0 ;
  assign y2310 = ~n5309 ;
  assign y2311 = ~n5310 ;
  assign y2312 = ~n5311 ;
  assign y2313 = ~n5312 ;
  assign y2314 = ~n5321 ;
  assign y2315 = ~1'b0 ;
  assign y2316 = ~n5322 ;
  assign y2317 = n5324 ;
  assign y2318 = ~n5329 ;
  assign y2319 = n5331 ;
  assign y2320 = n5333 ;
  assign y2321 = ~1'b0 ;
  assign y2322 = ~n5337 ;
  assign y2323 = ~n5341 ;
  assign y2324 = ~n5342 ;
  assign y2325 = n5344 ;
  assign y2326 = n5346 ;
  assign y2327 = ~n5355 ;
  assign y2328 = ~n5356 ;
  assign y2329 = n5357 ;
  assign y2330 = n5361 ;
  assign y2331 = ~1'b0 ;
  assign y2332 = n5364 ;
  assign y2333 = ~n5365 ;
  assign y2334 = ~n5366 ;
  assign y2335 = n5368 ;
  assign y2336 = n5372 ;
  assign y2337 = ~n5374 ;
  assign y2338 = n5376 ;
  assign y2339 = ~n5378 ;
  assign y2340 = n5381 ;
  assign y2341 = n44 ;
  assign y2342 = ~1'b0 ;
  assign y2343 = ~n5384 ;
  assign y2344 = n5386 ;
  assign y2345 = ~n5391 ;
  assign y2346 = ~n5392 ;
  assign y2347 = ~1'b0 ;
  assign y2348 = n45 ;
  assign y2349 = ~1'b0 ;
  assign y2350 = ~1'b0 ;
  assign y2351 = n5394 ;
  assign y2352 = ~n5396 ;
  assign y2353 = n5399 ;
  assign y2354 = ~n5402 ;
  assign y2355 = n5417 ;
  assign y2356 = ~n5421 ;
  assign y2357 = ~n5430 ;
  assign y2358 = ~n5433 ;
  assign y2359 = ~n5435 ;
  assign y2360 = n5436 ;
  assign y2361 = n5437 ;
  assign y2362 = n5440 ;
  assign y2363 = n2674 ;
  assign y2364 = n2391 ;
  assign y2365 = ~1'b0 ;
  assign y2366 = ~1'b0 ;
  assign y2367 = n5442 ;
  assign y2368 = n1904 ;
  assign y2369 = n5446 ;
  assign y2370 = n5461 ;
  assign y2371 = 1'b0 ;
  assign y2372 = n5468 ;
  assign y2373 = n892 ;
  assign y2374 = ~n5469 ;
  assign y2375 = n455 ;
  assign y2376 = n5479 ;
  assign y2377 = n5481 ;
  assign y2378 = n5486 ;
  assign y2379 = n5491 ;
  assign y2380 = n5493 ;
  assign y2381 = ~1'b0 ;
  assign y2382 = ~n5495 ;
  assign y2383 = n4681 ;
  assign y2384 = ~n5498 ;
  assign y2385 = ~n1766 ;
  assign y2386 = n615 ;
  assign y2387 = ~n5506 ;
  assign y2388 = ~n5508 ;
  assign y2389 = ~n5512 ;
  assign y2390 = ~n5513 ;
  assign y2391 = ~1'b0 ;
  assign y2392 = ~1'b0 ;
  assign y2393 = n5533 ;
  assign y2394 = ~1'b0 ;
  assign y2395 = n5534 ;
  assign y2396 = 1'b0 ;
  assign y2397 = ~n5536 ;
  assign y2398 = ~1'b0 ;
  assign y2399 = ~1'b0 ;
  assign y2400 = ~n5540 ;
  assign y2401 = ~n5550 ;
  assign y2402 = ~1'b0 ;
  assign y2403 = 1'b0 ;
  assign y2404 = n5552 ;
  assign y2405 = ~n5556 ;
  assign y2406 = n5562 ;
  assign y2407 = ~1'b0 ;
  assign y2408 = n5563 ;
  assign y2409 = n5564 ;
  assign y2410 = ~n3563 ;
  assign y2411 = n5568 ;
  assign y2412 = n5570 ;
  assign y2413 = ~n5571 ;
  assign y2414 = ~n5573 ;
  assign y2415 = ~1'b0 ;
  assign y2416 = ~n5576 ;
  assign y2417 = n5585 ;
  assign y2418 = n5589 ;
  assign y2419 = n5595 ;
  assign y2420 = ~n5601 ;
  assign y2421 = n5604 ;
  assign y2422 = n5610 ;
  assign y2423 = ~1'b0 ;
  assign y2424 = ~1'b0 ;
  assign y2425 = ~n5615 ;
  assign y2426 = n5622 ;
  assign y2427 = ~n5623 ;
  assign y2428 = n5625 ;
  assign y2429 = n2190 ;
  assign y2430 = ~n5627 ;
  assign y2431 = ~1'b0 ;
  assign y2432 = n5628 ;
  assign y2433 = n5631 ;
  assign y2434 = n5632 ;
  assign y2435 = ~1'b0 ;
  assign y2436 = n5635 ;
  assign y2437 = ~1'b0 ;
  assign y2438 = ~n5641 ;
  assign y2439 = ~n5650 ;
  assign y2440 = ~n5653 ;
  assign y2441 = ~n5655 ;
  assign y2442 = ~1'b0 ;
  assign y2443 = ~n5658 ;
  assign y2444 = ~n1169 ;
  assign y2445 = n5662 ;
  assign y2446 = ~1'b0 ;
  assign y2447 = ~1'b0 ;
  assign y2448 = ~n5663 ;
  assign y2449 = n5668 ;
  assign y2450 = n5679 ;
  assign y2451 = ~n5688 ;
  assign y2452 = ~n4976 ;
  assign y2453 = n5690 ;
  assign y2454 = n5693 ;
  assign y2455 = ~n5697 ;
  assign y2456 = ~n5704 ;
  assign y2457 = 1'b0 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = n5708 ;
  assign y2460 = ~n5709 ;
  assign y2461 = 1'b0 ;
  assign y2462 = ~1'b0 ;
  assign y2463 = n5712 ;
  assign y2464 = ~n5719 ;
  assign y2465 = ~n5725 ;
  assign y2466 = n5730 ;
  assign y2467 = ~1'b0 ;
  assign y2468 = ~n5734 ;
  assign y2469 = 1'b0 ;
  assign y2470 = ~n5736 ;
  assign y2471 = n5738 ;
  assign y2472 = n5741 ;
  assign y2473 = n5743 ;
  assign y2474 = ~1'b0 ;
  assign y2475 = ~1'b0 ;
  assign y2476 = n5744 ;
  assign y2477 = ~1'b0 ;
  assign y2478 = n2019 ;
  assign y2479 = 1'b0 ;
  assign y2480 = ~n5745 ;
  assign y2481 = ~1'b0 ;
  assign y2482 = n5747 ;
  assign y2483 = ~1'b0 ;
  assign y2484 = n5750 ;
  assign y2485 = n5753 ;
  assign y2486 = ~n5757 ;
  assign y2487 = ~1'b0 ;
  assign y2488 = ~n5758 ;
  assign y2489 = ~n5764 ;
  assign y2490 = n5771 ;
  assign y2491 = ~n5778 ;
  assign y2492 = ~n5781 ;
  assign y2493 = ~n5785 ;
  assign y2494 = ~1'b0 ;
  assign y2495 = ~n5786 ;
  assign y2496 = ~n5788 ;
  assign y2497 = ~n5790 ;
  assign y2498 = ~n5791 ;
  assign y2499 = ~n5796 ;
  assign y2500 = n5799 ;
  assign y2501 = ~1'b0 ;
  assign y2502 = n5803 ;
  assign y2503 = n5804 ;
  assign y2504 = n5806 ;
  assign y2505 = ~1'b0 ;
  assign y2506 = ~n5808 ;
  assign y2507 = ~n5813 ;
  assign y2508 = ~n5815 ;
  assign y2509 = ~n5823 ;
  assign y2510 = ~n5824 ;
  assign y2511 = ~1'b0 ;
  assign y2512 = ~n5830 ;
  assign y2513 = ~n5836 ;
  assign y2514 = n5837 ;
  assign y2515 = ~n5844 ;
  assign y2516 = ~n5847 ;
  assign y2517 = ~1'b0 ;
  assign y2518 = ~n5850 ;
  assign y2519 = ~n5851 ;
  assign y2520 = n5854 ;
  assign y2521 = ~n5858 ;
  assign y2522 = ~n5860 ;
  assign y2523 = n5861 ;
  assign y2524 = ~1'b0 ;
  assign y2525 = ~n5862 ;
  assign y2526 = ~n5864 ;
  assign y2527 = n5867 ;
  assign y2528 = ~1'b0 ;
  assign y2529 = ~1'b0 ;
  assign y2530 = ~n5868 ;
  assign y2531 = ~n5872 ;
  assign y2532 = n5877 ;
  assign y2533 = n5879 ;
  assign y2534 = ~n5882 ;
  assign y2535 = n5888 ;
  assign y2536 = n5896 ;
  assign y2537 = n5902 ;
  assign y2538 = ~n99 ;
  assign y2539 = ~1'b0 ;
  assign y2540 = ~1'b0 ;
  assign y2541 = n5903 ;
  assign y2542 = n5904 ;
  assign y2543 = n4147 ;
  assign y2544 = ~n5907 ;
  assign y2545 = n5911 ;
  assign y2546 = ~n5912 ;
  assign y2547 = ~1'b0 ;
  assign y2548 = n5914 ;
  assign y2549 = n5915 ;
  assign y2550 = n5916 ;
  assign y2551 = n5920 ;
  assign y2552 = ~n5923 ;
  assign y2553 = n5925 ;
  assign y2554 = ~1'b0 ;
  assign y2555 = ~n5927 ;
  assign y2556 = n5928 ;
  assign y2557 = n5931 ;
  assign y2558 = n5932 ;
  assign y2559 = ~n5933 ;
  assign y2560 = ~n5941 ;
  assign y2561 = ~1'b0 ;
  assign y2562 = n3717 ;
  assign y2563 = 1'b0 ;
  assign y2564 = ~n5948 ;
  assign y2565 = ~n5949 ;
  assign y2566 = n5953 ;
  assign y2567 = ~n5955 ;
  assign y2568 = n5958 ;
  assign y2569 = ~n5959 ;
  assign y2570 = ~n5963 ;
  assign y2571 = ~1'b0 ;
  assign y2572 = ~1'b0 ;
  assign y2573 = ~1'b0 ;
  assign y2574 = n5969 ;
  assign y2575 = ~n5972 ;
  assign y2576 = ~1'b0 ;
  assign y2577 = ~n5975 ;
  assign y2578 = ~n5978 ;
  assign y2579 = n5979 ;
  assign y2580 = n5982 ;
  assign y2581 = n5988 ;
  assign y2582 = ~n5995 ;
  assign y2583 = ~n5996 ;
  assign y2584 = ~1'b0 ;
  assign y2585 = n5997 ;
  assign y2586 = ~n5998 ;
  assign y2587 = ~n6003 ;
  assign y2588 = n6004 ;
  assign y2589 = 1'b0 ;
  assign y2590 = ~1'b0 ;
  assign y2591 = n6005 ;
  assign y2592 = n6010 ;
  assign y2593 = ~n6014 ;
  assign y2594 = ~n6016 ;
  assign y2595 = ~n6019 ;
  assign y2596 = ~n6020 ;
  assign y2597 = ~n6022 ;
  assign y2598 = 1'b0 ;
  assign y2599 = n4803 ;
  assign y2600 = ~1'b0 ;
  assign y2601 = ~1'b0 ;
  assign y2602 = ~n6026 ;
  assign y2603 = n6027 ;
  assign y2604 = n6030 ;
  assign y2605 = ~n6034 ;
  assign y2606 = n6040 ;
  assign y2607 = ~n6042 ;
  assign y2608 = ~n6043 ;
  assign y2609 = ~1'b0 ;
  assign y2610 = n6049 ;
  assign y2611 = ~n6050 ;
  assign y2612 = ~n1348 ;
  assign y2613 = ~n6060 ;
  assign y2614 = ~n6064 ;
  assign y2615 = ~1'b0 ;
  assign y2616 = ~n6069 ;
  assign y2617 = ~n6074 ;
  assign y2618 = ~n6075 ;
  assign y2619 = n6080 ;
  assign y2620 = ~1'b0 ;
  assign y2621 = ~n6082 ;
  assign y2622 = ~1'b0 ;
  assign y2623 = n4545 ;
  assign y2624 = ~n6089 ;
  assign y2625 = n6091 ;
  assign y2626 = 1'b0 ;
  assign y2627 = ~n6093 ;
  assign y2628 = n6094 ;
  assign y2629 = ~n6096 ;
  assign y2630 = n6097 ;
  assign y2631 = ~1'b0 ;
  assign y2632 = n6098 ;
  assign y2633 = n6100 ;
  assign y2634 = n6101 ;
  assign y2635 = n6107 ;
  assign y2636 = ~1'b0 ;
  assign y2637 = ~n6116 ;
  assign y2638 = ~n6121 ;
  assign y2639 = ~n6122 ;
  assign y2640 = n6129 ;
  assign y2641 = n6131 ;
  assign y2642 = ~n6134 ;
  assign y2643 = ~n6135 ;
  assign y2644 = ~n6138 ;
  assign y2645 = n6147 ;
  assign y2646 = ~1'b0 ;
  assign y2647 = ~1'b0 ;
  assign y2648 = n6149 ;
  assign y2649 = ~n6155 ;
  assign y2650 = ~n6159 ;
  assign y2651 = ~n6160 ;
  assign y2652 = ~1'b0 ;
  assign y2653 = n6163 ;
  assign y2654 = ~1'b0 ;
  assign y2655 = ~1'b0 ;
  assign y2656 = ~1'b0 ;
  assign y2657 = n6167 ;
  assign y2658 = 1'b0 ;
  assign y2659 = 1'b0 ;
  assign y2660 = n1540 ;
  assign y2661 = ~n6168 ;
  assign y2662 = ~1'b0 ;
  assign y2663 = ~n6171 ;
  assign y2664 = ~1'b0 ;
  assign y2665 = n6173 ;
  assign y2666 = ~n6174 ;
  assign y2667 = n6176 ;
  assign y2668 = n3985 ;
  assign y2669 = ~n6178 ;
  assign y2670 = ~n6182 ;
  assign y2671 = ~n6183 ;
  assign y2672 = n6186 ;
  assign y2673 = ~n6188 ;
  assign y2674 = ~n6191 ;
  assign y2675 = n6193 ;
  assign y2676 = ~n6198 ;
  assign y2677 = n6199 ;
  assign y2678 = ~n6204 ;
  assign y2679 = ~n6206 ;
  assign y2680 = n1170 ;
  assign y2681 = ~n6210 ;
  assign y2682 = ~n6211 ;
  assign y2683 = ~1'b0 ;
  assign y2684 = n6212 ;
  assign y2685 = n6214 ;
  assign y2686 = ~n6218 ;
  assign y2687 = ~n3345 ;
  assign y2688 = ~1'b0 ;
  assign y2689 = ~n6219 ;
  assign y2690 = n6222 ;
  assign y2691 = ~1'b0 ;
  assign y2692 = ~n6223 ;
  assign y2693 = ~1'b0 ;
  assign y2694 = n6224 ;
  assign y2695 = ~n6225 ;
  assign y2696 = ~1'b0 ;
  assign y2697 = ~n6227 ;
  assign y2698 = n6229 ;
  assign y2699 = n6231 ;
  assign y2700 = ~1'b0 ;
  assign y2701 = ~1'b0 ;
  assign y2702 = ~1'b0 ;
  assign y2703 = ~1'b0 ;
  assign y2704 = n3517 ;
  assign y2705 = ~n6236 ;
  assign y2706 = n6239 ;
  assign y2707 = n6242 ;
  assign y2708 = ~n6251 ;
  assign y2709 = ~n6253 ;
  assign y2710 = n6254 ;
  assign y2711 = n6259 ;
  assign y2712 = n6267 ;
  assign y2713 = ~n6272 ;
  assign y2714 = ~n5400 ;
  assign y2715 = n6273 ;
  assign y2716 = ~1'b0 ;
  assign y2717 = ~n6274 ;
  assign y2718 = ~1'b0 ;
  assign y2719 = ~1'b0 ;
  assign y2720 = ~1'b0 ;
  assign y2721 = n6275 ;
  assign y2722 = n6282 ;
  assign y2723 = n6285 ;
  assign y2724 = ~1'b0 ;
  assign y2725 = ~1'b0 ;
  assign y2726 = n6291 ;
  assign y2727 = ~1'b0 ;
  assign y2728 = ~n6293 ;
  assign y2729 = 1'b0 ;
  assign y2730 = ~n2375 ;
  assign y2731 = ~n6294 ;
  assign y2732 = ~n6296 ;
  assign y2733 = ~1'b0 ;
  assign y2734 = ~1'b0 ;
  assign y2735 = ~1'b0 ;
  assign y2736 = ~1'b0 ;
  assign y2737 = n6299 ;
  assign y2738 = ~1'b0 ;
  assign y2739 = ~n6301 ;
  assign y2740 = ~n6307 ;
  assign y2741 = ~n6308 ;
  assign y2742 = n6310 ;
  assign y2743 = n6313 ;
  assign y2744 = n6317 ;
  assign y2745 = ~1'b0 ;
  assign y2746 = ~n6319 ;
  assign y2747 = n6324 ;
  assign y2748 = n6328 ;
  assign y2749 = ~n6330 ;
  assign y2750 = ~n6332 ;
  assign y2751 = ~n6335 ;
  assign y2752 = n6336 ;
  assign y2753 = n6340 ;
  assign y2754 = ~1'b0 ;
  assign y2755 = n4195 ;
  assign y2756 = ~n4877 ;
  assign y2757 = ~n6343 ;
  assign y2758 = ~n4937 ;
  assign y2759 = ~1'b0 ;
  assign y2760 = ~1'b0 ;
  assign y2761 = n6345 ;
  assign y2762 = ~n6346 ;
  assign y2763 = ~n6351 ;
  assign y2764 = n6352 ;
  assign y2765 = n6360 ;
  assign y2766 = ~n6366 ;
  assign y2767 = ~n6370 ;
  assign y2768 = ~n6375 ;
  assign y2769 = n3926 ;
  assign y2770 = ~1'b0 ;
  assign y2771 = ~1'b0 ;
  assign y2772 = 1'b0 ;
  assign y2773 = 1'b0 ;
  assign y2774 = n6376 ;
  assign y2775 = ~n6377 ;
  assign y2776 = n3784 ;
  assign y2777 = ~n6379 ;
  assign y2778 = ~n6381 ;
  assign y2779 = n2502 ;
  assign y2780 = n6382 ;
  assign y2781 = ~n6383 ;
  assign y2782 = ~1'b0 ;
  assign y2783 = n6385 ;
  assign y2784 = n6386 ;
  assign y2785 = ~n6387 ;
  assign y2786 = ~1'b0 ;
  assign y2787 = n6388 ;
  assign y2788 = ~n6390 ;
  assign y2789 = n6398 ;
  assign y2790 = ~n6403 ;
  assign y2791 = n6406 ;
  assign y2792 = ~n6407 ;
  assign y2793 = n6408 ;
  assign y2794 = ~n6411 ;
  assign y2795 = ~n926 ;
  assign y2796 = n6415 ;
  assign y2797 = n6417 ;
  assign y2798 = ~n3812 ;
  assign y2799 = ~1'b0 ;
  assign y2800 = ~1'b0 ;
  assign y2801 = ~1'b0 ;
  assign y2802 = 1'b0 ;
  assign y2803 = ~1'b0 ;
  assign y2804 = n6418 ;
  assign y2805 = ~n6420 ;
  assign y2806 = n6421 ;
  assign y2807 = n6422 ;
  assign y2808 = ~1'b0 ;
  assign y2809 = ~n6423 ;
  assign y2810 = ~1'b0 ;
  assign y2811 = ~1'b0 ;
  assign y2812 = ~1'b0 ;
  assign y2813 = ~1'b0 ;
  assign y2814 = n6431 ;
  assign y2815 = n6433 ;
  assign y2816 = n6441 ;
  assign y2817 = ~1'b0 ;
  assign y2818 = ~1'b0 ;
  assign y2819 = ~1'b0 ;
  assign y2820 = ~n6444 ;
  assign y2821 = ~1'b0 ;
  assign y2822 = n6446 ;
  assign y2823 = n6449 ;
  assign y2824 = n6450 ;
  assign y2825 = n6452 ;
  assign y2826 = ~n6454 ;
  assign y2827 = n6455 ;
  assign y2828 = ~n4376 ;
  assign y2829 = ~1'b0 ;
  assign y2830 = ~1'b0 ;
  assign y2831 = ~1'b0 ;
  assign y2832 = ~1'b0 ;
  assign y2833 = n6457 ;
  assign y2834 = ~n6464 ;
  assign y2835 = ~1'b0 ;
  assign y2836 = ~n6473 ;
  assign y2837 = ~n6478 ;
  assign y2838 = 1'b0 ;
  assign y2839 = n2334 ;
  assign y2840 = n6480 ;
  assign y2841 = ~n6482 ;
  assign y2842 = ~1'b0 ;
  assign y2843 = n6488 ;
  assign y2844 = ~n6495 ;
  assign y2845 = 1'b0 ;
  assign y2846 = ~n6496 ;
  assign y2847 = ~1'b0 ;
  assign y2848 = 1'b0 ;
  assign y2849 = ~1'b0 ;
  assign y2850 = ~1'b0 ;
  assign y2851 = ~1'b0 ;
  assign y2852 = ~1'b0 ;
  assign y2853 = n6497 ;
  assign y2854 = ~1'b0 ;
  assign y2855 = ~n6498 ;
  assign y2856 = n6500 ;
  assign y2857 = ~n6501 ;
  assign y2858 = n6506 ;
  assign y2859 = n6508 ;
  assign y2860 = ~n6509 ;
  assign y2861 = ~1'b0 ;
  assign y2862 = n6511 ;
  assign y2863 = ~1'b0 ;
  assign y2864 = 1'b0 ;
  assign y2865 = n6521 ;
  assign y2866 = n6523 ;
  assign y2867 = n6524 ;
  assign y2868 = n6526 ;
  assign y2869 = n6527 ;
  assign y2870 = n2784 ;
  assign y2871 = n6531 ;
  assign y2872 = n6532 ;
  assign y2873 = ~n6547 ;
  assign y2874 = ~n6549 ;
  assign y2875 = ~n6550 ;
  assign y2876 = ~n6552 ;
  assign y2877 = ~1'b0 ;
  assign y2878 = ~1'b0 ;
  assign y2879 = n6554 ;
  assign y2880 = ~n6556 ;
  assign y2881 = ~n6557 ;
  assign y2882 = n6561 ;
  assign y2883 = ~n6569 ;
  assign y2884 = ~n6575 ;
  assign y2885 = n6581 ;
  assign y2886 = ~n6582 ;
  assign y2887 = ~n6587 ;
  assign y2888 = n6593 ;
  assign y2889 = n6596 ;
  assign y2890 = n5415 ;
  assign y2891 = ~1'b0 ;
  assign y2892 = ~1'b0 ;
  assign y2893 = n6600 ;
  assign y2894 = n6601 ;
  assign y2895 = ~n6605 ;
  assign y2896 = ~n6606 ;
  assign y2897 = ~n6613 ;
  assign y2898 = n6615 ;
  assign y2899 = ~n6618 ;
  assign y2900 = ~n6622 ;
  assign y2901 = n6627 ;
  assign y2902 = n6628 ;
  assign y2903 = ~n6629 ;
  assign y2904 = n6630 ;
  assign y2905 = n6632 ;
  assign y2906 = ~1'b0 ;
  assign y2907 = ~n6636 ;
  assign y2908 = ~n6639 ;
  assign y2909 = n6640 ;
  assign y2910 = ~n6641 ;
  assign y2911 = n6650 ;
  assign y2912 = ~n6652 ;
  assign y2913 = n6658 ;
  assign y2914 = n6659 ;
  assign y2915 = ~1'b0 ;
  assign y2916 = ~1'b0 ;
  assign y2917 = n6660 ;
  assign y2918 = ~1'b0 ;
  assign y2919 = ~n5854 ;
  assign y2920 = n6661 ;
  assign y2921 = ~1'b0 ;
  assign y2922 = n6662 ;
  assign y2923 = n6666 ;
  assign y2924 = ~n6667 ;
  assign y2925 = ~1'b0 ;
  assign y2926 = ~1'b0 ;
  assign y2927 = n6670 ;
  assign y2928 = n6671 ;
  assign y2929 = ~1'b0 ;
  assign y2930 = n6673 ;
  assign y2931 = ~n6676 ;
  assign y2932 = ~n6681 ;
  assign y2933 = n6683 ;
  assign y2934 = ~n6686 ;
  assign y2935 = ~n6687 ;
  assign y2936 = ~n6690 ;
  assign y2937 = ~n6695 ;
  assign y2938 = ~n6702 ;
  assign y2939 = ~1'b0 ;
  assign y2940 = n6703 ;
  assign y2941 = ~1'b0 ;
  assign y2942 = ~n6707 ;
  assign y2943 = n6709 ;
  assign y2944 = n6710 ;
  assign y2945 = ~n6716 ;
  assign y2946 = ~n6722 ;
  assign y2947 = ~n6723 ;
  assign y2948 = n1064 ;
  assign y2949 = ~1'b0 ;
  assign y2950 = n6725 ;
  assign y2951 = ~n6729 ;
  assign y2952 = ~1'b0 ;
  assign y2953 = ~n6731 ;
  assign y2954 = n6732 ;
  assign y2955 = ~1'b0 ;
  assign y2956 = n6739 ;
  assign y2957 = n6746 ;
  assign y2958 = ~n6747 ;
  assign y2959 = ~1'b0 ;
  assign y2960 = ~n6748 ;
  assign y2961 = ~n6754 ;
  assign y2962 = n6766 ;
  assign y2963 = n6767 ;
  assign y2964 = ~n54 ;
  assign y2965 = ~n6768 ;
  assign y2966 = ~1'b0 ;
  assign y2967 = ~n6771 ;
  assign y2968 = 1'b0 ;
  assign y2969 = n6776 ;
  assign y2970 = ~n6779 ;
  assign y2971 = n6781 ;
  assign y2972 = n6784 ;
  assign y2973 = ~n6787 ;
  assign y2974 = n6792 ;
  assign y2975 = ~n6796 ;
  assign y2976 = n6801 ;
  assign y2977 = n6806 ;
  assign y2978 = ~n6819 ;
  assign y2979 = n6820 ;
  assign y2980 = ~1'b0 ;
  assign y2981 = n6821 ;
  assign y2982 = ~n6823 ;
  assign y2983 = n6829 ;
  assign y2984 = ~n6831 ;
  assign y2985 = n6839 ;
  assign y2986 = n4599 ;
  assign y2987 = ~n6841 ;
  assign y2988 = ~n6844 ;
  assign y2989 = n6846 ;
  assign y2990 = n6848 ;
  assign y2991 = ~n6849 ;
  assign y2992 = n6851 ;
  assign y2993 = ~1'b0 ;
  assign y2994 = ~1'b0 ;
  assign y2995 = ~n6852 ;
  assign y2996 = n6853 ;
  assign y2997 = ~n6858 ;
  assign y2998 = n6865 ;
  assign y2999 = ~n6872 ;
  assign y3000 = ~n6873 ;
  assign y3001 = n6874 ;
  assign y3002 = ~n6878 ;
  assign y3003 = ~n6882 ;
  assign y3004 = ~1'b0 ;
  assign y3005 = ~n6883 ;
  assign y3006 = ~1'b0 ;
  assign y3007 = n6885 ;
  assign y3008 = ~n6042 ;
  assign y3009 = ~1'b0 ;
  assign y3010 = ~n6886 ;
  assign y3011 = n6888 ;
  assign y3012 = n6889 ;
  assign y3013 = n6893 ;
  assign y3014 = ~1'b0 ;
  assign y3015 = n6898 ;
  assign y3016 = n6901 ;
  assign y3017 = ~n6902 ;
  assign y3018 = n6903 ;
  assign y3019 = n6906 ;
  assign y3020 = ~1'b0 ;
  assign y3021 = n6910 ;
  assign y3022 = n1105 ;
  assign y3023 = ~n6915 ;
  assign y3024 = n6916 ;
  assign y3025 = ~n6922 ;
  assign y3026 = ~n6923 ;
  assign y3027 = n6924 ;
  assign y3028 = n6925 ;
  assign y3029 = n6938 ;
  assign y3030 = ~1'b0 ;
  assign y3031 = n6941 ;
  assign y3032 = ~n6942 ;
  assign y3033 = ~1'b0 ;
  assign y3034 = ~1'b0 ;
  assign y3035 = n2859 ;
  assign y3036 = ~n6945 ;
  assign y3037 = n6948 ;
  assign y3038 = ~n6954 ;
  assign y3039 = ~1'b0 ;
  assign y3040 = ~1'b0 ;
  assign y3041 = ~n6955 ;
  assign y3042 = n6958 ;
  assign y3043 = ~n285 ;
  assign y3044 = n6962 ;
  assign y3045 = ~n6965 ;
  assign y3046 = n6968 ;
  assign y3047 = ~n6969 ;
  assign y3048 = ~n6973 ;
  assign y3049 = n6977 ;
  assign y3050 = n6978 ;
  assign y3051 = ~n6979 ;
  assign y3052 = ~1'b0 ;
  assign y3053 = ~1'b0 ;
  assign y3054 = n6981 ;
  assign y3055 = n6988 ;
  assign y3056 = ~1'b0 ;
  assign y3057 = ~n6992 ;
  assign y3058 = ~n7000 ;
  assign y3059 = ~1'b0 ;
  assign y3060 = ~1'b0 ;
  assign y3061 = n7005 ;
  assign y3062 = ~1'b0 ;
  assign y3063 = ~1'b0 ;
  assign y3064 = ~n7008 ;
  assign y3065 = n7010 ;
  assign y3066 = n7014 ;
  assign y3067 = ~1'b0 ;
  assign y3068 = n5722 ;
  assign y3069 = ~n7021 ;
  assign y3070 = n7023 ;
  assign y3071 = ~1'b0 ;
  assign y3072 = ~n7033 ;
  assign y3073 = n7035 ;
  assign y3074 = ~n7039 ;
  assign y3075 = ~n7040 ;
  assign y3076 = n7041 ;
  assign y3077 = ~1'b0 ;
  assign y3078 = ~1'b0 ;
  assign y3079 = ~1'b0 ;
  assign y3080 = ~1'b0 ;
  assign y3081 = n7043 ;
  assign y3082 = ~n7046 ;
  assign y3083 = n7047 ;
  assign y3084 = ~1'b0 ;
  assign y3085 = n7054 ;
  assign y3086 = ~n7056 ;
  assign y3087 = ~1'b0 ;
  assign y3088 = 1'b0 ;
  assign y3089 = ~1'b0 ;
  assign y3090 = n7060 ;
  assign y3091 = ~n7064 ;
  assign y3092 = ~n7067 ;
  assign y3093 = n7072 ;
  assign y3094 = ~n7074 ;
  assign y3095 = n7076 ;
  assign y3096 = n3679 ;
  assign y3097 = n7077 ;
  assign y3098 = n7078 ;
  assign y3099 = n7080 ;
  assign y3100 = n5533 ;
  assign y3101 = ~n7086 ;
  assign y3102 = ~n3245 ;
  assign y3103 = ~1'b0 ;
  assign y3104 = ~1'b0 ;
  assign y3105 = n7091 ;
  assign y3106 = ~n7098 ;
  assign y3107 = ~1'b0 ;
  assign y3108 = ~n7102 ;
  assign y3109 = ~1'b0 ;
  assign y3110 = ~1'b0 ;
  assign y3111 = ~n7103 ;
  assign y3112 = n7114 ;
  assign y3113 = ~1'b0 ;
  assign y3114 = ~n7118 ;
  assign y3115 = ~n1835 ;
  assign y3116 = n7119 ;
  assign y3117 = ~1'b0 ;
  assign y3118 = n7120 ;
  assign y3119 = n7125 ;
  assign y3120 = n7134 ;
  assign y3121 = ~n7135 ;
  assign y3122 = n7138 ;
  assign y3123 = ~1'b0 ;
  assign y3124 = ~n7140 ;
  assign y3125 = n7142 ;
  assign y3126 = ~n7146 ;
  assign y3127 = ~1'b0 ;
  assign y3128 = ~1'b0 ;
  assign y3129 = ~n7149 ;
  assign y3130 = 1'b0 ;
  assign y3131 = n7150 ;
  assign y3132 = ~n7158 ;
  assign y3133 = ~n3626 ;
  assign y3134 = ~n7161 ;
  assign y3135 = ~1'b0 ;
  assign y3136 = ~n7165 ;
  assign y3137 = ~n7167 ;
  assign y3138 = ~1'b0 ;
  assign y3139 = ~1'b0 ;
  assign y3140 = ~1'b0 ;
  assign y3141 = ~n7174 ;
  assign y3142 = n7180 ;
  assign y3143 = ~n7182 ;
  assign y3144 = ~n7185 ;
  assign y3145 = ~n7188 ;
  assign y3146 = ~1'b0 ;
  assign y3147 = ~n7189 ;
  assign y3148 = n7193 ;
  assign y3149 = ~n7194 ;
  assign y3150 = ~n7195 ;
  assign y3151 = ~1'b0 ;
  assign y3152 = n7196 ;
  assign y3153 = ~n7208 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = n7213 ;
  assign y3156 = ~n7214 ;
  assign y3157 = ~1'b0 ;
  assign y3158 = n7216 ;
  assign y3159 = n7218 ;
  assign y3160 = ~n7219 ;
  assign y3161 = ~n7221 ;
  assign y3162 = ~n7223 ;
  assign y3163 = ~1'b0 ;
  assign y3164 = n7225 ;
  assign y3165 = ~1'b0 ;
  assign y3166 = ~1'b0 ;
  assign y3167 = n7226 ;
  assign y3168 = n1616 ;
  assign y3169 = ~1'b0 ;
  assign y3170 = ~n7230 ;
  assign y3171 = ~1'b0 ;
  assign y3172 = n7231 ;
  assign y3173 = ~1'b0 ;
  assign y3174 = ~1'b0 ;
  assign y3175 = ~1'b0 ;
  assign y3176 = n7235 ;
  assign y3177 = n7239 ;
  assign y3178 = ~1'b0 ;
  assign y3179 = ~1'b0 ;
  assign y3180 = n7243 ;
  assign y3181 = ~1'b0 ;
  assign y3182 = ~n7250 ;
  assign y3183 = ~n7251 ;
  assign y3184 = n7252 ;
  assign y3185 = ~n7253 ;
  assign y3186 = ~1'b0 ;
  assign y3187 = ~1'b0 ;
  assign y3188 = ~1'b0 ;
  assign y3189 = ~1'b0 ;
  assign y3190 = n7255 ;
  assign y3191 = ~n7259 ;
  assign y3192 = ~1'b0 ;
  assign y3193 = n7260 ;
  assign y3194 = n3248 ;
  assign y3195 = ~1'b0 ;
  assign y3196 = n7264 ;
  assign y3197 = ~n7267 ;
  assign y3198 = ~n7268 ;
  assign y3199 = n7269 ;
  assign y3200 = 1'b0 ;
  assign y3201 = ~n7271 ;
  assign y3202 = n4002 ;
  assign y3203 = ~n7278 ;
  assign y3204 = ~1'b0 ;
  assign y3205 = n7280 ;
  assign y3206 = ~1'b0 ;
  assign y3207 = n7288 ;
  assign y3208 = ~n7292 ;
  assign y3209 = n7293 ;
  assign y3210 = ~n7295 ;
  assign y3211 = ~1'b0 ;
  assign y3212 = n5997 ;
  assign y3213 = ~n7296 ;
  assign y3214 = ~1'b0 ;
  assign y3215 = n7297 ;
  assign y3216 = ~n6699 ;
  assign y3217 = n7298 ;
  assign y3218 = ~n7302 ;
  assign y3219 = n7303 ;
  assign y3220 = n7307 ;
  assign y3221 = ~1'b0 ;
  assign y3222 = n7314 ;
  assign y3223 = ~n7318 ;
  assign y3224 = ~1'b0 ;
  assign y3225 = n7324 ;
  assign y3226 = n7328 ;
  assign y3227 = ~n7330 ;
  assign y3228 = n7334 ;
  assign y3229 = ~n7345 ;
  assign y3230 = n7349 ;
  assign y3231 = n7350 ;
  assign y3232 = n7370 ;
  assign y3233 = ~1'b0 ;
  assign y3234 = ~n5022 ;
  assign y3235 = n7371 ;
  assign y3236 = ~n7376 ;
  assign y3237 = ~n7377 ;
  assign y3238 = ~1'b0 ;
  assign y3239 = n7380 ;
  assign y3240 = ~n7386 ;
  assign y3241 = ~n7388 ;
  assign y3242 = ~1'b0 ;
  assign y3243 = ~n7391 ;
  assign y3244 = n7397 ;
  assign y3245 = ~n6253 ;
  assign y3246 = ~1'b0 ;
  assign y3247 = n7401 ;
  assign y3248 = ~n7404 ;
  assign y3249 = n7414 ;
  assign y3250 = n7417 ;
  assign y3251 = ~1'b0 ;
  assign y3252 = n7419 ;
  assign y3253 = ~n7423 ;
  assign y3254 = n7426 ;
  assign y3255 = ~1'b0 ;
  assign y3256 = n7427 ;
  assign y3257 = n7428 ;
  assign y3258 = n7430 ;
  assign y3259 = ~1'b0 ;
  assign y3260 = ~n7432 ;
  assign y3261 = ~n7433 ;
  assign y3262 = n7436 ;
  assign y3263 = n7438 ;
  assign y3264 = ~n7446 ;
  assign y3265 = ~n7447 ;
  assign y3266 = n7451 ;
  assign y3267 = ~n7459 ;
  assign y3268 = ~n7464 ;
  assign y3269 = ~n7465 ;
  assign y3270 = n7469 ;
  assign y3271 = ~n7470 ;
  assign y3272 = ~1'b0 ;
  assign y3273 = ~n7475 ;
  assign y3274 = n7478 ;
  assign y3275 = ~n7483 ;
  assign y3276 = ~n7484 ;
  assign y3277 = n7487 ;
  assign y3278 = n7488 ;
  assign y3279 = ~n7493 ;
  assign y3280 = ~n7495 ;
  assign y3281 = n4992 ;
  assign y3282 = ~1'b0 ;
  assign y3283 = ~n7498 ;
  assign y3284 = 1'b0 ;
  assign y3285 = ~n7499 ;
  assign y3286 = n7505 ;
  assign y3287 = ~n7506 ;
  assign y3288 = ~n7508 ;
  assign y3289 = ~1'b0 ;
  assign y3290 = ~n7512 ;
  assign y3291 = n7514 ;
  assign y3292 = ~n7520 ;
  assign y3293 = n7525 ;
  assign y3294 = n7526 ;
  assign y3295 = ~1'b0 ;
  assign y3296 = n7527 ;
  assign y3297 = ~n6010 ;
  assign y3298 = ~1'b0 ;
  assign y3299 = n7530 ;
  assign y3300 = ~n7531 ;
  assign y3301 = ~1'b0 ;
  assign y3302 = ~n7534 ;
  assign y3303 = n2678 ;
  assign y3304 = n7540 ;
  assign y3305 = ~1'b0 ;
  assign y3306 = ~1'b0 ;
  assign y3307 = n7543 ;
  assign y3308 = n7544 ;
  assign y3309 = n7550 ;
  assign y3310 = ~n7551 ;
  assign y3311 = ~n7554 ;
  assign y3312 = ~1'b0 ;
  assign y3313 = ~n7556 ;
  assign y3314 = ~n5329 ;
  assign y3315 = n7561 ;
  assign y3316 = n7563 ;
  assign y3317 = ~n7568 ;
  assign y3318 = ~1'b0 ;
  assign y3319 = n7569 ;
  assign y3320 = ~n7572 ;
  assign y3321 = ~n7574 ;
  assign y3322 = ~1'b0 ;
  assign y3323 = ~n7586 ;
  assign y3324 = ~n7588 ;
  assign y3325 = ~1'b0 ;
  assign y3326 = ~1'b0 ;
  assign y3327 = ~1'b0 ;
  assign y3328 = ~1'b0 ;
  assign y3329 = n7590 ;
  assign y3330 = n7594 ;
  assign y3331 = n7605 ;
  assign y3332 = ~n7610 ;
  assign y3333 = ~n7612 ;
  assign y3334 = n7613 ;
  assign y3335 = ~n7614 ;
  assign y3336 = n7617 ;
  assign y3337 = n7620 ;
  assign y3338 = ~1'b0 ;
  assign y3339 = n7626 ;
  assign y3340 = ~1'b0 ;
  assign y3341 = ~n7627 ;
  assign y3342 = n3195 ;
  assign y3343 = 1'b0 ;
  assign y3344 = 1'b0 ;
  assign y3345 = n7629 ;
  assign y3346 = ~1'b0 ;
  assign y3347 = ~1'b0 ;
  assign y3348 = n7630 ;
  assign y3349 = ~n7631 ;
  assign y3350 = ~1'b0 ;
  assign y3351 = n7633 ;
  assign y3352 = n7635 ;
  assign y3353 = n7639 ;
  assign y3354 = n7644 ;
  assign y3355 = ~n7652 ;
  assign y3356 = n7653 ;
  assign y3357 = n7654 ;
  assign y3358 = ~n7656 ;
  assign y3359 = ~n7659 ;
  assign y3360 = ~n7661 ;
  assign y3361 = n7674 ;
  assign y3362 = ~n7676 ;
  assign y3363 = n7682 ;
  assign y3364 = n4212 ;
  assign y3365 = ~1'b0 ;
  assign y3366 = ~n7686 ;
  assign y3367 = ~n7687 ;
  assign y3368 = ~1'b0 ;
  assign y3369 = ~1'b0 ;
  assign y3370 = n7690 ;
  assign y3371 = n6229 ;
  assign y3372 = ~n7697 ;
  assign y3373 = n7704 ;
  assign y3374 = n7705 ;
  assign y3375 = ~n7715 ;
  assign y3376 = ~n7717 ;
  assign y3377 = ~n7718 ;
  assign y3378 = ~n7722 ;
  assign y3379 = 1'b0 ;
  assign y3380 = ~n7726 ;
  assign y3381 = n7728 ;
  assign y3382 = ~n7730 ;
  assign y3383 = ~n7734 ;
  assign y3384 = n3313 ;
  assign y3385 = ~n7735 ;
  assign y3386 = ~n7737 ;
  assign y3387 = ~n7741 ;
  assign y3388 = n7746 ;
  assign y3389 = n7754 ;
  assign y3390 = ~n7755 ;
  assign y3391 = ~n3460 ;
  assign y3392 = ~n7757 ;
  assign y3393 = ~1'b0 ;
  assign y3394 = n7759 ;
  assign y3395 = n7760 ;
  assign y3396 = ~1'b0 ;
  assign y3397 = ~1'b0 ;
  assign y3398 = ~1'b0 ;
  assign y3399 = n7766 ;
  assign y3400 = n7767 ;
  assign y3401 = ~1'b0 ;
  assign y3402 = n7773 ;
  assign y3403 = n7775 ;
  assign y3404 = n7776 ;
  assign y3405 = ~1'b0 ;
  assign y3406 = ~n7782 ;
  assign y3407 = ~1'b0 ;
  assign y3408 = ~n7785 ;
  assign y3409 = n7787 ;
  assign y3410 = ~1'b0 ;
  assign y3411 = n7791 ;
  assign y3412 = n7795 ;
  assign y3413 = ~1'b0 ;
  assign y3414 = ~1'b0 ;
  assign y3415 = ~n7799 ;
  assign y3416 = n7801 ;
  assign y3417 = ~1'b0 ;
  assign y3418 = ~n1787 ;
  assign y3419 = ~1'b0 ;
  assign y3420 = ~n7802 ;
  assign y3421 = ~n7810 ;
  assign y3422 = ~n7812 ;
  assign y3423 = n7815 ;
  assign y3424 = ~1'b0 ;
  assign y3425 = ~1'b0 ;
  assign y3426 = n7822 ;
  assign y3427 = n7823 ;
  assign y3428 = ~1'b0 ;
  assign y3429 = ~1'b0 ;
  assign y3430 = ~n7825 ;
  assign y3431 = ~n7830 ;
  assign y3432 = ~1'b0 ;
  assign y3433 = ~1'b0 ;
  assign y3434 = n4093 ;
  assign y3435 = n7832 ;
  assign y3436 = n7834 ;
  assign y3437 = ~n7846 ;
  assign y3438 = n7848 ;
  assign y3439 = n7851 ;
  assign y3440 = n7856 ;
  assign y3441 = ~1'b0 ;
  assign y3442 = ~n7859 ;
  assign y3443 = ~1'b0 ;
  assign y3444 = ~n7863 ;
  assign y3445 = n7866 ;
  assign y3446 = n7867 ;
  assign y3447 = ~n7869 ;
  assign y3448 = ~1'b0 ;
  assign y3449 = n7874 ;
  assign y3450 = n7875 ;
  assign y3451 = ~1'b0 ;
  assign y3452 = ~n7878 ;
  assign y3453 = ~1'b0 ;
  assign y3454 = ~1'b0 ;
  assign y3455 = n7881 ;
  assign y3456 = ~n7882 ;
  assign y3457 = 1'b0 ;
  assign y3458 = n7885 ;
  assign y3459 = ~1'b0 ;
  assign y3460 = ~n7888 ;
  assign y3461 = n7891 ;
  assign y3462 = n7892 ;
  assign y3463 = ~1'b0 ;
  assign y3464 = ~n1435 ;
  assign y3465 = ~1'b0 ;
  assign y3466 = n7896 ;
  assign y3467 = ~1'b0 ;
  assign y3468 = ~n7904 ;
  assign y3469 = ~n7906 ;
  assign y3470 = ~1'b0 ;
  assign y3471 = n7907 ;
  assign y3472 = n7912 ;
  assign y3473 = ~n7916 ;
  assign y3474 = n7923 ;
  assign y3475 = ~n5301 ;
  assign y3476 = ~n7927 ;
  assign y3477 = ~n7930 ;
  assign y3478 = ~n7931 ;
  assign y3479 = n7932 ;
  assign y3480 = n7933 ;
  assign y3481 = ~n7938 ;
  assign y3482 = ~1'b0 ;
  assign y3483 = ~n7939 ;
  assign y3484 = ~n7941 ;
  assign y3485 = n7943 ;
  assign y3486 = n7944 ;
  assign y3487 = ~n7945 ;
  assign y3488 = ~n7947 ;
  assign y3489 = n7949 ;
  assign y3490 = n7952 ;
  assign y3491 = n6485 ;
  assign y3492 = n7954 ;
  assign y3493 = n5683 ;
  assign y3494 = n7970 ;
  assign y3495 = n7974 ;
  assign y3496 = n7975 ;
  assign y3497 = n7976 ;
  assign y3498 = 1'b0 ;
  assign y3499 = ~n398 ;
  assign y3500 = n7978 ;
  assign y3501 = ~n7980 ;
  assign y3502 = n7982 ;
  assign y3503 = ~n7987 ;
  assign y3504 = n7994 ;
  assign y3505 = ~n7997 ;
  assign y3506 = ~n8001 ;
  assign y3507 = ~n4285 ;
  assign y3508 = ~n8010 ;
  assign y3509 = ~n8015 ;
  assign y3510 = ~1'b0 ;
  assign y3511 = ~n8016 ;
  assign y3512 = ~n8018 ;
  assign y3513 = n8021 ;
  assign y3514 = n8023 ;
  assign y3515 = ~n8027 ;
  assign y3516 = ~1'b0 ;
  assign y3517 = n8028 ;
  assign y3518 = ~n6607 ;
  assign y3519 = n8029 ;
  assign y3520 = n8031 ;
  assign y3521 = ~n8033 ;
  assign y3522 = ~n1026 ;
  assign y3523 = n8034 ;
  assign y3524 = ~n8045 ;
  assign y3525 = ~n8054 ;
  assign y3526 = n8055 ;
  assign y3527 = ~n7535 ;
  assign y3528 = n8056 ;
  assign y3529 = ~1'b0 ;
  assign y3530 = ~1'b0 ;
  assign y3531 = ~1'b0 ;
  assign y3532 = n8058 ;
  assign y3533 = ~n8065 ;
  assign y3534 = n8067 ;
  assign y3535 = 1'b0 ;
  assign y3536 = ~n8071 ;
  assign y3537 = ~1'b0 ;
  assign y3538 = n8076 ;
  assign y3539 = n8079 ;
  assign y3540 = n8080 ;
  assign y3541 = ~n8082 ;
  assign y3542 = 1'b0 ;
  assign y3543 = ~1'b0 ;
  assign y3544 = ~1'b0 ;
  assign y3545 = n8083 ;
  assign y3546 = ~n8084 ;
  assign y3547 = ~n8085 ;
  assign y3548 = n8086 ;
  assign y3549 = n8088 ;
  assign y3550 = ~n8089 ;
  assign y3551 = ~n8090 ;
  assign y3552 = ~1'b0 ;
  assign y3553 = ~1'b0 ;
  assign y3554 = ~n879 ;
  assign y3555 = 1'b0 ;
  assign y3556 = n8093 ;
  assign y3557 = ~1'b0 ;
  assign y3558 = n8094 ;
  assign y3559 = n8095 ;
  assign y3560 = 1'b0 ;
  assign y3561 = n8098 ;
  assign y3562 = ~n8103 ;
  assign y3563 = ~n8108 ;
  assign y3564 = ~n8109 ;
  assign y3565 = n8112 ;
  assign y3566 = 1'b0 ;
  assign y3567 = ~n8113 ;
  assign y3568 = n8120 ;
  assign y3569 = ~n8122 ;
  assign y3570 = ~n469 ;
  assign y3571 = ~n8123 ;
  assign y3572 = ~n4216 ;
  assign y3573 = ~1'b0 ;
  assign y3574 = n8125 ;
  assign y3575 = ~n8126 ;
  assign y3576 = ~n8128 ;
  assign y3577 = ~n8134 ;
  assign y3578 = ~1'b0 ;
  assign y3579 = ~n8135 ;
  assign y3580 = ~n8137 ;
  assign y3581 = ~n8138 ;
  assign y3582 = ~n8140 ;
  assign y3583 = ~n8147 ;
  assign y3584 = n8149 ;
  assign y3585 = n8153 ;
  assign y3586 = ~n8158 ;
  assign y3587 = n8162 ;
  assign y3588 = ~n8166 ;
  assign y3589 = n8167 ;
  assign y3590 = n8172 ;
  assign y3591 = n8173 ;
  assign y3592 = n8175 ;
  assign y3593 = n8176 ;
  assign y3594 = ~n8181 ;
  assign y3595 = ~1'b0 ;
  assign y3596 = n2196 ;
  assign y3597 = ~1'b0 ;
  assign y3598 = n8182 ;
  assign y3599 = n8184 ;
  assign y3600 = 1'b0 ;
  assign y3601 = n8185 ;
  assign y3602 = n8187 ;
  assign y3603 = n8191 ;
  assign y3604 = ~n8197 ;
  assign y3605 = ~1'b0 ;
  assign y3606 = ~n8201 ;
  assign y3607 = n8204 ;
  assign y3608 = ~n8205 ;
  assign y3609 = n8208 ;
  assign y3610 = ~n8211 ;
  assign y3611 = n8212 ;
  assign y3612 = ~n8214 ;
  assign y3613 = n8216 ;
  assign y3614 = n8225 ;
  assign y3615 = n8226 ;
  assign y3616 = n4055 ;
  assign y3617 = ~n8228 ;
  assign y3618 = n8231 ;
  assign y3619 = n8236 ;
  assign y3620 = n8239 ;
  assign y3621 = n8241 ;
  assign y3622 = ~1'b0 ;
  assign y3623 = n8242 ;
  assign y3624 = ~n8244 ;
  assign y3625 = ~1'b0 ;
  assign y3626 = n8245 ;
  assign y3627 = n8247 ;
  assign y3628 = ~1'b0 ;
  assign y3629 = ~1'b0 ;
  assign y3630 = ~n8248 ;
  assign y3631 = n8254 ;
  assign y3632 = n8258 ;
  assign y3633 = ~n8262 ;
  assign y3634 = ~1'b0 ;
  assign y3635 = ~n8266 ;
  assign y3636 = ~1'b0 ;
  assign y3637 = n8268 ;
  assign y3638 = ~n8269 ;
  assign y3639 = n8271 ;
  assign y3640 = ~1'b0 ;
  assign y3641 = ~n8275 ;
  assign y3642 = ~1'b0 ;
  assign y3643 = ~n8277 ;
  assign y3644 = n8279 ;
  assign y3645 = n8281 ;
  assign y3646 = n8284 ;
  assign y3647 = ~n8291 ;
  assign y3648 = ~1'b0 ;
  assign y3649 = ~1'b0 ;
  assign y3650 = n8298 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = ~1'b0 ;
  assign y3653 = ~1'b0 ;
  assign y3654 = ~n8306 ;
  assign y3655 = n8308 ;
  assign y3656 = n8310 ;
  assign y3657 = ~1'b0 ;
  assign y3658 = ~n8311 ;
  assign y3659 = ~n8312 ;
  assign y3660 = ~1'b0 ;
  assign y3661 = n8314 ;
  assign y3662 = n865 ;
  assign y3663 = n4014 ;
  assign y3664 = n8316 ;
  assign y3665 = ~n8318 ;
  assign y3666 = n8327 ;
  assign y3667 = ~n8330 ;
  assign y3668 = ~1'b0 ;
  assign y3669 = n8331 ;
  assign y3670 = n8333 ;
  assign y3671 = ~n8334 ;
  assign y3672 = n8337 ;
  assign y3673 = n8343 ;
  assign y3674 = ~n8348 ;
  assign y3675 = n8353 ;
  assign y3676 = ~1'b0 ;
  assign y3677 = ~1'b0 ;
  assign y3678 = n8354 ;
  assign y3679 = ~n5876 ;
  assign y3680 = ~1'b0 ;
  assign y3681 = ~1'b0 ;
  assign y3682 = ~n8356 ;
  assign y3683 = ~1'b0 ;
  assign y3684 = ~n8357 ;
  assign y3685 = ~n8361 ;
  assign y3686 = ~n8364 ;
  assign y3687 = n8367 ;
  assign y3688 = n8369 ;
  assign y3689 = ~n8374 ;
  assign y3690 = ~1'b0 ;
  assign y3691 = ~n8378 ;
  assign y3692 = n8385 ;
  assign y3693 = n8387 ;
  assign y3694 = ~1'b0 ;
  assign y3695 = ~n8392 ;
  assign y3696 = ~n8395 ;
  assign y3697 = ~n8401 ;
  assign y3698 = ~1'b0 ;
  assign y3699 = ~1'b0 ;
  assign y3700 = ~n3039 ;
  assign y3701 = n8403 ;
  assign y3702 = n8413 ;
  assign y3703 = ~n8416 ;
  assign y3704 = ~n8421 ;
  assign y3705 = n8427 ;
  assign y3706 = ~n8429 ;
  assign y3707 = ~n8431 ;
  assign y3708 = ~n8434 ;
  assign y3709 = ~1'b0 ;
  assign y3710 = ~1'b0 ;
  assign y3711 = ~1'b0 ;
  assign y3712 = ~1'b0 ;
  assign y3713 = ~1'b0 ;
  assign y3714 = ~1'b0 ;
  assign y3715 = n694 ;
  assign y3716 = ~1'b0 ;
  assign y3717 = ~n8435 ;
  assign y3718 = ~1'b0 ;
  assign y3719 = ~1'b0 ;
  assign y3720 = n8438 ;
  assign y3721 = ~1'b0 ;
  assign y3722 = ~n8442 ;
  assign y3723 = ~n8450 ;
  assign y3724 = ~n8451 ;
  assign y3725 = ~1'b0 ;
  assign y3726 = ~1'b0 ;
  assign y3727 = ~1'b0 ;
  assign y3728 = ~n8455 ;
  assign y3729 = n8457 ;
  assign y3730 = n8460 ;
  assign y3731 = ~n8465 ;
  assign y3732 = ~n8472 ;
  assign y3733 = n8483 ;
  assign y3734 = n8496 ;
  assign y3735 = n8508 ;
  assign y3736 = ~1'b0 ;
  assign y3737 = ~n8509 ;
  assign y3738 = ~n8514 ;
  assign y3739 = ~n8519 ;
  assign y3740 = ~1'b0 ;
  assign y3741 = ~1'b0 ;
  assign y3742 = ~1'b0 ;
  assign y3743 = n1272 ;
  assign y3744 = ~n8522 ;
  assign y3745 = n8523 ;
  assign y3746 = n8524 ;
  assign y3747 = n8526 ;
  assign y3748 = ~n8528 ;
  assign y3749 = n8536 ;
  assign y3750 = n8537 ;
  assign y3751 = ~n8541 ;
  assign y3752 = n8544 ;
  assign y3753 = ~n8547 ;
  assign y3754 = n8549 ;
  assign y3755 = n8551 ;
  assign y3756 = n1400 ;
  assign y3757 = ~n8554 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = n8556 ;
  assign y3760 = ~n8557 ;
  assign y3761 = ~1'b0 ;
  assign y3762 = ~n8562 ;
  assign y3763 = ~n8565 ;
  assign y3764 = n8571 ;
  assign y3765 = ~1'b0 ;
  assign y3766 = ~n8574 ;
  assign y3767 = n8575 ;
  assign y3768 = ~n8577 ;
  assign y3769 = ~n8581 ;
  assign y3770 = n8586 ;
  assign y3771 = n8590 ;
  assign y3772 = n8592 ;
  assign y3773 = ~n8600 ;
  assign y3774 = n8601 ;
  assign y3775 = n8605 ;
  assign y3776 = n8606 ;
  assign y3777 = ~n8612 ;
  assign y3778 = n8615 ;
  assign y3779 = ~n8616 ;
  assign y3780 = ~n8628 ;
  assign y3781 = ~n8629 ;
  assign y3782 = ~1'b0 ;
  assign y3783 = ~n8635 ;
  assign y3784 = ~1'b0 ;
  assign y3785 = n8636 ;
  assign y3786 = ~n8639 ;
  assign y3787 = ~n8654 ;
  assign y3788 = ~1'b0 ;
  assign y3789 = ~1'b0 ;
  assign y3790 = ~n8656 ;
  assign y3791 = n8660 ;
  assign y3792 = n8661 ;
  assign y3793 = ~n7468 ;
  assign y3794 = n8662 ;
  assign y3795 = ~1'b0 ;
  assign y3796 = n8663 ;
  assign y3797 = n8671 ;
  assign y3798 = ~n8672 ;
  assign y3799 = n8673 ;
  assign y3800 = n8674 ;
  assign y3801 = ~n8678 ;
  assign y3802 = ~1'b0 ;
  assign y3803 = ~1'b0 ;
  assign y3804 = ~1'b0 ;
  assign y3805 = ~n8681 ;
  assign y3806 = ~1'b0 ;
  assign y3807 = ~n8682 ;
  assign y3808 = ~n7505 ;
  assign y3809 = n8684 ;
  assign y3810 = ~n8691 ;
  assign y3811 = n8696 ;
  assign y3812 = ~n23 ;
  assign y3813 = n8701 ;
  assign y3814 = n8704 ;
  assign y3815 = ~n8712 ;
  assign y3816 = ~n8717 ;
  assign y3817 = n8719 ;
  assign y3818 = ~n8724 ;
  assign y3819 = ~1'b0 ;
  assign y3820 = ~n8725 ;
  assign y3821 = n8727 ;
  assign y3822 = ~1'b0 ;
  assign y3823 = n8728 ;
  assign y3824 = n8743 ;
  assign y3825 = ~n8745 ;
  assign y3826 = ~1'b0 ;
  assign y3827 = ~n8747 ;
  assign y3828 = 1'b0 ;
  assign y3829 = n8758 ;
  assign y3830 = ~n8763 ;
  assign y3831 = ~n8764 ;
  assign y3832 = n8765 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = n8769 ;
  assign y3835 = ~1'b0 ;
  assign y3836 = ~n8772 ;
  assign y3837 = ~n8774 ;
  assign y3838 = n8775 ;
  assign y3839 = ~n2418 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = ~n8777 ;
  assign y3842 = ~n7240 ;
  assign y3843 = ~n8783 ;
  assign y3844 = n8787 ;
  assign y3845 = n8795 ;
  assign y3846 = n8797 ;
  assign y3847 = ~1'b0 ;
  assign y3848 = n8798 ;
  assign y3849 = n8800 ;
  assign y3850 = ~1'b0 ;
  assign y3851 = ~n8807 ;
  assign y3852 = ~n8810 ;
  assign y3853 = ~n8812 ;
  assign y3854 = ~1'b0 ;
  assign y3855 = ~n8813 ;
  assign y3856 = ~n8820 ;
  assign y3857 = ~n8821 ;
  assign y3858 = ~n8822 ;
  assign y3859 = ~1'b0 ;
  assign y3860 = ~n8824 ;
  assign y3861 = ~n8826 ;
  assign y3862 = n8828 ;
  assign y3863 = n8835 ;
  assign y3864 = n8845 ;
  assign y3865 = ~n8850 ;
  assign y3866 = ~n8852 ;
  assign y3867 = n8859 ;
  assign y3868 = n8860 ;
  assign y3869 = n8861 ;
  assign y3870 = n8866 ;
  assign y3871 = ~1'b0 ;
  assign y3872 = ~n6167 ;
  assign y3873 = ~n8868 ;
  assign y3874 = n8872 ;
  assign y3875 = n8876 ;
  assign y3876 = ~1'b0 ;
  assign y3877 = n8877 ;
  assign y3878 = ~n8878 ;
  assign y3879 = ~1'b0 ;
  assign y3880 = ~1'b0 ;
  assign y3881 = ~n8881 ;
  assign y3882 = n8884 ;
  assign y3883 = ~n8885 ;
  assign y3884 = ~1'b0 ;
  assign y3885 = ~n8888 ;
  assign y3886 = ~1'b0 ;
  assign y3887 = ~1'b0 ;
  assign y3888 = ~1'b0 ;
  assign y3889 = n1932 ;
  assign y3890 = n8890 ;
  assign y3891 = n184 ;
  assign y3892 = ~n8893 ;
  assign y3893 = ~n8895 ;
  assign y3894 = ~n8902 ;
  assign y3895 = n8909 ;
  assign y3896 = n4548 ;
  assign y3897 = ~n8910 ;
  assign y3898 = ~n8913 ;
  assign y3899 = n8921 ;
  assign y3900 = ~n8923 ;
  assign y3901 = n8925 ;
  assign y3902 = ~n8926 ;
  assign y3903 = ~n6711 ;
  assign y3904 = n8927 ;
  assign y3905 = ~n8931 ;
  assign y3906 = ~n8933 ;
  assign y3907 = n8936 ;
  assign y3908 = ~n8937 ;
  assign y3909 = n8703 ;
  assign y3910 = n8939 ;
  assign y3911 = ~n8945 ;
  assign y3912 = ~n8948 ;
  assign y3913 = ~n8950 ;
  assign y3914 = n8958 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = ~1'b0 ;
  assign y3917 = ~1'b0 ;
  assign y3918 = n8965 ;
  assign y3919 = n8973 ;
  assign y3920 = ~1'b0 ;
  assign y3921 = ~n8977 ;
  assign y3922 = n8979 ;
  assign y3923 = n8986 ;
  assign y3924 = ~1'b0 ;
  assign y3925 = ~n8988 ;
  assign y3926 = ~1'b0 ;
  assign y3927 = ~n8991 ;
  assign y3928 = n8994 ;
  assign y3929 = n9000 ;
  assign y3930 = ~1'b0 ;
  assign y3931 = ~n9003 ;
  assign y3932 = ~1'b0 ;
  assign y3933 = ~n9006 ;
  assign y3934 = n9009 ;
  assign y3935 = ~1'b0 ;
  assign y3936 = ~n711 ;
  assign y3937 = n9026 ;
  assign y3938 = n9027 ;
  assign y3939 = ~n9034 ;
  assign y3940 = n9041 ;
  assign y3941 = ~n9042 ;
  assign y3942 = n9043 ;
  assign y3943 = n9049 ;
  assign y3944 = ~n9051 ;
  assign y3945 = ~n9054 ;
  assign y3946 = n9057 ;
  assign y3947 = n9059 ;
  assign y3948 = ~1'b0 ;
  assign y3949 = ~1'b0 ;
  assign y3950 = ~1'b0 ;
  assign y3951 = n9060 ;
  assign y3952 = n9063 ;
  assign y3953 = n9066 ;
  assign y3954 = ~n9070 ;
  assign y3955 = ~n9074 ;
  assign y3956 = ~1'b0 ;
  assign y3957 = 1'b0 ;
  assign y3958 = ~1'b0 ;
  assign y3959 = ~n9083 ;
  assign y3960 = ~n9084 ;
  assign y3961 = ~1'b0 ;
  assign y3962 = n9087 ;
  assign y3963 = ~n9095 ;
  assign y3964 = n9096 ;
  assign y3965 = ~n9099 ;
  assign y3966 = n9108 ;
  assign y3967 = n9111 ;
  assign y3968 = n9113 ;
  assign y3969 = ~1'b0 ;
  assign y3970 = ~n9118 ;
  assign y3971 = n9119 ;
  assign y3972 = ~n9124 ;
  assign y3973 = ~n9125 ;
  assign y3974 = ~n9130 ;
  assign y3975 = ~n9137 ;
  assign y3976 = ~n9139 ;
  assign y3977 = ~n9142 ;
  assign y3978 = ~n9143 ;
  assign y3979 = ~1'b0 ;
  assign y3980 = ~1'b0 ;
  assign y3981 = ~n9145 ;
  assign y3982 = ~n9148 ;
  assign y3983 = ~n9150 ;
  assign y3984 = ~n9152 ;
  assign y3985 = n9156 ;
  assign y3986 = ~n9158 ;
  assign y3987 = n9159 ;
  assign y3988 = n9161 ;
  assign y3989 = n542 ;
  assign y3990 = ~1'b0 ;
  assign y3991 = ~n9164 ;
  assign y3992 = ~1'b0 ;
  assign y3993 = n9168 ;
  assign y3994 = ~n9171 ;
  assign y3995 = n9173 ;
  assign y3996 = ~1'b0 ;
  assign y3997 = n9175 ;
  assign y3998 = n9176 ;
  assign y3999 = n9179 ;
  assign y4000 = ~1'b0 ;
  assign y4001 = n9181 ;
  assign y4002 = ~n9189 ;
  assign y4003 = ~n9192 ;
  assign y4004 = n9193 ;
  assign y4005 = n9197 ;
  assign y4006 = ~n9204 ;
  assign y4007 = ~1'b0 ;
  assign y4008 = ~n9215 ;
  assign y4009 = n9216 ;
  assign y4010 = n9221 ;
  assign y4011 = ~n9223 ;
  assign y4012 = ~1'b0 ;
  assign y4013 = n1751 ;
  assign y4014 = ~1'b0 ;
  assign y4015 = n9226 ;
  assign y4016 = n9230 ;
  assign y4017 = ~n9232 ;
  assign y4018 = ~n9236 ;
  assign y4019 = ~n9238 ;
  assign y4020 = ~n9240 ;
  assign y4021 = n9248 ;
  assign y4022 = 1'b0 ;
  assign y4023 = ~n9255 ;
  assign y4024 = n9257 ;
  assign y4025 = ~n6739 ;
  assign y4026 = ~n9267 ;
  assign y4027 = ~n213 ;
  assign y4028 = n9269 ;
  assign y4029 = ~n9273 ;
  assign y4030 = ~1'b0 ;
  assign y4031 = ~n9274 ;
  assign y4032 = 1'b0 ;
  assign y4033 = ~1'b0 ;
  assign y4034 = ~1'b0 ;
  assign y4035 = n9275 ;
  assign y4036 = n9276 ;
  assign y4037 = ~1'b0 ;
  assign y4038 = ~n9278 ;
  assign y4039 = ~n9283 ;
  assign y4040 = ~n9284 ;
  assign y4041 = n9293 ;
  assign y4042 = n9299 ;
  assign y4043 = ~1'b0 ;
  assign y4044 = n9304 ;
  assign y4045 = ~1'b0 ;
  assign y4046 = ~1'b0 ;
  assign y4047 = 1'b0 ;
  assign y4048 = ~n9306 ;
  assign y4049 = ~1'b0 ;
  assign y4050 = ~n9311 ;
  assign y4051 = ~1'b0 ;
  assign y4052 = ~n9312 ;
  assign y4053 = n5716 ;
  assign y4054 = ~n9313 ;
  assign y4055 = n9315 ;
  assign y4056 = ~1'b0 ;
  assign y4057 = n9320 ;
  assign y4058 = ~n9323 ;
  assign y4059 = ~n9324 ;
  assign y4060 = ~1'b0 ;
  assign y4061 = n9325 ;
  assign y4062 = ~n9326 ;
  assign y4063 = n9328 ;
  assign y4064 = n9331 ;
  assign y4065 = ~n9333 ;
  assign y4066 = ~n9334 ;
  assign y4067 = ~n9337 ;
  assign y4068 = n9340 ;
  assign y4069 = n9347 ;
  assign y4070 = ~n6193 ;
  assign y4071 = n9351 ;
  assign y4072 = ~n9353 ;
  assign y4073 = ~n9354 ;
  assign y4074 = ~n9355 ;
  assign y4075 = ~n9357 ;
  assign y4076 = ~1'b0 ;
  assign y4077 = ~n9361 ;
  assign y4078 = ~1'b0 ;
  assign y4079 = ~1'b0 ;
  assign y4080 = n9363 ;
  assign y4081 = ~n9367 ;
  assign y4082 = ~n9371 ;
  assign y4083 = ~1'b0 ;
  assign y4084 = n9372 ;
  assign y4085 = ~n9379 ;
  assign y4086 = ~n9384 ;
  assign y4087 = ~1'b0 ;
  assign y4088 = ~1'b0 ;
  assign y4089 = n9386 ;
  assign y4090 = ~n9391 ;
  assign y4091 = n9392 ;
  assign y4092 = ~n9395 ;
  assign y4093 = ~1'b0 ;
  assign y4094 = ~n9399 ;
  assign y4095 = n9401 ;
  assign y4096 = n9402 ;
  assign y4097 = ~n9409 ;
  assign y4098 = ~1'b0 ;
  assign y4099 = n9415 ;
  assign y4100 = n9418 ;
  assign y4101 = ~1'b0 ;
  assign y4102 = ~1'b0 ;
  assign y4103 = ~1'b0 ;
  assign y4104 = ~1'b0 ;
  assign y4105 = n9422 ;
  assign y4106 = ~n9423 ;
  assign y4107 = n9424 ;
  assign y4108 = ~n9425 ;
  assign y4109 = ~1'b0 ;
  assign y4110 = n9430 ;
  assign y4111 = n9432 ;
  assign y4112 = ~n9435 ;
  assign y4113 = n9436 ;
  assign y4114 = ~1'b0 ;
  assign y4115 = ~n9438 ;
  assign y4116 = n9439 ;
  assign y4117 = ~n9441 ;
  assign y4118 = n9443 ;
  assign y4119 = ~1'b0 ;
  assign y4120 = n9449 ;
  assign y4121 = ~1'b0 ;
  assign y4122 = 1'b0 ;
  assign y4123 = ~n9451 ;
  assign y4124 = n9454 ;
  assign y4125 = n9457 ;
  assign y4126 = ~n9460 ;
  assign y4127 = n9467 ;
  assign y4128 = n9478 ;
  assign y4129 = ~1'b0 ;
  assign y4130 = n9481 ;
  assign y4131 = ~n9483 ;
  assign y4132 = ~n9484 ;
  assign y4133 = ~1'b0 ;
  assign y4134 = n9485 ;
  assign y4135 = n9493 ;
  assign y4136 = ~n9501 ;
  assign y4137 = ~1'b0 ;
  assign y4138 = ~n9503 ;
  assign y4139 = ~n9504 ;
  assign y4140 = ~1'b0 ;
  assign y4141 = ~n9506 ;
  assign y4142 = ~1'b0 ;
  assign y4143 = ~1'b0 ;
  assign y4144 = ~n9522 ;
  assign y4145 = n9526 ;
  assign y4146 = ~1'b0 ;
  assign y4147 = ~1'b0 ;
  assign y4148 = n9527 ;
  assign y4149 = n9528 ;
  assign y4150 = n9529 ;
  assign y4151 = ~n9530 ;
  assign y4152 = ~n9533 ;
  assign y4153 = n9543 ;
  assign y4154 = ~1'b0 ;
  assign y4155 = ~n9545 ;
  assign y4156 = ~n9548 ;
  assign y4157 = ~1'b0 ;
  assign y4158 = ~n9553 ;
  assign y4159 = n9557 ;
  assign y4160 = ~1'b0 ;
  assign y4161 = ~n9162 ;
  assign y4162 = ~n9562 ;
  assign y4163 = ~n9563 ;
  assign y4164 = n9568 ;
  assign y4165 = n9578 ;
  assign y4166 = n9584 ;
  assign y4167 = n4262 ;
  assign y4168 = n9586 ;
  assign y4169 = n9589 ;
  assign y4170 = ~n9594 ;
  assign y4171 = ~1'b0 ;
  assign y4172 = n9596 ;
  assign y4173 = n9597 ;
  assign y4174 = n5673 ;
  assign y4175 = ~n9598 ;
  assign y4176 = ~1'b0 ;
  assign y4177 = ~1'b0 ;
  assign y4178 = n9600 ;
  assign y4179 = ~1'b0 ;
  assign y4180 = ~1'b0 ;
  assign y4181 = ~1'b0 ;
  assign y4182 = ~1'b0 ;
  assign y4183 = ~1'b0 ;
  assign y4184 = n9605 ;
  assign y4185 = n9613 ;
  assign y4186 = ~n9614 ;
  assign y4187 = ~n9616 ;
  assign y4188 = ~n9619 ;
  assign y4189 = ~n9625 ;
  assign y4190 = ~n9626 ;
  assign y4191 = ~n9627 ;
  assign y4192 = ~1'b0 ;
  assign y4193 = ~n9633 ;
  assign y4194 = ~n9634 ;
  assign y4195 = n9636 ;
  assign y4196 = ~n9639 ;
  assign y4197 = ~n9640 ;
  assign y4198 = ~1'b0 ;
  assign y4199 = ~n9643 ;
  assign y4200 = ~n9644 ;
  assign y4201 = ~n9645 ;
  assign y4202 = ~n9646 ;
  assign y4203 = ~1'b0 ;
  assign y4204 = 1'b0 ;
  assign y4205 = ~n9647 ;
  assign y4206 = n9652 ;
  assign y4207 = ~n9653 ;
  assign y4208 = ~n9656 ;
  assign y4209 = ~n9661 ;
  assign y4210 = ~n9663 ;
  assign y4211 = n9664 ;
  assign y4212 = ~n9669 ;
  assign y4213 = ~1'b0 ;
  assign y4214 = ~n9673 ;
  assign y4215 = ~1'b0 ;
  assign y4216 = ~1'b0 ;
  assign y4217 = ~1'b0 ;
  assign y4218 = n9676 ;
  assign y4219 = ~1'b0 ;
  assign y4220 = n9679 ;
  assign y4221 = n9680 ;
  assign y4222 = ~1'b0 ;
  assign y4223 = ~1'b0 ;
  assign y4224 = ~1'b0 ;
  assign y4225 = ~n9681 ;
  assign y4226 = ~1'b0 ;
  assign y4227 = n9686 ;
  assign y4228 = ~n9687 ;
  assign y4229 = ~1'b0 ;
  assign y4230 = ~1'b0 ;
  assign y4231 = n9694 ;
  assign y4232 = n9698 ;
  assign y4233 = ~1'b0 ;
  assign y4234 = n9699 ;
  assign y4235 = n2873 ;
  assign y4236 = ~1'b0 ;
  assign y4237 = n9700 ;
  assign y4238 = ~n9703 ;
  assign y4239 = ~n9705 ;
  assign y4240 = n9706 ;
  assign y4241 = n9712 ;
  assign y4242 = n9715 ;
  assign y4243 = ~n9716 ;
  assign y4244 = n9722 ;
  assign y4245 = ~1'b0 ;
  assign y4246 = ~n9723 ;
  assign y4247 = ~n9724 ;
  assign y4248 = ~1'b0 ;
  assign y4249 = n9729 ;
  assign y4250 = ~1'b0 ;
  assign y4251 = n9730 ;
  assign y4252 = ~n9737 ;
  assign y4253 = ~n9741 ;
  assign y4254 = ~1'b0 ;
  assign y4255 = n8912 ;
  assign y4256 = ~n9746 ;
  assign y4257 = n9750 ;
  assign y4258 = n9760 ;
  assign y4259 = ~n9761 ;
  assign y4260 = ~n6451 ;
  assign y4261 = ~1'b0 ;
  assign y4262 = n9764 ;
  assign y4263 = ~n9766 ;
  assign y4264 = ~1'b0 ;
  assign y4265 = ~1'b0 ;
  assign y4266 = n7391 ;
  assign y4267 = n9768 ;
  assign y4268 = ~n9772 ;
  assign y4269 = n9779 ;
  assign y4270 = n9780 ;
  assign y4271 = ~n9782 ;
  assign y4272 = ~n9789 ;
  assign y4273 = ~n9790 ;
  assign y4274 = ~n9793 ;
  assign y4275 = ~n9794 ;
  assign y4276 = n9798 ;
  assign y4277 = ~1'b0 ;
  assign y4278 = ~1'b0 ;
  assign y4279 = ~n9801 ;
  assign y4280 = ~n9802 ;
  assign y4281 = ~n9804 ;
  assign y4282 = n9805 ;
  assign y4283 = ~n9806 ;
  assign y4284 = ~1'b0 ;
  assign y4285 = n9808 ;
  assign y4286 = ~n9813 ;
  assign y4287 = ~n4126 ;
  assign y4288 = n9817 ;
  assign y4289 = n9818 ;
  assign y4290 = n9819 ;
  assign y4291 = ~1'b0 ;
  assign y4292 = ~1'b0 ;
  assign y4293 = ~1'b0 ;
  assign y4294 = ~n9820 ;
  assign y4295 = n9823 ;
  assign y4296 = ~n9826 ;
  assign y4297 = ~1'b0 ;
  assign y4298 = ~n9827 ;
  assign y4299 = n9829 ;
  assign y4300 = n9830 ;
  assign y4301 = ~n9838 ;
  assign y4302 = ~n9841 ;
  assign y4303 = ~1'b0 ;
  assign y4304 = n3949 ;
  assign y4305 = ~n9847 ;
  assign y4306 = n9862 ;
  assign y4307 = ~n9863 ;
  assign y4308 = n191 ;
  assign y4309 = n9869 ;
  assign y4310 = ~n9875 ;
  assign y4311 = ~n9880 ;
  assign y4312 = ~1'b0 ;
  assign y4313 = ~n9882 ;
  assign y4314 = 1'b0 ;
  assign y4315 = ~n9884 ;
  assign y4316 = n9893 ;
  assign y4317 = n9894 ;
  assign y4318 = ~n9896 ;
  assign y4319 = n9904 ;
  assign y4320 = ~n9905 ;
  assign y4321 = ~1'b0 ;
  assign y4322 = ~n9907 ;
  assign y4323 = ~n9911 ;
  assign y4324 = ~n9915 ;
  assign y4325 = ~n9917 ;
  assign y4326 = ~1'b0 ;
  assign y4327 = ~1'b0 ;
  assign y4328 = ~1'b0 ;
  assign y4329 = ~1'b0 ;
  assign y4330 = ~1'b0 ;
  assign y4331 = n9920 ;
  assign y4332 = ~n9926 ;
  assign y4333 = ~n9932 ;
  assign y4334 = ~n9934 ;
  assign y4335 = ~n9937 ;
  assign y4336 = ~1'b0 ;
  assign y4337 = ~1'b0 ;
  assign y4338 = ~1'b0 ;
  assign y4339 = ~n9938 ;
  assign y4340 = ~n9942 ;
  assign y4341 = n9948 ;
  assign y4342 = n9950 ;
  assign y4343 = ~n9954 ;
  assign y4344 = ~1'b0 ;
  assign y4345 = n9958 ;
  assign y4346 = ~1'b0 ;
  assign y4347 = ~1'b0 ;
  assign y4348 = ~1'b0 ;
  assign y4349 = ~n9961 ;
  assign y4350 = ~n9964 ;
  assign y4351 = ~1'b0 ;
  assign y4352 = ~n9966 ;
  assign y4353 = ~n9968 ;
  assign y4354 = ~n1402 ;
  assign y4355 = n9972 ;
  assign y4356 = n9979 ;
  assign y4357 = ~n9982 ;
  assign y4358 = ~1'b0 ;
  assign y4359 = ~1'b0 ;
  assign y4360 = n9983 ;
  assign y4361 = ~1'b0 ;
  assign y4362 = n9987 ;
  assign y4363 = ~n9991 ;
  assign y4364 = ~n9995 ;
  assign y4365 = ~n9996 ;
  assign y4366 = ~n9998 ;
  assign y4367 = ~1'b0 ;
  assign y4368 = 1'b0 ;
  assign y4369 = ~n10003 ;
  assign y4370 = ~n10005 ;
  assign y4371 = n10010 ;
  assign y4372 = ~n10014 ;
  assign y4373 = ~n10020 ;
  assign y4374 = n10021 ;
  assign y4375 = ~n10027 ;
  assign y4376 = 1'b0 ;
  assign y4377 = n10031 ;
  assign y4378 = n10033 ;
  assign y4379 = n10037 ;
  assign y4380 = n10048 ;
  assign y4381 = ~1'b0 ;
  assign y4382 = ~n10049 ;
  assign y4383 = ~1'b0 ;
  assign y4384 = n10050 ;
  assign y4385 = ~1'b0 ;
  assign y4386 = n10051 ;
  assign y4387 = ~n10055 ;
  assign y4388 = ~n10056 ;
  assign y4389 = n10058 ;
  assign y4390 = n10059 ;
  assign y4391 = n10063 ;
  assign y4392 = 1'b0 ;
  assign y4393 = ~1'b0 ;
  assign y4394 = n10066 ;
  assign y4395 = ~1'b0 ;
  assign y4396 = n10072 ;
  assign y4397 = ~1'b0 ;
  assign y4398 = ~n10074 ;
  assign y4399 = n10077 ;
  assign y4400 = ~1'b0 ;
  assign y4401 = ~1'b0 ;
  assign y4402 = ~n10078 ;
  assign y4403 = ~1'b0 ;
  assign y4404 = ~n10082 ;
  assign y4405 = ~1'b0 ;
  assign y4406 = n10085 ;
  assign y4407 = n10086 ;
  assign y4408 = n10087 ;
  assign y4409 = ~1'b0 ;
  assign y4410 = ~n10091 ;
  assign y4411 = ~1'b0 ;
  assign y4412 = ~1'b0 ;
  assign y4413 = ~1'b0 ;
  assign y4414 = n10094 ;
  assign y4415 = ~n10096 ;
  assign y4416 = n10102 ;
  assign y4417 = n10106 ;
  assign y4418 = ~1'b0 ;
  assign y4419 = n6670 ;
  assign y4420 = ~n10111 ;
  assign y4421 = ~n10115 ;
  assign y4422 = ~n10122 ;
  assign y4423 = ~n10130 ;
  assign y4424 = ~n10135 ;
  assign y4425 = ~n10140 ;
  assign y4426 = ~n10143 ;
  assign y4427 = ~n10151 ;
  assign y4428 = ~n10153 ;
  assign y4429 = n10154 ;
  assign y4430 = n10161 ;
  assign y4431 = ~1'b0 ;
  assign y4432 = n5281 ;
  assign y4433 = n10169 ;
  assign y4434 = ~n8740 ;
  assign y4435 = n10173 ;
  assign y4436 = ~1'b0 ;
  assign y4437 = n10177 ;
  assign y4438 = ~1'b0 ;
  assign y4439 = ~n10178 ;
  assign y4440 = ~1'b0 ;
  assign y4441 = ~n10183 ;
  assign y4442 = n10186 ;
  assign y4443 = ~1'b0 ;
  assign y4444 = n10190 ;
  assign y4445 = ~1'b0 ;
  assign y4446 = n10195 ;
  assign y4447 = ~1'b0 ;
  assign y4448 = ~n10196 ;
  assign y4449 = ~1'b0 ;
  assign y4450 = ~n10204 ;
  assign y4451 = ~n10209 ;
  assign y4452 = n10210 ;
  assign y4453 = 1'b0 ;
  assign y4454 = ~n10212 ;
  assign y4455 = n10213 ;
  assign y4456 = n10217 ;
  assign y4457 = ~n10218 ;
  assign y4458 = n10221 ;
  assign y4459 = ~1'b0 ;
  assign y4460 = ~1'b0 ;
  assign y4461 = ~n10226 ;
  assign y4462 = ~1'b0 ;
  assign y4463 = n10228 ;
  assign y4464 = ~n10230 ;
  assign y4465 = ~1'b0 ;
  assign y4466 = n10231 ;
  assign y4467 = ~1'b0 ;
  assign y4468 = ~1'b0 ;
  assign y4469 = ~1'b0 ;
  assign y4470 = ~n10232 ;
  assign y4471 = n10233 ;
  assign y4472 = ~n10236 ;
  assign y4473 = ~n10238 ;
  assign y4474 = ~1'b0 ;
  assign y4475 = ~n10244 ;
  assign y4476 = ~n10245 ;
  assign y4477 = ~1'b0 ;
  assign y4478 = ~1'b0 ;
  assign y4479 = n10247 ;
  assign y4480 = n10249 ;
  assign y4481 = ~1'b0 ;
  assign y4482 = n10252 ;
  assign y4483 = ~n10254 ;
  assign y4484 = ~1'b0 ;
  assign y4485 = n10256 ;
  assign y4486 = ~n10258 ;
  assign y4487 = ~n10261 ;
  assign y4488 = ~1'b0 ;
  assign y4489 = ~n10266 ;
  assign y4490 = ~1'b0 ;
  assign y4491 = n10269 ;
  assign y4492 = n10270 ;
  assign y4493 = ~n10272 ;
  assign y4494 = ~n10273 ;
  assign y4495 = ~1'b0 ;
  assign y4496 = ~n8941 ;
  assign y4497 = n10274 ;
  assign y4498 = ~n10276 ;
  assign y4499 = n10279 ;
  assign y4500 = ~n10292 ;
  assign y4501 = ~1'b0 ;
  assign y4502 = ~1'b0 ;
  assign y4503 = ~1'b0 ;
  assign y4504 = n10294 ;
  assign y4505 = n10297 ;
  assign y4506 = ~1'b0 ;
  assign y4507 = n10301 ;
  assign y4508 = ~n10305 ;
  assign y4509 = n10308 ;
  assign y4510 = ~n10311 ;
  assign y4511 = ~n10312 ;
  assign y4512 = n7363 ;
  assign y4513 = ~n10318 ;
  assign y4514 = ~1'b0 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = ~n10322 ;
  assign y4517 = ~n10325 ;
  assign y4518 = ~n10329 ;
  assign y4519 = ~n10330 ;
  assign y4520 = ~n1410 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = n10335 ;
  assign y4523 = ~1'b0 ;
  assign y4524 = ~n10337 ;
  assign y4525 = n10340 ;
  assign y4526 = n10342 ;
  assign y4527 = ~n10343 ;
  assign y4528 = ~n10344 ;
  assign y4529 = ~1'b0 ;
  assign y4530 = ~1'b0 ;
  assign y4531 = n10345 ;
  assign y4532 = n4578 ;
  assign y4533 = ~n10346 ;
  assign y4534 = ~n4059 ;
  assign y4535 = n10347 ;
  assign y4536 = n10352 ;
  assign y4537 = ~n10361 ;
  assign y4538 = ~1'b0 ;
  assign y4539 = ~1'b0 ;
  assign y4540 = ~n10368 ;
  assign y4541 = ~n10371 ;
  assign y4542 = ~1'b0 ;
  assign y4543 = ~n10372 ;
  assign y4544 = n23 ;
  assign y4545 = n10373 ;
  assign y4546 = ~1'b0 ;
  assign y4547 = ~1'b0 ;
  assign y4548 = n10375 ;
  assign y4549 = n10378 ;
  assign y4550 = n10381 ;
  assign y4551 = ~n7672 ;
  assign y4552 = ~1'b0 ;
  assign y4553 = n10383 ;
  assign y4554 = ~1'b0 ;
  assign y4555 = n10384 ;
  assign y4556 = n352 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = n10387 ;
  assign y4559 = n10392 ;
  assign y4560 = ~1'b0 ;
  assign y4561 = n10393 ;
  assign y4562 = n10394 ;
  assign y4563 = n10395 ;
  assign y4564 = n10396 ;
  assign y4565 = ~n10398 ;
  assign y4566 = n10400 ;
  assign y4567 = ~n10404 ;
  assign y4568 = ~n10406 ;
  assign y4569 = ~n10416 ;
  assign y4570 = ~n8088 ;
  assign y4571 = n5339 ;
  assign y4572 = ~1'b0 ;
  assign y4573 = n10417 ;
  assign y4574 = ~n10418 ;
  assign y4575 = ~n10421 ;
  assign y4576 = ~n10423 ;
  assign y4577 = ~1'b0 ;
  assign y4578 = ~1'b0 ;
  assign y4579 = n10432 ;
  assign y4580 = ~n10433 ;
  assign y4581 = n10435 ;
  assign y4582 = ~n10440 ;
  assign y4583 = ~1'b0 ;
  assign y4584 = ~n10443 ;
  assign y4585 = ~1'b0 ;
  assign y4586 = ~1'b0 ;
  assign y4587 = ~n10446 ;
  assign y4588 = ~n10448 ;
  assign y4589 = n10450 ;
  assign y4590 = ~1'b0 ;
  assign y4591 = ~1'b0 ;
  assign y4592 = ~n10457 ;
  assign y4593 = ~n10461 ;
  assign y4594 = ~1'b0 ;
  assign y4595 = ~1'b0 ;
  assign y4596 = n10464 ;
  assign y4597 = ~n10472 ;
  assign y4598 = ~n3181 ;
  assign y4599 = n10473 ;
  assign y4600 = n10478 ;
  assign y4601 = n10480 ;
  assign y4602 = ~n10482 ;
  assign y4603 = n10484 ;
  assign y4604 = ~n10487 ;
  assign y4605 = ~1'b0 ;
  assign y4606 = ~1'b0 ;
  assign y4607 = n10490 ;
  assign y4608 = ~n10491 ;
  assign y4609 = ~1'b0 ;
  assign y4610 = ~n10492 ;
  assign y4611 = ~1'b0 ;
  assign y4612 = ~1'b0 ;
  assign y4613 = n10496 ;
  assign y4614 = n10498 ;
  assign y4615 = ~n10499 ;
  assign y4616 = n10500 ;
  assign y4617 = n10501 ;
  assign y4618 = ~1'b0 ;
  assign y4619 = ~n10503 ;
  assign y4620 = ~1'b0 ;
  assign y4621 = ~n10514 ;
  assign y4622 = ~n10521 ;
  assign y4623 = n10523 ;
  assign y4624 = n10528 ;
  assign y4625 = n10532 ;
  assign y4626 = ~n10539 ;
  assign y4627 = ~n10550 ;
  assign y4628 = ~n10557 ;
  assign y4629 = ~1'b0 ;
  assign y4630 = ~n10559 ;
  assign y4631 = n10562 ;
  assign y4632 = ~n10565 ;
  assign y4633 = ~n10567 ;
  assign y4634 = n10568 ;
  assign y4635 = ~n10572 ;
  assign y4636 = ~n10577 ;
  assign y4637 = n9631 ;
  assign y4638 = n10582 ;
  assign y4639 = n8043 ;
  assign y4640 = ~1'b0 ;
  assign y4641 = n10585 ;
  assign y4642 = ~1'b0 ;
  assign y4643 = ~1'b0 ;
  assign y4644 = n10586 ;
  assign y4645 = n10588 ;
  assign y4646 = ~n10591 ;
  assign y4647 = ~1'b0 ;
  assign y4648 = ~n10592 ;
  assign y4649 = ~1'b0 ;
  assign y4650 = n8170 ;
  assign y4651 = ~n10593 ;
  assign y4652 = n10594 ;
  assign y4653 = n5016 ;
  assign y4654 = n543 ;
  assign y4655 = ~1'b0 ;
  assign y4656 = ~n10596 ;
  assign y4657 = ~1'b0 ;
  assign y4658 = ~n10599 ;
  assign y4659 = ~n10600 ;
  assign y4660 = n10621 ;
  assign y4661 = ~n10623 ;
  assign y4662 = ~n10624 ;
  assign y4663 = ~n10630 ;
  assign y4664 = ~1'b0 ;
  assign y4665 = ~1'b0 ;
  assign y4666 = n10631 ;
  assign y4667 = n2044 ;
  assign y4668 = n10635 ;
  assign y4669 = n10643 ;
  assign y4670 = n10646 ;
  assign y4671 = n10648 ;
  assign y4672 = n10650 ;
  assign y4673 = ~n10654 ;
  assign y4674 = ~1'b0 ;
  assign y4675 = ~1'b0 ;
  assign y4676 = ~n10658 ;
  assign y4677 = ~1'b0 ;
  assign y4678 = n10664 ;
  assign y4679 = ~n10665 ;
  assign y4680 = n10667 ;
  assign y4681 = n10668 ;
  assign y4682 = n10670 ;
  assign y4683 = ~n10673 ;
  assign y4684 = n10675 ;
  assign y4685 = n1487 ;
  assign y4686 = ~n9921 ;
  assign y4687 = ~1'b0 ;
  assign y4688 = ~1'b0 ;
  assign y4689 = ~n10677 ;
  assign y4690 = n10684 ;
  assign y4691 = ~1'b0 ;
  assign y4692 = ~n10685 ;
  assign y4693 = ~n10688 ;
  assign y4694 = ~n5930 ;
  assign y4695 = ~1'b0 ;
  assign y4696 = ~n10708 ;
  assign y4697 = n10712 ;
  assign y4698 = ~n10717 ;
  assign y4699 = n10720 ;
  assign y4700 = n5713 ;
  assign y4701 = ~n10722 ;
  assign y4702 = ~n10724 ;
  assign y4703 = ~n10726 ;
  assign y4704 = n10733 ;
  assign y4705 = n10747 ;
  assign y4706 = ~1'b0 ;
  assign y4707 = n10748 ;
  assign y4708 = n10749 ;
  assign y4709 = ~1'b0 ;
  assign y4710 = ~n10751 ;
  assign y4711 = ~1'b0 ;
  assign y4712 = n10753 ;
  assign y4713 = ~n10348 ;
  assign y4714 = n10754 ;
  assign y4715 = ~n10756 ;
  assign y4716 = ~n10764 ;
  assign y4717 = n10765 ;
  assign y4718 = n10769 ;
  assign y4719 = ~1'b0 ;
  assign y4720 = n10772 ;
  assign y4721 = n10773 ;
  assign y4722 = n10775 ;
  assign y4723 = ~1'b0 ;
  assign y4724 = n1891 ;
  assign y4725 = ~n10781 ;
  assign y4726 = ~1'b0 ;
  assign y4727 = ~n10783 ;
  assign y4728 = ~n5501 ;
  assign y4729 = n10791 ;
  assign y4730 = ~n10792 ;
  assign y4731 = n10795 ;
  assign y4732 = n10797 ;
  assign y4733 = ~1'b0 ;
  assign y4734 = ~n10802 ;
  assign y4735 = ~n10803 ;
  assign y4736 = 1'b0 ;
  assign y4737 = ~n10807 ;
  assign y4738 = n10809 ;
  assign y4739 = ~1'b0 ;
  assign y4740 = n10811 ;
  assign y4741 = ~n10815 ;
  assign y4742 = ~n10817 ;
  assign y4743 = n10819 ;
  assign y4744 = n10822 ;
  assign y4745 = n10824 ;
  assign y4746 = ~n10827 ;
  assign y4747 = ~n3758 ;
  assign y4748 = ~1'b0 ;
  assign y4749 = ~n10833 ;
  assign y4750 = ~n10836 ;
  assign y4751 = ~1'b0 ;
  assign y4752 = ~1'b0 ;
  assign y4753 = ~1'b0 ;
  assign y4754 = ~n10842 ;
  assign y4755 = n10848 ;
  assign y4756 = ~n10857 ;
  assign y4757 = ~1'b0 ;
  assign y4758 = ~n4549 ;
  assign y4759 = ~1'b0 ;
  assign y4760 = n10859 ;
  assign y4761 = ~1'b0 ;
  assign y4762 = ~n10861 ;
  assign y4763 = ~1'b0 ;
  assign y4764 = ~n10863 ;
  assign y4765 = ~1'b0 ;
  assign y4766 = n10870 ;
  assign y4767 = ~n10872 ;
  assign y4768 = n10873 ;
  assign y4769 = n10878 ;
  assign y4770 = ~n10886 ;
  assign y4771 = ~n10894 ;
  assign y4772 = ~1'b0 ;
  assign y4773 = ~n10897 ;
  assign y4774 = ~n10352 ;
  assign y4775 = n10898 ;
  assign y4776 = ~1'b0 ;
  assign y4777 = ~1'b0 ;
  assign y4778 = ~n10899 ;
  assign y4779 = ~n5740 ;
  assign y4780 = n10900 ;
  assign y4781 = ~1'b0 ;
  assign y4782 = n1771 ;
  assign y4783 = n10902 ;
  assign y4784 = ~1'b0 ;
  assign y4785 = ~n4275 ;
  assign y4786 = ~n10907 ;
  assign y4787 = ~n10913 ;
  assign y4788 = ~1'b0 ;
  assign y4789 = n1414 ;
  assign y4790 = n10920 ;
  assign y4791 = ~n10924 ;
  assign y4792 = ~n10928 ;
  assign y4793 = ~n10930 ;
  assign y4794 = ~n10933 ;
  assign y4795 = ~1'b0 ;
  assign y4796 = 1'b0 ;
  assign y4797 = n10934 ;
  assign y4798 = ~n10935 ;
  assign y4799 = ~n10938 ;
  assign y4800 = ~n10940 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = ~1'b0 ;
  assign y4803 = ~1'b0 ;
  assign y4804 = ~n10941 ;
  assign y4805 = ~n10948 ;
  assign y4806 = ~1'b0 ;
  assign y4807 = n10957 ;
  assign y4808 = ~n1105 ;
  assign y4809 = ~n10958 ;
  assign y4810 = ~1'b0 ;
  assign y4811 = n10959 ;
  assign y4812 = ~n10963 ;
  assign y4813 = ~1'b0 ;
  assign y4814 = n10966 ;
  assign y4815 = n3840 ;
  assign y4816 = n10967 ;
  assign y4817 = 1'b0 ;
  assign y4818 = ~n10969 ;
  assign y4819 = ~n10971 ;
  assign y4820 = ~1'b0 ;
  assign y4821 = ~n10973 ;
  assign y4822 = ~n10974 ;
  assign y4823 = ~n10975 ;
  assign y4824 = n10976 ;
  assign y4825 = n10977 ;
  assign y4826 = ~n10978 ;
  assign y4827 = ~n10981 ;
  assign y4828 = ~1'b0 ;
  assign y4829 = ~1'b0 ;
  assign y4830 = ~n10982 ;
  assign y4831 = ~n10986 ;
  assign y4832 = ~1'b0 ;
  assign y4833 = ~1'b0 ;
  assign y4834 = n10987 ;
  assign y4835 = ~n10990 ;
  assign y4836 = n8536 ;
  assign y4837 = n10995 ;
  assign y4838 = ~n10997 ;
  assign y4839 = 1'b0 ;
  assign y4840 = n11003 ;
  assign y4841 = ~n11004 ;
  assign y4842 = n11006 ;
  assign y4843 = ~n11018 ;
  assign y4844 = ~n11022 ;
  assign y4845 = ~n11028 ;
  assign y4846 = n11029 ;
  assign y4847 = n4050 ;
  assign y4848 = n11033 ;
  assign y4849 = n11037 ;
  assign y4850 = 1'b0 ;
  assign y4851 = ~n11038 ;
  assign y4852 = n11041 ;
  assign y4853 = n11045 ;
  assign y4854 = ~n11048 ;
  assign y4855 = ~1'b0 ;
  assign y4856 = 1'b0 ;
  assign y4857 = ~n11050 ;
  assign y4858 = ~n11052 ;
  assign y4859 = ~1'b0 ;
  assign y4860 = n11057 ;
  assign y4861 = ~n11071 ;
  assign y4862 = ~1'b0 ;
  assign y4863 = ~1'b0 ;
  assign y4864 = n11073 ;
  assign y4865 = ~n11074 ;
  assign y4866 = n11076 ;
  assign y4867 = n11078 ;
  assign y4868 = ~n11086 ;
  assign y4869 = n11091 ;
  assign y4870 = ~n11094 ;
  assign y4871 = ~1'b0 ;
  assign y4872 = ~1'b0 ;
  assign y4873 = n11098 ;
  assign y4874 = ~1'b0 ;
  assign y4875 = ~n11101 ;
  assign y4876 = n11104 ;
  assign y4877 = ~1'b0 ;
  assign y4878 = ~n11115 ;
  assign y4879 = ~n11116 ;
  assign y4880 = ~n11118 ;
  assign y4881 = ~1'b0 ;
  assign y4882 = n1084 ;
  assign y4883 = ~n11119 ;
  assign y4884 = ~n11124 ;
  assign y4885 = n11129 ;
  assign y4886 = n9863 ;
  assign y4887 = ~n11134 ;
  assign y4888 = ~1'b0 ;
  assign y4889 = ~n11136 ;
  assign y4890 = n11145 ;
  assign y4891 = ~1'b0 ;
  assign y4892 = n11147 ;
  assign y4893 = ~n11153 ;
  assign y4894 = ~1'b0 ;
  assign y4895 = 1'b0 ;
  assign y4896 = n11157 ;
  assign y4897 = n7544 ;
  assign y4898 = n11159 ;
  assign y4899 = ~1'b0 ;
  assign y4900 = ~1'b0 ;
  assign y4901 = ~1'b0 ;
  assign y4902 = n11163 ;
  assign y4903 = ~1'b0 ;
  assign y4904 = ~1'b0 ;
  assign y4905 = ~n11169 ;
  assign y4906 = ~n11171 ;
  assign y4907 = n11172 ;
  assign y4908 = n11173 ;
  assign y4909 = n11178 ;
  assign y4910 = n11180 ;
  assign y4911 = ~n11184 ;
  assign y4912 = n11187 ;
  assign y4913 = n11188 ;
  assign y4914 = ~n11189 ;
  assign y4915 = n11199 ;
  assign y4916 = ~n11211 ;
  assign y4917 = n3156 ;
  assign y4918 = ~1'b0 ;
  assign y4919 = n11216 ;
  assign y4920 = ~n11218 ;
  assign y4921 = n11220 ;
  assign y4922 = ~n11221 ;
  assign y4923 = ~1'b0 ;
  assign y4924 = ~n11222 ;
  assign y4925 = ~1'b0 ;
  assign y4926 = ~1'b0 ;
  assign y4927 = ~n11226 ;
  assign y4928 = ~n11229 ;
  assign y4929 = n11230 ;
  assign y4930 = ~n11231 ;
  assign y4931 = n11233 ;
  assign y4932 = n4830 ;
  assign y4933 = ~n11235 ;
  assign y4934 = n11238 ;
  assign y4935 = n11239 ;
  assign y4936 = ~n11250 ;
  assign y4937 = ~n11251 ;
  assign y4938 = ~n11256 ;
  assign y4939 = ~n11269 ;
  assign y4940 = n11273 ;
  assign y4941 = ~1'b0 ;
  assign y4942 = ~n11274 ;
  assign y4943 = ~1'b0 ;
  assign y4944 = ~n11275 ;
  assign y4945 = ~n11279 ;
  assign y4946 = n11282 ;
  assign y4947 = ~1'b0 ;
  assign y4948 = n11292 ;
  assign y4949 = ~n11294 ;
  assign y4950 = n11295 ;
  assign y4951 = ~n11296 ;
  assign y4952 = ~n11301 ;
  assign y4953 = ~1'b0 ;
  assign y4954 = ~1'b0 ;
  assign y4955 = n11304 ;
  assign y4956 = ~n6804 ;
  assign y4957 = ~1'b0 ;
  assign y4958 = ~n11305 ;
  assign y4959 = 1'b0 ;
  assign y4960 = ~n11307 ;
  assign y4961 = n575 ;
  assign y4962 = ~n11311 ;
  assign y4963 = 1'b0 ;
  assign y4964 = n11312 ;
  assign y4965 = ~1'b0 ;
  assign y4966 = n11316 ;
  assign y4967 = n11320 ;
  assign y4968 = ~1'b0 ;
  assign y4969 = ~1'b0 ;
  assign y4970 = n11323 ;
  assign y4971 = ~n601 ;
  assign y4972 = ~n11325 ;
  assign y4973 = n11327 ;
  assign y4974 = ~n11332 ;
  assign y4975 = ~n11333 ;
  assign y4976 = ~1'b0 ;
  assign y4977 = ~1'b0 ;
  assign y4978 = ~1'b0 ;
  assign y4979 = ~1'b0 ;
  assign y4980 = ~1'b0 ;
  assign y4981 = ~1'b0 ;
  assign y4982 = n11337 ;
  assign y4983 = n11340 ;
  assign y4984 = n11346 ;
  assign y4985 = n11352 ;
  assign y4986 = ~n11353 ;
  assign y4987 = ~1'b0 ;
  assign y4988 = ~1'b0 ;
  assign y4989 = ~1'b0 ;
  assign y4990 = ~n11355 ;
  assign y4991 = 1'b0 ;
  assign y4992 = n11357 ;
  assign y4993 = n11367 ;
  assign y4994 = n11373 ;
  assign y4995 = n3043 ;
  assign y4996 = n11379 ;
  assign y4997 = ~1'b0 ;
  assign y4998 = n11381 ;
  assign y4999 = ~1'b0 ;
  assign y5000 = ~1'b0 ;
  assign y5001 = n11382 ;
  assign y5002 = ~1'b0 ;
  assign y5003 = ~n11385 ;
  assign y5004 = n11386 ;
  assign y5005 = n11399 ;
  assign y5006 = n2597 ;
  assign y5007 = n11402 ;
  assign y5008 = ~1'b0 ;
  assign y5009 = n11403 ;
  assign y5010 = ~1'b0 ;
  assign y5011 = ~n11406 ;
  assign y5012 = ~n11410 ;
  assign y5013 = ~n11413 ;
  assign y5014 = ~1'b0 ;
  assign y5015 = n11418 ;
  assign y5016 = ~n11419 ;
  assign y5017 = ~n11420 ;
  assign y5018 = n11422 ;
  assign y5019 = n11433 ;
  assign y5020 = n11442 ;
  assign y5021 = ~1'b0 ;
  assign y5022 = ~1'b0 ;
  assign y5023 = n11443 ;
  assign y5024 = n11446 ;
  assign y5025 = n11456 ;
  assign y5026 = ~1'b0 ;
  assign y5027 = n11458 ;
  assign y5028 = n11462 ;
  assign y5029 = n11467 ;
  assign y5030 = ~n11469 ;
  assign y5031 = n11470 ;
  assign y5032 = ~1'b0 ;
  assign y5033 = ~1'b0 ;
  assign y5034 = ~1'b0 ;
  assign y5035 = ~1'b0 ;
  assign y5036 = ~n11472 ;
  assign y5037 = ~1'b0 ;
  assign y5038 = ~n11475 ;
  assign y5039 = n11483 ;
  assign y5040 = n11490 ;
  assign y5041 = n11491 ;
  assign y5042 = ~1'b0 ;
  assign y5043 = ~n11494 ;
  assign y5044 = n11497 ;
  assign y5045 = 1'b0 ;
  assign y5046 = n6657 ;
  assign y5047 = n11498 ;
  assign y5048 = ~n11502 ;
  assign y5049 = n11503 ;
  assign y5050 = ~n11505 ;
  assign y5051 = ~n11507 ;
  assign y5052 = ~n11511 ;
  assign y5053 = n11513 ;
  assign y5054 = ~1'b0 ;
  assign y5055 = n8171 ;
  assign y5056 = n11514 ;
  assign y5057 = ~n11517 ;
  assign y5058 = ~1'b0 ;
  assign y5059 = ~n11521 ;
  assign y5060 = ~1'b0 ;
  assign y5061 = ~1'b0 ;
  assign y5062 = ~n11523 ;
  assign y5063 = ~n11528 ;
  assign y5064 = ~n11529 ;
  assign y5065 = ~1'b0 ;
  assign y5066 = n10775 ;
  assign y5067 = ~n11535 ;
  assign y5068 = ~1'b0 ;
  assign y5069 = ~n11536 ;
  assign y5070 = ~n11538 ;
  assign y5071 = n11540 ;
  assign y5072 = ~1'b0 ;
  assign y5073 = ~n11542 ;
  assign y5074 = ~n11543 ;
  assign y5075 = ~n11546 ;
  assign y5076 = ~1'b0 ;
  assign y5077 = ~n11549 ;
  assign y5078 = ~n11551 ;
  assign y5079 = ~1'b0 ;
  assign y5080 = ~n381 ;
  assign y5081 = ~1'b0 ;
  assign y5082 = ~n11554 ;
  assign y5083 = n4447 ;
  assign y5084 = ~1'b0 ;
  assign y5085 = n11559 ;
  assign y5086 = n11562 ;
  assign y5087 = ~n3066 ;
  assign y5088 = ~n11564 ;
  assign y5089 = ~1'b0 ;
  assign y5090 = ~n11566 ;
  assign y5091 = ~n11567 ;
  assign y5092 = ~1'b0 ;
  assign y5093 = ~n11568 ;
  assign y5094 = ~1'b0 ;
  assign y5095 = ~1'b0 ;
  assign y5096 = ~1'b0 ;
  assign y5097 = n11569 ;
  assign y5098 = ~n11572 ;
  assign y5099 = ~n11573 ;
  assign y5100 = n11574 ;
  assign y5101 = ~n11583 ;
  assign y5102 = ~n11591 ;
  assign y5103 = ~1'b0 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = n4892 ;
  assign y5106 = ~n10163 ;
  assign y5107 = ~1'b0 ;
  assign y5108 = n11593 ;
  assign y5109 = n11594 ;
  assign y5110 = ~n11595 ;
  assign y5111 = n11597 ;
  assign y5112 = n11599 ;
  assign y5113 = ~n11602 ;
  assign y5114 = 1'b0 ;
  assign y5115 = ~n11606 ;
  assign y5116 = n4057 ;
  assign y5117 = ~1'b0 ;
  assign y5118 = n11607 ;
  assign y5119 = n11609 ;
  assign y5120 = ~n11612 ;
  assign y5121 = n11614 ;
  assign y5122 = n11617 ;
  assign y5123 = ~n11620 ;
  assign y5124 = ~1'b0 ;
  assign y5125 = ~n7106 ;
  assign y5126 = ~n11622 ;
  assign y5127 = ~n11624 ;
  assign y5128 = ~1'b0 ;
  assign y5129 = n11631 ;
  assign y5130 = ~1'b0 ;
  assign y5131 = ~n11640 ;
  assign y5132 = ~n11643 ;
  assign y5133 = n11644 ;
  assign y5134 = ~n113 ;
  assign y5135 = ~1'b0 ;
  assign y5136 = n11650 ;
  assign y5137 = n11652 ;
  assign y5138 = n8024 ;
  assign y5139 = ~n11657 ;
  assign y5140 = ~n11662 ;
  assign y5141 = ~n11666 ;
  assign y5142 = ~n11678 ;
  assign y5143 = ~n11689 ;
  assign y5144 = ~n11691 ;
  assign y5145 = ~n11697 ;
  assign y5146 = n11698 ;
  assign y5147 = n11700 ;
  assign y5148 = n11704 ;
  assign y5149 = n11707 ;
  assign y5150 = ~n11711 ;
  assign y5151 = ~n11712 ;
  assign y5152 = ~n11713 ;
  assign y5153 = ~n11715 ;
  assign y5154 = n11717 ;
  assign y5155 = ~n11720 ;
  assign y5156 = ~1'b0 ;
  assign y5157 = n11723 ;
  assign y5158 = ~1'b0 ;
  assign y5159 = ~n11727 ;
  assign y5160 = ~1'b0 ;
  assign y5161 = 1'b0 ;
  assign y5162 = ~n11729 ;
  assign y5163 = ~1'b0 ;
  assign y5164 = 1'b0 ;
  assign y5165 = ~n11731 ;
  assign y5166 = n11733 ;
  assign y5167 = ~n11734 ;
  assign y5168 = ~1'b0 ;
  assign y5169 = ~n11735 ;
  assign y5170 = n11738 ;
  assign y5171 = ~n11743 ;
  assign y5172 = n11744 ;
  assign y5173 = ~n11746 ;
  assign y5174 = ~1'b0 ;
  assign y5175 = 1'b0 ;
  assign y5176 = ~n11750 ;
  assign y5177 = n11752 ;
  assign y5178 = ~n11753 ;
  assign y5179 = ~n11544 ;
  assign y5180 = n11762 ;
  assign y5181 = n11773 ;
  assign y5182 = ~1'b0 ;
  assign y5183 = n11778 ;
  assign y5184 = n1586 ;
  assign y5185 = ~1'b0 ;
  assign y5186 = n11780 ;
  assign y5187 = ~1'b0 ;
  assign y5188 = ~n11788 ;
  assign y5189 = n2631 ;
  assign y5190 = ~n11792 ;
  assign y5191 = ~1'b0 ;
  assign y5192 = n11794 ;
  assign y5193 = ~n11307 ;
  assign y5194 = ~1'b0 ;
  assign y5195 = n11798 ;
  assign y5196 = ~1'b0 ;
  assign y5197 = ~1'b0 ;
  assign y5198 = n11803 ;
  assign y5199 = ~n11805 ;
  assign y5200 = ~1'b0 ;
  assign y5201 = n11808 ;
  assign y5202 = ~n11812 ;
  assign y5203 = n11813 ;
  assign y5204 = ~n11818 ;
  assign y5205 = ~n11820 ;
  assign y5206 = ~n11825 ;
  assign y5207 = n11834 ;
  assign y5208 = ~1'b0 ;
  assign y5209 = ~1'b0 ;
  assign y5210 = n11836 ;
  assign y5211 = n11841 ;
  assign y5212 = n11846 ;
  assign y5213 = n11847 ;
  assign y5214 = 1'b0 ;
  assign y5215 = ~n11848 ;
  assign y5216 = ~1'b0 ;
  assign y5217 = n11850 ;
  assign y5218 = n11853 ;
  assign y5219 = ~1'b0 ;
  assign y5220 = ~n11854 ;
  assign y5221 = ~1'b0 ;
  assign y5222 = ~1'b0 ;
  assign y5223 = n11862 ;
  assign y5224 = n11864 ;
  assign y5225 = ~n11865 ;
  assign y5226 = ~n11872 ;
  assign y5227 = n11873 ;
  assign y5228 = n11877 ;
  assign y5229 = n11879 ;
  assign y5230 = n11880 ;
  assign y5231 = ~n11881 ;
  assign y5232 = ~1'b0 ;
  assign y5233 = ~1'b0 ;
  assign y5234 = ~n11890 ;
  assign y5235 = ~n11893 ;
  assign y5236 = n11894 ;
  assign y5237 = n11898 ;
  assign y5238 = ~1'b0 ;
  assign y5239 = n11911 ;
  assign y5240 = ~n11916 ;
  assign y5241 = n11919 ;
  assign y5242 = n11928 ;
  assign y5243 = ~n11938 ;
  assign y5244 = ~1'b0 ;
  assign y5245 = ~n11941 ;
  assign y5246 = ~1'b0 ;
  assign y5247 = ~n11943 ;
  assign y5248 = n11949 ;
  assign y5249 = n11950 ;
  assign y5250 = n11954 ;
  assign y5251 = ~n11955 ;
  assign y5252 = ~1'b0 ;
  assign y5253 = n11957 ;
  assign y5254 = ~n11963 ;
  assign y5255 = ~1'b0 ;
  assign y5256 = n11964 ;
  assign y5257 = n11966 ;
  assign y5258 = ~n11967 ;
  assign y5259 = ~1'b0 ;
  assign y5260 = n11968 ;
  assign y5261 = n11971 ;
  assign y5262 = ~n11973 ;
  assign y5263 = n11980 ;
  assign y5264 = n11987 ;
  assign y5265 = ~1'b0 ;
  assign y5266 = n4992 ;
  assign y5267 = n10829 ;
  assign y5268 = ~1'b0 ;
  assign y5269 = n11988 ;
  assign y5270 = n11996 ;
  assign y5271 = n11997 ;
  assign y5272 = ~1'b0 ;
  assign y5273 = ~n11998 ;
  assign y5274 = n12000 ;
  assign y5275 = ~1'b0 ;
  assign y5276 = n12004 ;
  assign y5277 = ~n12005 ;
  assign y5278 = ~n12008 ;
  assign y5279 = ~1'b0 ;
  assign y5280 = n12010 ;
  assign y5281 = ~n12014 ;
  assign y5282 = ~1'b0 ;
  assign y5283 = ~1'b0 ;
  assign y5284 = ~n12016 ;
  assign y5285 = n12021 ;
  assign y5286 = n12022 ;
  assign y5287 = ~n12025 ;
  assign y5288 = n12028 ;
  assign y5289 = ~n12034 ;
  assign y5290 = ~n12038 ;
  assign y5291 = ~1'b0 ;
  assign y5292 = ~n12048 ;
  assign y5293 = ~1'b0 ;
  assign y5294 = ~n12051 ;
  assign y5295 = ~n12057 ;
  assign y5296 = n12058 ;
  assign y5297 = n12061 ;
  assign y5298 = ~1'b0 ;
  assign y5299 = n12062 ;
  assign y5300 = n12063 ;
  assign y5301 = ~n12065 ;
  assign y5302 = ~1'b0 ;
  assign y5303 = ~n12068 ;
  assign y5304 = ~n12070 ;
  assign y5305 = ~1'b0 ;
  assign y5306 = ~n12073 ;
  assign y5307 = n12076 ;
  assign y5308 = n12080 ;
  assign y5309 = ~n12082 ;
  assign y5310 = n12086 ;
  assign y5311 = ~n12088 ;
  assign y5312 = ~n12095 ;
  assign y5313 = ~1'b0 ;
  assign y5314 = ~n12099 ;
  assign y5315 = ~1'b0 ;
  assign y5316 = ~1'b0 ;
  assign y5317 = ~n12100 ;
  assign y5318 = ~1'b0 ;
  assign y5319 = ~n12101 ;
  assign y5320 = n12102 ;
  assign y5321 = ~n12106 ;
  assign y5322 = ~n12107 ;
  assign y5323 = ~n12108 ;
  assign y5324 = ~1'b0 ;
  assign y5325 = n12112 ;
  assign y5326 = ~n12115 ;
  assign y5327 = n12116 ;
  assign y5328 = ~n12124 ;
  assign y5329 = n12128 ;
  assign y5330 = ~n12133 ;
  assign y5331 = n12135 ;
  assign y5332 = ~1'b0 ;
  assign y5333 = n12138 ;
  assign y5334 = ~n7790 ;
  assign y5335 = n12142 ;
  assign y5336 = ~n12112 ;
  assign y5337 = ~n12150 ;
  assign y5338 = ~n12151 ;
  assign y5339 = ~1'b0 ;
  assign y5340 = n12153 ;
  assign y5341 = ~n12162 ;
  assign y5342 = n12164 ;
  assign y5343 = ~1'b0 ;
  assign y5344 = ~n12171 ;
  assign y5345 = ~n12173 ;
  assign y5346 = ~n12174 ;
  assign y5347 = ~n12177 ;
  assign y5348 = ~n12178 ;
  assign y5349 = ~n12180 ;
  assign y5350 = ~n12183 ;
  assign y5351 = n12186 ;
  assign y5352 = ~n12187 ;
  assign y5353 = ~1'b0 ;
  assign y5354 = ~1'b0 ;
  assign y5355 = n12190 ;
  assign y5356 = ~1'b0 ;
  assign y5357 = n12192 ;
  assign y5358 = n12194 ;
  assign y5359 = 1'b0 ;
  assign y5360 = n2319 ;
  assign y5361 = ~n7295 ;
  assign y5362 = n12196 ;
  assign y5363 = ~n8962 ;
  assign y5364 = n12199 ;
  assign y5365 = ~n12200 ;
  assign y5366 = ~n6433 ;
  assign y5367 = ~n12204 ;
  assign y5368 = ~1'b0 ;
  assign y5369 = ~n12208 ;
  assign y5370 = ~n12211 ;
  assign y5371 = n12212 ;
  assign y5372 = ~1'b0 ;
  assign y5373 = ~n12213 ;
  assign y5374 = n8815 ;
  assign y5375 = ~n12217 ;
  assign y5376 = n12219 ;
  assign y5377 = n12224 ;
  assign y5378 = ~n12225 ;
  assign y5379 = n12229 ;
  assign y5380 = n12231 ;
  assign y5381 = 1'b0 ;
  assign y5382 = ~n10459 ;
  assign y5383 = ~n12233 ;
  assign y5384 = ~1'b0 ;
  assign y5385 = ~n12234 ;
  assign y5386 = ~n12235 ;
  assign y5387 = ~1'b0 ;
  assign y5388 = n12243 ;
  assign y5389 = ~1'b0 ;
  assign y5390 = n12245 ;
  assign y5391 = ~n12249 ;
  assign y5392 = ~n12253 ;
  assign y5393 = n12257 ;
  assign y5394 = ~n12258 ;
  assign y5395 = ~1'b0 ;
  assign y5396 = ~n10537 ;
  assign y5397 = ~n12262 ;
  assign y5398 = ~1'b0 ;
  assign y5399 = n12267 ;
  assign y5400 = ~1'b0 ;
  assign y5401 = ~1'b0 ;
  assign y5402 = ~1'b0 ;
  assign y5403 = n12269 ;
  assign y5404 = ~n5024 ;
  assign y5405 = ~1'b0 ;
  assign y5406 = ~1'b0 ;
  assign y5407 = n12271 ;
  assign y5408 = ~n12276 ;
  assign y5409 = n12279 ;
  assign y5410 = ~n12283 ;
  assign y5411 = ~n12284 ;
  assign y5412 = n12287 ;
  assign y5413 = ~n12288 ;
  assign y5414 = ~n12293 ;
  assign y5415 = n12296 ;
  assign y5416 = ~1'b0 ;
  assign y5417 = ~n12301 ;
  assign y5418 = n12305 ;
  assign y5419 = n12313 ;
  assign y5420 = ~1'b0 ;
  assign y5421 = n12320 ;
  assign y5422 = n12321 ;
  assign y5423 = ~n12322 ;
  assign y5424 = n12328 ;
  assign y5425 = n11764 ;
  assign y5426 = ~1'b0 ;
  assign y5427 = ~n12333 ;
  assign y5428 = 1'b0 ;
  assign y5429 = n12340 ;
  assign y5430 = ~1'b0 ;
  assign y5431 = ~n12342 ;
  assign y5432 = n12343 ;
  assign y5433 = n12349 ;
  assign y5434 = n12351 ;
  assign y5435 = n12362 ;
  assign y5436 = ~n12363 ;
  assign y5437 = n12364 ;
  assign y5438 = ~n12366 ;
  assign y5439 = ~n12372 ;
  assign y5440 = ~1'b0 ;
  assign y5441 = ~n12374 ;
  assign y5442 = ~n12378 ;
  assign y5443 = n12379 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = ~1'b0 ;
  assign y5446 = n12384 ;
  assign y5447 = n12385 ;
  assign y5448 = n12388 ;
  assign y5449 = ~n12390 ;
  assign y5450 = n12391 ;
  assign y5451 = n12395 ;
  assign y5452 = ~n12399 ;
  assign y5453 = 1'b0 ;
  assign y5454 = n12400 ;
  assign y5455 = ~1'b0 ;
  assign y5456 = ~1'b0 ;
  assign y5457 = ~n12403 ;
  assign y5458 = 1'b0 ;
  assign y5459 = ~n12405 ;
  assign y5460 = n12406 ;
  assign y5461 = n10453 ;
  assign y5462 = ~n12410 ;
  assign y5463 = 1'b0 ;
  assign y5464 = ~n12414 ;
  assign y5465 = n12416 ;
  assign y5466 = ~n12422 ;
  assign y5467 = ~n7008 ;
  assign y5468 = n12432 ;
  assign y5469 = n12433 ;
  assign y5470 = ~n12437 ;
  assign y5471 = n12439 ;
  assign y5472 = n5932 ;
  assign y5473 = ~n12442 ;
  assign y5474 = ~1'b0 ;
  assign y5475 = ~n12444 ;
  assign y5476 = n12447 ;
  assign y5477 = n12452 ;
  assign y5478 = ~n12459 ;
  assign y5479 = 1'b0 ;
  assign y5480 = ~n12463 ;
  assign y5481 = n12465 ;
  assign y5482 = ~n12477 ;
  assign y5483 = ~1'b0 ;
  assign y5484 = ~n12478 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = ~n12480 ;
  assign y5487 = n12481 ;
  assign y5488 = n9453 ;
  assign y5489 = ~1'b0 ;
  assign y5490 = ~n12482 ;
  assign y5491 = ~n12487 ;
  assign y5492 = ~n12488 ;
  assign y5493 = ~n10129 ;
  assign y5494 = ~n12489 ;
  assign y5495 = n12490 ;
  assign y5496 = n12495 ;
  assign y5497 = n12497 ;
  assign y5498 = ~1'b0 ;
  assign y5499 = n976 ;
  assign y5500 = ~n12504 ;
  assign y5501 = ~1'b0 ;
  assign y5502 = n12510 ;
  assign y5503 = n11974 ;
  assign y5504 = ~1'b0 ;
  assign y5505 = ~1'b0 ;
  assign y5506 = n12514 ;
  assign y5507 = n12525 ;
  assign y5508 = ~n12531 ;
  assign y5509 = n12535 ;
  assign y5510 = ~n12537 ;
  assign y5511 = n12539 ;
  assign y5512 = ~1'b0 ;
  assign y5513 = n12540 ;
  assign y5514 = n12545 ;
  assign y5515 = n12549 ;
  assign y5516 = ~1'b0 ;
  assign y5517 = n12551 ;
  assign y5518 = ~n12554 ;
  assign y5519 = n12556 ;
  assign y5520 = n12557 ;
  assign y5521 = ~1'b0 ;
  assign y5522 = ~n12564 ;
  assign y5523 = ~n12568 ;
  assign y5524 = ~1'b0 ;
  assign y5525 = ~n12573 ;
  assign y5526 = n12575 ;
  assign y5527 = ~n12581 ;
  assign y5528 = n12585 ;
  assign y5529 = n12587 ;
  assign y5530 = ~n12590 ;
  assign y5531 = n12593 ;
  assign y5532 = ~n12249 ;
  assign y5533 = ~n12597 ;
  assign y5534 = n12600 ;
  assign y5535 = n12601 ;
  assign y5536 = n12604 ;
  assign y5537 = n12607 ;
  assign y5538 = n12608 ;
  assign y5539 = ~n12610 ;
  assign y5540 = ~n12616 ;
  assign y5541 = n12617 ;
  assign y5542 = n12618 ;
  assign y5543 = ~n12623 ;
  assign y5544 = ~n12629 ;
  assign y5545 = n12630 ;
  assign y5546 = ~n12633 ;
  assign y5547 = n12637 ;
  assign y5548 = ~n12638 ;
  assign y5549 = ~1'b0 ;
  assign y5550 = ~1'b0 ;
  assign y5551 = n12639 ;
  assign y5552 = ~1'b0 ;
  assign y5553 = n12642 ;
  assign y5554 = ~n12645 ;
  assign y5555 = ~n12652 ;
  assign y5556 = n12654 ;
  assign y5557 = ~n12657 ;
  assign y5558 = ~n12659 ;
  assign y5559 = n12661 ;
  assign y5560 = ~n12665 ;
  assign y5561 = ~1'b0 ;
  assign y5562 = ~1'b0 ;
  assign y5563 = 1'b0 ;
  assign y5564 = n12671 ;
  assign y5565 = n12674 ;
  assign y5566 = ~1'b0 ;
  assign y5567 = n12678 ;
  assign y5568 = n12679 ;
  assign y5569 = ~1'b0 ;
  assign y5570 = ~n12680 ;
  assign y5571 = n12683 ;
  assign y5572 = n12684 ;
  assign y5573 = ~1'b0 ;
  assign y5574 = ~1'b0 ;
  assign y5575 = n12685 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = ~n12687 ;
  assign y5578 = n12688 ;
  assign y5579 = n12691 ;
  assign y5580 = ~n12694 ;
  assign y5581 = ~n12695 ;
  assign y5582 = n12697 ;
  assign y5583 = ~1'b0 ;
  assign y5584 = n12698 ;
  assign y5585 = ~n12701 ;
  assign y5586 = ~1'b0 ;
  assign y5587 = ~1'b0 ;
  assign y5588 = ~n12702 ;
  assign y5589 = n12709 ;
  assign y5590 = n12712 ;
  assign y5591 = n12713 ;
  assign y5592 = ~1'b0 ;
  assign y5593 = ~n12717 ;
  assign y5594 = n2449 ;
  assign y5595 = ~n12718 ;
  assign y5596 = ~n12722 ;
  assign y5597 = ~n12723 ;
  assign y5598 = ~1'b0 ;
  assign y5599 = ~1'b0 ;
  assign y5600 = n12727 ;
  assign y5601 = n12730 ;
  assign y5602 = ~n3773 ;
  assign y5603 = ~n12732 ;
  assign y5604 = ~n12737 ;
  assign y5605 = ~n4769 ;
  assign y5606 = n12744 ;
  assign y5607 = n12745 ;
  assign y5608 = ~n523 ;
  assign y5609 = n12746 ;
  assign y5610 = n1807 ;
  assign y5611 = ~1'b0 ;
  assign y5612 = ~1'b0 ;
  assign y5613 = ~n12747 ;
  assign y5614 = n12750 ;
  assign y5615 = ~1'b0 ;
  assign y5616 = n11345 ;
  assign y5617 = n12752 ;
  assign y5618 = ~n12755 ;
  assign y5619 = ~1'b0 ;
  assign y5620 = ~n12758 ;
  assign y5621 = n12759 ;
  assign y5622 = n3067 ;
  assign y5623 = ~1'b0 ;
  assign y5624 = ~n12768 ;
  assign y5625 = ~1'b0 ;
  assign y5626 = ~n12777 ;
  assign y5627 = ~1'b0 ;
  assign y5628 = n12787 ;
  assign y5629 = ~n12788 ;
  assign y5630 = ~1'b0 ;
  assign y5631 = n12793 ;
  assign y5632 = ~1'b0 ;
  assign y5633 = ~n12797 ;
  assign y5634 = n12800 ;
  assign y5635 = n12802 ;
  assign y5636 = ~1'b0 ;
  assign y5637 = ~n12805 ;
  assign y5638 = n12807 ;
  assign y5639 = n12808 ;
  assign y5640 = ~n12817 ;
  assign y5641 = ~n12818 ;
  assign y5642 = ~n5342 ;
  assign y5643 = ~1'b0 ;
  assign y5644 = ~1'b0 ;
  assign y5645 = ~1'b0 ;
  assign y5646 = n12820 ;
  assign y5647 = ~1'b0 ;
  assign y5648 = ~1'b0 ;
  assign y5649 = ~1'b0 ;
  assign y5650 = n12822 ;
  assign y5651 = n12823 ;
  assign y5652 = ~n12828 ;
  assign y5653 = ~n12833 ;
  assign y5654 = n12836 ;
  assign y5655 = ~n12839 ;
  assign y5656 = n12845 ;
  assign y5657 = n12847 ;
  assign y5658 = ~n12850 ;
  assign y5659 = ~n12851 ;
  assign y5660 = n12857 ;
  assign y5661 = n12860 ;
  assign y5662 = n12864 ;
  assign y5663 = ~1'b0 ;
  assign y5664 = n12870 ;
  assign y5665 = ~1'b0 ;
  assign y5666 = ~n12873 ;
  assign y5667 = n12874 ;
  assign y5668 = n9439 ;
  assign y5669 = ~1'b0 ;
  assign y5670 = 1'b0 ;
  assign y5671 = ~n12875 ;
  assign y5672 = ~n12878 ;
  assign y5673 = n12884 ;
  assign y5674 = n12886 ;
  assign y5675 = n12889 ;
  assign y5676 = ~n12893 ;
  assign y5677 = n12906 ;
  assign y5678 = n12909 ;
  assign y5679 = ~1'b0 ;
  assign y5680 = n12920 ;
  assign y5681 = n12921 ;
  assign y5682 = ~n12925 ;
  assign y5683 = 1'b0 ;
  assign y5684 = ~n12927 ;
  assign y5685 = n12928 ;
  assign y5686 = ~n12929 ;
  assign y5687 = ~n12932 ;
  assign y5688 = ~n12934 ;
  assign y5689 = ~1'b0 ;
  assign y5690 = ~1'b0 ;
  assign y5691 = n12938 ;
  assign y5692 = n12942 ;
  assign y5693 = ~1'b0 ;
  assign y5694 = ~n12943 ;
  assign y5695 = ~n12574 ;
  assign y5696 = ~n12950 ;
  assign y5697 = n12956 ;
  assign y5698 = n12957 ;
  assign y5699 = n12960 ;
  assign y5700 = 1'b0 ;
  assign y5701 = n12963 ;
  assign y5702 = n12965 ;
  assign y5703 = ~n12967 ;
  assign y5704 = n4339 ;
  assign y5705 = ~n12975 ;
  assign y5706 = ~1'b0 ;
  assign y5707 = ~n12980 ;
  assign y5708 = ~n12983 ;
  assign y5709 = ~1'b0 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = ~n12985 ;
  assign y5712 = ~1'b0 ;
  assign y5713 = n12986 ;
  assign y5714 = ~n12988 ;
  assign y5715 = n12989 ;
  assign y5716 = n12088 ;
  assign y5717 = n12992 ;
  assign y5718 = ~n12998 ;
  assign y5719 = ~n12999 ;
  assign y5720 = n13006 ;
  assign y5721 = 1'b0 ;
  assign y5722 = ~n13010 ;
  assign y5723 = ~n13011 ;
  assign y5724 = ~n13017 ;
  assign y5725 = ~n13019 ;
  assign y5726 = ~n13021 ;
  assign y5727 = ~n13023 ;
  assign y5728 = ~1'b0 ;
  assign y5729 = ~n13028 ;
  assign y5730 = ~1'b0 ;
  assign y5731 = n13035 ;
  assign y5732 = ~n13038 ;
  assign y5733 = n13042 ;
  assign y5734 = ~1'b0 ;
  assign y5735 = ~n13047 ;
  assign y5736 = ~1'b0 ;
  assign y5737 = ~n13051 ;
  assign y5738 = ~1'b0 ;
  assign y5739 = ~n13063 ;
  assign y5740 = ~1'b0 ;
  assign y5741 = n13064 ;
  assign y5742 = ~1'b0 ;
  assign y5743 = ~1'b0 ;
  assign y5744 = ~n13071 ;
  assign y5745 = ~n13080 ;
  assign y5746 = n13084 ;
  assign y5747 = ~1'b0 ;
  assign y5748 = n13089 ;
  assign y5749 = ~n13090 ;
  assign y5750 = n13093 ;
  assign y5751 = ~n13096 ;
  assign y5752 = ~n13097 ;
  assign y5753 = ~n13106 ;
  assign y5754 = ~n13108 ;
  assign y5755 = n13110 ;
  assign y5756 = ~n13114 ;
  assign y5757 = n13116 ;
  assign y5758 = ~1'b0 ;
  assign y5759 = n13117 ;
  assign y5760 = ~n13119 ;
  assign y5761 = ~1'b0 ;
  assign y5762 = ~1'b0 ;
  assign y5763 = ~n13122 ;
  assign y5764 = ~n13127 ;
  assign y5765 = n13129 ;
  assign y5766 = ~n13137 ;
  assign y5767 = n13138 ;
  assign y5768 = ~n13139 ;
  assign y5769 = ~n13141 ;
  assign y5770 = n13145 ;
  assign y5771 = n13147 ;
  assign y5772 = n12779 ;
  assign y5773 = n13148 ;
  assign y5774 = n13149 ;
  assign y5775 = 1'b0 ;
  assign y5776 = ~n13154 ;
  assign y5777 = n13158 ;
  assign y5778 = ~n13160 ;
  assign y5779 = n13162 ;
  assign y5780 = ~n13164 ;
  assign y5781 = 1'b0 ;
  assign y5782 = n13170 ;
  assign y5783 = ~n13174 ;
  assign y5784 = ~1'b0 ;
  assign y5785 = n13179 ;
  assign y5786 = n13182 ;
  assign y5787 = n13193 ;
  assign y5788 = n13195 ;
  assign y5789 = ~n13196 ;
  assign y5790 = ~1'b0 ;
  assign y5791 = ~n13197 ;
  assign y5792 = ~n13199 ;
  assign y5793 = ~1'b0 ;
  assign y5794 = n13201 ;
  assign y5795 = ~1'b0 ;
  assign y5796 = n13202 ;
  assign y5797 = n13208 ;
  assign y5798 = n13211 ;
  assign y5799 = ~1'b0 ;
  assign y5800 = ~n13213 ;
  assign y5801 = ~n13217 ;
  assign y5802 = n13223 ;
  assign y5803 = ~n13231 ;
  assign y5804 = ~n13232 ;
  assign y5805 = ~1'b0 ;
  assign y5806 = 1'b0 ;
  assign y5807 = n13237 ;
  assign y5808 = ~1'b0 ;
  assign y5809 = n13238 ;
  assign y5810 = ~n13242 ;
  assign y5811 = n13247 ;
  assign y5812 = ~1'b0 ;
  assign y5813 = ~n13249 ;
  assign y5814 = ~n13251 ;
  assign y5815 = n13261 ;
  assign y5816 = ~1'b0 ;
  assign y5817 = ~n10379 ;
  assign y5818 = n13262 ;
  assign y5819 = ~1'b0 ;
  assign y5820 = ~n13266 ;
  assign y5821 = n13268 ;
  assign y5822 = ~1'b0 ;
  assign y5823 = n13272 ;
  assign y5824 = n13280 ;
  assign y5825 = n5311 ;
  assign y5826 = ~1'b0 ;
  assign y5827 = ~n9120 ;
  assign y5828 = n13282 ;
  assign y5829 = ~1'b0 ;
  assign y5830 = n13285 ;
  assign y5831 = n5144 ;
  assign y5832 = ~n13289 ;
  assign y5833 = ~1'b0 ;
  assign y5834 = n177 ;
  assign y5835 = n13293 ;
  assign y5836 = ~n13300 ;
  assign y5837 = ~n13303 ;
  assign y5838 = n13307 ;
  assign y5839 = ~n6167 ;
  assign y5840 = ~1'b0 ;
  assign y5841 = n13308 ;
  assign y5842 = n13312 ;
  assign y5843 = n13317 ;
  assign y5844 = ~n13322 ;
  assign y5845 = ~1'b0 ;
  assign y5846 = ~n13327 ;
  assign y5847 = n13332 ;
  assign y5848 = ~n13335 ;
  assign y5849 = n13337 ;
  assign y5850 = ~n13340 ;
  assign y5851 = ~n13342 ;
  assign y5852 = n13343 ;
  assign y5853 = ~n13348 ;
  assign y5854 = n13352 ;
  assign y5855 = ~n13354 ;
  assign y5856 = 1'b0 ;
  assign y5857 = ~n13364 ;
  assign y5858 = ~n13365 ;
  assign y5859 = ~1'b0 ;
  assign y5860 = ~n13370 ;
  assign y5861 = n13372 ;
  assign y5862 = n13380 ;
  assign y5863 = ~n13385 ;
  assign y5864 = n13388 ;
  assign y5865 = n8907 ;
  assign y5866 = n13390 ;
  assign y5867 = ~1'b0 ;
  assign y5868 = n13393 ;
  assign y5869 = n13394 ;
  assign y5870 = ~1'b0 ;
  assign y5871 = ~1'b0 ;
  assign y5872 = ~n13399 ;
  assign y5873 = ~1'b0 ;
  assign y5874 = ~1'b0 ;
  assign y5875 = ~1'b0 ;
  assign y5876 = ~1'b0 ;
  assign y5877 = n12002 ;
  assign y5878 = ~n13407 ;
  assign y5879 = ~1'b0 ;
  assign y5880 = n13408 ;
  assign y5881 = n13413 ;
  assign y5882 = 1'b0 ;
  assign y5883 = ~1'b0 ;
  assign y5884 = ~n13418 ;
  assign y5885 = n13422 ;
  assign y5886 = ~n13426 ;
  assign y5887 = ~1'b0 ;
  assign y5888 = ~1'b0 ;
  assign y5889 = ~1'b0 ;
  assign y5890 = n13427 ;
  assign y5891 = n13428 ;
  assign y5892 = ~1'b0 ;
  assign y5893 = n13432 ;
  assign y5894 = n11219 ;
  assign y5895 = n13433 ;
  assign y5896 = ~n13435 ;
  assign y5897 = ~1'b0 ;
  assign y5898 = ~1'b0 ;
  assign y5899 = ~1'b0 ;
  assign y5900 = n13442 ;
  assign y5901 = n13443 ;
  assign y5902 = n13445 ;
  assign y5903 = ~n1805 ;
  assign y5904 = ~n13449 ;
  assign y5905 = n13451 ;
  assign y5906 = ~1'b0 ;
  assign y5907 = ~1'b0 ;
  assign y5908 = ~n13453 ;
  assign y5909 = n13456 ;
  assign y5910 = ~n13457 ;
  assign y5911 = n13459 ;
  assign y5912 = ~n13461 ;
  assign y5913 = ~n9226 ;
  assign y5914 = ~n13462 ;
  assign y5915 = ~n13465 ;
  assign y5916 = ~n13467 ;
  assign y5917 = n13470 ;
  assign y5918 = n13475 ;
  assign y5919 = ~1'b0 ;
  assign y5920 = ~1'b0 ;
  assign y5921 = ~1'b0 ;
  assign y5922 = 1'b0 ;
  assign y5923 = ~1'b0 ;
  assign y5924 = n6142 ;
  assign y5925 = n13486 ;
  assign y5926 = ~n13488 ;
  assign y5927 = n13489 ;
  assign y5928 = n13490 ;
  assign y5929 = n13498 ;
  assign y5930 = ~1'b0 ;
  assign y5931 = ~n13504 ;
  assign y5932 = ~n13508 ;
  assign y5933 = n13513 ;
  assign y5934 = ~1'b0 ;
  assign y5935 = ~1'b0 ;
  assign y5936 = n13516 ;
  assign y5937 = ~1'b0 ;
  assign y5938 = ~1'b0 ;
  assign y5939 = ~1'b0 ;
  assign y5940 = ~n9072 ;
  assign y5941 = 1'b0 ;
  assign y5942 = ~1'b0 ;
  assign y5943 = n13517 ;
  assign y5944 = n13520 ;
  assign y5945 = n13521 ;
  assign y5946 = ~n13524 ;
  assign y5947 = ~1'b0 ;
  assign y5948 = n13526 ;
  assign y5949 = ~n13530 ;
  assign y5950 = ~1'b0 ;
  assign y5951 = n13533 ;
  assign y5952 = n13538 ;
  assign y5953 = ~n13541 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = n13542 ;
  assign y5956 = n13544 ;
  assign y5957 = ~n13545 ;
  assign y5958 = ~n13547 ;
  assign y5959 = ~n13548 ;
  assign y5960 = ~n13549 ;
  assign y5961 = ~n11551 ;
  assign y5962 = ~n13552 ;
  assign y5963 = ~1'b0 ;
  assign y5964 = n7047 ;
  assign y5965 = ~1'b0 ;
  assign y5966 = ~n13554 ;
  assign y5967 = ~1'b0 ;
  assign y5968 = ~n13556 ;
  assign y5969 = n13557 ;
  assign y5970 = ~1'b0 ;
  assign y5971 = ~n13560 ;
  assign y5972 = n13561 ;
  assign y5973 = ~n13563 ;
  assign y5974 = ~n13565 ;
  assign y5975 = ~n13569 ;
  assign y5976 = ~n13572 ;
  assign y5977 = n13574 ;
  assign y5978 = ~n13578 ;
  assign y5979 = ~n13582 ;
  assign y5980 = ~1'b0 ;
  assign y5981 = n13583 ;
  assign y5982 = ~1'b0 ;
  assign y5983 = ~n13585 ;
  assign y5984 = n13586 ;
  assign y5985 = ~n13593 ;
  assign y5986 = n13595 ;
  assign y5987 = n13597 ;
  assign y5988 = ~1'b0 ;
  assign y5989 = n13603 ;
  assign y5990 = ~n13607 ;
  assign y5991 = ~n13608 ;
  assign y5992 = n13609 ;
  assign y5993 = ~n13614 ;
  assign y5994 = n13617 ;
  assign y5995 = n13619 ;
  assign y5996 = ~n13625 ;
  assign y5997 = ~n13626 ;
  assign y5998 = ~n13629 ;
  assign y5999 = ~n13634 ;
  assign y6000 = n13637 ;
  assign y6001 = ~1'b0 ;
  assign y6002 = n13642 ;
  assign y6003 = n13648 ;
  assign y6004 = n13649 ;
  assign y6005 = ~n13651 ;
  assign y6006 = ~n13654 ;
  assign y6007 = ~n13658 ;
  assign y6008 = ~1'b0 ;
  assign y6009 = n13660 ;
  assign y6010 = ~n13661 ;
  assign y6011 = n13665 ;
  assign y6012 = n13667 ;
  assign y6013 = ~n13668 ;
  assign y6014 = ~n13671 ;
  assign y6015 = ~1'b0 ;
  assign y6016 = n13673 ;
  assign y6017 = ~n13678 ;
  assign y6018 = ~1'b0 ;
  assign y6019 = ~1'b0 ;
  assign y6020 = ~n13679 ;
  assign y6021 = n3784 ;
  assign y6022 = n13688 ;
  assign y6023 = n9221 ;
  assign y6024 = n13694 ;
  assign y6025 = ~n13698 ;
  assign y6026 = n13699 ;
  assign y6027 = ~n13702 ;
  assign y6028 = ~n13706 ;
  assign y6029 = ~1'b0 ;
  assign y6030 = n13713 ;
  assign y6031 = ~1'b0 ;
  assign y6032 = ~n13714 ;
  assign y6033 = ~1'b0 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = ~1'b0 ;
  assign y6036 = n13719 ;
  assign y6037 = n13720 ;
  assign y6038 = ~n13727 ;
  assign y6039 = n13733 ;
  assign y6040 = ~n13735 ;
  assign y6041 = n13736 ;
  assign y6042 = n13741 ;
  assign y6043 = ~1'b0 ;
  assign y6044 = ~n13747 ;
  assign y6045 = ~1'b0 ;
  assign y6046 = ~n13748 ;
  assign y6047 = ~n13749 ;
  assign y6048 = ~1'b0 ;
  assign y6049 = ~n13757 ;
  assign y6050 = n13760 ;
  assign y6051 = ~n13761 ;
  assign y6052 = n13762 ;
  assign y6053 = ~n13768 ;
  assign y6054 = n13770 ;
  assign y6055 = ~n13775 ;
  assign y6056 = n13777 ;
  assign y6057 = n6455 ;
  assign y6058 = ~1'b0 ;
  assign y6059 = n13783 ;
  assign y6060 = ~n13785 ;
  assign y6061 = n13806 ;
  assign y6062 = 1'b0 ;
  assign y6063 = ~1'b0 ;
  assign y6064 = ~n2946 ;
  assign y6065 = n13808 ;
  assign y6066 = n13810 ;
  assign y6067 = n13812 ;
  assign y6068 = n13813 ;
  assign y6069 = ~1'b0 ;
  assign y6070 = n13817 ;
  assign y6071 = ~1'b0 ;
  assign y6072 = n13818 ;
  assign y6073 = n13441 ;
  assign y6074 = ~n13819 ;
  assign y6075 = n13829 ;
  assign y6076 = n13842 ;
  assign y6077 = ~n13845 ;
  assign y6078 = ~n13846 ;
  assign y6079 = n13849 ;
  assign y6080 = n13850 ;
  assign y6081 = ~n13853 ;
  assign y6082 = ~n13858 ;
  assign y6083 = n13859 ;
  assign y6084 = ~1'b0 ;
  assign y6085 = ~1'b0 ;
  assign y6086 = ~1'b0 ;
  assign y6087 = ~n13862 ;
  assign y6088 = n13870 ;
  assign y6089 = ~n13873 ;
  assign y6090 = ~n13878 ;
  assign y6091 = ~n13884 ;
  assign y6092 = ~1'b0 ;
  assign y6093 = ~n13887 ;
  assign y6094 = ~1'b0 ;
  assign y6095 = ~n13895 ;
  assign y6096 = n9125 ;
  assign y6097 = n13900 ;
  assign y6098 = n13902 ;
  assign y6099 = ~n13903 ;
  assign y6100 = ~1'b0 ;
  assign y6101 = n13907 ;
  assign y6102 = n13913 ;
  assign y6103 = n13914 ;
  assign y6104 = ~1'b0 ;
  assign y6105 = ~n13916 ;
  assign y6106 = n13920 ;
  assign y6107 = ~n13931 ;
  assign y6108 = ~1'b0 ;
  assign y6109 = n13934 ;
  assign y6110 = ~1'b0 ;
  assign y6111 = n13941 ;
  assign y6112 = n13942 ;
  assign y6113 = ~n12421 ;
  assign y6114 = ~1'b0 ;
  assign y6115 = n13951 ;
  assign y6116 = 1'b0 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = ~n13954 ;
  assign y6119 = n13962 ;
  assign y6120 = n13963 ;
  assign y6121 = ~n13965 ;
  assign y6122 = n13970 ;
  assign y6123 = n13979 ;
  assign y6124 = ~1'b0 ;
  assign y6125 = ~n13982 ;
  assign y6126 = ~1'b0 ;
  assign y6127 = ~n13990 ;
  assign y6128 = ~n13991 ;
  assign y6129 = ~n13995 ;
  assign y6130 = n13999 ;
  assign y6131 = n14001 ;
  assign y6132 = n14005 ;
  assign y6133 = n14007 ;
  assign y6134 = n14009 ;
  assign y6135 = n517 ;
  assign y6136 = ~n14014 ;
  assign y6137 = ~1'b0 ;
  assign y6138 = ~n14019 ;
  assign y6139 = ~1'b0 ;
  assign y6140 = ~1'b0 ;
  assign y6141 = ~n14024 ;
  assign y6142 = ~1'b0 ;
  assign y6143 = ~n14035 ;
  assign y6144 = n14037 ;
  assign y6145 = ~n14043 ;
  assign y6146 = n14047 ;
  assign y6147 = ~n14048 ;
  assign y6148 = ~n14054 ;
  assign y6149 = n14063 ;
  assign y6150 = n8659 ;
  assign y6151 = ~n14065 ;
  assign y6152 = ~1'b0 ;
  assign y6153 = ~1'b0 ;
  assign y6154 = n14068 ;
  assign y6155 = ~n14080 ;
  assign y6156 = n14088 ;
  assign y6157 = n14091 ;
  assign y6158 = n14094 ;
  assign y6159 = ~n14098 ;
  assign y6160 = ~n14100 ;
  assign y6161 = ~1'b0 ;
  assign y6162 = n14104 ;
  assign y6163 = ~n14109 ;
  assign y6164 = ~n14110 ;
  assign y6165 = ~n14121 ;
  assign y6166 = n14125 ;
  assign y6167 = ~n14127 ;
  assign y6168 = n14135 ;
  assign y6169 = ~1'b0 ;
  assign y6170 = ~1'b0 ;
  assign y6171 = n8885 ;
  assign y6172 = ~n14139 ;
  assign y6173 = ~n14144 ;
  assign y6174 = ~n14150 ;
  assign y6175 = n14151 ;
  assign y6176 = ~1'b0 ;
  assign y6177 = n14152 ;
  assign y6178 = n14153 ;
  assign y6179 = n14157 ;
  assign y6180 = n14158 ;
  assign y6181 = ~n14159 ;
  assign y6182 = ~1'b0 ;
  assign y6183 = n14161 ;
  assign y6184 = ~1'b0 ;
  assign y6185 = ~1'b0 ;
  assign y6186 = ~1'b0 ;
  assign y6187 = ~n14162 ;
  assign y6188 = ~1'b0 ;
  assign y6189 = ~n14164 ;
  assign y6190 = n14166 ;
  assign y6191 = n14172 ;
  assign y6192 = ~n14173 ;
  assign y6193 = n14175 ;
  assign y6194 = ~n8881 ;
  assign y6195 = n14178 ;
  assign y6196 = ~n14179 ;
  assign y6197 = n14181 ;
  assign y6198 = n14189 ;
  assign y6199 = ~n14193 ;
  assign y6200 = n14198 ;
  assign y6201 = n14208 ;
  assign y6202 = ~1'b0 ;
  assign y6203 = n14212 ;
  assign y6204 = ~n14214 ;
  assign y6205 = n14216 ;
  assign y6206 = ~1'b0 ;
  assign y6207 = ~n14218 ;
  assign y6208 = ~n3282 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = n14220 ;
  assign y6211 = n14226 ;
  assign y6212 = n14227 ;
  assign y6213 = n12698 ;
  assign y6214 = 1'b0 ;
  assign y6215 = n14236 ;
  assign y6216 = ~n14239 ;
  assign y6217 = n1043 ;
  assign y6218 = n14241 ;
  assign y6219 = n14243 ;
  assign y6220 = ~n14249 ;
  assign y6221 = ~n14251 ;
  assign y6222 = ~1'b0 ;
  assign y6223 = ~1'b0 ;
  assign y6224 = ~n14252 ;
  assign y6225 = n14254 ;
  assign y6226 = n14255 ;
  assign y6227 = n14257 ;
  assign y6228 = n14259 ;
  assign y6229 = ~n7354 ;
  assign y6230 = ~n14261 ;
  assign y6231 = ~n14263 ;
  assign y6232 = n13992 ;
  assign y6233 = n14264 ;
  assign y6234 = n9716 ;
  assign y6235 = ~1'b0 ;
  assign y6236 = ~1'b0 ;
  assign y6237 = n14266 ;
  assign y6238 = ~n3908 ;
  assign y6239 = n14270 ;
  assign y6240 = ~n14275 ;
  assign y6241 = ~n14278 ;
  assign y6242 = ~1'b0 ;
  assign y6243 = ~n14281 ;
  assign y6244 = ~1'b0 ;
  assign y6245 = n14287 ;
  assign y6246 = n14288 ;
  assign y6247 = ~1'b0 ;
  assign y6248 = n12402 ;
  assign y6249 = ~n14290 ;
  assign y6250 = ~1'b0 ;
  assign y6251 = ~1'b0 ;
  assign y6252 = n14293 ;
  assign y6253 = ~n14296 ;
  assign y6254 = n14298 ;
  assign y6255 = n14301 ;
  assign y6256 = n14303 ;
  assign y6257 = ~n14307 ;
  assign y6258 = ~n14310 ;
  assign y6259 = n14313 ;
  assign y6260 = ~n14316 ;
  assign y6261 = n14323 ;
  assign y6262 = n14324 ;
  assign y6263 = ~n14326 ;
  assign y6264 = ~n14329 ;
  assign y6265 = ~n14333 ;
  assign y6266 = n14335 ;
  assign y6267 = ~n14337 ;
  assign y6268 = ~n14342 ;
  assign y6269 = n14343 ;
  assign y6270 = ~n14344 ;
  assign y6271 = ~n14348 ;
  assign y6272 = ~1'b0 ;
  assign y6273 = ~n14351 ;
  assign y6274 = ~1'b0 ;
  assign y6275 = ~n14356 ;
  assign y6276 = n14364 ;
  assign y6277 = n14366 ;
  assign y6278 = n14367 ;
  assign y6279 = ~1'b0 ;
  assign y6280 = n14371 ;
  assign y6281 = ~n14374 ;
  assign y6282 = ~n14377 ;
  assign y6283 = n14378 ;
  assign y6284 = ~n9043 ;
  assign y6285 = ~1'b0 ;
  assign y6286 = ~1'b0 ;
  assign y6287 = 1'b0 ;
  assign y6288 = ~n14381 ;
  assign y6289 = n14383 ;
  assign y6290 = ~n14385 ;
  assign y6291 = ~n14391 ;
  assign y6292 = ~1'b0 ;
  assign y6293 = n14393 ;
  assign y6294 = n14399 ;
  assign y6295 = ~n14405 ;
  assign y6296 = ~n14407 ;
  assign y6297 = ~n14409 ;
  assign y6298 = ~n14411 ;
  assign y6299 = n14413 ;
  assign y6300 = 1'b0 ;
  assign y6301 = n14415 ;
  assign y6302 = ~1'b0 ;
  assign y6303 = ~n14421 ;
  assign y6304 = ~1'b0 ;
  assign y6305 = ~n14422 ;
  assign y6306 = ~1'b0 ;
  assign y6307 = n14427 ;
  assign y6308 = ~1'b0 ;
  assign y6309 = ~n14428 ;
  assign y6310 = n14433 ;
  assign y6311 = ~n4160 ;
  assign y6312 = n9879 ;
  assign y6313 = n14434 ;
  assign y6314 = ~n14439 ;
  assign y6315 = ~1'b0 ;
  assign y6316 = n14440 ;
  assign y6317 = ~1'b0 ;
  assign y6318 = n1746 ;
  assign y6319 = ~1'b0 ;
  assign y6320 = n14441 ;
  assign y6321 = ~1'b0 ;
  assign y6322 = n14442 ;
  assign y6323 = ~n14447 ;
  assign y6324 = ~n14449 ;
  assign y6325 = ~1'b0 ;
  assign y6326 = ~n14454 ;
  assign y6327 = ~n14458 ;
  assign y6328 = ~1'b0 ;
  assign y6329 = n14459 ;
  assign y6330 = ~n14462 ;
  assign y6331 = ~n14464 ;
  assign y6332 = ~1'b0 ;
  assign y6333 = ~1'b0 ;
  assign y6334 = n14465 ;
  assign y6335 = ~n14473 ;
  assign y6336 = ~1'b0 ;
  assign y6337 = n14477 ;
  assign y6338 = n14478 ;
  assign y6339 = ~1'b0 ;
  assign y6340 = n14480 ;
  assign y6341 = n14482 ;
  assign y6342 = ~n14483 ;
  assign y6343 = n14485 ;
  assign y6344 = ~n14488 ;
  assign y6345 = n14492 ;
  assign y6346 = n14498 ;
  assign y6347 = n14499 ;
  assign y6348 = n14503 ;
  assign y6349 = 1'b0 ;
  assign y6350 = n14504 ;
  assign y6351 = ~n14506 ;
  assign y6352 = n14512 ;
  assign y6353 = ~n14517 ;
  assign y6354 = ~1'b0 ;
  assign y6355 = ~1'b0 ;
  assign y6356 = ~n14518 ;
  assign y6357 = 1'b0 ;
  assign y6358 = ~1'b0 ;
  assign y6359 = ~n14522 ;
  assign y6360 = ~1'b0 ;
  assign y6361 = ~1'b0 ;
  assign y6362 = ~1'b0 ;
  assign y6363 = ~n14527 ;
  assign y6364 = n14529 ;
  assign y6365 = ~1'b0 ;
  assign y6366 = ~1'b0 ;
  assign y6367 = n14531 ;
  assign y6368 = n14533 ;
  assign y6369 = ~n14539 ;
  assign y6370 = n14542 ;
  assign y6371 = ~n14543 ;
  assign y6372 = ~1'b0 ;
  assign y6373 = ~1'b0 ;
  assign y6374 = n14544 ;
  assign y6375 = ~n14545 ;
  assign y6376 = ~n14550 ;
  assign y6377 = ~1'b0 ;
  assign y6378 = ~1'b0 ;
  assign y6379 = n14554 ;
  assign y6380 = ~1'b0 ;
  assign y6381 = n14560 ;
  assign y6382 = ~n14565 ;
  assign y6383 = ~1'b0 ;
  assign y6384 = n14566 ;
  assign y6385 = ~n14567 ;
  assign y6386 = ~n14575 ;
  assign y6387 = n14583 ;
  assign y6388 = ~n14584 ;
  assign y6389 = ~1'b0 ;
  assign y6390 = ~1'b0 ;
  assign y6391 = n14585 ;
  assign y6392 = n14589 ;
  assign y6393 = n14590 ;
  assign y6394 = n14592 ;
  assign y6395 = ~1'b0 ;
  assign y6396 = n14605 ;
  assign y6397 = n14619 ;
  assign y6398 = ~1'b0 ;
  assign y6399 = ~n416 ;
  assign y6400 = ~n14620 ;
  assign y6401 = ~1'b0 ;
  assign y6402 = ~n14634 ;
  assign y6403 = ~n14635 ;
  assign y6404 = n14636 ;
  assign y6405 = ~n14640 ;
  assign y6406 = n10001 ;
  assign y6407 = ~n14642 ;
  assign y6408 = n9773 ;
  assign y6409 = ~n14645 ;
  assign y6410 = n14650 ;
  assign y6411 = n14653 ;
  assign y6412 = n14656 ;
  assign y6413 = n14657 ;
  assign y6414 = ~n14658 ;
  assign y6415 = ~1'b0 ;
  assign y6416 = ~n14662 ;
  assign y6417 = ~n14663 ;
  assign y6418 = ~n14664 ;
  assign y6419 = ~n14670 ;
  assign y6420 = n14671 ;
  assign y6421 = n14684 ;
  assign y6422 = n14686 ;
  assign y6423 = ~1'b0 ;
  assign y6424 = ~n14687 ;
  assign y6425 = n14688 ;
  assign y6426 = n14694 ;
  assign y6427 = ~n14695 ;
  assign y6428 = n14696 ;
  assign y6429 = ~n14698 ;
  assign y6430 = ~n14701 ;
  assign y6431 = n14703 ;
  assign y6432 = ~1'b0 ;
  assign y6433 = n14710 ;
  assign y6434 = ~1'b0 ;
  assign y6435 = ~n14711 ;
  assign y6436 = ~n14714 ;
  assign y6437 = n14718 ;
  assign y6438 = n14723 ;
  assign y6439 = ~n14725 ;
  assign y6440 = ~1'b0 ;
  assign y6441 = n14729 ;
  assign y6442 = ~n4913 ;
  assign y6443 = ~n14734 ;
  assign y6444 = n14741 ;
  assign y6445 = n14743 ;
  assign y6446 = ~n14749 ;
  assign y6447 = ~n14750 ;
  assign y6448 = n14753 ;
  assign y6449 = ~1'b0 ;
  assign y6450 = n14758 ;
  assign y6451 = ~n14764 ;
  assign y6452 = ~n14765 ;
  assign y6453 = ~n14768 ;
  assign y6454 = n14771 ;
  assign y6455 = n8030 ;
  assign y6456 = ~n14772 ;
  assign y6457 = ~1'b0 ;
  assign y6458 = ~1'b0 ;
  assign y6459 = n14774 ;
  assign y6460 = ~n14777 ;
  assign y6461 = n12622 ;
  assign y6462 = ~n14779 ;
  assign y6463 = ~1'b0 ;
  assign y6464 = n14786 ;
  assign y6465 = ~1'b0 ;
  assign y6466 = n14788 ;
  assign y6467 = n14790 ;
  assign y6468 = n2047 ;
  assign y6469 = ~n14794 ;
  assign y6470 = ~1'b0 ;
  assign y6471 = n14797 ;
  assign y6472 = ~1'b0 ;
  assign y6473 = n14798 ;
  assign y6474 = ~n14799 ;
  assign y6475 = ~1'b0 ;
  assign y6476 = n14801 ;
  assign y6477 = n14803 ;
  assign y6478 = ~n14812 ;
  assign y6479 = n14817 ;
  assign y6480 = ~1'b0 ;
  assign y6481 = ~n14818 ;
  assign y6482 = ~n14840 ;
  assign y6483 = n14841 ;
  assign y6484 = n14842 ;
  assign y6485 = ~1'b0 ;
  assign y6486 = ~1'b0 ;
  assign y6487 = n14843 ;
  assign y6488 = n14846 ;
  assign y6489 = ~1'b0 ;
  assign y6490 = ~n14847 ;
  assign y6491 = ~n14849 ;
  assign y6492 = ~n1910 ;
  assign y6493 = ~n14851 ;
  assign y6494 = n14855 ;
  assign y6495 = ~n14856 ;
  assign y6496 = ~n14862 ;
  assign y6497 = ~n14867 ;
  assign y6498 = ~n14870 ;
  assign y6499 = ~1'b0 ;
  assign y6500 = n14871 ;
  assign y6501 = n14879 ;
  assign y6502 = n14883 ;
  assign y6503 = n14887 ;
  assign y6504 = ~1'b0 ;
  assign y6505 = n14892 ;
  assign y6506 = ~1'b0 ;
  assign y6507 = n1311 ;
  assign y6508 = ~1'b0 ;
  assign y6509 = n14895 ;
  assign y6510 = n1251 ;
  assign y6511 = ~n14897 ;
  assign y6512 = ~1'b0 ;
  assign y6513 = n14902 ;
  assign y6514 = ~n14905 ;
  assign y6515 = n14906 ;
  assign y6516 = ~1'b0 ;
  assign y6517 = n14909 ;
  assign y6518 = n14913 ;
  assign y6519 = ~n14922 ;
  assign y6520 = ~n1139 ;
  assign y6521 = n14925 ;
  assign y6522 = 1'b0 ;
  assign y6523 = ~1'b0 ;
  assign y6524 = ~n14929 ;
  assign y6525 = ~n14930 ;
  assign y6526 = ~n14931 ;
  assign y6527 = ~n14932 ;
  assign y6528 = n14934 ;
  assign y6529 = n14938 ;
  assign y6530 = ~n14939 ;
  assign y6531 = ~n14941 ;
  assign y6532 = ~n14943 ;
  assign y6533 = n14950 ;
  assign y6534 = 1'b0 ;
  assign y6535 = ~1'b0 ;
  assign y6536 = ~n14951 ;
  assign y6537 = ~n14954 ;
  assign y6538 = ~1'b0 ;
  assign y6539 = ~1'b0 ;
  assign y6540 = ~n14956 ;
  assign y6541 = n14958 ;
  assign y6542 = ~n14960 ;
  assign y6543 = n14969 ;
  assign y6544 = ~1'b0 ;
  assign y6545 = ~n14970 ;
  assign y6546 = ~n14974 ;
  assign y6547 = ~n14987 ;
  assign y6548 = ~n14990 ;
  assign y6549 = n11662 ;
  assign y6550 = n14991 ;
  assign y6551 = n12465 ;
  assign y6552 = ~1'b0 ;
  assign y6553 = n14996 ;
  assign y6554 = ~n12111 ;
  assign y6555 = n15020 ;
  assign y6556 = n15021 ;
  assign y6557 = ~n15022 ;
  assign y6558 = ~1'b0 ;
  assign y6559 = n15025 ;
  assign y6560 = n15027 ;
  assign y6561 = n15028 ;
  assign y6562 = n15030 ;
  assign y6563 = n15031 ;
  assign y6564 = n15032 ;
  assign y6565 = ~n15034 ;
  assign y6566 = n15036 ;
  assign y6567 = ~1'b0 ;
  assign y6568 = ~n15044 ;
  assign y6569 = ~n15046 ;
  assign y6570 = n15048 ;
  assign y6571 = n6188 ;
  assign y6572 = 1'b0 ;
  assign y6573 = ~n15049 ;
  assign y6574 = n15050 ;
  assign y6575 = ~n15055 ;
  assign y6576 = ~n15060 ;
  assign y6577 = ~1'b0 ;
  assign y6578 = ~n15063 ;
  assign y6579 = ~n15064 ;
  assign y6580 = ~n15068 ;
  assign y6581 = ~n15071 ;
  assign y6582 = ~n15075 ;
  assign y6583 = n15079 ;
  assign y6584 = ~n15085 ;
  assign y6585 = ~n15096 ;
  assign y6586 = ~1'b0 ;
  assign y6587 = n15100 ;
  assign y6588 = ~n15101 ;
  assign y6589 = ~n15102 ;
  assign y6590 = n15106 ;
  assign y6591 = n15107 ;
  assign y6592 = n6965 ;
  assign y6593 = ~n4180 ;
  assign y6594 = n15111 ;
  assign y6595 = ~n15115 ;
  assign y6596 = n15118 ;
  assign y6597 = ~1'b0 ;
  assign y6598 = ~1'b0 ;
  assign y6599 = n15124 ;
  assign y6600 = n15129 ;
  assign y6601 = ~n15133 ;
  assign y6602 = n15140 ;
  assign y6603 = n15142 ;
  assign y6604 = ~n15145 ;
  assign y6605 = n15146 ;
  assign y6606 = ~n15153 ;
  assign y6607 = ~n10752 ;
  assign y6608 = ~1'b0 ;
  assign y6609 = n15157 ;
  assign y6610 = ~n15160 ;
  assign y6611 = ~n15165 ;
  assign y6612 = ~1'b0 ;
  assign y6613 = ~1'b0 ;
  assign y6614 = ~1'b0 ;
  assign y6615 = n15166 ;
  assign y6616 = ~n10703 ;
  assign y6617 = n15170 ;
  assign y6618 = ~1'b0 ;
  assign y6619 = ~n15175 ;
  assign y6620 = ~n14775 ;
  assign y6621 = ~1'b0 ;
  assign y6622 = ~1'b0 ;
  assign y6623 = ~n15176 ;
  assign y6624 = ~1'b0 ;
  assign y6625 = n15177 ;
  assign y6626 = ~n15180 ;
  assign y6627 = n15181 ;
  assign y6628 = ~1'b0 ;
  assign y6629 = n15183 ;
  assign y6630 = n15187 ;
  assign y6631 = n15193 ;
  assign y6632 = n15194 ;
  assign y6633 = n15195 ;
  assign y6634 = ~n15197 ;
  assign y6635 = n15200 ;
  assign y6636 = ~n15201 ;
  assign y6637 = ~n15205 ;
  assign y6638 = n2667 ;
  assign y6639 = ~1'b0 ;
  assign y6640 = ~1'b0 ;
  assign y6641 = ~1'b0 ;
  assign y6642 = n15206 ;
  assign y6643 = ~n15208 ;
  assign y6644 = ~n15209 ;
  assign y6645 = ~n15210 ;
  assign y6646 = ~n15224 ;
  assign y6647 = ~1'b0 ;
  assign y6648 = ~1'b0 ;
  assign y6649 = ~n5101 ;
  assign y6650 = ~n4536 ;
  assign y6651 = ~n15225 ;
  assign y6652 = n15227 ;
  assign y6653 = n11134 ;
  assign y6654 = ~1'b0 ;
  assign y6655 = n15228 ;
  assign y6656 = ~1'b0 ;
  assign y6657 = n15229 ;
  assign y6658 = ~n15230 ;
  assign y6659 = ~1'b0 ;
  assign y6660 = ~n15232 ;
  assign y6661 = ~n15233 ;
  assign y6662 = ~n15237 ;
  assign y6663 = ~n15240 ;
  assign y6664 = ~1'b0 ;
  assign y6665 = n15241 ;
  assign y6666 = n15243 ;
  assign y6667 = ~1'b0 ;
  assign y6668 = ~1'b0 ;
  assign y6669 = ~1'b0 ;
  assign y6670 = ~n15251 ;
  assign y6671 = ~n15252 ;
  assign y6672 = n15257 ;
  assign y6673 = n15258 ;
  assign y6674 = n15262 ;
  assign y6675 = ~n15264 ;
  assign y6676 = ~1'b0 ;
  assign y6677 = n15269 ;
  assign y6678 = n15274 ;
  assign y6679 = ~n15280 ;
  assign y6680 = ~1'b0 ;
  assign y6681 = ~1'b0 ;
  assign y6682 = ~n15282 ;
  assign y6683 = n928 ;
  assign y6684 = ~n15287 ;
  assign y6685 = ~n15290 ;
  assign y6686 = ~n15291 ;
  assign y6687 = ~1'b0 ;
  assign y6688 = ~1'b0 ;
  assign y6689 = ~n15292 ;
  assign y6690 = n15296 ;
  assign y6691 = ~1'b0 ;
  assign y6692 = ~n5273 ;
  assign y6693 = ~n15299 ;
  assign y6694 = ~n15304 ;
  assign y6695 = ~1'b0 ;
  assign y6696 = ~1'b0 ;
  assign y6697 = ~n15309 ;
  assign y6698 = ~n12040 ;
  assign y6699 = ~n15311 ;
  assign y6700 = ~1'b0 ;
  assign y6701 = ~n15313 ;
  assign y6702 = ~1'b0 ;
  assign y6703 = ~n15314 ;
  assign y6704 = ~1'b0 ;
  assign y6705 = n15319 ;
  assign y6706 = ~n15323 ;
  assign y6707 = ~n15326 ;
  assign y6708 = n15327 ;
  assign y6709 = ~1'b0 ;
  assign y6710 = ~n15328 ;
  assign y6711 = n8325 ;
  assign y6712 = n572 ;
  assign y6713 = n15331 ;
  assign y6714 = ~1'b0 ;
  assign y6715 = n15333 ;
  assign y6716 = n15335 ;
  assign y6717 = ~n15337 ;
  assign y6718 = ~n15343 ;
  assign y6719 = n15353 ;
  assign y6720 = ~1'b0 ;
  assign y6721 = ~n15355 ;
  assign y6722 = n15360 ;
  assign y6723 = n15364 ;
  assign y6724 = 1'b0 ;
  assign y6725 = ~n15366 ;
  assign y6726 = ~n15375 ;
  assign y6727 = n15379 ;
  assign y6728 = n15381 ;
  assign y6729 = ~1'b0 ;
  assign y6730 = n15383 ;
  assign y6731 = ~n15394 ;
  assign y6732 = ~1'b0 ;
  assign y6733 = ~n15399 ;
  assign y6734 = ~n15401 ;
  assign y6735 = ~1'b0 ;
  assign y6736 = n15404 ;
  assign y6737 = n15405 ;
  assign y6738 = ~n15406 ;
  assign y6739 = ~1'b0 ;
  assign y6740 = ~1'b0 ;
  assign y6741 = n14674 ;
  assign y6742 = n15407 ;
  assign y6743 = n6050 ;
  assign y6744 = ~n15410 ;
  assign y6745 = ~n15416 ;
  assign y6746 = ~n3449 ;
  assign y6747 = ~n15418 ;
  assign y6748 = n15420 ;
  assign y6749 = ~1'b0 ;
  assign y6750 = ~1'b0 ;
  assign y6751 = n15423 ;
  assign y6752 = ~n15428 ;
  assign y6753 = n15431 ;
  assign y6754 = ~n15436 ;
  assign y6755 = ~n15441 ;
  assign y6756 = ~1'b0 ;
  assign y6757 = n15446 ;
  assign y6758 = ~n15450 ;
  assign y6759 = ~1'b0 ;
  assign y6760 = ~n15455 ;
  assign y6761 = ~n15456 ;
  assign y6762 = n15457 ;
  assign y6763 = ~1'b0 ;
  assign y6764 = n15462 ;
  assign y6765 = n15464 ;
  assign y6766 = ~1'b0 ;
  assign y6767 = n15466 ;
  assign y6768 = n9360 ;
  assign y6769 = n15468 ;
  assign y6770 = ~n15473 ;
  assign y6771 = ~1'b0 ;
  assign y6772 = ~n15475 ;
  assign y6773 = ~1'b0 ;
  assign y6774 = ~n15477 ;
  assign y6775 = ~n15478 ;
  assign y6776 = ~n15479 ;
  assign y6777 = ~n15481 ;
  assign y6778 = ~n15487 ;
  assign y6779 = ~n15489 ;
  assign y6780 = n10129 ;
  assign y6781 = ~n15492 ;
  assign y6782 = ~1'b0 ;
  assign y6783 = ~n15495 ;
  assign y6784 = ~n12018 ;
  assign y6785 = n9621 ;
  assign y6786 = ~n15497 ;
  assign y6787 = ~n15498 ;
  assign y6788 = ~n15501 ;
  assign y6789 = ~n15503 ;
  assign y6790 = n15505 ;
  assign y6791 = ~1'b0 ;
  assign y6792 = ~n15507 ;
  assign y6793 = ~n15513 ;
  assign y6794 = ~1'b0 ;
  assign y6795 = n15518 ;
  assign y6796 = ~n15520 ;
  assign y6797 = ~n15522 ;
  assign y6798 = ~1'b0 ;
  assign y6799 = ~1'b0 ;
  assign y6800 = ~1'b0 ;
  assign y6801 = n15523 ;
  assign y6802 = ~n15525 ;
  assign y6803 = n15527 ;
  assign y6804 = ~1'b0 ;
  assign y6805 = ~n15528 ;
  assign y6806 = ~1'b0 ;
  assign y6807 = ~n4675 ;
  assign y6808 = ~1'b0 ;
  assign y6809 = ~n15529 ;
  assign y6810 = n15533 ;
  assign y6811 = 1'b0 ;
  assign y6812 = ~n15534 ;
  assign y6813 = n15537 ;
  assign y6814 = n15546 ;
  assign y6815 = ~n15550 ;
  assign y6816 = n15554 ;
  assign y6817 = ~n15557 ;
  assign y6818 = n15558 ;
  assign y6819 = ~1'b0 ;
  assign y6820 = ~1'b0 ;
  assign y6821 = n15560 ;
  assign y6822 = ~n15565 ;
  assign y6823 = ~n15566 ;
  assign y6824 = ~1'b0 ;
  assign y6825 = ~n15571 ;
  assign y6826 = ~n15573 ;
  assign y6827 = n15574 ;
  assign y6828 = n15579 ;
  assign y6829 = n15581 ;
  assign y6830 = n15582 ;
  assign y6831 = n15585 ;
  assign y6832 = n15589 ;
  assign y6833 = n15590 ;
  assign y6834 = ~1'b0 ;
  assign y6835 = ~n15592 ;
  assign y6836 = ~1'b0 ;
  assign y6837 = ~n15604 ;
  assign y6838 = ~n15608 ;
  assign y6839 = ~1'b0 ;
  assign y6840 = n15613 ;
  assign y6841 = n9462 ;
  assign y6842 = n15621 ;
  assign y6843 = n15624 ;
  assign y6844 = 1'b0 ;
  assign y6845 = ~1'b0 ;
  assign y6846 = ~n15628 ;
  assign y6847 = ~n15637 ;
  assign y6848 = n15640 ;
  assign y6849 = ~1'b0 ;
  assign y6850 = ~n15647 ;
  assign y6851 = n15650 ;
  assign y6852 = ~1'b0 ;
  assign y6853 = ~n15651 ;
  assign y6854 = ~1'b0 ;
  assign y6855 = ~1'b0 ;
  assign y6856 = n15652 ;
  assign y6857 = n15653 ;
  assign y6858 = n15660 ;
  assign y6859 = n15663 ;
  assign y6860 = n15666 ;
  assign y6861 = ~1'b0 ;
  assign y6862 = n15669 ;
  assign y6863 = ~1'b0 ;
  assign y6864 = ~n5458 ;
  assign y6865 = ~1'b0 ;
  assign y6866 = ~n15671 ;
  assign y6867 = ~n15672 ;
  assign y6868 = ~n15678 ;
  assign y6869 = ~1'b0 ;
  assign y6870 = ~1'b0 ;
  assign y6871 = ~1'b0 ;
  assign y6872 = ~1'b0 ;
  assign y6873 = ~1'b0 ;
  assign y6874 = n15679 ;
  assign y6875 = ~n15680 ;
  assign y6876 = ~n15683 ;
  assign y6877 = ~n15684 ;
  assign y6878 = n15685 ;
  assign y6879 = n15692 ;
  assign y6880 = n15695 ;
  assign y6881 = n8656 ;
  assign y6882 = n15696 ;
  assign y6883 = ~1'b0 ;
  assign y6884 = ~n15704 ;
  assign y6885 = ~n14719 ;
  assign y6886 = ~n15716 ;
  assign y6887 = ~1'b0 ;
  assign y6888 = ~1'b0 ;
  assign y6889 = ~1'b0 ;
  assign y6890 = n15724 ;
  assign y6891 = ~n6123 ;
  assign y6892 = n15728 ;
  assign y6893 = ~n15730 ;
  assign y6894 = n15733 ;
  assign y6895 = 1'b0 ;
  assign y6896 = ~n15739 ;
  assign y6897 = ~1'b0 ;
  assign y6898 = n15741 ;
  assign y6899 = ~1'b0 ;
  assign y6900 = ~n15742 ;
  assign y6901 = ~n15748 ;
  assign y6902 = ~n15749 ;
  assign y6903 = n15752 ;
  assign y6904 = n15754 ;
  assign y6905 = n15759 ;
  assign y6906 = ~1'b0 ;
  assign y6907 = n3252 ;
  assign y6908 = n15765 ;
  assign y6909 = ~n15770 ;
  assign y6910 = ~n15775 ;
  assign y6911 = n15777 ;
  assign y6912 = n15784 ;
  assign y6913 = ~n15785 ;
  assign y6914 = n15789 ;
  assign y6915 = n15792 ;
  assign y6916 = ~n15796 ;
  assign y6917 = ~n15797 ;
  assign y6918 = ~n15803 ;
  assign y6919 = n15807 ;
  assign y6920 = ~n9043 ;
  assign y6921 = ~n15809 ;
  assign y6922 = ~1'b0 ;
  assign y6923 = ~1'b0 ;
  assign y6924 = ~n15813 ;
  assign y6925 = n15815 ;
  assign y6926 = n15816 ;
  assign y6927 = ~1'b0 ;
  assign y6928 = ~1'b0 ;
  assign y6929 = ~1'b0 ;
  assign y6930 = n15817 ;
  assign y6931 = ~1'b0 ;
  assign y6932 = n15820 ;
  assign y6933 = ~n15833 ;
  assign y6934 = ~n15835 ;
  assign y6935 = n15836 ;
  assign y6936 = n15839 ;
  assign y6937 = n15843 ;
  assign y6938 = n15845 ;
  assign y6939 = n15846 ;
  assign y6940 = n9879 ;
  assign y6941 = ~n15852 ;
  assign y6942 = n15857 ;
  assign y6943 = n15861 ;
  assign y6944 = ~1'b0 ;
  assign y6945 = ~n15863 ;
  assign y6946 = ~n15864 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = n3098 ;
  assign y6949 = ~n15871 ;
  assign y6950 = ~n15876 ;
  assign y6951 = ~n15879 ;
  assign y6952 = ~n15880 ;
  assign y6953 = ~n15882 ;
  assign y6954 = ~n15884 ;
  assign y6955 = ~1'b0 ;
  assign y6956 = ~n15886 ;
  assign y6957 = ~n15890 ;
  assign y6958 = ~1'b0 ;
  assign y6959 = n15895 ;
  assign y6960 = ~n15897 ;
  assign y6961 = ~n15910 ;
  assign y6962 = ~n15911 ;
  assign y6963 = n15912 ;
  assign y6964 = ~n15916 ;
  assign y6965 = n15918 ;
  assign y6966 = ~n15919 ;
  assign y6967 = ~1'b0 ;
  assign y6968 = ~n15921 ;
  assign y6969 = ~1'b0 ;
  assign y6970 = ~1'b0 ;
  assign y6971 = ~n15925 ;
  assign y6972 = ~n15926 ;
  assign y6973 = n15930 ;
  assign y6974 = ~n15931 ;
  assign y6975 = ~n15936 ;
  assign y6976 = ~n15937 ;
  assign y6977 = n15943 ;
  assign y6978 = n15949 ;
  assign y6979 = n15952 ;
  assign y6980 = n15955 ;
  assign y6981 = ~1'b0 ;
  assign y6982 = ~1'b0 ;
  assign y6983 = ~n15959 ;
  assign y6984 = ~n15960 ;
  assign y6985 = ~1'b0 ;
  assign y6986 = n15962 ;
  assign y6987 = ~1'b0 ;
  assign y6988 = n15966 ;
  assign y6989 = n15967 ;
  assign y6990 = ~n1761 ;
  assign y6991 = ~n15971 ;
  assign y6992 = ~1'b0 ;
  assign y6993 = n15972 ;
  assign y6994 = ~n15973 ;
  assign y6995 = ~n15976 ;
  assign y6996 = n6245 ;
  assign y6997 = ~1'b0 ;
  assign y6998 = ~n9081 ;
  assign y6999 = n15977 ;
  assign y7000 = n15981 ;
  assign y7001 = ~n15984 ;
  assign y7002 = n15988 ;
  assign y7003 = n15989 ;
  assign y7004 = n15990 ;
  assign y7005 = n3455 ;
  assign y7006 = ~n15991 ;
  assign y7007 = ~1'b0 ;
  assign y7008 = n7505 ;
  assign y7009 = ~1'b0 ;
  assign y7010 = ~n15994 ;
  assign y7011 = n15995 ;
  assign y7012 = ~1'b0 ;
  assign y7013 = ~1'b0 ;
  assign y7014 = ~1'b0 ;
  assign y7015 = ~1'b0 ;
  assign y7016 = ~n15996 ;
  assign y7017 = ~n15997 ;
  assign y7018 = n16000 ;
  assign y7019 = n16004 ;
  assign y7020 = ~n16005 ;
  assign y7021 = ~n16006 ;
  assign y7022 = ~n16008 ;
  assign y7023 = n16011 ;
  assign y7024 = n16014 ;
  assign y7025 = ~n16019 ;
  assign y7026 = ~1'b0 ;
  assign y7027 = n16023 ;
  assign y7028 = ~n15876 ;
  assign y7029 = n16024 ;
  assign y7030 = ~1'b0 ;
  assign y7031 = ~1'b0 ;
  assign y7032 = n16027 ;
  assign y7033 = ~n16030 ;
  assign y7034 = 1'b0 ;
  assign y7035 = n16032 ;
  assign y7036 = ~n16033 ;
  assign y7037 = n16035 ;
  assign y7038 = ~n16036 ;
  assign y7039 = ~n16041 ;
  assign y7040 = ~1'b0 ;
  assign y7041 = n16046 ;
  assign y7042 = ~n16050 ;
  assign y7043 = ~1'b0 ;
  assign y7044 = n3906 ;
  assign y7045 = n16053 ;
  assign y7046 = n16058 ;
  assign y7047 = ~n16059 ;
  assign y7048 = n16060 ;
  assign y7049 = ~n16063 ;
  assign y7050 = ~1'b0 ;
  assign y7051 = n16065 ;
  assign y7052 = n13011 ;
  assign y7053 = ~n11852 ;
  assign y7054 = ~1'b0 ;
  assign y7055 = n16066 ;
  assign y7056 = ~1'b0 ;
  assign y7057 = ~1'b0 ;
  assign y7058 = n16067 ;
  assign y7059 = n9715 ;
  assign y7060 = n16071 ;
  assign y7061 = n16075 ;
  assign y7062 = n16077 ;
  assign y7063 = ~n16081 ;
  assign y7064 = n16087 ;
  assign y7065 = ~1'b0 ;
  assign y7066 = n16091 ;
  assign y7067 = n16093 ;
  assign y7068 = ~n16096 ;
  assign y7069 = n16097 ;
  assign y7070 = ~n16098 ;
  assign y7071 = n16102 ;
  assign y7072 = ~n16104 ;
  assign y7073 = ~n16106 ;
  assign y7074 = ~n16117 ;
  assign y7075 = ~n16122 ;
  assign y7076 = n10138 ;
  assign y7077 = ~n16123 ;
  assign y7078 = ~n16126 ;
  assign y7079 = n16127 ;
  assign y7080 = n16130 ;
  assign y7081 = ~1'b0 ;
  assign y7082 = n16133 ;
  assign y7083 = n16140 ;
  assign y7084 = n16146 ;
  assign y7085 = ~1'b0 ;
  assign y7086 = ~n11260 ;
  assign y7087 = ~1'b0 ;
  assign y7088 = n16154 ;
  assign y7089 = ~n16157 ;
  assign y7090 = n16166 ;
  assign y7091 = ~n16170 ;
  assign y7092 = ~1'b0 ;
  assign y7093 = ~n8480 ;
  assign y7094 = ~1'b0 ;
  assign y7095 = n16171 ;
  assign y7096 = 1'b0 ;
  assign y7097 = n16181 ;
  assign y7098 = n16182 ;
  assign y7099 = ~n16186 ;
  assign y7100 = ~1'b0 ;
  assign y7101 = ~n16194 ;
  assign y7102 = n16195 ;
  assign y7103 = n16196 ;
  assign y7104 = ~1'b0 ;
  assign y7105 = 1'b0 ;
  assign y7106 = n16198 ;
  assign y7107 = ~1'b0 ;
  assign y7108 = n16199 ;
  assign y7109 = ~n16201 ;
  assign y7110 = ~n16203 ;
  assign y7111 = ~1'b0 ;
  assign y7112 = n16205 ;
  assign y7113 = ~n16208 ;
  assign y7114 = ~n16210 ;
  assign y7115 = ~1'b0 ;
  assign y7116 = n16218 ;
  assign y7117 = n16219 ;
  assign y7118 = ~n16225 ;
  assign y7119 = n16226 ;
  assign y7120 = ~n16230 ;
  assign y7121 = n11832 ;
  assign y7122 = ~1'b0 ;
  assign y7123 = n16231 ;
  assign y7124 = ~n16232 ;
  assign y7125 = 1'b0 ;
  assign y7126 = n16235 ;
  assign y7127 = ~n16238 ;
  assign y7128 = n16240 ;
  assign y7129 = ~n16244 ;
  assign y7130 = ~n16250 ;
  assign y7131 = 1'b0 ;
  assign y7132 = ~1'b0 ;
  assign y7133 = n16255 ;
  assign y7134 = n16256 ;
  assign y7135 = n16259 ;
  assign y7136 = ~1'b0 ;
  assign y7137 = ~1'b0 ;
  assign y7138 = n16260 ;
  assign y7139 = ~1'b0 ;
  assign y7140 = n16262 ;
  assign y7141 = ~n16264 ;
  assign y7142 = ~n16273 ;
  assign y7143 = n16274 ;
  assign y7144 = ~n16277 ;
  assign y7145 = n16278 ;
  assign y7146 = ~n16279 ;
  assign y7147 = ~n16280 ;
  assign y7148 = n16286 ;
  assign y7149 = ~n16290 ;
  assign y7150 = ~1'b0 ;
  assign y7151 = n16291 ;
  assign y7152 = ~n16293 ;
  assign y7153 = ~1'b0 ;
  assign y7154 = ~n16296 ;
  assign y7155 = n16299 ;
  assign y7156 = ~1'b0 ;
  assign y7157 = ~1'b0 ;
  assign y7158 = ~1'b0 ;
  assign y7159 = ~n14194 ;
  assign y7160 = ~1'b0 ;
  assign y7161 = ~1'b0 ;
  assign y7162 = n16302 ;
  assign y7163 = n16304 ;
  assign y7164 = n16311 ;
  assign y7165 = n16314 ;
  assign y7166 = ~1'b0 ;
  assign y7167 = n16317 ;
  assign y7168 = ~n16318 ;
  assign y7169 = ~n16327 ;
  assign y7170 = ~1'b0 ;
  assign y7171 = ~n16328 ;
  assign y7172 = n16330 ;
  assign y7173 = n16332 ;
  assign y7174 = n16336 ;
  assign y7175 = ~n16341 ;
  assign y7176 = n16342 ;
  assign y7177 = ~n11656 ;
  assign y7178 = ~1'b0 ;
  assign y7179 = ~n16343 ;
  assign y7180 = n16350 ;
  assign y7181 = ~n12421 ;
  assign y7182 = ~n16353 ;
  assign y7183 = ~1'b0 ;
  assign y7184 = ~1'b0 ;
  assign y7185 = ~1'b0 ;
  assign y7186 = ~1'b0 ;
  assign y7187 = ~n16357 ;
  assign y7188 = n16360 ;
  assign y7189 = 1'b0 ;
  assign y7190 = ~n16362 ;
  assign y7191 = ~n16365 ;
  assign y7192 = ~n5872 ;
  assign y7193 = ~1'b0 ;
  assign y7194 = ~n16366 ;
  assign y7195 = ~1'b0 ;
  assign y7196 = ~1'b0 ;
  assign y7197 = ~1'b0 ;
  assign y7198 = ~n11998 ;
  assign y7199 = n16367 ;
  assign y7200 = ~1'b0 ;
  assign y7201 = ~n16373 ;
  assign y7202 = ~n16374 ;
  assign y7203 = ~n16376 ;
  assign y7204 = ~n16381 ;
  assign y7205 = n16383 ;
  assign y7206 = ~1'b0 ;
  assign y7207 = n9075 ;
  assign y7208 = n16385 ;
  assign y7209 = ~n16391 ;
  assign y7210 = n16393 ;
  assign y7211 = n16394 ;
  assign y7212 = n16396 ;
  assign y7213 = ~1'b0 ;
  assign y7214 = n16398 ;
  assign y7215 = ~1'b0 ;
  assign y7216 = n16399 ;
  assign y7217 = ~n16400 ;
  assign y7218 = ~1'b0 ;
  assign y7219 = n16404 ;
  assign y7220 = ~1'b0 ;
  assign y7221 = ~1'b0 ;
  assign y7222 = ~n16406 ;
  assign y7223 = ~n16413 ;
  assign y7224 = ~1'b0 ;
  assign y7225 = ~1'b0 ;
  assign y7226 = ~n16417 ;
  assign y7227 = n16420 ;
  assign y7228 = n16421 ;
  assign y7229 = n16425 ;
  assign y7230 = ~n16428 ;
  assign y7231 = ~1'b0 ;
  assign y7232 = n16430 ;
  assign y7233 = n16439 ;
  assign y7234 = ~1'b0 ;
  assign y7235 = ~n16444 ;
  assign y7236 = n16447 ;
  assign y7237 = ~n2689 ;
  assign y7238 = ~n16451 ;
  assign y7239 = n16452 ;
  assign y7240 = ~n16457 ;
  assign y7241 = n16459 ;
  assign y7242 = ~1'b0 ;
  assign y7243 = ~n16461 ;
  assign y7244 = n16465 ;
  assign y7245 = ~1'b0 ;
  assign y7246 = n16468 ;
  assign y7247 = n16470 ;
  assign y7248 = ~n16477 ;
  assign y7249 = n16483 ;
  assign y7250 = ~n16484 ;
  assign y7251 = ~1'b0 ;
  assign y7252 = ~1'b0 ;
  assign y7253 = ~n16487 ;
  assign y7254 = ~1'b0 ;
  assign y7255 = ~1'b0 ;
  assign y7256 = ~1'b0 ;
  assign y7257 = ~n16496 ;
  assign y7258 = n16497 ;
  assign y7259 = ~n16502 ;
  assign y7260 = n16505 ;
  assign y7261 = ~1'b0 ;
  assign y7262 = ~n16510 ;
  assign y7263 = ~n16511 ;
  assign y7264 = ~n16513 ;
  assign y7265 = ~n16516 ;
  assign y7266 = n16517 ;
  assign y7267 = ~1'b0 ;
  assign y7268 = n16523 ;
  assign y7269 = n16526 ;
  assign y7270 = n16531 ;
  assign y7271 = ~n16538 ;
  assign y7272 = n16539 ;
  assign y7273 = n16542 ;
  assign y7274 = ~1'b0 ;
  assign y7275 = 1'b0 ;
  assign y7276 = ~n4004 ;
  assign y7277 = n16544 ;
  assign y7278 = ~1'b0 ;
  assign y7279 = n16548 ;
  assign y7280 = n16549 ;
  assign y7281 = n16552 ;
  assign y7282 = n16560 ;
  assign y7283 = n16563 ;
  assign y7284 = ~n16568 ;
  assign y7285 = n16571 ;
  assign y7286 = ~1'b0 ;
  assign y7287 = n16572 ;
  assign y7288 = n16573 ;
  assign y7289 = n16574 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = ~1'b0 ;
  assign y7292 = ~1'b0 ;
  assign y7293 = ~1'b0 ;
  assign y7294 = ~1'b0 ;
  assign y7295 = n16575 ;
  assign y7296 = ~1'b0 ;
  assign y7297 = ~n16578 ;
  assign y7298 = ~n16580 ;
  assign y7299 = ~1'b0 ;
  assign y7300 = n7218 ;
  assign y7301 = ~1'b0 ;
  assign y7302 = ~1'b0 ;
  assign y7303 = ~n15993 ;
  assign y7304 = ~1'b0 ;
  assign y7305 = ~n16585 ;
  assign y7306 = ~n16587 ;
  assign y7307 = n16589 ;
  assign y7308 = ~n16599 ;
  assign y7309 = ~n16603 ;
  assign y7310 = 1'b0 ;
  assign y7311 = n16610 ;
  assign y7312 = n16611 ;
  assign y7313 = ~1'b0 ;
  assign y7314 = n16612 ;
  assign y7315 = n16614 ;
  assign y7316 = ~n16618 ;
  assign y7317 = 1'b0 ;
  assign y7318 = n16623 ;
  assign y7319 = n16624 ;
  assign y7320 = ~1'b0 ;
  assign y7321 = n16625 ;
  assign y7322 = ~n16627 ;
  assign y7323 = n16629 ;
  assign y7324 = ~n16632 ;
  assign y7325 = ~1'b0 ;
  assign y7326 = ~n16635 ;
  assign y7327 = n16636 ;
  assign y7328 = ~1'b0 ;
  assign y7329 = ~n16640 ;
  assign y7330 = ~n16642 ;
  assign y7331 = ~1'b0 ;
  assign y7332 = n16651 ;
  assign y7333 = ~n16653 ;
  assign y7334 = n16658 ;
  assign y7335 = ~1'b0 ;
  assign y7336 = ~n16663 ;
  assign y7337 = n16666 ;
  assign y7338 = ~n16668 ;
  assign y7339 = ~n16669 ;
  assign y7340 = ~n16687 ;
  assign y7341 = ~n8605 ;
  assign y7342 = ~n16689 ;
  assign y7343 = ~n16704 ;
  assign y7344 = n16706 ;
  assign y7345 = ~n16707 ;
  assign y7346 = ~1'b0 ;
  assign y7347 = ~n16709 ;
  assign y7348 = ~n16711 ;
  assign y7349 = ~n16717 ;
  assign y7350 = n39 ;
  assign y7351 = n16720 ;
  assign y7352 = 1'b0 ;
  assign y7353 = n1654 ;
  assign y7354 = ~n16723 ;
  assign y7355 = ~n8950 ;
  assign y7356 = ~1'b0 ;
  assign y7357 = ~1'b0 ;
  assign y7358 = ~1'b0 ;
  assign y7359 = ~1'b0 ;
  assign y7360 = ~n16726 ;
  assign y7361 = ~1'b0 ;
  assign y7362 = ~n16730 ;
  assign y7363 = n16736 ;
  assign y7364 = ~n16748 ;
  assign y7365 = ~1'b0 ;
  assign y7366 = ~n16749 ;
  assign y7367 = ~1'b0 ;
  assign y7368 = n16751 ;
  assign y7369 = ~n16753 ;
  assign y7370 = ~n16759 ;
  assign y7371 = ~1'b0 ;
  assign y7372 = n16762 ;
  assign y7373 = ~n16763 ;
  assign y7374 = ~n5335 ;
  assign y7375 = n16768 ;
  assign y7376 = n16772 ;
  assign y7377 = ~1'b0 ;
  assign y7378 = n16774 ;
  assign y7379 = n16778 ;
  assign y7380 = ~n16780 ;
  assign y7381 = ~n16786 ;
  assign y7382 = ~1'b0 ;
  assign y7383 = ~1'b0 ;
  assign y7384 = ~n16789 ;
  assign y7385 = ~n16797 ;
  assign y7386 = ~1'b0 ;
  assign y7387 = ~1'b0 ;
  assign y7388 = ~1'b0 ;
  assign y7389 = ~1'b0 ;
  assign y7390 = n16798 ;
  assign y7391 = n16805 ;
  assign y7392 = ~1'b0 ;
  assign y7393 = ~n16810 ;
  assign y7394 = ~n16811 ;
  assign y7395 = ~n4805 ;
  assign y7396 = ~n16812 ;
  assign y7397 = ~1'b0 ;
  assign y7398 = n2879 ;
  assign y7399 = ~1'b0 ;
  assign y7400 = ~n16813 ;
  assign y7401 = ~n16814 ;
  assign y7402 = ~n16818 ;
  assign y7403 = ~1'b0 ;
  assign y7404 = ~n16819 ;
  assign y7405 = n16821 ;
  assign y7406 = n16825 ;
  assign y7407 = ~n16735 ;
  assign y7408 = n16827 ;
  assign y7409 = ~n16829 ;
  assign y7410 = ~n16835 ;
  assign y7411 = ~1'b0 ;
  assign y7412 = ~n16836 ;
  assign y7413 = n16838 ;
  assign y7414 = ~1'b0 ;
  assign y7415 = n16840 ;
  assign y7416 = ~n16846 ;
  assign y7417 = n16854 ;
  assign y7418 = n16855 ;
  assign y7419 = n16859 ;
  assign y7420 = n16863 ;
  assign y7421 = ~n14188 ;
  assign y7422 = n16864 ;
  assign y7423 = n16867 ;
  assign y7424 = ~n16868 ;
  assign y7425 = ~1'b0 ;
  assign y7426 = ~1'b0 ;
  assign y7427 = ~n16873 ;
  assign y7428 = n16877 ;
  assign y7429 = ~1'b0 ;
  assign y7430 = n16878 ;
  assign y7431 = ~n16879 ;
  assign y7432 = ~1'b0 ;
  assign y7433 = ~1'b0 ;
  assign y7434 = ~1'b0 ;
  assign y7435 = n16881 ;
  assign y7436 = ~n16882 ;
  assign y7437 = n16885 ;
  assign y7438 = ~n16888 ;
  assign y7439 = ~n16890 ;
  assign y7440 = ~1'b0 ;
  assign y7441 = n16891 ;
  assign y7442 = ~n16893 ;
  assign y7443 = n16894 ;
  assign y7444 = ~n16898 ;
  assign y7445 = ~n16903 ;
  assign y7446 = n16904 ;
  assign y7447 = n16906 ;
  assign y7448 = ~n16907 ;
  assign y7449 = ~n16911 ;
  assign y7450 = n16913 ;
  assign y7451 = ~n16918 ;
  assign y7452 = ~n16920 ;
  assign y7453 = n16927 ;
  assign y7454 = ~n16931 ;
  assign y7455 = n16936 ;
  assign y7456 = ~n16938 ;
  assign y7457 = ~n16942 ;
  assign y7458 = ~1'b0 ;
  assign y7459 = ~1'b0 ;
  assign y7460 = ~n16946 ;
  assign y7461 = n16950 ;
  assign y7462 = n16951 ;
  assign y7463 = ~1'b0 ;
  assign y7464 = n16953 ;
  assign y7465 = n16955 ;
  assign y7466 = ~1'b0 ;
  assign y7467 = ~n16959 ;
  assign y7468 = n16961 ;
  assign y7469 = ~n16963 ;
  assign y7470 = n16965 ;
  assign y7471 = ~n16967 ;
  assign y7472 = ~1'b0 ;
  assign y7473 = n16971 ;
  assign y7474 = n16976 ;
  assign y7475 = ~1'b0 ;
  assign y7476 = ~n16982 ;
  assign y7477 = ~n16983 ;
  assign y7478 = ~1'b0 ;
  assign y7479 = n16988 ;
  assign y7480 = ~1'b0 ;
  assign y7481 = ~n16993 ;
  assign y7482 = ~n16997 ;
  assign y7483 = n17000 ;
  assign y7484 = ~1'b0 ;
  assign y7485 = ~n17003 ;
  assign y7486 = ~1'b0 ;
  assign y7487 = ~n17010 ;
  assign y7488 = n17012 ;
  assign y7489 = ~n17014 ;
  assign y7490 = ~n17015 ;
  assign y7491 = n17016 ;
  assign y7492 = ~1'b0 ;
  assign y7493 = ~n17027 ;
  assign y7494 = n17029 ;
  assign y7495 = n17031 ;
  assign y7496 = ~n17041 ;
  assign y7497 = n17042 ;
  assign y7498 = ~1'b0 ;
  assign y7499 = ~n17045 ;
  assign y7500 = ~n17051 ;
  assign y7501 = ~1'b0 ;
  assign y7502 = ~1'b0 ;
  assign y7503 = n17053 ;
  assign y7504 = ~n17057 ;
  assign y7505 = n17058 ;
  assign y7506 = ~n17060 ;
  assign y7507 = ~n17065 ;
  assign y7508 = ~1'b0 ;
  assign y7509 = ~1'b0 ;
  assign y7510 = n17070 ;
  assign y7511 = n17081 ;
  assign y7512 = n17083 ;
  assign y7513 = n17085 ;
  assign y7514 = ~n17088 ;
  assign y7515 = ~n16269 ;
  assign y7516 = n17092 ;
  assign y7517 = n17094 ;
  assign y7518 = ~1'b0 ;
  assign y7519 = ~1'b0 ;
  assign y7520 = ~n17095 ;
  assign y7521 = ~1'b0 ;
  assign y7522 = ~n17097 ;
  assign y7523 = ~n17100 ;
  assign y7524 = n17102 ;
  assign y7525 = n17108 ;
  assign y7526 = ~1'b0 ;
  assign y7527 = n17109 ;
  assign y7528 = ~1'b0 ;
  assign y7529 = n4454 ;
  assign y7530 = ~n17113 ;
  assign y7531 = ~1'b0 ;
  assign y7532 = n17118 ;
  assign y7533 = ~n17121 ;
  assign y7534 = n17125 ;
  assign y7535 = ~n17133 ;
  assign y7536 = ~n17135 ;
  assign y7537 = ~n17137 ;
  assign y7538 = ~1'b0 ;
  assign y7539 = ~1'b0 ;
  assign y7540 = ~1'b0 ;
  assign y7541 = ~1'b0 ;
  assign y7542 = ~1'b0 ;
  assign y7543 = ~n17139 ;
  assign y7544 = ~1'b0 ;
  assign y7545 = n17140 ;
  assign y7546 = ~n17142 ;
  assign y7547 = ~n17143 ;
  assign y7548 = ~n17145 ;
  assign y7549 = n17150 ;
  assign y7550 = ~1'b0 ;
  assign y7551 = ~1'b0 ;
  assign y7552 = ~n17151 ;
  assign y7553 = n17158 ;
  assign y7554 = ~n17160 ;
  assign y7555 = n17165 ;
  assign y7556 = ~n17168 ;
  assign y7557 = ~n17171 ;
  assign y7558 = ~1'b0 ;
  assign y7559 = ~1'b0 ;
  assign y7560 = ~n17174 ;
  assign y7561 = n17175 ;
  assign y7562 = n17177 ;
  assign y7563 = ~n17179 ;
  assign y7564 = ~n17180 ;
  assign y7565 = ~n17181 ;
  assign y7566 = 1'b0 ;
  assign y7567 = ~1'b0 ;
  assign y7568 = ~n17182 ;
  assign y7569 = 1'b0 ;
  assign y7570 = n17187 ;
  assign y7571 = ~n17192 ;
  assign y7572 = n17196 ;
  assign y7573 = n937 ;
  assign y7574 = n17201 ;
  assign y7575 = n14779 ;
  assign y7576 = ~1'b0 ;
  assign y7577 = n17202 ;
  assign y7578 = ~n17212 ;
  assign y7579 = n6083 ;
  assign y7580 = ~n17216 ;
  assign y7581 = ~n17217 ;
  assign y7582 = ~1'b0 ;
  assign y7583 = ~1'b0 ;
  assign y7584 = n17218 ;
  assign y7585 = ~n17222 ;
  assign y7586 = ~1'b0 ;
  assign y7587 = ~1'b0 ;
  assign y7588 = 1'b0 ;
  assign y7589 = n17223 ;
  assign y7590 = ~n17228 ;
  assign y7591 = ~1'b0 ;
  assign y7592 = ~1'b0 ;
  assign y7593 = n17229 ;
  assign y7594 = ~n17233 ;
  assign y7595 = n17237 ;
  assign y7596 = ~n17239 ;
  assign y7597 = n17240 ;
  assign y7598 = ~n17226 ;
  assign y7599 = n17242 ;
  assign y7600 = n17244 ;
  assign y7601 = ~1'b0 ;
  assign y7602 = ~n17245 ;
  assign y7603 = n17250 ;
  assign y7604 = n17252 ;
  assign y7605 = n17256 ;
  assign y7606 = ~n17258 ;
  assign y7607 = ~1'b0 ;
  assign y7608 = ~1'b0 ;
  assign y7609 = ~n11231 ;
  assign y7610 = ~n17259 ;
  assign y7611 = n17262 ;
  assign y7612 = n17264 ;
  assign y7613 = ~n17266 ;
  assign y7614 = ~n17270 ;
  assign y7615 = n17272 ;
  assign y7616 = n17274 ;
  assign y7617 = n17275 ;
  assign y7618 = n17277 ;
  assign y7619 = n17280 ;
  assign y7620 = 1'b0 ;
  assign y7621 = n17289 ;
  assign y7622 = ~n17296 ;
  assign y7623 = ~1'b0 ;
  assign y7624 = ~n17297 ;
  assign y7625 = ~n17299 ;
  assign y7626 = n17301 ;
  assign y7627 = n17302 ;
  assign y7628 = ~1'b0 ;
  assign y7629 = n17307 ;
  assign y7630 = n17308 ;
  assign y7631 = n17309 ;
  assign y7632 = n17311 ;
  assign y7633 = n17316 ;
  assign y7634 = n17323 ;
  assign y7635 = ~1'b0 ;
  assign y7636 = n17324 ;
  assign y7637 = n17327 ;
  assign y7638 = ~n17329 ;
  assign y7639 = ~n17334 ;
  assign y7640 = n17335 ;
  assign y7641 = n14659 ;
  assign y7642 = ~n17338 ;
  assign y7643 = ~n17342 ;
  assign y7644 = ~1'b0 ;
  assign y7645 = n17343 ;
  assign y7646 = n17355 ;
  assign y7647 = n17356 ;
  assign y7648 = ~n17357 ;
  assign y7649 = ~n17360 ;
  assign y7650 = ~n17365 ;
  assign y7651 = n4463 ;
  assign y7652 = ~n17367 ;
  assign y7653 = ~1'b0 ;
  assign y7654 = 1'b0 ;
  assign y7655 = ~1'b0 ;
  assign y7656 = n17373 ;
  assign y7657 = n17374 ;
  assign y7658 = n17376 ;
  assign y7659 = n17378 ;
  assign y7660 = ~1'b0 ;
  assign y7661 = n17383 ;
  assign y7662 = ~n791 ;
  assign y7663 = ~n17387 ;
  assign y7664 = n4944 ;
  assign y7665 = ~n17392 ;
  assign y7666 = n17396 ;
  assign y7667 = ~1'b0 ;
  assign y7668 = ~n17401 ;
  assign y7669 = ~1'b0 ;
  assign y7670 = ~n17402 ;
  assign y7671 = n17403 ;
  assign y7672 = ~n17404 ;
  assign y7673 = n17411 ;
  assign y7674 = ~1'b0 ;
  assign y7675 = ~n17415 ;
  assign y7676 = ~n17416 ;
  assign y7677 = ~n17418 ;
  assign y7678 = ~1'b0 ;
  assign y7679 = ~1'b0 ;
  assign y7680 = n17420 ;
  assign y7681 = ~1'b0 ;
  assign y7682 = n17428 ;
  assign y7683 = ~n17432 ;
  assign y7684 = ~n17434 ;
  assign y7685 = n17440 ;
  assign y7686 = ~n17449 ;
  assign y7687 = ~n17451 ;
  assign y7688 = n17462 ;
  assign y7689 = n17463 ;
  assign y7690 = ~n17466 ;
  assign y7691 = ~n17467 ;
  assign y7692 = n17468 ;
  assign y7693 = ~1'b0 ;
  assign y7694 = ~n17469 ;
  assign y7695 = ~n3090 ;
  assign y7696 = ~n17472 ;
  assign y7697 = ~n17484 ;
  assign y7698 = n11573 ;
  assign y7699 = ~n17487 ;
  assign y7700 = n17488 ;
  assign y7701 = n17491 ;
  assign y7702 = ~n17493 ;
  assign y7703 = n15618 ;
  assign y7704 = ~1'b0 ;
  assign y7705 = ~1'b0 ;
  assign y7706 = ~n17500 ;
  assign y7707 = n17502 ;
  assign y7708 = ~n17503 ;
  assign y7709 = n17505 ;
  assign y7710 = ~n17508 ;
  assign y7711 = ~n17511 ;
  assign y7712 = ~n962 ;
  assign y7713 = ~n17513 ;
  assign y7714 = ~1'b0 ;
  assign y7715 = ~1'b0 ;
  assign y7716 = n17514 ;
  assign y7717 = ~n17516 ;
  assign y7718 = n17523 ;
  assign y7719 = ~1'b0 ;
  assign y7720 = ~1'b0 ;
  assign y7721 = n17524 ;
  assign y7722 = n15308 ;
  assign y7723 = n17526 ;
  assign y7724 = ~n17536 ;
  assign y7725 = ~n17539 ;
  assign y7726 = n17541 ;
  assign y7727 = n17544 ;
  assign y7728 = ~1'b0 ;
  assign y7729 = ~n17546 ;
  assign y7730 = n17548 ;
  assign y7731 = ~n17550 ;
  assign y7732 = ~1'b0 ;
  assign y7733 = ~1'b0 ;
  assign y7734 = ~1'b0 ;
  assign y7735 = ~n17551 ;
  assign y7736 = ~n17552 ;
  assign y7737 = ~1'b0 ;
  assign y7738 = ~n17560 ;
  assign y7739 = ~1'b0 ;
  assign y7740 = n17561 ;
  assign y7741 = ~n17564 ;
  assign y7742 = ~n17565 ;
  assign y7743 = ~n17569 ;
  assign y7744 = ~1'b0 ;
  assign y7745 = ~1'b0 ;
  assign y7746 = ~1'b0 ;
  assign y7747 = n17572 ;
  assign y7748 = ~1'b0 ;
  assign y7749 = n17574 ;
  assign y7750 = n17578 ;
  assign y7751 = ~1'b0 ;
  assign y7752 = n17580 ;
  assign y7753 = ~n17583 ;
  assign y7754 = n17585 ;
  assign y7755 = n17587 ;
  assign y7756 = n17594 ;
  assign y7757 = ~n7614 ;
  assign y7758 = ~1'b0 ;
  assign y7759 = ~n17607 ;
  assign y7760 = ~n17610 ;
  assign y7761 = ~1'b0 ;
  assign y7762 = ~n17613 ;
  assign y7763 = ~1'b0 ;
  assign y7764 = n17617 ;
  assign y7765 = ~n17622 ;
  assign y7766 = ~n17623 ;
  assign y7767 = ~n17627 ;
  assign y7768 = ~n17628 ;
  assign y7769 = n17632 ;
  assign y7770 = ~n17633 ;
  assign y7771 = ~n17634 ;
  assign y7772 = ~n17635 ;
  assign y7773 = ~n17644 ;
  assign y7774 = ~1'b0 ;
  assign y7775 = n17645 ;
  assign y7776 = n17646 ;
  assign y7777 = ~n17648 ;
  assign y7778 = n17649 ;
  assign y7779 = ~1'b0 ;
  assign y7780 = ~1'b0 ;
  assign y7781 = ~1'b0 ;
  assign y7782 = n17653 ;
  assign y7783 = ~n17655 ;
  assign y7784 = ~1'b0 ;
  assign y7785 = ~1'b0 ;
  assign y7786 = ~n3039 ;
  assign y7787 = ~1'b0 ;
  assign y7788 = n17656 ;
  assign y7789 = ~1'b0 ;
  assign y7790 = n17664 ;
  assign y7791 = n17665 ;
  assign y7792 = ~n17673 ;
  assign y7793 = ~n17674 ;
  assign y7794 = n17676 ;
  assign y7795 = ~1'b0 ;
  assign y7796 = n17679 ;
  assign y7797 = ~n11636 ;
  assign y7798 = n17682 ;
  assign y7799 = ~n17685 ;
  assign y7800 = ~1'b0 ;
  assign y7801 = ~n8077 ;
  assign y7802 = ~n17690 ;
  assign y7803 = 1'b0 ;
  assign y7804 = n17698 ;
  assign y7805 = ~n17700 ;
  assign y7806 = n17704 ;
  assign y7807 = n17706 ;
  assign y7808 = ~n17708 ;
  assign y7809 = ~1'b0 ;
  assign y7810 = n17714 ;
  assign y7811 = n17717 ;
  assign y7812 = n17720 ;
  assign y7813 = ~1'b0 ;
  assign y7814 = ~1'b0 ;
  assign y7815 = ~1'b0 ;
  assign y7816 = ~n17722 ;
  assign y7817 = n17724 ;
  assign y7818 = ~1'b0 ;
  assign y7819 = ~1'b0 ;
  assign y7820 = ~n17729 ;
  assign y7821 = ~1'b0 ;
  assign y7822 = ~n17738 ;
  assign y7823 = 1'b0 ;
  assign y7824 = ~n17739 ;
  assign y7825 = ~1'b0 ;
  assign y7826 = n17741 ;
  assign y7827 = n17744 ;
  assign y7828 = ~1'b0 ;
  assign y7829 = n17752 ;
  assign y7830 = ~1'b0 ;
  assign y7831 = ~1'b0 ;
  assign y7832 = ~n17756 ;
  assign y7833 = ~n17763 ;
  assign y7834 = ~1'b0 ;
  assign y7835 = ~1'b0 ;
  assign y7836 = ~n17765 ;
  assign y7837 = ~n17767 ;
  assign y7838 = n17768 ;
  assign y7839 = n17769 ;
  assign y7840 = ~1'b0 ;
  assign y7841 = ~1'b0 ;
  assign y7842 = ~1'b0 ;
  assign y7843 = ~n17770 ;
  assign y7844 = ~1'b0 ;
  assign y7845 = n17776 ;
  assign y7846 = ~1'b0 ;
  assign y7847 = ~1'b0 ;
  assign y7848 = ~n17778 ;
  assign y7849 = ~1'b0 ;
  assign y7850 = n17782 ;
  assign y7851 = ~n17783 ;
  assign y7852 = n17791 ;
  assign y7853 = n17797 ;
  assign y7854 = ~1'b0 ;
  assign y7855 = n17798 ;
  assign y7856 = 1'b0 ;
  assign y7857 = ~n17802 ;
  assign y7858 = n17807 ;
  assign y7859 = ~1'b0 ;
  assign y7860 = ~1'b0 ;
  assign y7861 = n17811 ;
  assign y7862 = n17812 ;
  assign y7863 = ~1'b0 ;
  assign y7864 = ~n2612 ;
  assign y7865 = ~1'b0 ;
  assign y7866 = ~n17814 ;
  assign y7867 = ~n17827 ;
  assign y7868 = n17830 ;
  assign y7869 = n17832 ;
  assign y7870 = ~n17833 ;
  assign y7871 = n17834 ;
  assign y7872 = ~1'b0 ;
  assign y7873 = n7506 ;
  assign y7874 = ~n17835 ;
  assign y7875 = ~1'b0 ;
  assign y7876 = ~n17837 ;
  assign y7877 = n17839 ;
  assign y7878 = ~n17843 ;
  assign y7879 = ~n17844 ;
  assign y7880 = n17845 ;
  assign y7881 = ~n17846 ;
  assign y7882 = n17848 ;
  assign y7883 = ~n17857 ;
  assign y7884 = ~n17859 ;
  assign y7885 = n17862 ;
  assign y7886 = ~n17864 ;
  assign y7887 = n17865 ;
  assign y7888 = ~n17868 ;
  assign y7889 = ~n17873 ;
  assign y7890 = 1'b0 ;
  assign y7891 = n1118 ;
  assign y7892 = n17875 ;
  assign y7893 = ~n17883 ;
  assign y7894 = ~n17886 ;
  assign y7895 = ~n17891 ;
  assign y7896 = ~n17897 ;
  assign y7897 = ~n17898 ;
  assign y7898 = n17899 ;
  assign y7899 = n17901 ;
  assign y7900 = n17903 ;
  assign y7901 = ~1'b0 ;
  assign y7902 = n17904 ;
  assign y7903 = ~n2885 ;
  assign y7904 = ~n17906 ;
  assign y7905 = n17907 ;
  assign y7906 = n17910 ;
  assign y7907 = ~1'b0 ;
  assign y7908 = n17912 ;
  assign y7909 = n17916 ;
  assign y7910 = ~1'b0 ;
  assign y7911 = n17917 ;
  assign y7912 = n17923 ;
  assign y7913 = ~n17927 ;
  assign y7914 = ~n17928 ;
  assign y7915 = ~n17929 ;
  assign y7916 = ~n15886 ;
  assign y7917 = n17930 ;
  assign y7918 = n17938 ;
  assign y7919 = ~n17945 ;
  assign y7920 = ~1'b0 ;
  assign y7921 = n17946 ;
  assign y7922 = n17947 ;
  assign y7923 = n17948 ;
  assign y7924 = n571 ;
  assign y7925 = n17949 ;
  assign y7926 = ~n17950 ;
  assign y7927 = ~n17959 ;
  assign y7928 = ~n17963 ;
  assign y7929 = ~n11618 ;
  assign y7930 = ~n17965 ;
  assign y7931 = ~n17977 ;
  assign y7932 = n17979 ;
  assign y7933 = ~1'b0 ;
  assign y7934 = 1'b0 ;
  assign y7935 = n17980 ;
  assign y7936 = ~n17981 ;
  assign y7937 = ~1'b0 ;
  assign y7938 = ~n17983 ;
  assign y7939 = ~1'b0 ;
  assign y7940 = ~n17985 ;
  assign y7941 = ~1'b0 ;
  assign y7942 = n17989 ;
  assign y7943 = ~n17990 ;
  assign y7944 = n17995 ;
  assign y7945 = ~n17996 ;
  assign y7946 = ~1'b0 ;
  assign y7947 = ~n17997 ;
  assign y7948 = n17998 ;
  assign y7949 = ~n18000 ;
  assign y7950 = n18001 ;
  assign y7951 = ~1'b0 ;
  assign y7952 = ~1'b0 ;
  assign y7953 = n18005 ;
  assign y7954 = ~1'b0 ;
  assign y7955 = n18006 ;
  assign y7956 = ~n18012 ;
  assign y7957 = ~n18014 ;
  assign y7958 = ~1'b0 ;
  assign y7959 = ~n18015 ;
  assign y7960 = n18017 ;
  assign y7961 = ~n18023 ;
  assign y7962 = n18025 ;
  assign y7963 = n18027 ;
  assign y7964 = ~1'b0 ;
  assign y7965 = n18029 ;
  assign y7966 = n18030 ;
  assign y7967 = ~n18033 ;
  assign y7968 = n18034 ;
  assign y7969 = ~1'b0 ;
  assign y7970 = ~n18047 ;
  assign y7971 = n18051 ;
  assign y7972 = ~1'b0 ;
  assign y7973 = ~1'b0 ;
  assign y7974 = ~1'b0 ;
  assign y7975 = ~n18053 ;
  assign y7976 = ~1'b0 ;
  assign y7977 = ~n14711 ;
  assign y7978 = ~1'b0 ;
  assign y7979 = ~1'b0 ;
  assign y7980 = ~1'b0 ;
  assign y7981 = ~n6010 ;
  assign y7982 = ~1'b0 ;
  assign y7983 = n18057 ;
  assign y7984 = n18059 ;
  assign y7985 = ~1'b0 ;
  assign y7986 = n18060 ;
  assign y7987 = n18061 ;
  assign y7988 = n10222 ;
  assign y7989 = n18062 ;
  assign y7990 = n18063 ;
  assign y7991 = ~n18065 ;
  assign y7992 = ~n18066 ;
  assign y7993 = ~1'b0 ;
  assign y7994 = ~1'b0 ;
  assign y7995 = ~1'b0 ;
  assign y7996 = ~1'b0 ;
  assign y7997 = n18069 ;
  assign y7998 = n18072 ;
  assign y7999 = n18073 ;
  assign y8000 = n18079 ;
  assign y8001 = n18084 ;
  assign y8002 = ~n18090 ;
  assign y8003 = n18092 ;
  assign y8004 = n18093 ;
  assign y8005 = ~1'b0 ;
  assign y8006 = n18095 ;
  assign y8007 = ~n11982 ;
  assign y8008 = n18096 ;
  assign y8009 = n18097 ;
  assign y8010 = n18098 ;
  assign y8011 = ~1'b0 ;
  assign y8012 = ~n18102 ;
  assign y8013 = ~n16664 ;
  assign y8014 = ~n18104 ;
  assign y8015 = n18110 ;
  assign y8016 = n18118 ;
  assign y8017 = n18119 ;
  assign y8018 = ~n11969 ;
  assign y8019 = ~n18127 ;
  assign y8020 = ~1'b0 ;
  assign y8021 = ~1'b0 ;
  assign y8022 = ~1'b0 ;
  assign y8023 = ~n18129 ;
  assign y8024 = n18132 ;
  assign y8025 = n18134 ;
  assign y8026 = ~n18142 ;
  assign y8027 = ~n18145 ;
  assign y8028 = ~1'b0 ;
  assign y8029 = n18147 ;
  assign y8030 = ~n18148 ;
  assign y8031 = ~n18151 ;
  assign y8032 = n18152 ;
  assign y8033 = n18153 ;
  assign y8034 = ~n18154 ;
  assign y8035 = ~1'b0 ;
  assign y8036 = ~n18157 ;
  assign y8037 = n18160 ;
  assign y8038 = n18166 ;
  assign y8039 = ~n18169 ;
  assign y8040 = n18172 ;
  assign y8041 = ~1'b0 ;
  assign y8042 = ~1'b0 ;
  assign y8043 = n18175 ;
  assign y8044 = ~n18180 ;
  assign y8045 = n18188 ;
  assign y8046 = ~n18193 ;
  assign y8047 = n18195 ;
  assign y8048 = n18198 ;
  assign y8049 = n18202 ;
  assign y8050 = ~n18205 ;
  assign y8051 = ~1'b0 ;
  assign y8052 = ~n18207 ;
  assign y8053 = n18208 ;
  assign y8054 = n18211 ;
  assign y8055 = n18213 ;
  assign y8056 = n10433 ;
  assign y8057 = ~n18218 ;
  assign y8058 = ~n18220 ;
  assign y8059 = ~n18223 ;
  assign y8060 = ~n18224 ;
  assign y8061 = ~n18226 ;
  assign y8062 = ~n18227 ;
  assign y8063 = ~n18228 ;
  assign y8064 = ~n18231 ;
  assign y8065 = n18237 ;
  assign y8066 = ~1'b0 ;
  assign y8067 = ~1'b0 ;
  assign y8068 = ~1'b0 ;
  assign y8069 = ~1'b0 ;
  assign y8070 = n3120 ;
  assign y8071 = ~n18241 ;
  assign y8072 = n18243 ;
  assign y8073 = ~1'b0 ;
  assign y8074 = ~1'b0 ;
  assign y8075 = n18248 ;
  assign y8076 = ~n18249 ;
  assign y8077 = ~n18250 ;
  assign y8078 = ~1'b0 ;
  assign y8079 = ~n18255 ;
  assign y8080 = ~n18256 ;
  assign y8081 = ~n13197 ;
  assign y8082 = ~n18260 ;
  assign y8083 = ~n18264 ;
  assign y8084 = ~n18265 ;
  assign y8085 = ~1'b0 ;
  assign y8086 = n18266 ;
  assign y8087 = ~1'b0 ;
  assign y8088 = ~n18272 ;
  assign y8089 = n18274 ;
  assign y8090 = ~n4949 ;
  assign y8091 = ~1'b0 ;
  assign y8092 = ~1'b0 ;
  assign y8093 = ~n18282 ;
  assign y8094 = ~1'b0 ;
  assign y8095 = ~n18284 ;
  assign y8096 = ~n18291 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = n18157 ;
  assign y8099 = ~n18292 ;
  assign y8100 = n18299 ;
  assign y8101 = n18301 ;
  assign y8102 = ~n18304 ;
  assign y8103 = n18305 ;
  assign y8104 = ~1'b0 ;
  assign y8105 = ~1'b0 ;
  assign y8106 = ~n18314 ;
  assign y8107 = ~1'b0 ;
  assign y8108 = n18316 ;
  assign y8109 = n18320 ;
  assign y8110 = ~n18324 ;
  assign y8111 = ~1'b0 ;
  assign y8112 = ~n18325 ;
  assign y8113 = ~n18326 ;
  assign y8114 = ~n18327 ;
  assign y8115 = ~1'b0 ;
  assign y8116 = ~n18331 ;
  assign y8117 = ~n18333 ;
  assign y8118 = n18338 ;
  assign y8119 = ~1'b0 ;
  assign y8120 = n18341 ;
  assign y8121 = ~1'b0 ;
  assign y8122 = ~n18346 ;
  assign y8123 = n18347 ;
  assign y8124 = ~1'b0 ;
  assign y8125 = ~1'b0 ;
  assign y8126 = ~n18348 ;
  assign y8127 = ~1'b0 ;
  assign y8128 = n18349 ;
  assign y8129 = n18350 ;
  assign y8130 = ~1'b0 ;
  assign y8131 = ~1'b0 ;
  assign y8132 = ~n2677 ;
  assign y8133 = ~1'b0 ;
  assign y8134 = ~n18356 ;
  assign y8135 = ~n18359 ;
  assign y8136 = n18360 ;
  assign y8137 = ~n18361 ;
  assign y8138 = n18363 ;
  assign y8139 = 1'b0 ;
  assign y8140 = n18365 ;
  assign y8141 = ~1'b0 ;
  assign y8142 = ~n18369 ;
  assign y8143 = ~1'b0 ;
  assign y8144 = ~1'b0 ;
  assign y8145 = n2387 ;
  assign y8146 = ~1'b0 ;
  assign y8147 = ~n18373 ;
  assign y8148 = ~n18374 ;
  assign y8149 = ~n18375 ;
  assign y8150 = ~1'b0 ;
  assign y8151 = ~n18378 ;
  assign y8152 = ~n18383 ;
  assign y8153 = ~1'b0 ;
  assign y8154 = n18384 ;
  assign y8155 = n18386 ;
  assign y8156 = n18388 ;
  assign y8157 = ~n18390 ;
  assign y8158 = n18391 ;
  assign y8159 = ~n18394 ;
  assign y8160 = n18395 ;
  assign y8161 = ~n18396 ;
  assign y8162 = ~n18402 ;
  assign y8163 = n18408 ;
  assign y8164 = ~n18410 ;
  assign y8165 = ~n18414 ;
  assign y8166 = ~n18416 ;
  assign y8167 = n18417 ;
  assign y8168 = ~1'b0 ;
  assign y8169 = n18419 ;
  assign y8170 = n18420 ;
  assign y8171 = ~n18426 ;
  assign y8172 = ~n18430 ;
  assign y8173 = ~n6524 ;
  assign y8174 = ~1'b0 ;
  assign y8175 = n18431 ;
  assign y8176 = ~n18435 ;
  assign y8177 = n18436 ;
  assign y8178 = ~1'b0 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = ~1'b0 ;
  assign y8181 = n18447 ;
  assign y8182 = ~n9479 ;
  assign y8183 = ~n18459 ;
  assign y8184 = n18465 ;
  assign y8185 = n18467 ;
  assign y8186 = ~n18469 ;
  assign y8187 = ~1'b0 ;
  assign y8188 = ~n18473 ;
  assign y8189 = ~1'b0 ;
  assign y8190 = ~1'b0 ;
  assign y8191 = n18475 ;
  assign y8192 = ~n18476 ;
  assign y8193 = ~1'b0 ;
  assign y8194 = ~1'b0 ;
  assign y8195 = ~n4436 ;
  assign y8196 = ~n18479 ;
  assign y8197 = ~n18480 ;
  assign y8198 = n18485 ;
  assign y8199 = ~1'b0 ;
  assign y8200 = ~n18487 ;
  assign y8201 = n18492 ;
  assign y8202 = n18493 ;
  assign y8203 = n18495 ;
  assign y8204 = ~1'b0 ;
  assign y8205 = ~1'b0 ;
  assign y8206 = n18496 ;
  assign y8207 = n18497 ;
  assign y8208 = ~n18501 ;
  assign y8209 = ~n18513 ;
  assign y8210 = ~1'b0 ;
  assign y8211 = n18514 ;
  assign y8212 = n18518 ;
  assign y8213 = n18520 ;
  assign y8214 = ~1'b0 ;
  assign y8215 = n18525 ;
  assign y8216 = n18531 ;
  assign y8217 = ~n18536 ;
  assign y8218 = n18538 ;
  assign y8219 = ~n18539 ;
  assign y8220 = n18542 ;
  assign y8221 = n18547 ;
  assign y8222 = ~n18550 ;
  assign y8223 = n18552 ;
  assign y8224 = ~1'b0 ;
  assign y8225 = n18555 ;
  assign y8226 = ~1'b0 ;
  assign y8227 = ~n18560 ;
  assign y8228 = 1'b0 ;
  assign y8229 = n18563 ;
  assign y8230 = ~1'b0 ;
  assign y8231 = n18566 ;
  assign y8232 = ~n18578 ;
  assign y8233 = ~1'b0 ;
  assign y8234 = ~n18586 ;
  assign y8235 = ~1'b0 ;
  assign y8236 = ~n18591 ;
  assign y8237 = ~n18593 ;
  assign y8238 = ~n18594 ;
  assign y8239 = ~1'b0 ;
  assign y8240 = ~n18596 ;
  assign y8241 = n18597 ;
  assign y8242 = ~n18602 ;
  assign y8243 = ~n18608 ;
  assign y8244 = n18609 ;
  assign y8245 = ~1'b0 ;
  assign y8246 = ~n18613 ;
  assign y8247 = n18614 ;
  assign y8248 = ~n18628 ;
  assign y8249 = ~1'b0 ;
  assign y8250 = ~1'b0 ;
  assign y8251 = ~n18637 ;
  assign y8252 = ~1'b0 ;
  assign y8253 = ~1'b0 ;
  assign y8254 = ~n18638 ;
  assign y8255 = ~n18640 ;
  assign y8256 = ~1'b0 ;
  assign y8257 = n18642 ;
  assign y8258 = ~n18645 ;
  assign y8259 = n18646 ;
  assign y8260 = ~n18651 ;
  assign y8261 = n18654 ;
  assign y8262 = n18655 ;
  assign y8263 = ~1'b0 ;
  assign y8264 = n18658 ;
  assign y8265 = ~1'b0 ;
  assign y8266 = ~n18660 ;
  assign y8267 = 1'b0 ;
  assign y8268 = ~1'b0 ;
  assign y8269 = ~1'b0 ;
  assign y8270 = ~n13384 ;
  assign y8271 = n18664 ;
  assign y8272 = n18667 ;
  assign y8273 = ~1'b0 ;
  assign y8274 = n18668 ;
  assign y8275 = ~1'b0 ;
  assign y8276 = ~n18671 ;
  assign y8277 = ~n18672 ;
  assign y8278 = n18674 ;
  assign y8279 = ~1'b0 ;
  assign y8280 = ~n18677 ;
  assign y8281 = ~1'b0 ;
  assign y8282 = ~n18683 ;
  assign y8283 = n18687 ;
  assign y8284 = ~1'b0 ;
  assign y8285 = ~n18688 ;
  assign y8286 = n18689 ;
  assign y8287 = ~1'b0 ;
  assign y8288 = n18701 ;
  assign y8289 = ~1'b0 ;
  assign y8290 = ~n18706 ;
  assign y8291 = ~n18707 ;
  assign y8292 = ~n18710 ;
  assign y8293 = ~1'b0 ;
  assign y8294 = n18712 ;
  assign y8295 = ~n18717 ;
  assign y8296 = ~n18721 ;
  assign y8297 = ~n18725 ;
  assign y8298 = ~n18726 ;
  assign y8299 = ~1'b0 ;
  assign y8300 = ~n18731 ;
  assign y8301 = n18732 ;
  assign y8302 = ~n18736 ;
  assign y8303 = ~1'b0 ;
  assign y8304 = n18757 ;
  assign y8305 = ~n15956 ;
  assign y8306 = ~n18758 ;
  assign y8307 = n18759 ;
  assign y8308 = ~n18763 ;
  assign y8309 = ~n18764 ;
  assign y8310 = ~1'b0 ;
  assign y8311 = n18765 ;
  assign y8312 = ~n18766 ;
  assign y8313 = ~n18768 ;
  assign y8314 = ~n18771 ;
  assign y8315 = ~n18777 ;
  assign y8316 = n18787 ;
  assign y8317 = n18788 ;
  assign y8318 = ~n18789 ;
  assign y8319 = ~n18791 ;
  assign y8320 = n18792 ;
  assign y8321 = n18793 ;
  assign y8322 = ~n18796 ;
  assign y8323 = ~1'b0 ;
  assign y8324 = 1'b0 ;
  assign y8325 = n18797 ;
  assign y8326 = ~n18800 ;
  assign y8327 = ~n18802 ;
  assign y8328 = ~n18803 ;
  assign y8329 = ~1'b0 ;
  assign y8330 = ~n18808 ;
  assign y8331 = ~1'b0 ;
  assign y8332 = ~1'b0 ;
  assign y8333 = ~n18818 ;
  assign y8334 = ~1'b0 ;
  assign y8335 = n18822 ;
  assign y8336 = n18823 ;
  assign y8337 = ~n18824 ;
  assign y8338 = n18829 ;
  assign y8339 = ~1'b0 ;
  assign y8340 = ~1'b0 ;
  assign y8341 = n18840 ;
  assign y8342 = ~n18846 ;
  assign y8343 = ~n18848 ;
  assign y8344 = ~n18849 ;
  assign y8345 = ~1'b0 ;
  assign y8346 = ~1'b0 ;
  assign y8347 = ~1'b0 ;
  assign y8348 = n18858 ;
  assign y8349 = n18862 ;
  assign y8350 = ~n18870 ;
  assign y8351 = 1'b0 ;
  assign y8352 = n18873 ;
  assign y8353 = n18874 ;
  assign y8354 = n18879 ;
  assign y8355 = 1'b0 ;
  assign y8356 = ~1'b0 ;
  assign y8357 = n18880 ;
  assign y8358 = ~1'b0 ;
  assign y8359 = n18885 ;
  assign y8360 = n4067 ;
  assign y8361 = ~1'b0 ;
  assign y8362 = ~n18890 ;
  assign y8363 = ~n18893 ;
  assign y8364 = ~n18894 ;
  assign y8365 = ~n18895 ;
  assign y8366 = n18896 ;
  assign y8367 = ~n18899 ;
  assign y8368 = ~n18905 ;
  assign y8369 = ~n18910 ;
  assign y8370 = n18913 ;
  assign y8371 = n18914 ;
  assign y8372 = ~1'b0 ;
  assign y8373 = n18917 ;
  assign y8374 = ~n18921 ;
  assign y8375 = ~n18929 ;
  assign y8376 = n18930 ;
  assign y8377 = ~1'b0 ;
  assign y8378 = ~n18931 ;
  assign y8379 = n5897 ;
  assign y8380 = n18932 ;
  assign y8381 = ~1'b0 ;
  assign y8382 = ~n18933 ;
  assign y8383 = n18941 ;
  assign y8384 = n18943 ;
  assign y8385 = ~n18944 ;
  assign y8386 = ~1'b0 ;
  assign y8387 = n18947 ;
  assign y8388 = 1'b0 ;
  assign y8389 = ~n18952 ;
  assign y8390 = ~1'b0 ;
  assign y8391 = n18957 ;
  assign y8392 = n18959 ;
  assign y8393 = ~n18966 ;
  assign y8394 = n18969 ;
  assign y8395 = ~1'b0 ;
  assign y8396 = ~1'b0 ;
  assign y8397 = n18974 ;
  assign y8398 = ~n18975 ;
  assign y8399 = n18976 ;
  assign y8400 = ~n18989 ;
  assign y8401 = ~n18990 ;
  assign y8402 = n6139 ;
  assign y8403 = ~n18991 ;
  assign y8404 = ~1'b0 ;
  assign y8405 = ~n18992 ;
  assign y8406 = ~1'b0 ;
  assign y8407 = ~1'b0 ;
  assign y8408 = ~n8936 ;
  assign y8409 = ~n18997 ;
  assign y8410 = ~n18999 ;
  assign y8411 = ~n19009 ;
  assign y8412 = n19010 ;
  assign y8413 = n19016 ;
  assign y8414 = ~n7468 ;
  assign y8415 = n19017 ;
  assign y8416 = ~n19018 ;
  assign y8417 = ~n19021 ;
  assign y8418 = n19022 ;
  assign y8419 = n19023 ;
  assign y8420 = ~1'b0 ;
  assign y8421 = ~1'b0 ;
  assign y8422 = n19024 ;
  assign y8423 = n19026 ;
  assign y8424 = ~n19028 ;
  assign y8425 = ~n19029 ;
  assign y8426 = ~1'b0 ;
  assign y8427 = ~1'b0 ;
  assign y8428 = ~n19034 ;
  assign y8429 = n11919 ;
  assign y8430 = n19039 ;
  assign y8431 = n19042 ;
  assign y8432 = ~1'b0 ;
  assign y8433 = 1'b0 ;
  assign y8434 = ~n19045 ;
  assign y8435 = ~1'b0 ;
  assign y8436 = ~n19047 ;
  assign y8437 = ~n19051 ;
  assign y8438 = ~n19053 ;
  assign y8439 = n19055 ;
  assign y8440 = ~n19057 ;
  assign y8441 = n19062 ;
  assign y8442 = ~1'b0 ;
  assign y8443 = ~n19064 ;
  assign y8444 = n19065 ;
  assign y8445 = ~n19066 ;
  assign y8446 = ~1'b0 ;
  assign y8447 = ~n19068 ;
  assign y8448 = ~1'b0 ;
  assign y8449 = ~n19071 ;
  assign y8450 = ~1'b0 ;
  assign y8451 = ~1'b0 ;
  assign y8452 = n19072 ;
  assign y8453 = ~n15799 ;
  assign y8454 = ~n19074 ;
  assign y8455 = n19077 ;
  assign y8456 = ~1'b0 ;
  assign y8457 = ~n19080 ;
  assign y8458 = ~n19083 ;
  assign y8459 = n19084 ;
  assign y8460 = ~n19086 ;
  assign y8461 = n19090 ;
  assign y8462 = ~n19094 ;
  assign y8463 = ~1'b0 ;
  assign y8464 = ~1'b0 ;
  assign y8465 = ~n19095 ;
  assign y8466 = n19096 ;
  assign y8467 = ~n19098 ;
  assign y8468 = n19099 ;
  assign y8469 = ~n19100 ;
  assign y8470 = ~n19101 ;
  assign y8471 = ~n19104 ;
  assign y8472 = ~1'b0 ;
  assign y8473 = ~n19105 ;
  assign y8474 = ~1'b0 ;
  assign y8475 = ~n19109 ;
  assign y8476 = ~n19139 ;
  assign y8477 = ~1'b0 ;
  assign y8478 = ~1'b0 ;
  assign y8479 = n19140 ;
  assign y8480 = 1'b0 ;
  assign y8481 = n19141 ;
  assign y8482 = ~n11973 ;
  assign y8483 = ~n19143 ;
  assign y8484 = ~n576 ;
  assign y8485 = ~n19144 ;
  assign y8486 = n19147 ;
  assign y8487 = n19152 ;
  assign y8488 = ~1'b0 ;
  assign y8489 = ~n19155 ;
  assign y8490 = ~n19158 ;
  assign y8491 = n19161 ;
  assign y8492 = n19163 ;
  assign y8493 = ~1'b0 ;
  assign y8494 = ~n19167 ;
  assign y8495 = n19175 ;
  assign y8496 = ~n19181 ;
  assign y8497 = n19182 ;
  assign y8498 = n19183 ;
  assign y8499 = n19185 ;
  assign y8500 = ~1'b0 ;
  assign y8501 = ~1'b0 ;
  assign y8502 = ~n3923 ;
  assign y8503 = ~n19190 ;
  assign y8504 = ~1'b0 ;
  assign y8505 = n19193 ;
  assign y8506 = n19194 ;
  assign y8507 = n19195 ;
  assign y8508 = n19198 ;
  assign y8509 = n19199 ;
  assign y8510 = n19200 ;
  assign y8511 = n19205 ;
  assign y8512 = n19214 ;
  assign y8513 = ~1'b0 ;
  assign y8514 = ~n19218 ;
  assign y8515 = n19223 ;
  assign y8516 = ~1'b0 ;
  assign y8517 = n19226 ;
  assign y8518 = n14385 ;
  assign y8519 = n19229 ;
  assign y8520 = 1'b0 ;
  assign y8521 = n3825 ;
  assign y8522 = n5706 ;
  assign y8523 = ~1'b0 ;
  assign y8524 = n19232 ;
  assign y8525 = n19235 ;
  assign y8526 = ~n19242 ;
  assign y8527 = ~n19244 ;
  assign y8528 = ~n19245 ;
  assign y8529 = n19250 ;
  assign y8530 = n19260 ;
  assign y8531 = n19261 ;
  assign y8532 = ~1'b0 ;
  assign y8533 = ~n19265 ;
  assign y8534 = n19268 ;
  assign y8535 = ~n19269 ;
  assign y8536 = n19272 ;
  assign y8537 = n19273 ;
  assign y8538 = ~n19281 ;
  assign y8539 = ~n19285 ;
  assign y8540 = ~n19288 ;
  assign y8541 = ~n19296 ;
  assign y8542 = 1'b0 ;
  assign y8543 = n17851 ;
  assign y8544 = n9230 ;
  assign y8545 = 1'b0 ;
  assign y8546 = ~n19297 ;
  assign y8547 = ~n19298 ;
  assign y8548 = n19302 ;
  assign y8549 = ~n19308 ;
  assign y8550 = ~1'b0 ;
  assign y8551 = ~n19309 ;
  assign y8552 = ~n19315 ;
  assign y8553 = 1'b0 ;
  assign y8554 = ~n19316 ;
  assign y8555 = ~n19319 ;
  assign y8556 = n19320 ;
  assign y8557 = n19321 ;
  assign y8558 = ~n19327 ;
  assign y8559 = n19330 ;
  assign y8560 = n19332 ;
  assign y8561 = ~1'b0 ;
  assign y8562 = ~n19337 ;
  assign y8563 = ~n19340 ;
  assign y8564 = ~n19341 ;
  assign y8565 = ~n19342 ;
  assign y8566 = ~1'b0 ;
  assign y8567 = n19351 ;
  assign y8568 = ~1'b0 ;
  assign y8569 = ~1'b0 ;
  assign y8570 = ~n19352 ;
  assign y8571 = ~n19353 ;
  assign y8572 = ~n19355 ;
  assign y8573 = n19358 ;
  assign y8574 = n19359 ;
  assign y8575 = ~1'b0 ;
  assign y8576 = ~n19365 ;
  assign y8577 = n19370 ;
  assign y8578 = ~n19371 ;
  assign y8579 = ~n19379 ;
  assign y8580 = n19383 ;
  assign y8581 = ~1'b0 ;
  assign y8582 = ~1'b0 ;
  assign y8583 = ~n19384 ;
  assign y8584 = ~1'b0 ;
  assign y8585 = ~1'b0 ;
  assign y8586 = ~n19390 ;
  assign y8587 = ~n19393 ;
  assign y8588 = n19396 ;
  assign y8589 = n19402 ;
  assign y8590 = n19405 ;
  assign y8591 = ~1'b0 ;
  assign y8592 = 1'b0 ;
  assign y8593 = ~n19409 ;
  assign y8594 = ~1'b0 ;
  assign y8595 = n19411 ;
  assign y8596 = n19412 ;
  assign y8597 = ~n19413 ;
  assign y8598 = ~n19414 ;
  assign y8599 = 1'b0 ;
  assign y8600 = 1'b0 ;
  assign y8601 = ~n19417 ;
  assign y8602 = n19421 ;
  assign y8603 = n7896 ;
  assign y8604 = n19422 ;
  assign y8605 = ~n19425 ;
  assign y8606 = ~n19427 ;
  assign y8607 = n19431 ;
  assign y8608 = n19435 ;
  assign y8609 = ~1'b0 ;
  assign y8610 = ~1'b0 ;
  assign y8611 = n9298 ;
  assign y8612 = ~1'b0 ;
  assign y8613 = ~n19441 ;
  assign y8614 = ~1'b0 ;
  assign y8615 = n19444 ;
  assign y8616 = n19446 ;
  assign y8617 = ~n19448 ;
  assign y8618 = n19451 ;
  assign y8619 = n5244 ;
  assign y8620 = ~n1951 ;
  assign y8621 = ~1'b0 ;
  assign y8622 = ~n19461 ;
  assign y8623 = n19467 ;
  assign y8624 = ~1'b0 ;
  assign y8625 = ~n19468 ;
  assign y8626 = ~1'b0 ;
  assign y8627 = ~1'b0 ;
  assign y8628 = ~1'b0 ;
  assign y8629 = n19470 ;
  assign y8630 = ~n19472 ;
  assign y8631 = n19477 ;
  assign y8632 = ~1'b0 ;
  assign y8633 = ~n19478 ;
  assign y8634 = n774 ;
  assign y8635 = n19480 ;
  assign y8636 = ~1'b0 ;
  assign y8637 = ~n19483 ;
  assign y8638 = n19487 ;
  assign y8639 = ~n19489 ;
  assign y8640 = ~1'b0 ;
  assign y8641 = ~n19493 ;
  assign y8642 = n19494 ;
  assign y8643 = ~n19496 ;
  assign y8644 = ~1'b0 ;
  assign y8645 = ~n19499 ;
  assign y8646 = n19506 ;
  assign y8647 = ~n19507 ;
  assign y8648 = n19510 ;
  assign y8649 = ~n19513 ;
  assign y8650 = ~n19515 ;
  assign y8651 = ~n19521 ;
  assign y8652 = ~1'b0 ;
  assign y8653 = n19523 ;
  assign y8654 = n19524 ;
  assign y8655 = ~1'b0 ;
  assign y8656 = n19528 ;
  assign y8657 = ~n19532 ;
  assign y8658 = n19543 ;
  assign y8659 = 1'b0 ;
  assign y8660 = ~1'b0 ;
  assign y8661 = n19547 ;
  assign y8662 = n19548 ;
  assign y8663 = ~1'b0 ;
  assign y8664 = ~n19551 ;
  assign y8665 = 1'b0 ;
  assign y8666 = ~1'b0 ;
  assign y8667 = n19555 ;
  assign y8668 = ~n19559 ;
  assign y8669 = ~1'b0 ;
  assign y8670 = ~1'b0 ;
  assign y8671 = ~1'b0 ;
  assign y8672 = ~n19565 ;
  assign y8673 = ~1'b0 ;
  assign y8674 = ~n19567 ;
  assign y8675 = ~1'b0 ;
  assign y8676 = ~n1818 ;
  assign y8677 = ~n19578 ;
  assign y8678 = ~1'b0 ;
  assign y8679 = ~1'b0 ;
  assign y8680 = n19579 ;
  assign y8681 = n19587 ;
  assign y8682 = n19588 ;
  assign y8683 = ~n19591 ;
  assign y8684 = ~1'b0 ;
  assign y8685 = n19592 ;
  assign y8686 = n19593 ;
  assign y8687 = n11111 ;
  assign y8688 = n19594 ;
  assign y8689 = ~1'b0 ;
  assign y8690 = ~1'b0 ;
  assign y8691 = ~n19597 ;
  assign y8692 = ~1'b0 ;
  assign y8693 = ~n19605 ;
  assign y8694 = n19607 ;
  assign y8695 = ~n19610 ;
  assign y8696 = ~1'b0 ;
  assign y8697 = n19611 ;
  assign y8698 = n19615 ;
  assign y8699 = n19619 ;
  assign y8700 = ~n19623 ;
  assign y8701 = n19625 ;
  assign y8702 = ~1'b0 ;
  assign y8703 = ~n19629 ;
  assign y8704 = ~1'b0 ;
  assign y8705 = n19632 ;
  assign y8706 = ~1'b0 ;
  assign y8707 = ~n19633 ;
  assign y8708 = n19634 ;
  assign y8709 = ~n19638 ;
  assign y8710 = ~n19642 ;
  assign y8711 = 1'b0 ;
  assign y8712 = ~n19648 ;
  assign y8713 = n19652 ;
  assign y8714 = ~1'b0 ;
  assign y8715 = n19655 ;
  assign y8716 = ~1'b0 ;
  assign y8717 = ~n19656 ;
  assign y8718 = ~1'b0 ;
  assign y8719 = ~n19666 ;
  assign y8720 = ~n19667 ;
  assign y8721 = n19668 ;
  assign y8722 = ~n19670 ;
  assign y8723 = ~n19673 ;
  assign y8724 = ~1'b0 ;
  assign y8725 = ~n19675 ;
  assign y8726 = ~1'b0 ;
  assign y8727 = ~n19679 ;
  assign y8728 = n6261 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = ~1'b0 ;
  assign y8731 = ~n19684 ;
  assign y8732 = ~n19697 ;
  assign y8733 = n19700 ;
  assign y8734 = ~n19705 ;
  assign y8735 = ~1'b0 ;
  assign y8736 = n19706 ;
  assign y8737 = ~n19709 ;
  assign y8738 = n19712 ;
  assign y8739 = ~1'b0 ;
  assign y8740 = ~n19713 ;
  assign y8741 = n9507 ;
  assign y8742 = ~1'b0 ;
  assign y8743 = ~n19715 ;
  assign y8744 = ~n19719 ;
  assign y8745 = ~n19726 ;
  assign y8746 = ~n19732 ;
  assign y8747 = ~n19733 ;
  assign y8748 = ~n19734 ;
  assign y8749 = ~1'b0 ;
  assign y8750 = ~1'b0 ;
  assign y8751 = n19737 ;
  assign y8752 = ~1'b0 ;
  assign y8753 = ~1'b0 ;
  assign y8754 = ~n19739 ;
  assign y8755 = ~1'b0 ;
  assign y8756 = n6126 ;
  assign y8757 = ~n19748 ;
  assign y8758 = ~1'b0 ;
  assign y8759 = n19749 ;
  assign y8760 = ~n19750 ;
  assign y8761 = ~1'b0 ;
  assign y8762 = ~1'b0 ;
  assign y8763 = ~n19756 ;
  assign y8764 = ~n19763 ;
  assign y8765 = ~n19767 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = ~1'b0 ;
  assign y8768 = n19771 ;
  assign y8769 = n19772 ;
  assign y8770 = 1'b0 ;
  assign y8771 = ~n19776 ;
  assign y8772 = ~1'b0 ;
  assign y8773 = n19781 ;
  assign y8774 = ~1'b0 ;
  assign y8775 = ~1'b0 ;
  assign y8776 = ~n19782 ;
  assign y8777 = ~n19783 ;
  assign y8778 = n19785 ;
  assign y8779 = ~n19788 ;
  assign y8780 = ~1'b0 ;
  assign y8781 = n19790 ;
  assign y8782 = ~1'b0 ;
  assign y8783 = ~n19792 ;
  assign y8784 = ~1'b0 ;
  assign y8785 = ~1'b0 ;
  assign y8786 = n19795 ;
  assign y8787 = n19800 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = n19803 ;
  assign y8790 = ~n19805 ;
  assign y8791 = ~n2621 ;
  assign y8792 = n19811 ;
  assign y8793 = ~n19812 ;
  assign y8794 = ~n19813 ;
  assign y8795 = 1'b0 ;
  assign y8796 = ~n19817 ;
  assign y8797 = ~n19819 ;
  assign y8798 = ~1'b0 ;
  assign y8799 = ~n19824 ;
  assign y8800 = n19828 ;
  assign y8801 = n19829 ;
  assign y8802 = ~n19835 ;
  assign y8803 = ~n19839 ;
  assign y8804 = ~1'b0 ;
  assign y8805 = n19840 ;
  assign y8806 = ~n19842 ;
  assign y8807 = ~n19843 ;
  assign y8808 = n19847 ;
  assign y8809 = n19848 ;
  assign y8810 = ~1'b0 ;
  assign y8811 = ~n19850 ;
  assign y8812 = ~1'b0 ;
  assign y8813 = ~1'b0 ;
  assign y8814 = n19857 ;
  assign y8815 = n19860 ;
  assign y8816 = n19861 ;
  assign y8817 = ~n19862 ;
  assign y8818 = n968 ;
  assign y8819 = ~n19865 ;
  assign y8820 = n19869 ;
  assign y8821 = ~n19874 ;
  assign y8822 = ~1'b0 ;
  assign y8823 = n19876 ;
  assign y8824 = n19879 ;
  assign y8825 = n19881 ;
  assign y8826 = n19883 ;
  assign y8827 = n19889 ;
  assign y8828 = ~n6152 ;
  assign y8829 = n19890 ;
  assign y8830 = ~n19892 ;
  assign y8831 = ~1'b0 ;
  assign y8832 = ~1'b0 ;
  assign y8833 = ~n19897 ;
  assign y8834 = ~1'b0 ;
  assign y8835 = ~1'b0 ;
  assign y8836 = ~n19898 ;
  assign y8837 = ~n19899 ;
  assign y8838 = n19905 ;
  assign y8839 = ~n19911 ;
  assign y8840 = ~n19913 ;
  assign y8841 = ~n19915 ;
  assign y8842 = ~1'b0 ;
  assign y8843 = n19922 ;
  assign y8844 = ~n19924 ;
  assign y8845 = n19927 ;
  assign y8846 = ~n19938 ;
  assign y8847 = ~n5837 ;
  assign y8848 = n15218 ;
  assign y8849 = ~n19943 ;
  assign y8850 = n19948 ;
  assign y8851 = ~1'b0 ;
  assign y8852 = n19950 ;
  assign y8853 = ~n19954 ;
  assign y8854 = ~n19955 ;
  assign y8855 = ~1'b0 ;
  assign y8856 = n19957 ;
  assign y8857 = n19958 ;
  assign y8858 = ~n19213 ;
  assign y8859 = n19969 ;
  assign y8860 = n19976 ;
  assign y8861 = ~n19981 ;
  assign y8862 = n19982 ;
  assign y8863 = ~1'b0 ;
  assign y8864 = ~n19984 ;
  assign y8865 = ~n19989 ;
  assign y8866 = ~1'b0 ;
  assign y8867 = n19991 ;
  assign y8868 = n19994 ;
  assign y8869 = ~n19995 ;
  assign y8870 = ~1'b0 ;
  assign y8871 = n19997 ;
  assign y8872 = n20000 ;
  assign y8873 = n20001 ;
  assign y8874 = ~n17712 ;
  assign y8875 = ~1'b0 ;
  assign y8876 = ~n20005 ;
  assign y8877 = ~1'b0 ;
  assign y8878 = n20007 ;
  assign y8879 = ~1'b0 ;
  assign y8880 = ~n18570 ;
  assign y8881 = ~1'b0 ;
  assign y8882 = ~n20017 ;
  assign y8883 = ~n20018 ;
  assign y8884 = ~n16419 ;
  assign y8885 = n20026 ;
  assign y8886 = n14296 ;
  assign y8887 = ~1'b0 ;
  assign y8888 = ~1'b0 ;
  assign y8889 = ~1'b0 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = n20030 ;
  assign y8892 = 1'b0 ;
  assign y8893 = n10942 ;
  assign y8894 = ~n20035 ;
  assign y8895 = ~n20039 ;
  assign y8896 = ~n20041 ;
  assign y8897 = ~1'b0 ;
  assign y8898 = n20045 ;
  assign y8899 = n20046 ;
  assign y8900 = ~n20047 ;
  assign y8901 = n20048 ;
  assign y8902 = n20052 ;
  assign y8903 = ~n20055 ;
  assign y8904 = ~1'b0 ;
  assign y8905 = ~n20057 ;
  assign y8906 = ~n20060 ;
  assign y8907 = ~n20064 ;
  assign y8908 = ~n20067 ;
  assign y8909 = 1'b0 ;
  assign y8910 = n20069 ;
  assign y8911 = n20074 ;
  assign y8912 = n20075 ;
  assign y8913 = n20078 ;
  assign y8914 = ~n20081 ;
  assign y8915 = n20085 ;
  assign y8916 = ~n20086 ;
  assign y8917 = ~n20087 ;
  assign y8918 = n20094 ;
  assign y8919 = ~1'b0 ;
  assign y8920 = n20095 ;
  assign y8921 = ~1'b0 ;
  assign y8922 = ~1'b0 ;
  assign y8923 = n20099 ;
  assign y8924 = n20101 ;
  assign y8925 = n20103 ;
  assign y8926 = n17755 ;
  assign y8927 = n20106 ;
  assign y8928 = ~n20107 ;
  assign y8929 = ~n20109 ;
  assign y8930 = ~1'b0 ;
  assign y8931 = ~1'b0 ;
  assign y8932 = n20110 ;
  assign y8933 = ~n20118 ;
  assign y8934 = ~1'b0 ;
  assign y8935 = ~n20121 ;
  assign y8936 = n20122 ;
  assign y8937 = n20125 ;
  assign y8938 = n20127 ;
  assign y8939 = n20128 ;
  assign y8940 = ~n20132 ;
  assign y8941 = ~1'b0 ;
  assign y8942 = ~1'b0 ;
  assign y8943 = n20135 ;
  assign y8944 = n20137 ;
  assign y8945 = ~n20139 ;
  assign y8946 = n20144 ;
  assign y8947 = ~n12281 ;
  assign y8948 = n20146 ;
  assign y8949 = ~1'b0 ;
  assign y8950 = ~n20147 ;
  assign y8951 = ~1'b0 ;
  assign y8952 = ~1'b0 ;
  assign y8953 = ~n20149 ;
  assign y8954 = ~n20151 ;
  assign y8955 = ~1'b0 ;
  assign y8956 = ~1'b0 ;
  assign y8957 = ~n20153 ;
  assign y8958 = ~n20158 ;
  assign y8959 = n20161 ;
  assign y8960 = n9809 ;
  assign y8961 = ~n20163 ;
  assign y8962 = n20166 ;
  assign y8963 = n20167 ;
  assign y8964 = ~n20175 ;
  assign y8965 = n20183 ;
  assign y8966 = ~1'b0 ;
  assign y8967 = ~n20185 ;
  assign y8968 = n20189 ;
  assign y8969 = ~1'b0 ;
  assign y8970 = ~n20193 ;
  assign y8971 = ~n20197 ;
  assign y8972 = n20198 ;
  assign y8973 = n20203 ;
  assign y8974 = n20204 ;
  assign y8975 = ~1'b0 ;
  assign y8976 = ~n20206 ;
  assign y8977 = n13481 ;
  assign y8978 = n20210 ;
  assign y8979 = n20213 ;
  assign y8980 = n20215 ;
  assign y8981 = ~n10313 ;
  assign y8982 = 1'b0 ;
  assign y8983 = ~1'b0 ;
  assign y8984 = ~n20216 ;
  assign y8985 = ~n20220 ;
  assign y8986 = ~1'b0 ;
  assign y8987 = n20222 ;
  assign y8988 = ~n20224 ;
  assign y8989 = ~n20225 ;
  assign y8990 = n20226 ;
  assign y8991 = n20228 ;
  assign y8992 = ~n20232 ;
  assign y8993 = n20233 ;
  assign y8994 = ~n20240 ;
  assign y8995 = ~1'b0 ;
  assign y8996 = n20247 ;
  assign y8997 = ~n20251 ;
  assign y8998 = ~1'b0 ;
  assign y8999 = ~n20252 ;
  assign y9000 = ~1'b0 ;
  assign y9001 = ~1'b0 ;
  assign y9002 = ~1'b0 ;
  assign y9003 = n20254 ;
  assign y9004 = n20256 ;
  assign y9005 = ~n20258 ;
  assign y9006 = ~n20260 ;
  assign y9007 = ~1'b0 ;
  assign y9008 = ~n20263 ;
  assign y9009 = n20269 ;
  assign y9010 = ~1'b0 ;
  assign y9011 = n20271 ;
  assign y9012 = n20272 ;
  assign y9013 = n20273 ;
  assign y9014 = n20274 ;
  assign y9015 = ~n20276 ;
  assign y9016 = ~1'b0 ;
  assign y9017 = n20279 ;
  assign y9018 = ~1'b0 ;
  assign y9019 = 1'b0 ;
  assign y9020 = ~n20282 ;
  assign y9021 = ~n20283 ;
  assign y9022 = n20291 ;
  assign y9023 = ~1'b0 ;
  assign y9024 = n20297 ;
  assign y9025 = ~n20298 ;
  assign y9026 = n20302 ;
  assign y9027 = ~n20305 ;
  assign y9028 = ~n20317 ;
  assign y9029 = 1'b0 ;
  assign y9030 = n20320 ;
  assign y9031 = 1'b0 ;
  assign y9032 = ~n473 ;
  assign y9033 = ~1'b0 ;
  assign y9034 = ~n20321 ;
  assign y9035 = ~n20324 ;
  assign y9036 = ~n20326 ;
  assign y9037 = ~1'b0 ;
  assign y9038 = n20328 ;
  assign y9039 = ~1'b0 ;
  assign y9040 = n8427 ;
  assign y9041 = ~n20329 ;
  assign y9042 = ~n20335 ;
  assign y9043 = ~1'b0 ;
  assign y9044 = ~n20337 ;
  assign y9045 = n20340 ;
  assign y9046 = ~1'b0 ;
  assign y9047 = ~n20341 ;
  assign y9048 = ~n1996 ;
  assign y9049 = ~n20345 ;
  assign y9050 = ~n20350 ;
  assign y9051 = ~1'b0 ;
  assign y9052 = n20353 ;
  assign y9053 = ~n20358 ;
  assign y9054 = ~n20360 ;
  assign y9055 = ~1'b0 ;
  assign y9056 = n20362 ;
  assign y9057 = ~n20366 ;
  assign y9058 = ~n20370 ;
  assign y9059 = ~1'b0 ;
  assign y9060 = ~1'b0 ;
  assign y9061 = ~n16297 ;
  assign y9062 = n10350 ;
  assign y9063 = n20372 ;
  assign y9064 = ~n7087 ;
  assign y9065 = ~1'b0 ;
  assign y9066 = 1'b0 ;
  assign y9067 = ~n20375 ;
  assign y9068 = ~n20381 ;
  assign y9069 = ~1'b0 ;
  assign y9070 = n20385 ;
  assign y9071 = ~n20386 ;
  assign y9072 = 1'b0 ;
  assign y9073 = ~n20403 ;
  assign y9074 = ~1'b0 ;
  assign y9075 = n20404 ;
  assign y9076 = n20405 ;
  assign y9077 = ~1'b0 ;
  assign y9078 = ~n705 ;
  assign y9079 = ~n20406 ;
  assign y9080 = n20409 ;
  assign y9081 = ~n20412 ;
  assign y9082 = ~n20416 ;
  assign y9083 = n20421 ;
  assign y9084 = n20422 ;
  assign y9085 = n4315 ;
  assign y9086 = ~n12701 ;
  assign y9087 = n20430 ;
  assign y9088 = n20433 ;
  assign y9089 = n20437 ;
  assign y9090 = ~n20439 ;
  assign y9091 = ~1'b0 ;
  assign y9092 = ~1'b0 ;
  assign y9093 = n20441 ;
  assign y9094 = n20448 ;
  assign y9095 = ~n20449 ;
  assign y9096 = ~1'b0 ;
  assign y9097 = n20450 ;
  assign y9098 = ~n20453 ;
  assign y9099 = ~n20455 ;
  assign y9100 = n17887 ;
  assign y9101 = ~n20456 ;
  assign y9102 = n20458 ;
  assign y9103 = n20462 ;
  assign y9104 = ~n20464 ;
  assign y9105 = n20466 ;
  assign y9106 = ~n20470 ;
  assign y9107 = ~n20473 ;
  assign y9108 = ~n20476 ;
  assign y9109 = n20477 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = n20490 ;
  assign y9112 = n4804 ;
  assign y9113 = n20501 ;
  assign y9114 = ~1'b0 ;
  assign y9115 = ~n20505 ;
  assign y9116 = n20507 ;
  assign y9117 = ~1'b0 ;
  assign y9118 = ~n20510 ;
  assign y9119 = ~n2695 ;
  assign y9120 = n20511 ;
  assign y9121 = ~1'b0 ;
  assign y9122 = n20513 ;
  assign y9123 = ~n20514 ;
  assign y9124 = ~n14798 ;
  assign y9125 = n20515 ;
  assign y9126 = 1'b0 ;
  assign y9127 = ~1'b0 ;
  assign y9128 = n20517 ;
  assign y9129 = ~1'b0 ;
  assign y9130 = ~n20518 ;
  assign y9131 = ~1'b0 ;
  assign y9132 = ~n20522 ;
  assign y9133 = n20528 ;
  assign y9134 = ~n20531 ;
  assign y9135 = n20533 ;
  assign y9136 = ~1'b0 ;
  assign y9137 = n20536 ;
  assign y9138 = ~n20537 ;
  assign y9139 = n20538 ;
  assign y9140 = ~1'b0 ;
  assign y9141 = n20546 ;
  assign y9142 = ~n1261 ;
  assign y9143 = n20548 ;
  assign y9144 = ~1'b0 ;
  assign y9145 = ~n8054 ;
  assign y9146 = ~1'b0 ;
  assign y9147 = n20550 ;
  assign y9148 = ~1'b0 ;
  assign y9149 = ~1'b0 ;
  assign y9150 = ~1'b0 ;
  assign y9151 = ~1'b0 ;
  assign y9152 = ~n20551 ;
  assign y9153 = n20554 ;
  assign y9154 = ~n20557 ;
  assign y9155 = n20561 ;
  assign y9156 = ~n20566 ;
  assign y9157 = ~n20571 ;
  assign y9158 = ~n20576 ;
  assign y9159 = ~n20578 ;
  assign y9160 = n20583 ;
  assign y9161 = ~1'b0 ;
  assign y9162 = ~1'b0 ;
  assign y9163 = ~1'b0 ;
  assign y9164 = ~1'b0 ;
  assign y9165 = ~1'b0 ;
  assign y9166 = ~n20585 ;
  assign y9167 = n20586 ;
  assign y9168 = ~n20590 ;
  assign y9169 = ~n20592 ;
  assign y9170 = n9621 ;
  assign y9171 = n20594 ;
  assign y9172 = ~1'b0 ;
  assign y9173 = ~1'b0 ;
  assign y9174 = ~n10745 ;
  assign y9175 = ~1'b0 ;
  assign y9176 = n20605 ;
  assign y9177 = ~n20609 ;
  assign y9178 = ~1'b0 ;
  assign y9179 = n18907 ;
  assign y9180 = ~1'b0 ;
  assign y9181 = ~1'b0 ;
  assign y9182 = ~n20611 ;
  assign y9183 = ~n20616 ;
  assign y9184 = ~n20623 ;
  assign y9185 = n20630 ;
  assign y9186 = ~n20631 ;
  assign y9187 = ~n20632 ;
  assign y9188 = n20635 ;
  assign y9189 = 1'b0 ;
  assign y9190 = ~1'b0 ;
  assign y9191 = n20644 ;
  assign y9192 = ~1'b0 ;
  assign y9193 = ~n20648 ;
  assign y9194 = n20649 ;
  assign y9195 = n20653 ;
  assign y9196 = ~n20654 ;
  assign y9197 = ~n20655 ;
  assign y9198 = ~n8143 ;
  assign y9199 = n10307 ;
  assign y9200 = n20656 ;
  assign y9201 = n20660 ;
  assign y9202 = ~1'b0 ;
  assign y9203 = ~1'b0 ;
  assign y9204 = ~n16251 ;
  assign y9205 = ~1'b0 ;
  assign y9206 = ~1'b0 ;
  assign y9207 = n20661 ;
  assign y9208 = ~n20667 ;
  assign y9209 = ~1'b0 ;
  assign y9210 = ~n20669 ;
  assign y9211 = ~n20674 ;
  assign y9212 = 1'b0 ;
  assign y9213 = n20677 ;
  assign y9214 = ~n20678 ;
  assign y9215 = n20681 ;
  assign y9216 = ~n18083 ;
  assign y9217 = ~n20682 ;
  assign y9218 = ~1'b0 ;
  assign y9219 = ~n20684 ;
  assign y9220 = n20686 ;
  assign y9221 = ~n20688 ;
  assign y9222 = n20689 ;
  assign y9223 = n20691 ;
  assign y9224 = n20693 ;
  assign y9225 = ~n20700 ;
  assign y9226 = n20702 ;
  assign y9227 = ~1'b0 ;
  assign y9228 = ~1'b0 ;
  assign y9229 = ~n20705 ;
  assign y9230 = n20711 ;
  assign y9231 = 1'b0 ;
  assign y9232 = ~1'b0 ;
  assign y9233 = ~n20712 ;
  assign y9234 = n20713 ;
  assign y9235 = ~n20715 ;
  assign y9236 = n20717 ;
  assign y9237 = ~n20719 ;
  assign y9238 = ~n20720 ;
  assign y9239 = ~n20722 ;
  assign y9240 = 1'b0 ;
  assign y9241 = ~n20731 ;
  assign y9242 = n20733 ;
  assign y9243 = n20736 ;
  assign y9244 = ~1'b0 ;
  assign y9245 = ~n20738 ;
  assign y9246 = n20742 ;
  assign y9247 = ~n20745 ;
  assign y9248 = n20747 ;
  assign y9249 = n20750 ;
  assign y9250 = ~n20751 ;
  assign y9251 = ~1'b0 ;
  assign y9252 = ~n20753 ;
  assign y9253 = ~n20754 ;
  assign y9254 = ~n20755 ;
  assign y9255 = n20756 ;
  assign y9256 = n20760 ;
  assign y9257 = ~1'b0 ;
  assign y9258 = ~1'b0 ;
  assign y9259 = ~1'b0 ;
  assign y9260 = n20762 ;
  assign y9261 = ~n12578 ;
  assign y9262 = ~n20763 ;
  assign y9263 = ~n20764 ;
  assign y9264 = ~n20765 ;
  assign y9265 = ~n20766 ;
  assign y9266 = ~1'b0 ;
  assign y9267 = ~n20767 ;
  assign y9268 = n20769 ;
  assign y9269 = 1'b0 ;
  assign y9270 = ~n20775 ;
  assign y9271 = ~n20783 ;
  assign y9272 = n20788 ;
  assign y9273 = n20792 ;
  assign y9274 = ~n20795 ;
  assign y9275 = ~n20799 ;
  assign y9276 = ~n20803 ;
  assign y9277 = ~n15324 ;
  assign y9278 = n20807 ;
  assign y9279 = n20809 ;
  assign y9280 = n20810 ;
  assign y9281 = ~1'b0 ;
  assign y9282 = ~n20813 ;
  assign y9283 = ~n20821 ;
  assign y9284 = n20822 ;
  assign y9285 = ~n7977 ;
  assign y9286 = ~n20824 ;
  assign y9287 = n20827 ;
  assign y9288 = n20832 ;
  assign y9289 = n20834 ;
  assign y9290 = ~1'b0 ;
  assign y9291 = n20836 ;
  assign y9292 = n4402 ;
  assign y9293 = n17738 ;
  assign y9294 = n20839 ;
  assign y9295 = ~n20840 ;
  assign y9296 = ~n20849 ;
  assign y9297 = ~1'b0 ;
  assign y9298 = 1'b0 ;
  assign y9299 = n20850 ;
  assign y9300 = ~1'b0 ;
  assign y9301 = n20852 ;
  assign y9302 = ~1'b0 ;
  assign y9303 = n20855 ;
  assign y9304 = ~1'b0 ;
  assign y9305 = ~n20863 ;
  assign y9306 = ~n20867 ;
  assign y9307 = n7031 ;
  assign y9308 = ~n20877 ;
  assign y9309 = ~1'b0 ;
  assign y9310 = ~1'b0 ;
  assign y9311 = n20878 ;
  assign y9312 = n20879 ;
  assign y9313 = n20882 ;
  assign y9314 = ~n20884 ;
  assign y9315 = ~1'b0 ;
  assign y9316 = ~1'b0 ;
  assign y9317 = n20886 ;
  assign y9318 = n20887 ;
  assign y9319 = ~1'b0 ;
  assign y9320 = n20888 ;
  assign y9321 = ~n20892 ;
  assign y9322 = ~n20893 ;
  assign y9323 = ~n9262 ;
  assign y9324 = n20895 ;
  assign y9325 = ~n20896 ;
  assign y9326 = ~n20897 ;
  assign y9327 = ~n20898 ;
  assign y9328 = n20899 ;
  assign y9329 = n20904 ;
  assign y9330 = ~n20905 ;
  assign y9331 = ~n20906 ;
  assign y9332 = ~n20909 ;
  assign y9333 = n20913 ;
  assign y9334 = ~n20915 ;
  assign y9335 = 1'b0 ;
  assign y9336 = n20919 ;
  assign y9337 = ~1'b0 ;
  assign y9338 = n20925 ;
  assign y9339 = n20929 ;
  assign y9340 = ~1'b0 ;
  assign y9341 = ~n20933 ;
  assign y9342 = ~1'b0 ;
  assign y9343 = n8175 ;
  assign y9344 = ~n20938 ;
  assign y9345 = ~1'b0 ;
  assign y9346 = n20942 ;
  assign y9347 = n20951 ;
  assign y9348 = n20953 ;
  assign y9349 = ~n20954 ;
  assign y9350 = n20955 ;
  assign y9351 = n20956 ;
  assign y9352 = ~n20957 ;
  assign y9353 = ~n20961 ;
  assign y9354 = ~n20965 ;
  assign y9355 = ~1'b0 ;
  assign y9356 = n20967 ;
  assign y9357 = n20968 ;
  assign y9358 = n20969 ;
  assign y9359 = ~n20971 ;
  assign y9360 = ~n20978 ;
  assign y9361 = n20983 ;
  assign y9362 = ~1'b0 ;
  assign y9363 = n20984 ;
  assign y9364 = ~n20985 ;
  assign y9365 = ~n20987 ;
  assign y9366 = n20988 ;
  assign y9367 = ~1'b0 ;
  assign y9368 = n10862 ;
  assign y9369 = ~1'b0 ;
  assign y9370 = n20989 ;
  assign y9371 = n20990 ;
  assign y9372 = n20993 ;
  assign y9373 = ~n20997 ;
  assign y9374 = ~n20998 ;
  assign y9375 = n21013 ;
  assign y9376 = n21015 ;
  assign y9377 = ~n21016 ;
  assign y9378 = ~1'b0 ;
  assign y9379 = ~1'b0 ;
  assign y9380 = ~n21022 ;
  assign y9381 = ~n21025 ;
  assign y9382 = n21030 ;
  assign y9383 = ~n21031 ;
  assign y9384 = n21033 ;
  assign y9385 = ~1'b0 ;
  assign y9386 = 1'b0 ;
  assign y9387 = ~1'b0 ;
  assign y9388 = n21040 ;
  assign y9389 = ~n21052 ;
  assign y9390 = n21056 ;
  assign y9391 = ~n21058 ;
  assign y9392 = ~1'b0 ;
  assign y9393 = n21061 ;
  assign y9394 = n21065 ;
  assign y9395 = ~n21066 ;
  assign y9396 = ~1'b0 ;
  assign y9397 = ~n21070 ;
  assign y9398 = n21072 ;
  assign y9399 = ~1'b0 ;
  assign y9400 = n21073 ;
  assign y9401 = n21074 ;
  assign y9402 = ~n21076 ;
  assign y9403 = ~n21077 ;
  assign y9404 = ~n21079 ;
  assign y9405 = n21084 ;
  assign y9406 = n21087 ;
  assign y9407 = n21090 ;
  assign y9408 = ~1'b0 ;
  assign y9409 = ~n21092 ;
  assign y9410 = n21113 ;
  assign y9411 = n21117 ;
  assign y9412 = ~1'b0 ;
  assign y9413 = ~n21120 ;
  assign y9414 = ~1'b0 ;
  assign y9415 = n21124 ;
  assign y9416 = ~n21128 ;
  assign y9417 = n21131 ;
  assign y9418 = ~1'b0 ;
  assign y9419 = ~n21135 ;
  assign y9420 = ~n21136 ;
  assign y9421 = ~1'b0 ;
  assign y9422 = ~n21142 ;
  assign y9423 = ~1'b0 ;
  assign y9424 = ~n21145 ;
  assign y9425 = n21146 ;
  assign y9426 = ~1'b0 ;
  assign y9427 = ~n21147 ;
  assign y9428 = n21149 ;
  assign y9429 = ~n21153 ;
  assign y9430 = ~1'b0 ;
  assign y9431 = n21156 ;
  assign y9432 = ~n21158 ;
  assign y9433 = ~n21161 ;
  assign y9434 = ~n21162 ;
  assign y9435 = ~1'b0 ;
  assign y9436 = ~n21166 ;
  assign y9437 = ~n21167 ;
  assign y9438 = ~n21174 ;
  assign y9439 = ~n21175 ;
  assign y9440 = ~1'b0 ;
  assign y9441 = ~n21178 ;
  assign y9442 = ~n21180 ;
  assign y9443 = ~n21181 ;
  assign y9444 = ~1'b0 ;
  assign y9445 = ~n21182 ;
  assign y9446 = ~n21191 ;
  assign y9447 = ~1'b0 ;
  assign y9448 = ~n21195 ;
  assign y9449 = ~n21196 ;
  assign y9450 = ~n21202 ;
  assign y9451 = n21204 ;
  assign y9452 = n21205 ;
  assign y9453 = n21208 ;
  assign y9454 = ~n21214 ;
  assign y9455 = n21217 ;
  assign y9456 = ~n21221 ;
  assign y9457 = ~n21222 ;
  assign y9458 = n15173 ;
  assign y9459 = n21223 ;
  assign y9460 = ~n21224 ;
  assign y9461 = ~n21232 ;
  assign y9462 = ~1'b0 ;
  assign y9463 = n21233 ;
  assign y9464 = ~n21234 ;
  assign y9465 = n21236 ;
  assign y9466 = n21240 ;
  assign y9467 = n21245 ;
  assign y9468 = n21246 ;
  assign y9469 = ~n21250 ;
  assign y9470 = n21261 ;
  assign y9471 = ~n21267 ;
  assign y9472 = n21269 ;
  assign y9473 = ~n21287 ;
  assign y9474 = ~n2787 ;
  assign y9475 = ~n21289 ;
  assign y9476 = ~n21292 ;
  assign y9477 = ~n21295 ;
  assign y9478 = ~n21296 ;
  assign y9479 = ~n21297 ;
  assign y9480 = ~n21302 ;
  assign y9481 = ~n21305 ;
  assign y9482 = ~n21307 ;
  assign y9483 = ~n21318 ;
  assign y9484 = ~1'b0 ;
  assign y9485 = ~n21319 ;
  assign y9486 = ~1'b0 ;
  assign y9487 = ~n2082 ;
  assign y9488 = ~1'b0 ;
  assign y9489 = ~n21329 ;
  assign y9490 = n21340 ;
  assign y9491 = ~1'b0 ;
  assign y9492 = ~1'b0 ;
  assign y9493 = ~n21342 ;
  assign y9494 = ~n21343 ;
  assign y9495 = ~n21344 ;
  assign y9496 = ~n21350 ;
  assign y9497 = ~1'b0 ;
  assign y9498 = ~1'b0 ;
  assign y9499 = ~n21353 ;
  assign y9500 = ~1'b0 ;
  assign y9501 = n21354 ;
  assign y9502 = n21357 ;
  assign y9503 = ~1'b0 ;
  assign y9504 = ~1'b0 ;
  assign y9505 = ~1'b0 ;
  assign y9506 = ~1'b0 ;
  assign y9507 = n21358 ;
  assign y9508 = ~n21360 ;
  assign y9509 = n21370 ;
  assign y9510 = n21375 ;
  assign y9511 = n21377 ;
  assign y9512 = ~n21380 ;
  assign y9513 = n4545 ;
  assign y9514 = n21381 ;
  assign y9515 = ~n21382 ;
  assign y9516 = ~n21383 ;
  assign y9517 = n21385 ;
  assign y9518 = ~1'b0 ;
  assign y9519 = ~1'b0 ;
  assign y9520 = ~n21390 ;
  assign y9521 = n21392 ;
  assign y9522 = ~n21396 ;
  assign y9523 = ~n21397 ;
  assign y9524 = ~n21400 ;
  assign y9525 = n21405 ;
  assign y9526 = ~1'b0 ;
  assign y9527 = ~1'b0 ;
  assign y9528 = n21407 ;
  assign y9529 = ~n21408 ;
  assign y9530 = ~n21412 ;
  assign y9531 = n21413 ;
  assign y9532 = ~n21416 ;
  assign y9533 = ~1'b0 ;
  assign y9534 = ~1'b0 ;
  assign y9535 = ~1'b0 ;
  assign y9536 = ~n21417 ;
  assign y9537 = ~1'b0 ;
  assign y9538 = n21421 ;
  assign y9539 = n21423 ;
  assign y9540 = ~1'b0 ;
  assign y9541 = n21427 ;
  assign y9542 = ~n21432 ;
  assign y9543 = n21439 ;
  assign y9544 = n21446 ;
  assign y9545 = ~1'b0 ;
  assign y9546 = ~n11666 ;
  assign y9547 = ~n21447 ;
  assign y9548 = ~n21448 ;
  assign y9549 = n21459 ;
  assign y9550 = ~1'b0 ;
  assign y9551 = ~1'b0 ;
  assign y9552 = n949 ;
  assign y9553 = 1'b0 ;
  assign y9554 = 1'b0 ;
  assign y9555 = ~1'b0 ;
  assign y9556 = n21462 ;
  assign y9557 = ~n21465 ;
  assign y9558 = n21467 ;
  assign y9559 = ~n21478 ;
  assign y9560 = n21480 ;
  assign y9561 = n21483 ;
  assign y9562 = ~n21489 ;
  assign y9563 = n21490 ;
  assign y9564 = 1'b0 ;
  assign y9565 = n13866 ;
  assign y9566 = n21497 ;
  assign y9567 = ~n21501 ;
  assign y9568 = ~1'b0 ;
  assign y9569 = ~1'b0 ;
  assign y9570 = ~1'b0 ;
  assign y9571 = ~n21503 ;
  assign y9572 = ~1'b0 ;
  assign y9573 = n21514 ;
  assign y9574 = n21517 ;
  assign y9575 = ~n1531 ;
  assign y9576 = ~n21521 ;
  assign y9577 = ~n21522 ;
  assign y9578 = n21525 ;
  assign y9579 = ~n21526 ;
  assign y9580 = ~n21529 ;
  assign y9581 = ~n11832 ;
  assign y9582 = ~n21530 ;
  assign y9583 = n21535 ;
  assign y9584 = ~n21539 ;
  assign y9585 = n21540 ;
  assign y9586 = n21541 ;
  assign y9587 = n21543 ;
  assign y9588 = n21544 ;
  assign y9589 = ~n21546 ;
  assign y9590 = ~n21557 ;
  assign y9591 = n21561 ;
  assign y9592 = ~n21564 ;
  assign y9593 = ~n21565 ;
  assign y9594 = ~n6713 ;
  assign y9595 = ~n21573 ;
  assign y9596 = n21574 ;
  assign y9597 = ~1'b0 ;
  assign y9598 = ~n21575 ;
  assign y9599 = n21576 ;
  assign y9600 = ~n21577 ;
  assign y9601 = n15680 ;
  assign y9602 = ~1'b0 ;
  assign y9603 = ~n21578 ;
  assign y9604 = n21579 ;
  assign y9605 = ~n21583 ;
  assign y9606 = ~1'b0 ;
  assign y9607 = ~n21584 ;
  assign y9608 = ~n21586 ;
  assign y9609 = ~n21589 ;
  assign y9610 = n21591 ;
  assign y9611 = ~n21593 ;
  assign y9612 = n21594 ;
  assign y9613 = n21595 ;
  assign y9614 = n21601 ;
  assign y9615 = ~n21605 ;
  assign y9616 = n21611 ;
  assign y9617 = n21612 ;
  assign y9618 = n21616 ;
  assign y9619 = n21617 ;
  assign y9620 = ~n21620 ;
  assign y9621 = n21625 ;
  assign y9622 = ~n21627 ;
  assign y9623 = ~n21628 ;
  assign y9624 = ~n21630 ;
  assign y9625 = n9014 ;
  assign y9626 = n21633 ;
  assign y9627 = ~n21636 ;
  assign y9628 = ~n21643 ;
  assign y9629 = n21646 ;
  assign y9630 = ~n21647 ;
  assign y9631 = n21655 ;
  assign y9632 = ~n21658 ;
  assign y9633 = ~n21660 ;
  assign y9634 = n21662 ;
  assign y9635 = n21663 ;
  assign y9636 = ~1'b0 ;
  assign y9637 = n21665 ;
  assign y9638 = ~n21669 ;
  assign y9639 = ~1'b0 ;
  assign y9640 = n21670 ;
  assign y9641 = ~1'b0 ;
  assign y9642 = ~1'b0 ;
  assign y9643 = ~n21672 ;
  assign y9644 = ~n21674 ;
  assign y9645 = n10212 ;
  assign y9646 = ~n21677 ;
  assign y9647 = ~1'b0 ;
  assign y9648 = n21681 ;
  assign y9649 = ~1'b0 ;
  assign y9650 = ~1'b0 ;
  assign y9651 = ~n21685 ;
  assign y9652 = ~n21690 ;
  assign y9653 = ~1'b0 ;
  assign y9654 = n21691 ;
  assign y9655 = ~n21695 ;
  assign y9656 = n21696 ;
  assign y9657 = ~n21697 ;
  assign y9658 = ~n21699 ;
  assign y9659 = ~n21700 ;
  assign y9660 = ~n21710 ;
  assign y9661 = ~1'b0 ;
  assign y9662 = ~n21712 ;
  assign y9663 = ~n21714 ;
  assign y9664 = ~n19973 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = ~n21718 ;
  assign y9667 = ~1'b0 ;
  assign y9668 = ~1'b0 ;
  assign y9669 = ~1'b0 ;
  assign y9670 = ~1'b0 ;
  assign y9671 = n21721 ;
  assign y9672 = ~n21725 ;
  assign y9673 = n21728 ;
  assign y9674 = ~1'b0 ;
  assign y9675 = n21737 ;
  assign y9676 = ~n16455 ;
  assign y9677 = n21738 ;
  assign y9678 = n21739 ;
  assign y9679 = ~1'b0 ;
  assign y9680 = ~1'b0 ;
  assign y9681 = ~n21740 ;
  assign y9682 = ~1'b0 ;
  assign y9683 = n21742 ;
  assign y9684 = ~n21743 ;
  assign y9685 = ~1'b0 ;
  assign y9686 = ~1'b0 ;
  assign y9687 = n21744 ;
  assign y9688 = ~n21747 ;
  assign y9689 = 1'b0 ;
  assign y9690 = ~n21748 ;
  assign y9691 = ~1'b0 ;
  assign y9692 = ~n21753 ;
  assign y9693 = n7061 ;
  assign y9694 = n15485 ;
  assign y9695 = ~n21754 ;
  assign y9696 = ~1'b0 ;
  assign y9697 = n21757 ;
  assign y9698 = ~n21760 ;
  assign y9699 = 1'b0 ;
  assign y9700 = n21761 ;
  assign y9701 = ~n21763 ;
  assign y9702 = 1'b0 ;
  assign y9703 = 1'b0 ;
  assign y9704 = n21764 ;
  assign y9705 = n21766 ;
  assign y9706 = ~1'b0 ;
  assign y9707 = n21768 ;
  assign y9708 = n21771 ;
  assign y9709 = ~n21773 ;
  assign y9710 = ~1'b0 ;
  assign y9711 = ~1'b0 ;
  assign y9712 = n21780 ;
  assign y9713 = ~n4447 ;
  assign y9714 = ~n21782 ;
  assign y9715 = ~n21785 ;
  assign y9716 = ~n21788 ;
  assign y9717 = ~1'b0 ;
  assign y9718 = ~n21790 ;
  assign y9719 = n21795 ;
  assign y9720 = ~1'b0 ;
  assign y9721 = ~1'b0 ;
  assign y9722 = ~n21797 ;
  assign y9723 = n21800 ;
  assign y9724 = n21802 ;
  assign y9725 = ~n21803 ;
  assign y9726 = ~n21804 ;
  assign y9727 = n21811 ;
  assign y9728 = n21814 ;
  assign y9729 = n21816 ;
  assign y9730 = ~1'b0 ;
  assign y9731 = ~1'b0 ;
  assign y9732 = ~1'b0 ;
  assign y9733 = n21825 ;
  assign y9734 = n21826 ;
  assign y9735 = ~n21828 ;
  assign y9736 = ~n21829 ;
  assign y9737 = ~n21835 ;
  assign y9738 = n21836 ;
  assign y9739 = ~n21842 ;
  assign y9740 = ~n21843 ;
  assign y9741 = n21844 ;
  assign y9742 = n21847 ;
  assign y9743 = n21850 ;
  assign y9744 = ~1'b0 ;
  assign y9745 = ~1'b0 ;
  assign y9746 = n21851 ;
  assign y9747 = n21854 ;
  assign y9748 = ~1'b0 ;
  assign y9749 = n12504 ;
  assign y9750 = ~n21856 ;
  assign y9751 = n21858 ;
  assign y9752 = n21864 ;
  assign y9753 = n21869 ;
  assign y9754 = ~n21872 ;
  assign y9755 = n21873 ;
  assign y9756 = ~1'b0 ;
  assign y9757 = n21876 ;
  assign y9758 = ~n4468 ;
  assign y9759 = ~1'b0 ;
  assign y9760 = n21877 ;
  assign y9761 = ~1'b0 ;
  assign y9762 = ~1'b0 ;
  assign y9763 = n21878 ;
  assign y9764 = n6415 ;
  assign y9765 = n21881 ;
  assign y9766 = ~1'b0 ;
  assign y9767 = ~1'b0 ;
  assign y9768 = n21884 ;
  assign y9769 = n21887 ;
  assign y9770 = ~n21889 ;
  assign y9771 = ~1'b0 ;
  assign y9772 = ~1'b0 ;
  assign y9773 = n21890 ;
  assign y9774 = n21892 ;
  assign y9775 = n21893 ;
  assign y9776 = n21899 ;
  assign y9777 = ~n21900 ;
  assign y9778 = n21908 ;
  assign y9779 = ~n21910 ;
  assign y9780 = ~1'b0 ;
  assign y9781 = n21911 ;
  assign y9782 = n21912 ;
  assign y9783 = ~n21915 ;
  assign y9784 = n21916 ;
  assign y9785 = ~1'b0 ;
  assign y9786 = ~1'b0 ;
  assign y9787 = ~1'b0 ;
  assign y9788 = n21919 ;
  assign y9789 = ~n21923 ;
  assign y9790 = ~1'b0 ;
  assign y9791 = n21925 ;
  assign y9792 = n21926 ;
  assign y9793 = ~n21931 ;
  assign y9794 = n21933 ;
  assign y9795 = n21938 ;
  assign y9796 = n21951 ;
  assign y9797 = ~1'b0 ;
  assign y9798 = ~1'b0 ;
  assign y9799 = ~1'b0 ;
  assign y9800 = n21952 ;
  assign y9801 = n21955 ;
  assign y9802 = n21957 ;
  assign y9803 = ~1'b0 ;
  assign y9804 = ~n21958 ;
  assign y9805 = ~n21960 ;
  assign y9806 = ~1'b0 ;
  assign y9807 = ~1'b0 ;
  assign y9808 = ~1'b0 ;
  assign y9809 = n21963 ;
  assign y9810 = ~n21969 ;
  assign y9811 = n21973 ;
  assign y9812 = ~1'b0 ;
  assign y9813 = n21974 ;
  assign y9814 = ~1'b0 ;
  assign y9815 = ~1'b0 ;
  assign y9816 = n21977 ;
  assign y9817 = n21978 ;
  assign y9818 = n21980 ;
  assign y9819 = n21981 ;
  assign y9820 = ~1'b0 ;
  assign y9821 = n21983 ;
  assign y9822 = ~n21986 ;
  assign y9823 = n21987 ;
  assign y9824 = n7280 ;
  assign y9825 = n21988 ;
  assign y9826 = n21989 ;
  assign y9827 = ~1'b0 ;
  assign y9828 = n21994 ;
  assign y9829 = n21998 ;
  assign y9830 = ~n22001 ;
  assign y9831 = ~1'b0 ;
  assign y9832 = ~1'b0 ;
  assign y9833 = ~1'b0 ;
  assign y9834 = ~1'b0 ;
  assign y9835 = n22007 ;
  assign y9836 = n22008 ;
  assign y9837 = ~1'b0 ;
  assign y9838 = ~1'b0 ;
  assign y9839 = ~n22014 ;
  assign y9840 = n22017 ;
  assign y9841 = n22019 ;
  assign y9842 = n22021 ;
  assign y9843 = 1'b0 ;
  assign y9844 = 1'b0 ;
  assign y9845 = ~1'b0 ;
  assign y9846 = ~n22022 ;
  assign y9847 = ~n22023 ;
  assign y9848 = ~n11971 ;
  assign y9849 = n22025 ;
  assign y9850 = ~1'b0 ;
  assign y9851 = ~n22026 ;
  assign y9852 = n22027 ;
  assign y9853 = ~n22029 ;
  assign y9854 = ~n22033 ;
  assign y9855 = ~n22037 ;
  assign y9856 = n22039 ;
  assign y9857 = ~n22040 ;
  assign y9858 = ~n22042 ;
  assign y9859 = ~n22044 ;
  assign y9860 = 1'b0 ;
  assign y9861 = n22047 ;
  assign y9862 = ~n22048 ;
  assign y9863 = n16661 ;
  assign y9864 = ~1'b0 ;
  assign y9865 = ~n22049 ;
  assign y9866 = ~1'b0 ;
  assign y9867 = n22054 ;
  assign y9868 = n22057 ;
  assign y9869 = ~n22059 ;
  assign y9870 = ~n22062 ;
  assign y9871 = ~n22064 ;
  assign y9872 = ~n13067 ;
  assign y9873 = ~1'b0 ;
  assign y9874 = ~n22066 ;
  assign y9875 = n22068 ;
  assign y9876 = n22070 ;
  assign y9877 = ~1'b0 ;
  assign y9878 = n22073 ;
  assign y9879 = ~1'b0 ;
  assign y9880 = ~n22074 ;
  assign y9881 = n22075 ;
  assign y9882 = ~n22083 ;
  assign y9883 = n8829 ;
  assign y9884 = n22092 ;
  assign y9885 = n22095 ;
  assign y9886 = ~n22100 ;
  assign y9887 = n22106 ;
  assign y9888 = ~1'b0 ;
  assign y9889 = n22112 ;
  assign y9890 = n14684 ;
  assign y9891 = n22113 ;
  assign y9892 = ~1'b0 ;
  assign y9893 = ~1'b0 ;
  assign y9894 = n22114 ;
  assign y9895 = n22118 ;
  assign y9896 = ~1'b0 ;
  assign y9897 = n22121 ;
  assign y9898 = ~n22123 ;
  assign y9899 = n22125 ;
  assign y9900 = ~n22129 ;
  assign y9901 = ~1'b0 ;
  assign y9902 = ~n22132 ;
  assign y9903 = ~n22137 ;
  assign y9904 = ~n22141 ;
  assign y9905 = ~1'b0 ;
  assign y9906 = ~1'b0 ;
  assign y9907 = n16246 ;
  assign y9908 = ~n22142 ;
  assign y9909 = ~n22143 ;
  assign y9910 = ~n22144 ;
  assign y9911 = ~n22145 ;
  assign y9912 = ~n22146 ;
  assign y9913 = ~n22147 ;
  assign y9914 = ~n22150 ;
  assign y9915 = ~n22151 ;
  assign y9916 = ~n22153 ;
  assign y9917 = ~1'b0 ;
  assign y9918 = ~n22160 ;
  assign y9919 = 1'b0 ;
  assign y9920 = ~1'b0 ;
  assign y9921 = n22163 ;
  assign y9922 = n22164 ;
  assign y9923 = n22165 ;
  assign y9924 = n22168 ;
  assign y9925 = ~n22174 ;
  assign y9926 = n8427 ;
  assign y9927 = ~1'b0 ;
  assign y9928 = ~n22175 ;
  assign y9929 = ~n22178 ;
  assign y9930 = ~n22182 ;
  assign y9931 = ~n22187 ;
  assign y9932 = ~1'b0 ;
  assign y9933 = ~n8622 ;
  assign y9934 = ~n22189 ;
  assign y9935 = ~1'b0 ;
  assign y9936 = n22198 ;
  assign y9937 = ~1'b0 ;
  assign y9938 = n22209 ;
  assign y9939 = n22215 ;
  assign y9940 = ~1'b0 ;
  assign y9941 = n22216 ;
  assign y9942 = ~1'b0 ;
  assign y9943 = ~n12909 ;
  assign y9944 = ~n13141 ;
  assign y9945 = n22222 ;
  assign y9946 = n22225 ;
  assign y9947 = ~1'b0 ;
  assign y9948 = ~n22232 ;
  assign y9949 = n22237 ;
  assign y9950 = ~1'b0 ;
  assign y9951 = n22240 ;
  assign y9952 = ~1'b0 ;
  assign y9953 = ~1'b0 ;
  assign y9954 = n22241 ;
  assign y9955 = n22243 ;
  assign y9956 = n22252 ;
  assign y9957 = ~n22255 ;
  assign y9958 = ~1'b0 ;
  assign y9959 = ~n22260 ;
  assign y9960 = n22265 ;
  assign y9961 = n22269 ;
  assign y9962 = n22270 ;
  assign y9963 = n22271 ;
  assign y9964 = ~n22272 ;
  assign y9965 = ~1'b0 ;
  assign y9966 = n22274 ;
  assign y9967 = n22275 ;
  assign y9968 = ~n22276 ;
  assign y9969 = n22278 ;
  assign y9970 = ~n22286 ;
  assign y9971 = n22287 ;
  assign y9972 = ~n22291 ;
  assign y9973 = ~n22293 ;
  assign y9974 = ~n22296 ;
  assign y9975 = n22303 ;
  assign y9976 = n22304 ;
  assign y9977 = ~1'b0 ;
  assign y9978 = ~n22310 ;
  assign y9979 = ~n22312 ;
  assign y9980 = ~1'b0 ;
  assign y9981 = n22318 ;
  assign y9982 = ~1'b0 ;
  assign y9983 = n10741 ;
  assign y9984 = ~n22323 ;
  assign y9985 = n22325 ;
  assign y9986 = n22330 ;
  assign y9987 = ~n22333 ;
  assign y9988 = ~1'b0 ;
  assign y9989 = ~1'b0 ;
  assign y9990 = ~n22342 ;
  assign y9991 = ~1'b0 ;
  assign y9992 = ~1'b0 ;
  assign y9993 = n22343 ;
  assign y9994 = ~n18911 ;
  assign y9995 = ~1'b0 ;
  assign y9996 = n22345 ;
  assign y9997 = ~n22346 ;
  assign y9998 = ~1'b0 ;
  assign y9999 = ~n22348 ;
  assign y10000 = ~n22352 ;
  assign y10001 = n22355 ;
  assign y10002 = n22365 ;
  assign y10003 = n22368 ;
  assign y10004 = ~1'b0 ;
  assign y10005 = ~n22373 ;
  assign y10006 = n22376 ;
  assign y10007 = ~n40 ;
  assign y10008 = ~1'b0 ;
  assign y10009 = ~n22379 ;
  assign y10010 = n22383 ;
  assign y10011 = ~1'b0 ;
  assign y10012 = n68 ;
  assign y10013 = n22386 ;
  assign y10014 = ~n22387 ;
  assign y10015 = ~n22388 ;
  assign y10016 = n22390 ;
  assign y10017 = ~n22392 ;
  assign y10018 = n22394 ;
  assign y10019 = n22395 ;
  assign y10020 = n22396 ;
  assign y10021 = n8684 ;
  assign y10022 = n22399 ;
  assign y10023 = ~1'b0 ;
  assign y10024 = n22400 ;
  assign y10025 = n22405 ;
  assign y10026 = ~1'b0 ;
  assign y10027 = ~n22407 ;
  assign y10028 = ~1'b0 ;
  assign y10029 = ~1'b0 ;
  assign y10030 = n22408 ;
  assign y10031 = n22417 ;
  assign y10032 = ~n22428 ;
  assign y10033 = n22429 ;
  assign y10034 = n22436 ;
  assign y10035 = ~n22438 ;
  assign y10036 = ~1'b0 ;
  assign y10037 = n7443 ;
  assign y10038 = n22440 ;
  assign y10039 = n22444 ;
  assign y10040 = ~1'b0 ;
  assign y10041 = n22445 ;
  assign y10042 = n22446 ;
  assign y10043 = ~1'b0 ;
  assign y10044 = n22448 ;
  assign y10045 = ~1'b0 ;
  assign y10046 = n22451 ;
  assign y10047 = ~n22452 ;
  assign y10048 = ~n22462 ;
  assign y10049 = ~1'b0 ;
  assign y10050 = ~1'b0 ;
  assign y10051 = ~n22465 ;
  assign y10052 = ~n22472 ;
  assign y10053 = n22475 ;
  assign y10054 = n22480 ;
  assign y10055 = n22481 ;
  assign y10056 = ~1'b0 ;
  assign y10057 = n22482 ;
  assign y10058 = n151 ;
  assign y10059 = ~n22485 ;
  assign y10060 = n22487 ;
  assign y10061 = n22490 ;
  assign y10062 = ~1'b0 ;
  assign y10063 = ~n1370 ;
  assign y10064 = n22499 ;
  assign y10065 = ~1'b0 ;
  assign y10066 = n22501 ;
  assign y10067 = ~n22502 ;
  assign y10068 = n7867 ;
  assign y10069 = ~n22511 ;
  assign y10070 = ~1'b0 ;
  assign y10071 = ~1'b0 ;
  assign y10072 = ~n22512 ;
  assign y10073 = ~1'b0 ;
  assign y10074 = ~n22514 ;
  assign y10075 = n22523 ;
  assign y10076 = ~n15912 ;
  assign y10077 = n22524 ;
  assign y10078 = ~n22526 ;
  assign y10079 = ~1'b0 ;
  assign y10080 = ~n22527 ;
  assign y10081 = n1036 ;
  assign y10082 = ~n22538 ;
  assign y10083 = ~1'b0 ;
  assign y10084 = ~n22540 ;
  assign y10085 = ~n22546 ;
  assign y10086 = ~1'b0 ;
  assign y10087 = ~1'b0 ;
  assign y10088 = ~1'b0 ;
  assign y10089 = ~1'b0 ;
  assign y10090 = n22551 ;
  assign y10091 = ~n22553 ;
  assign y10092 = n22554 ;
  assign y10093 = ~n22557 ;
  assign y10094 = ~n22561 ;
  assign y10095 = n22568 ;
  assign y10096 = ~1'b0 ;
  assign y10097 = ~n22571 ;
  assign y10098 = ~n3059 ;
  assign y10099 = n22577 ;
  assign y10100 = ~n22578 ;
  assign y10101 = ~1'b0 ;
  assign y10102 = ~1'b0 ;
  assign y10103 = ~n16730 ;
  assign y10104 = n22580 ;
  assign y10105 = ~n22583 ;
  assign y10106 = ~n22585 ;
  assign y10107 = n22586 ;
  assign y10108 = ~n9633 ;
  assign y10109 = n22588 ;
  assign y10110 = ~1'b0 ;
  assign y10111 = n22589 ;
  assign y10112 = ~n22590 ;
  assign y10113 = ~n22592 ;
  assign y10114 = ~n22594 ;
  assign y10115 = n22598 ;
  assign y10116 = ~n22602 ;
  assign y10117 = n22610 ;
  assign y10118 = n22611 ;
  assign y10119 = ~n22612 ;
  assign y10120 = ~n22615 ;
  assign y10121 = ~n22617 ;
  assign y10122 = ~1'b0 ;
  assign y10123 = ~1'b0 ;
  assign y10124 = ~n22620 ;
  assign y10125 = ~n22623 ;
  assign y10126 = ~n7468 ;
  assign y10127 = n22627 ;
  assign y10128 = ~1'b0 ;
  assign y10129 = ~n22628 ;
  assign y10130 = ~1'b0 ;
  assign y10131 = ~1'b0 ;
  assign y10132 = ~1'b0 ;
  assign y10133 = n22633 ;
  assign y10134 = ~n22634 ;
  assign y10135 = n22636 ;
  assign y10136 = n22638 ;
  assign y10137 = n22640 ;
  assign y10138 = n22641 ;
  assign y10139 = ~n22642 ;
  assign y10140 = n22644 ;
  assign y10141 = ~n22649 ;
  assign y10142 = ~n22652 ;
  assign y10143 = n22654 ;
  assign y10144 = n22656 ;
  assign y10145 = ~1'b0 ;
  assign y10146 = ~n22660 ;
  assign y10147 = n4860 ;
  assign y10148 = n22661 ;
  assign y10149 = n22666 ;
  assign y10150 = ~1'b0 ;
  assign y10151 = ~n22668 ;
  assign y10152 = ~n22669 ;
  assign y10153 = ~n22676 ;
  assign y10154 = ~n22681 ;
  assign y10155 = ~1'b0 ;
  assign y10156 = ~n22683 ;
  assign y10157 = n22687 ;
  assign y10158 = ~1'b0 ;
  assign y10159 = ~n11955 ;
  assign y10160 = ~n22688 ;
  assign y10161 = n22692 ;
  assign y10162 = ~n2225 ;
  assign y10163 = n22694 ;
  assign y10164 = ~n22699 ;
  assign y10165 = n5520 ;
  assign y10166 = n22702 ;
  assign y10167 = ~n22703 ;
  assign y10168 = n22704 ;
  assign y10169 = ~n22711 ;
  assign y10170 = ~n22714 ;
  assign y10171 = ~n22717 ;
  assign y10172 = ~1'b0 ;
  assign y10173 = ~1'b0 ;
  assign y10174 = ~1'b0 ;
  assign y10175 = ~n22721 ;
  assign y10176 = ~1'b0 ;
  assign y10177 = ~n22724 ;
  assign y10178 = n22728 ;
  assign y10179 = ~1'b0 ;
  assign y10180 = ~n22731 ;
  assign y10181 = n22738 ;
  assign y10182 = n22739 ;
  assign y10183 = n22741 ;
  assign y10184 = ~1'b0 ;
  assign y10185 = ~n22743 ;
  assign y10186 = ~n22753 ;
  assign y10187 = ~1'b0 ;
  assign y10188 = ~n22759 ;
  assign y10189 = ~1'b0 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = ~n22763 ;
  assign y10192 = n22765 ;
  assign y10193 = ~n22766 ;
  assign y10194 = n22770 ;
  assign y10195 = ~n22772 ;
  assign y10196 = ~n22773 ;
  assign y10197 = ~1'b0 ;
  assign y10198 = n11161 ;
  assign y10199 = n22774 ;
  assign y10200 = ~1'b0 ;
  assign y10201 = ~n7150 ;
  assign y10202 = ~n22780 ;
  assign y10203 = ~n22781 ;
  assign y10204 = n22785 ;
  assign y10205 = n22790 ;
  assign y10206 = n22791 ;
  assign y10207 = n22792 ;
  assign y10208 = ~1'b0 ;
  assign y10209 = ~n9919 ;
  assign y10210 = n22794 ;
  assign y10211 = ~n22798 ;
  assign y10212 = ~n22801 ;
  assign y10213 = ~1'b0 ;
  assign y10214 = n22802 ;
  assign y10215 = ~n22809 ;
  assign y10216 = ~1'b0 ;
  assign y10217 = n22810 ;
  assign y10218 = n22819 ;
  assign y10219 = ~1'b0 ;
  assign y10220 = n22821 ;
  assign y10221 = ~1'b0 ;
  assign y10222 = ~1'b0 ;
  assign y10223 = 1'b0 ;
  assign y10224 = n22825 ;
  assign y10225 = ~n22826 ;
  assign y10226 = n22828 ;
  assign y10227 = n22841 ;
  assign y10228 = ~n22843 ;
  assign y10229 = ~1'b0 ;
  assign y10230 = ~n22844 ;
  assign y10231 = n22848 ;
  assign y10232 = ~n22855 ;
  assign y10233 = ~n22856 ;
  assign y10234 = ~n22858 ;
  assign y10235 = ~1'b0 ;
  assign y10236 = n22865 ;
  assign y10237 = ~n22867 ;
  assign y10238 = n22871 ;
  assign y10239 = ~1'b0 ;
  assign y10240 = n22873 ;
  assign y10241 = n22876 ;
  assign y10242 = ~n16378 ;
  assign y10243 = ~n22884 ;
  assign y10244 = n22562 ;
  assign y10245 = ~n22887 ;
  assign y10246 = ~n22890 ;
  assign y10247 = ~n22894 ;
  assign y10248 = ~n22897 ;
  assign y10249 = ~1'b0 ;
  assign y10250 = ~1'b0 ;
  assign y10251 = ~n22899 ;
  assign y10252 = ~n22900 ;
  assign y10253 = n22902 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = ~n22905 ;
  assign y10256 = ~1'b0 ;
  assign y10257 = n22906 ;
  assign y10258 = ~1'b0 ;
  assign y10259 = n12994 ;
  assign y10260 = ~n22908 ;
  assign y10261 = ~n22909 ;
  assign y10262 = ~1'b0 ;
  assign y10263 = n22915 ;
  assign y10264 = n22920 ;
  assign y10265 = n22923 ;
  assign y10266 = ~n22924 ;
  assign y10267 = n22926 ;
  assign y10268 = n22931 ;
  assign y10269 = ~n22935 ;
  assign y10270 = ~n10673 ;
  assign y10271 = ~1'b0 ;
  assign y10272 = n22936 ;
  assign y10273 = ~1'b0 ;
  assign y10274 = n22938 ;
  assign y10275 = ~n22939 ;
  assign y10276 = n22940 ;
  assign y10277 = n22947 ;
  assign y10278 = n8349 ;
  assign y10279 = ~n22952 ;
  assign y10280 = ~n22956 ;
  assign y10281 = ~1'b0 ;
  assign y10282 = n22958 ;
  assign y10283 = ~n22962 ;
  assign y10284 = n22964 ;
  assign y10285 = ~n22972 ;
  assign y10286 = ~n22974 ;
  assign y10287 = n22975 ;
  assign y10288 = ~1'b0 ;
  assign y10289 = ~n22983 ;
  assign y10290 = ~1'b0 ;
  assign y10291 = ~n22989 ;
  assign y10292 = n22993 ;
  assign y10293 = n22995 ;
  assign y10294 = ~n22996 ;
  assign y10295 = ~1'b0 ;
  assign y10296 = ~n22998 ;
  assign y10297 = ~n23000 ;
  assign y10298 = ~n23003 ;
  assign y10299 = ~n23007 ;
  assign y10300 = ~1'b0 ;
  assign y10301 = ~n23013 ;
  assign y10302 = ~n23014 ;
  assign y10303 = ~n23015 ;
  assign y10304 = n23019 ;
  assign y10305 = n23022 ;
  assign y10306 = ~1'b0 ;
  assign y10307 = ~n23023 ;
  assign y10308 = n23026 ;
  assign y10309 = ~n23027 ;
  assign y10310 = n10849 ;
  assign y10311 = ~n151 ;
  assign y10312 = ~n23029 ;
  assign y10313 = n23030 ;
  assign y10314 = n23033 ;
  assign y10315 = ~1'b0 ;
  assign y10316 = ~n23038 ;
  assign y10317 = ~n23044 ;
  assign y10318 = n23046 ;
  assign y10319 = ~1'b0 ;
  assign y10320 = n2282 ;
  assign y10321 = n23049 ;
  assign y10322 = ~1'b0 ;
  assign y10323 = ~1'b0 ;
  assign y10324 = n23050 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = ~n23057 ;
  assign y10327 = 1'b0 ;
  assign y10328 = ~n23059 ;
  assign y10329 = n23060 ;
  assign y10330 = ~1'b0 ;
  assign y10331 = n23062 ;
  assign y10332 = ~n23063 ;
  assign y10333 = ~1'b0 ;
  assign y10334 = n23064 ;
  assign y10335 = n23065 ;
  assign y10336 = n23066 ;
  assign y10337 = n23067 ;
  assign y10338 = ~1'b0 ;
  assign y10339 = ~n23074 ;
  assign y10340 = ~n23076 ;
  assign y10341 = ~1'b0 ;
  assign y10342 = n23081 ;
  assign y10343 = ~n23083 ;
  assign y10344 = 1'b0 ;
  assign y10345 = ~n23087 ;
  assign y10346 = n23088 ;
  assign y10347 = ~1'b0 ;
  assign y10348 = n23096 ;
  assign y10349 = ~n23100 ;
  assign y10350 = ~n23101 ;
  assign y10351 = n23103 ;
  assign y10352 = n23105 ;
  assign y10353 = n23112 ;
  assign y10354 = n23120 ;
  assign y10355 = n23121 ;
  assign y10356 = ~1'b0 ;
  assign y10357 = ~n23124 ;
  assign y10358 = ~n23130 ;
  assign y10359 = ~n23131 ;
  assign y10360 = n23135 ;
  assign y10361 = ~1'b0 ;
  assign y10362 = n23136 ;
  assign y10363 = n23138 ;
  assign y10364 = ~1'b0 ;
  assign y10365 = ~n23142 ;
  assign y10366 = 1'b0 ;
  assign y10367 = n23144 ;
  assign y10368 = n23145 ;
  assign y10369 = ~n1138 ;
  assign y10370 = ~1'b0 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = ~1'b0 ;
  assign y10373 = ~1'b0 ;
  assign y10374 = ~1'b0 ;
  assign y10375 = ~1'b0 ;
  assign y10376 = n23147 ;
  assign y10377 = ~1'b0 ;
  assign y10378 = ~1'b0 ;
  assign y10379 = ~1'b0 ;
  assign y10380 = n12626 ;
  assign y10381 = n23148 ;
  assign y10382 = ~n23149 ;
  assign y10383 = n23151 ;
  assign y10384 = n23159 ;
  assign y10385 = ~1'b0 ;
  assign y10386 = ~1'b0 ;
  assign y10387 = n23161 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = n23162 ;
  assign y10390 = ~n23164 ;
  assign y10391 = ~1'b0 ;
  assign y10392 = ~1'b0 ;
  assign y10393 = n23165 ;
  assign y10394 = ~n23171 ;
  assign y10395 = ~n23173 ;
  assign y10396 = n23177 ;
  assign y10397 = ~n23179 ;
  assign y10398 = n23181 ;
  assign y10399 = ~n23185 ;
  assign y10400 = ~1'b0 ;
  assign y10401 = ~n23187 ;
  assign y10402 = n23189 ;
  assign y10403 = n23190 ;
  assign y10404 = ~1'b0 ;
  assign y10405 = ~n23191 ;
  assign y10406 = n1171 ;
  assign y10407 = ~n23195 ;
  assign y10408 = ~1'b0 ;
  assign y10409 = ~1'b0 ;
  assign y10410 = ~n23202 ;
  assign y10411 = ~n23204 ;
  assign y10412 = n23205 ;
  assign y10413 = n23208 ;
  assign y10414 = ~1'b0 ;
  assign y10415 = ~n23210 ;
  assign y10416 = n23211 ;
  assign y10417 = ~n23212 ;
  assign y10418 = n23216 ;
  assign y10419 = n23217 ;
  assign y10420 = n23222 ;
  assign y10421 = ~1'b0 ;
  assign y10422 = ~n23224 ;
  assign y10423 = n23225 ;
  assign y10424 = n23232 ;
  assign y10425 = ~n23234 ;
  assign y10426 = ~n23235 ;
  assign y10427 = ~n23237 ;
  assign y10428 = n23242 ;
  assign y10429 = ~n23250 ;
  assign y10430 = ~n23256 ;
  assign y10431 = ~n23259 ;
  assign y10432 = ~n23262 ;
  assign y10433 = n23267 ;
  assign y10434 = ~n23269 ;
  assign y10435 = ~n23271 ;
  assign y10436 = ~n23275 ;
  assign y10437 = ~1'b0 ;
  assign y10438 = n23278 ;
  assign y10439 = n23279 ;
  assign y10440 = ~n23288 ;
  assign y10441 = n23292 ;
  assign y10442 = n23295 ;
  assign y10443 = 1'b0 ;
  assign y10444 = n23296 ;
  assign y10445 = n23297 ;
  assign y10446 = n23300 ;
  assign y10447 = n23304 ;
  assign y10448 = ~1'b0 ;
  assign y10449 = ~1'b0 ;
  assign y10450 = ~n23305 ;
  assign y10451 = ~1'b0 ;
  assign y10452 = ~1'b0 ;
  assign y10453 = ~1'b0 ;
  assign y10454 = n23313 ;
  assign y10455 = ~n23314 ;
  assign y10456 = n23316 ;
  assign y10457 = n23318 ;
  assign y10458 = n23320 ;
  assign y10459 = n23326 ;
  assign y10460 = n23328 ;
  assign y10461 = ~n23330 ;
  assign y10462 = n10226 ;
  assign y10463 = n23337 ;
  assign y10464 = ~n23341 ;
  assign y10465 = n23342 ;
  assign y10466 = 1'b0 ;
  assign y10467 = ~n23343 ;
  assign y10468 = ~n23344 ;
  assign y10469 = ~1'b0 ;
  assign y10470 = n23345 ;
  assign y10471 = n23347 ;
  assign y10472 = ~1'b0 ;
  assign y10473 = ~x9 ;
  assign y10474 = ~n23349 ;
  assign y10475 = ~1'b0 ;
  assign y10476 = ~1'b0 ;
  assign y10477 = n23356 ;
  assign y10478 = n23357 ;
  assign y10479 = ~n23359 ;
  assign y10480 = ~n23361 ;
  assign y10481 = ~n23362 ;
  assign y10482 = n23366 ;
  assign y10483 = n5120 ;
  assign y10484 = n23369 ;
  assign y10485 = ~n23371 ;
  assign y10486 = n23375 ;
  assign y10487 = ~1'b0 ;
  assign y10488 = n23378 ;
  assign y10489 = n23380 ;
  assign y10490 = ~n23381 ;
  assign y10491 = ~n23382 ;
  assign y10492 = n23383 ;
  assign y10493 = ~1'b0 ;
  assign y10494 = ~n23384 ;
  assign y10495 = n23386 ;
  assign y10496 = ~1'b0 ;
  assign y10497 = ~1'b0 ;
  assign y10498 = ~n23387 ;
  assign y10499 = n23391 ;
  assign y10500 = ~1'b0 ;
  assign y10501 = n23394 ;
  assign y10502 = ~1'b0 ;
  assign y10503 = ~n23395 ;
  assign y10504 = n23398 ;
  assign y10505 = ~1'b0 ;
  assign y10506 = ~1'b0 ;
  assign y10507 = ~n23402 ;
  assign y10508 = ~1'b0 ;
  assign y10509 = ~1'b0 ;
  assign y10510 = n23404 ;
  assign y10511 = ~n23406 ;
  assign y10512 = n23410 ;
  assign y10513 = n23411 ;
  assign y10514 = ~1'b0 ;
  assign y10515 = ~n23416 ;
  assign y10516 = ~n23420 ;
  assign y10517 = n23424 ;
  assign y10518 = n23430 ;
  assign y10519 = ~1'b0 ;
  assign y10520 = ~n19083 ;
  assign y10521 = ~n23431 ;
  assign y10522 = ~n23435 ;
  assign y10523 = n23439 ;
  assign y10524 = ~1'b0 ;
  assign y10525 = ~1'b0 ;
  assign y10526 = ~n23442 ;
  assign y10527 = ~n23444 ;
  assign y10528 = n23448 ;
  assign y10529 = n23451 ;
  assign y10530 = n23454 ;
  assign y10531 = ~n23457 ;
  assign y10532 = n23463 ;
  assign y10533 = ~n23468 ;
  assign y10534 = n23469 ;
  assign y10535 = ~1'b0 ;
  assign y10536 = ~1'b0 ;
  assign y10537 = ~n23472 ;
  assign y10538 = ~n17245 ;
  assign y10539 = ~n23474 ;
  assign y10540 = ~1'b0 ;
  assign y10541 = ~n23477 ;
  assign y10542 = ~n23479 ;
  assign y10543 = ~n23481 ;
  assign y10544 = ~1'b0 ;
  assign y10545 = n23483 ;
  assign y10546 = ~n23485 ;
  assign y10547 = n23488 ;
  assign y10548 = n23489 ;
  assign y10549 = ~1'b0 ;
  assign y10550 = ~n23495 ;
  assign y10551 = ~n4465 ;
  assign y10552 = ~n23501 ;
  assign y10553 = n23507 ;
  assign y10554 = ~1'b0 ;
  assign y10555 = ~n23513 ;
  assign y10556 = ~1'b0 ;
  assign y10557 = n23516 ;
  assign y10558 = ~n23517 ;
  assign y10559 = ~n23519 ;
  assign y10560 = n23522 ;
  assign y10561 = n23524 ;
  assign y10562 = ~1'b0 ;
  assign y10563 = ~n23527 ;
  assign y10564 = n23528 ;
  assign y10565 = n23530 ;
  assign y10566 = n5120 ;
  assign y10567 = n23531 ;
  assign y10568 = ~n23535 ;
  assign y10569 = ~n23536 ;
  assign y10570 = ~n23554 ;
  assign y10571 = ~n23556 ;
  assign y10572 = ~1'b0 ;
  assign y10573 = ~n23562 ;
  assign y10574 = n392 ;
  assign y10575 = n23564 ;
  assign y10576 = ~n23568 ;
  assign y10577 = ~1'b0 ;
  assign y10578 = n23569 ;
  assign y10579 = n23570 ;
  assign y10580 = ~n23574 ;
  assign y10581 = ~1'b0 ;
  assign y10582 = n23576 ;
  assign y10583 = n23579 ;
  assign y10584 = ~n23581 ;
  assign y10585 = ~n2322 ;
  assign y10586 = n15119 ;
  assign y10587 = n2251 ;
  assign y10588 = ~1'b0 ;
  assign y10589 = n23582 ;
  assign y10590 = ~1'b0 ;
  assign y10591 = ~n23585 ;
  assign y10592 = n23591 ;
  assign y10593 = ~n5395 ;
  assign y10594 = ~n23595 ;
  assign y10595 = ~n23598 ;
  assign y10596 = ~n23600 ;
  assign y10597 = ~n23603 ;
  assign y10598 = ~1'b0 ;
  assign y10599 = n23605 ;
  assign y10600 = n23609 ;
  assign y10601 = n23620 ;
  assign y10602 = ~n23623 ;
  assign y10603 = ~n23626 ;
  assign y10604 = n23628 ;
  assign y10605 = ~1'b0 ;
  assign y10606 = ~n23629 ;
  assign y10607 = ~n23631 ;
  assign y10608 = ~n23633 ;
  assign y10609 = ~n23635 ;
  assign y10610 = n23638 ;
  assign y10611 = ~1'b0 ;
  assign y10612 = ~n23639 ;
  assign y10613 = n23640 ;
  assign y10614 = ~n23642 ;
  assign y10615 = ~n23644 ;
  assign y10616 = n23645 ;
  assign y10617 = ~n23647 ;
  assign y10618 = n23659 ;
  assign y10619 = ~n23661 ;
  assign y10620 = ~n23665 ;
  assign y10621 = ~n23667 ;
  assign y10622 = ~n23668 ;
  assign y10623 = ~n23669 ;
  assign y10624 = ~n18179 ;
  assign y10625 = n23678 ;
  assign y10626 = n23680 ;
  assign y10627 = n23681 ;
  assign y10628 = ~n23683 ;
  assign y10629 = n23685 ;
  assign y10630 = ~1'b0 ;
  assign y10631 = n23686 ;
  assign y10632 = n23689 ;
  assign y10633 = ~n23691 ;
  assign y10634 = n23695 ;
  assign y10635 = ~n23698 ;
  assign y10636 = ~n23702 ;
  assign y10637 = ~n23705 ;
  assign y10638 = ~n23707 ;
  assign y10639 = ~1'b0 ;
  assign y10640 = ~n23708 ;
  assign y10641 = n23709 ;
  assign y10642 = ~n23715 ;
  assign y10643 = n23716 ;
  assign y10644 = n23719 ;
  assign y10645 = ~n23723 ;
  assign y10646 = n23724 ;
  assign y10647 = n23726 ;
  assign y10648 = n23727 ;
  assign y10649 = ~n23730 ;
  assign y10650 = n23735 ;
  assign y10651 = n23736 ;
  assign y10652 = n23751 ;
  assign y10653 = n23752 ;
  assign y10654 = n23753 ;
  assign y10655 = ~1'b0 ;
  assign y10656 = ~1'b0 ;
  assign y10657 = n7255 ;
  assign y10658 = ~n23757 ;
  assign y10659 = n2620 ;
  assign y10660 = n23759 ;
  assign y10661 = ~n23763 ;
  assign y10662 = ~1'b0 ;
  assign y10663 = ~n23765 ;
  assign y10664 = n23767 ;
  assign y10665 = n23769 ;
  assign y10666 = ~1'b0 ;
  assign y10667 = n23771 ;
  assign y10668 = ~n23773 ;
  assign y10669 = ~1'b0 ;
  assign y10670 = ~n23774 ;
  assign y10671 = ~n23775 ;
  assign y10672 = n23779 ;
  assign y10673 = ~n23783 ;
  assign y10674 = ~1'b0 ;
  assign y10675 = ~n23785 ;
  assign y10676 = n23788 ;
  assign y10677 = ~n23798 ;
  assign y10678 = ~n23800 ;
  assign y10679 = ~1'b0 ;
  assign y10680 = ~n23803 ;
  assign y10681 = ~n23808 ;
  assign y10682 = n23813 ;
  assign y10683 = ~1'b0 ;
  assign y10684 = n23814 ;
  assign y10685 = ~n23818 ;
  assign y10686 = n23819 ;
  assign y10687 = ~n23822 ;
  assign y10688 = n23828 ;
  assign y10689 = 1'b0 ;
  assign y10690 = n23830 ;
  assign y10691 = n23831 ;
  assign y10692 = ~n23833 ;
  assign y10693 = ~1'b0 ;
  assign y10694 = ~1'b0 ;
  assign y10695 = ~n23837 ;
  assign y10696 = ~n23838 ;
  assign y10697 = n23845 ;
  assign y10698 = ~n23846 ;
  assign y10699 = ~n23848 ;
  assign y10700 = ~n23849 ;
  assign y10701 = 1'b0 ;
  assign y10702 = n23851 ;
  assign y10703 = ~n23854 ;
  assign y10704 = n23859 ;
  assign y10705 = ~n23862 ;
  assign y10706 = ~n23866 ;
  assign y10707 = n23867 ;
  assign y10708 = ~1'b0 ;
  assign y10709 = n23870 ;
  assign y10710 = 1'b0 ;
  assign y10711 = ~1'b0 ;
  assign y10712 = ~1'b0 ;
  assign y10713 = ~1'b0 ;
  assign y10714 = ~n23873 ;
  assign y10715 = ~n23875 ;
  assign y10716 = ~n23879 ;
  assign y10717 = n23881 ;
  assign y10718 = n23883 ;
  assign y10719 = n23888 ;
  assign y10720 = ~n23889 ;
  assign y10721 = n3731 ;
  assign y10722 = n23891 ;
  assign y10723 = n23894 ;
  assign y10724 = ~n23895 ;
  assign y10725 = ~1'b0 ;
  assign y10726 = ~1'b0 ;
  assign y10727 = ~n23897 ;
  assign y10728 = ~n23900 ;
  assign y10729 = n16177 ;
  assign y10730 = ~n23901 ;
  assign y10731 = ~1'b0 ;
  assign y10732 = ~n23902 ;
  assign y10733 = ~n23904 ;
  assign y10734 = ~n23907 ;
  assign y10735 = ~1'b0 ;
  assign y10736 = ~1'b0 ;
  assign y10737 = n23909 ;
  assign y10738 = ~n23911 ;
  assign y10739 = ~1'b0 ;
  assign y10740 = ~1'b0 ;
  assign y10741 = n23913 ;
  assign y10742 = ~n23914 ;
  assign y10743 = ~n23918 ;
  assign y10744 = n23926 ;
  assign y10745 = ~1'b0 ;
  assign y10746 = ~n23929 ;
  assign y10747 = ~n23930 ;
  assign y10748 = n23931 ;
  assign y10749 = n250 ;
  assign y10750 = n23937 ;
  assign y10751 = ~n11051 ;
  assign y10752 = n23938 ;
  assign y10753 = ~n23940 ;
  assign y10754 = n23950 ;
  assign y10755 = ~1'b0 ;
  assign y10756 = ~n23954 ;
  assign y10757 = n23955 ;
  assign y10758 = ~n23956 ;
  assign y10759 = n23959 ;
  assign y10760 = n23961 ;
  assign y10761 = n23966 ;
  assign y10762 = n23970 ;
  assign y10763 = ~1'b0 ;
  assign y10764 = n23971 ;
  assign y10765 = ~1'b0 ;
  assign y10766 = ~n23975 ;
  assign y10767 = ~n23979 ;
  assign y10768 = ~n23983 ;
  assign y10769 = n23984 ;
  assign y10770 = ~1'b0 ;
  assign y10771 = ~1'b0 ;
  assign y10772 = ~n23988 ;
  assign y10773 = n23989 ;
  assign y10774 = ~1'b0 ;
  assign y10775 = n23990 ;
  assign y10776 = ~1'b0 ;
  assign y10777 = n23994 ;
  assign y10778 = n23996 ;
  assign y10779 = ~1'b0 ;
  assign y10780 = ~1'b0 ;
  assign y10781 = ~n22177 ;
  assign y10782 = n23997 ;
  assign y10783 = ~1'b0 ;
  assign y10784 = ~n23999 ;
  assign y10785 = n24003 ;
  assign y10786 = n16021 ;
  assign y10787 = ~1'b0 ;
  assign y10788 = ~1'b0 ;
  assign y10789 = n24004 ;
  assign y10790 = n24005 ;
  assign y10791 = ~1'b0 ;
  assign y10792 = ~n24007 ;
  assign y10793 = ~1'b0 ;
  assign y10794 = ~n24010 ;
  assign y10795 = n24011 ;
  assign y10796 = ~1'b0 ;
  assign y10797 = n24013 ;
  assign y10798 = ~1'b0 ;
  assign y10799 = ~n19429 ;
  assign y10800 = n24014 ;
  assign y10801 = n24016 ;
  assign y10802 = ~n24019 ;
  assign y10803 = ~1'b0 ;
  assign y10804 = n24025 ;
  assign y10805 = ~1'b0 ;
  assign y10806 = ~1'b0 ;
  assign y10807 = n24026 ;
  assign y10808 = n624 ;
  assign y10809 = n24027 ;
  assign y10810 = ~n24029 ;
  assign y10811 = ~n469 ;
  assign y10812 = ~1'b0 ;
  assign y10813 = ~n24030 ;
  assign y10814 = ~n24032 ;
  assign y10815 = n24034 ;
  assign y10816 = ~n24035 ;
  assign y10817 = n24043 ;
  assign y10818 = n24045 ;
  assign y10819 = ~1'b0 ;
  assign y10820 = ~1'b0 ;
  assign y10821 = ~n24046 ;
  assign y10822 = ~n24047 ;
  assign y10823 = n13583 ;
  assign y10824 = n24049 ;
  assign y10825 = n24051 ;
  assign y10826 = n24053 ;
  assign y10827 = ~1'b0 ;
  assign y10828 = ~n24054 ;
  assign y10829 = n24055 ;
  assign y10830 = ~1'b0 ;
  assign y10831 = n24060 ;
  assign y10832 = ~1'b0 ;
  assign y10833 = n24062 ;
  assign y10834 = n24069 ;
  assign y10835 = n24073 ;
  assign y10836 = n24077 ;
  assign y10837 = ~1'b0 ;
  assign y10838 = ~n24081 ;
  assign y10839 = ~1'b0 ;
  assign y10840 = n24087 ;
  assign y10841 = ~n24090 ;
  assign y10842 = ~n24095 ;
  assign y10843 = n24096 ;
  assign y10844 = ~1'b0 ;
  assign y10845 = ~1'b0 ;
  assign y10846 = n24099 ;
  assign y10847 = ~n886 ;
  assign y10848 = n9830 ;
  assign y10849 = ~n24100 ;
  assign y10850 = ~1'b0 ;
  assign y10851 = ~n24104 ;
  assign y10852 = n24106 ;
  assign y10853 = n24109 ;
  assign y10854 = n24117 ;
  assign y10855 = ~n24119 ;
  assign y10856 = n24126 ;
  assign y10857 = n24128 ;
  assign y10858 = ~n24130 ;
  assign y10859 = ~n24134 ;
  assign y10860 = n24136 ;
  assign y10861 = n24145 ;
  assign y10862 = ~n24147 ;
  assign y10863 = ~1'b0 ;
  assign y10864 = ~n24151 ;
  assign y10865 = n24153 ;
  assign y10866 = n24163 ;
  assign y10867 = n24168 ;
  assign y10868 = n24171 ;
  assign y10869 = ~1'b0 ;
  assign y10870 = ~n24180 ;
  assign y10871 = ~1'b0 ;
  assign y10872 = ~1'b0 ;
  assign y10873 = ~1'b0 ;
  assign y10874 = n24182 ;
  assign y10875 = ~n24185 ;
  assign y10876 = n24186 ;
  assign y10877 = ~1'b0 ;
  assign y10878 = n24190 ;
  assign y10879 = n24192 ;
  assign y10880 = ~n24197 ;
  assign y10881 = n24199 ;
  assign y10882 = ~1'b0 ;
  assign y10883 = ~n24204 ;
  assign y10884 = ~n24207 ;
  assign y10885 = ~n24212 ;
  assign y10886 = ~n24219 ;
  assign y10887 = n24224 ;
  assign y10888 = n24230 ;
  assign y10889 = n24233 ;
  assign y10890 = n24239 ;
  assign y10891 = ~n24242 ;
  assign y10892 = ~n11038 ;
  assign y10893 = n24244 ;
  assign y10894 = n24247 ;
  assign y10895 = 1'b0 ;
  assign y10896 = n24254 ;
  assign y10897 = ~n24255 ;
  assign y10898 = ~n24260 ;
  assign y10899 = n24261 ;
  assign y10900 = n24265 ;
  assign y10901 = n24267 ;
  assign y10902 = ~n24272 ;
  assign y10903 = n24273 ;
  assign y10904 = ~1'b0 ;
  assign y10905 = ~n24274 ;
  assign y10906 = n18268 ;
  assign y10907 = ~n24281 ;
  assign y10908 = ~n8493 ;
  assign y10909 = n24283 ;
  assign y10910 = ~n19170 ;
  assign y10911 = ~1'b0 ;
  assign y10912 = ~1'b0 ;
  assign y10913 = ~n24286 ;
  assign y10914 = ~n24287 ;
  assign y10915 = n24289 ;
  assign y10916 = ~1'b0 ;
  assign y10917 = n23216 ;
  assign y10918 = ~1'b0 ;
  assign y10919 = n24291 ;
  assign y10920 = ~1'b0 ;
  assign y10921 = ~1'b0 ;
  assign y10922 = ~1'b0 ;
  assign y10923 = n24292 ;
  assign y10924 = n24298 ;
  assign y10925 = ~1'b0 ;
  assign y10926 = n24304 ;
  assign y10927 = ~n24312 ;
  assign y10928 = 1'b0 ;
  assign y10929 = ~1'b0 ;
  assign y10930 = ~1'b0 ;
  assign y10931 = n24316 ;
  assign y10932 = ~n24318 ;
  assign y10933 = 1'b0 ;
  assign y10934 = n24321 ;
  assign y10935 = ~1'b0 ;
  assign y10936 = n24324 ;
  assign y10937 = ~n24328 ;
  assign y10938 = n24330 ;
  assign y10939 = ~n24334 ;
  assign y10940 = n24340 ;
  assign y10941 = ~1'b0 ;
  assign y10942 = n24343 ;
  assign y10943 = n24345 ;
  assign y10944 = ~n24346 ;
  assign y10945 = n24347 ;
  assign y10946 = n24351 ;
  assign y10947 = ~n24353 ;
  assign y10948 = n24355 ;
  assign y10949 = n24358 ;
  assign y10950 = ~n24359 ;
  assign y10951 = ~n24360 ;
  assign y10952 = ~1'b0 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = n691 ;
  assign y10955 = ~1'b0 ;
  assign y10956 = ~1'b0 ;
  assign y10957 = ~n24364 ;
  assign y10958 = ~n24366 ;
  assign y10959 = n24367 ;
  assign y10960 = ~n24370 ;
  assign y10961 = ~n24372 ;
  assign y10962 = n24374 ;
  assign y10963 = n24376 ;
  assign y10964 = n24378 ;
  assign y10965 = ~n24382 ;
  assign y10966 = ~1'b0 ;
  assign y10967 = n24384 ;
  assign y10968 = ~n24385 ;
  assign y10969 = ~n18096 ;
  assign y10970 = n24388 ;
  assign y10971 = ~n24389 ;
  assign y10972 = ~n24392 ;
  assign y10973 = n24400 ;
  assign y10974 = ~1'b0 ;
  assign y10975 = n24402 ;
  assign y10976 = ~1'b0 ;
  assign y10977 = ~1'b0 ;
  assign y10978 = ~n24404 ;
  assign y10979 = n24406 ;
  assign y10980 = ~n24407 ;
  assign y10981 = n24410 ;
  assign y10982 = ~1'b0 ;
  assign y10983 = ~1'b0 ;
  assign y10984 = n181 ;
  assign y10985 = ~n24415 ;
  assign y10986 = ~n24419 ;
  assign y10987 = n24424 ;
  assign y10988 = ~1'b0 ;
  assign y10989 = n24425 ;
  assign y10990 = ~1'b0 ;
  assign y10991 = ~1'b0 ;
  assign y10992 = n24427 ;
  assign y10993 = ~n24430 ;
  assign y10994 = ~1'b0 ;
  assign y10995 = ~n24436 ;
  assign y10996 = ~n24439 ;
  assign y10997 = ~1'b0 ;
  assign y10998 = n24442 ;
  assign y10999 = ~n14460 ;
  assign y11000 = n24444 ;
  assign y11001 = ~n24446 ;
  assign y11002 = ~1'b0 ;
  assign y11003 = ~1'b0 ;
  assign y11004 = ~n24448 ;
  assign y11005 = ~n3383 ;
  assign y11006 = ~n24450 ;
  assign y11007 = ~1'b0 ;
  assign y11008 = n24451 ;
  assign y11009 = n24453 ;
  assign y11010 = ~1'b0 ;
  assign y11011 = ~1'b0 ;
  assign y11012 = ~n24454 ;
  assign y11013 = n12054 ;
  assign y11014 = n24457 ;
  assign y11015 = ~1'b0 ;
  assign y11016 = ~1'b0 ;
  assign y11017 = ~n24460 ;
  assign y11018 = ~1'b0 ;
  assign y11019 = n24467 ;
  assign y11020 = ~n24470 ;
  assign y11021 = n24473 ;
  assign y11022 = n24483 ;
  assign y11023 = 1'b0 ;
  assign y11024 = n24484 ;
  assign y11025 = n24488 ;
  assign y11026 = n24489 ;
  assign y11027 = ~n1962 ;
  assign y11028 = ~1'b0 ;
  assign y11029 = ~n24490 ;
  assign y11030 = n24494 ;
  assign y11031 = ~n2982 ;
  assign y11032 = n24495 ;
  assign y11033 = ~n24498 ;
  assign y11034 = n24501 ;
  assign y11035 = ~1'b0 ;
  assign y11036 = n20708 ;
  assign y11037 = ~1'b0 ;
  assign y11038 = ~n24504 ;
  assign y11039 = n24507 ;
  assign y11040 = ~n24509 ;
  assign y11041 = ~n24510 ;
  assign y11042 = n24511 ;
  assign y11043 = ~n24512 ;
  assign y11044 = ~n24515 ;
  assign y11045 = n24516 ;
  assign y11046 = ~n24517 ;
  assign y11047 = ~n24520 ;
  assign y11048 = n24522 ;
  assign y11049 = ~n24530 ;
  assign y11050 = ~1'b0 ;
  assign y11051 = n24534 ;
  assign y11052 = ~n24535 ;
  assign y11053 = ~n24538 ;
  assign y11054 = n24541 ;
  assign y11055 = ~n24546 ;
  assign y11056 = ~1'b0 ;
  assign y11057 = ~n24549 ;
  assign y11058 = 1'b0 ;
  assign y11059 = ~1'b0 ;
  assign y11060 = ~1'b0 ;
  assign y11061 = n24551 ;
  assign y11062 = ~n24556 ;
  assign y11063 = ~n24557 ;
  assign y11064 = ~1'b0 ;
  assign y11065 = n24560 ;
  assign y11066 = ~n24561 ;
  assign y11067 = ~1'b0 ;
  assign y11068 = ~1'b0 ;
  assign y11069 = ~n24563 ;
  assign y11070 = ~n24568 ;
  assign y11071 = ~n24576 ;
  assign y11072 = n24587 ;
  assign y11073 = ~n1185 ;
  assign y11074 = ~n24589 ;
  assign y11075 = n24591 ;
  assign y11076 = ~n24593 ;
  assign y11077 = n24595 ;
  assign y11078 = ~n24598 ;
  assign y11079 = ~n24599 ;
  assign y11080 = ~n24600 ;
  assign y11081 = n24604 ;
  assign y11082 = ~1'b0 ;
  assign y11083 = n24611 ;
  assign y11084 = ~n24615 ;
  assign y11085 = n20824 ;
  assign y11086 = n24618 ;
  assign y11087 = ~1'b0 ;
  assign y11088 = ~n24619 ;
  assign y11089 = n24621 ;
  assign y11090 = ~1'b0 ;
  assign y11091 = ~n24623 ;
  assign y11092 = n24625 ;
  assign y11093 = n24628 ;
  assign y11094 = n24636 ;
  assign y11095 = n24637 ;
  assign y11096 = n15209 ;
  assign y11097 = ~1'b0 ;
  assign y11098 = ~1'b0 ;
  assign y11099 = n24646 ;
  assign y11100 = ~n24651 ;
  assign y11101 = n24657 ;
  assign y11102 = ~n24660 ;
  assign y11103 = ~1'b0 ;
  assign y11104 = ~1'b0 ;
  assign y11105 = ~n24662 ;
  assign y11106 = ~1'b0 ;
  assign y11107 = ~n24668 ;
  assign y11108 = ~n24670 ;
  assign y11109 = ~n24672 ;
  assign y11110 = n24678 ;
  assign y11111 = ~1'b0 ;
  assign y11112 = ~1'b0 ;
  assign y11113 = n24683 ;
  assign y11114 = n24684 ;
  assign y11115 = n24686 ;
  assign y11116 = ~n24692 ;
  assign y11117 = n24695 ;
  assign y11118 = ~n24698 ;
  assign y11119 = n24700 ;
  assign y11120 = ~1'b0 ;
  assign y11121 = ~1'b0 ;
  assign y11122 = n24702 ;
  assign y11123 = ~1'b0 ;
  assign y11124 = ~n24706 ;
  assign y11125 = ~n24709 ;
  assign y11126 = ~n211 ;
  assign y11127 = ~n24711 ;
  assign y11128 = ~n16746 ;
  assign y11129 = ~n24712 ;
  assign y11130 = ~n24713 ;
  assign y11131 = ~n24715 ;
  assign y11132 = ~1'b0 ;
  assign y11133 = ~n24721 ;
  assign y11134 = 1'b0 ;
  assign y11135 = ~n24726 ;
  assign y11136 = n24728 ;
  assign y11137 = ~n24729 ;
  assign y11138 = ~1'b0 ;
  assign y11139 = n24731 ;
  assign y11140 = ~1'b0 ;
  assign y11141 = n24740 ;
  assign y11142 = ~1'b0 ;
  assign y11143 = ~n24742 ;
  assign y11144 = n24743 ;
  assign y11145 = 1'b0 ;
  assign y11146 = n24744 ;
  assign y11147 = ~n24746 ;
  assign y11148 = ~1'b0 ;
  assign y11149 = n24751 ;
  assign y11150 = n24752 ;
  assign y11151 = ~n24760 ;
  assign y11152 = n24763 ;
  assign y11153 = ~n24764 ;
  assign y11154 = ~1'b0 ;
  assign y11155 = ~n24765 ;
  assign y11156 = ~1'b0 ;
  assign y11157 = n24768 ;
  assign y11158 = ~1'b0 ;
  assign y11159 = ~1'b0 ;
  assign y11160 = n24771 ;
  assign y11161 = n5876 ;
  assign y11162 = ~1'b0 ;
  assign y11163 = n24773 ;
  assign y11164 = ~1'b0 ;
  assign y11165 = ~n24775 ;
  assign y11166 = n24776 ;
  assign y11167 = ~n24781 ;
  assign y11168 = ~1'b0 ;
  assign y11169 = n24782 ;
  assign y11170 = ~n24787 ;
  assign y11171 = ~n24792 ;
  assign y11172 = ~1'b0 ;
  assign y11173 = n24793 ;
  assign y11174 = n24802 ;
  assign y11175 = ~n24804 ;
  assign y11176 = ~n24808 ;
  assign y11177 = n11113 ;
  assign y11178 = n24811 ;
  assign y11179 = 1'b0 ;
  assign y11180 = ~n24814 ;
  assign y11181 = n24819 ;
  assign y11182 = ~n24821 ;
  assign y11183 = n24825 ;
  assign y11184 = 1'b0 ;
  assign y11185 = ~1'b0 ;
  assign y11186 = n24829 ;
  assign y11187 = 1'b0 ;
  assign y11188 = n24832 ;
  assign y11189 = n24598 ;
  assign y11190 = ~n24834 ;
  assign y11191 = ~1'b0 ;
  assign y11192 = ~n24839 ;
  assign y11193 = n24848 ;
  assign y11194 = ~n24850 ;
  assign y11195 = ~1'b0 ;
  assign y11196 = ~n24851 ;
  assign y11197 = n2306 ;
  assign y11198 = n24854 ;
  assign y11199 = ~n24859 ;
  assign y11200 = ~n24862 ;
  assign y11201 = ~1'b0 ;
  assign y11202 = ~n24863 ;
  assign y11203 = ~n24864 ;
  assign y11204 = ~1'b0 ;
  assign y11205 = ~1'b0 ;
  assign y11206 = n8569 ;
  assign y11207 = ~1'b0 ;
  assign y11208 = ~1'b0 ;
  assign y11209 = ~n3310 ;
  assign y11210 = n24871 ;
  assign y11211 = ~n21820 ;
  assign y11212 = n15483 ;
  assign y11213 = n24875 ;
  assign y11214 = ~1'b0 ;
  assign y11215 = ~n24881 ;
  assign y11216 = ~1'b0 ;
  assign y11217 = ~n24883 ;
  assign y11218 = ~n24887 ;
  assign y11219 = ~1'b0 ;
  assign y11220 = n24888 ;
  assign y11221 = ~n24896 ;
  assign y11222 = n24901 ;
  assign y11223 = ~1'b0 ;
  assign y11224 = n4226 ;
  assign y11225 = ~1'b0 ;
  assign y11226 = n24904 ;
  assign y11227 = n24909 ;
  assign y11228 = n24910 ;
  assign y11229 = n24911 ;
  assign y11230 = n24914 ;
  assign y11231 = ~1'b0 ;
  assign y11232 = ~1'b0 ;
  assign y11233 = ~1'b0 ;
  assign y11234 = ~n24917 ;
  assign y11235 = ~n24926 ;
  assign y11236 = ~n24933 ;
  assign y11237 = n24934 ;
  assign y11238 = n24943 ;
  assign y11239 = n24947 ;
  assign y11240 = n3781 ;
  assign y11241 = ~n24950 ;
  assign y11242 = ~1'b0 ;
  assign y11243 = n24951 ;
  assign y11244 = n24952 ;
  assign y11245 = ~n24953 ;
  assign y11246 = ~n24955 ;
  assign y11247 = ~n24957 ;
  assign y11248 = n24960 ;
  assign y11249 = ~1'b0 ;
  assign y11250 = n24963 ;
  assign y11251 = ~1'b0 ;
  assign y11252 = n24965 ;
  assign y11253 = n24966 ;
  assign y11254 = ~1'b0 ;
  assign y11255 = ~n24968 ;
  assign y11256 = ~n24975 ;
  assign y11257 = n24977 ;
  assign y11258 = n24986 ;
  assign y11259 = n7167 ;
  assign y11260 = ~1'b0 ;
  assign y11261 = n1922 ;
  assign y11262 = ~n24987 ;
  assign y11263 = ~n24988 ;
  assign y11264 = ~n24989 ;
  assign y11265 = n24993 ;
  assign y11266 = ~n24995 ;
  assign y11267 = ~n25001 ;
  assign y11268 = n25002 ;
  assign y11269 = ~n25004 ;
  assign y11270 = n25009 ;
  assign y11271 = ~1'b0 ;
  assign y11272 = n25010 ;
  assign y11273 = n25011 ;
  assign y11274 = ~n25013 ;
  assign y11275 = n25018 ;
  assign y11276 = n25020 ;
  assign y11277 = ~1'b0 ;
  assign y11278 = n25023 ;
  assign y11279 = ~n25025 ;
  assign y11280 = ~n10820 ;
  assign y11281 = n25026 ;
  assign y11282 = ~1'b0 ;
  assign y11283 = ~n25029 ;
  assign y11284 = n25034 ;
  assign y11285 = ~1'b0 ;
  assign y11286 = n25035 ;
  assign y11287 = ~n25036 ;
  assign y11288 = ~n25043 ;
  assign y11289 = n25044 ;
  assign y11290 = n25045 ;
  assign y11291 = ~n25048 ;
  assign y11292 = n25052 ;
  assign y11293 = n25056 ;
  assign y11294 = ~1'b0 ;
  assign y11295 = ~n25059 ;
  assign y11296 = ~1'b0 ;
  assign y11297 = n25065 ;
  assign y11298 = ~n25069 ;
  assign y11299 = n25071 ;
  assign y11300 = ~1'b0 ;
  assign y11301 = ~1'b0 ;
  assign y11302 = ~n25073 ;
  assign y11303 = ~n25082 ;
  assign y11304 = ~n25083 ;
  assign y11305 = ~n25086 ;
  assign y11306 = n25090 ;
  assign y11307 = ~1'b0 ;
  assign y11308 = ~1'b0 ;
  assign y11309 = n25093 ;
  assign y11310 = n25094 ;
  assign y11311 = n25096 ;
  assign y11312 = ~1'b0 ;
  assign y11313 = n25099 ;
  assign y11314 = ~1'b0 ;
  assign y11315 = ~1'b0 ;
  assign y11316 = n25105 ;
  assign y11317 = n25110 ;
  assign y11318 = ~1'b0 ;
  assign y11319 = 1'b0 ;
  assign y11320 = ~n25111 ;
  assign y11321 = ~1'b0 ;
  assign y11322 = n25113 ;
  assign y11323 = ~n25116 ;
  assign y11324 = n25117 ;
  assign y11325 = ~1'b0 ;
  assign y11326 = 1'b0 ;
  assign y11327 = ~n25120 ;
  assign y11328 = ~1'b0 ;
  assign y11329 = ~n25130 ;
  assign y11330 = ~n25137 ;
  assign y11331 = ~n25143 ;
  assign y11332 = n25151 ;
  assign y11333 = n25152 ;
  assign y11334 = n25153 ;
  assign y11335 = ~n25154 ;
  assign y11336 = n25160 ;
  assign y11337 = ~n25161 ;
  assign y11338 = ~1'b0 ;
  assign y11339 = ~1'b0 ;
  assign y11340 = ~n25162 ;
  assign y11341 = ~n25163 ;
  assign y11342 = ~n25164 ;
  assign y11343 = ~1'b0 ;
  assign y11344 = ~1'b0 ;
  assign y11345 = ~1'b0 ;
  assign y11346 = n25166 ;
  assign y11347 = ~1'b0 ;
  assign y11348 = n17377 ;
  assign y11349 = n25170 ;
  assign y11350 = ~n25171 ;
  assign y11351 = ~1'b0 ;
  assign y11352 = ~1'b0 ;
  assign y11353 = ~n25176 ;
  assign y11354 = ~n25179 ;
  assign y11355 = n25181 ;
  assign y11356 = ~n25185 ;
  assign y11357 = ~n25189 ;
  assign y11358 = n25193 ;
  assign y11359 = n25194 ;
  assign y11360 = n25197 ;
  assign y11361 = ~1'b0 ;
  assign y11362 = n25204 ;
  assign y11363 = ~n25209 ;
  assign y11364 = n25212 ;
  assign y11365 = ~1'b0 ;
  assign y11366 = n25213 ;
  assign y11367 = ~n25220 ;
  assign y11368 = n25221 ;
  assign y11369 = n25227 ;
  assign y11370 = ~n25230 ;
  assign y11371 = n25233 ;
  assign y11372 = n25236 ;
  assign y11373 = ~1'b0 ;
  assign y11374 = ~n25241 ;
  assign y11375 = ~n25243 ;
  assign y11376 = ~n25244 ;
  assign y11377 = n25248 ;
  assign y11378 = ~n25250 ;
  assign y11379 = n25253 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = ~n25255 ;
  assign y11382 = ~n25259 ;
  assign y11383 = ~1'b0 ;
  assign y11384 = n25263 ;
  assign y11385 = ~n25265 ;
  assign y11386 = ~n25268 ;
  assign y11387 = ~n15520 ;
  assign y11388 = ~n25271 ;
  assign y11389 = ~n25275 ;
  assign y11390 = n25278 ;
  assign y11391 = ~n13889 ;
  assign y11392 = ~n25281 ;
  assign y11393 = ~1'b0 ;
  assign y11394 = ~n25282 ;
  assign y11395 = ~n25285 ;
  assign y11396 = ~n25287 ;
  assign y11397 = ~1'b0 ;
  assign y11398 = n25294 ;
  assign y11399 = n25298 ;
  assign y11400 = ~n25300 ;
  assign y11401 = ~1'b0 ;
  assign y11402 = ~n25305 ;
  assign y11403 = ~1'b0 ;
  assign y11404 = n25308 ;
  assign y11405 = ~1'b0 ;
  assign y11406 = n25309 ;
  assign y11407 = n25310 ;
  assign y11408 = ~n25311 ;
  assign y11409 = n25338 ;
  assign y11410 = ~n25340 ;
  assign y11411 = ~n25342 ;
  assign y11412 = ~n25346 ;
  assign y11413 = ~n16790 ;
  assign y11414 = ~n25348 ;
  assign y11415 = ~1'b0 ;
  assign y11416 = ~n25349 ;
  assign y11417 = ~n25352 ;
  assign y11418 = n25353 ;
  assign y11419 = ~1'b0 ;
  assign y11420 = n25355 ;
  assign y11421 = n25357 ;
  assign y11422 = ~n25358 ;
  assign y11423 = ~1'b0 ;
  assign y11424 = n25368 ;
  assign y11425 = ~n25372 ;
  assign y11426 = n13057 ;
  assign y11427 = ~n25373 ;
  assign y11428 = ~1'b0 ;
  assign y11429 = ~1'b0 ;
  assign y11430 = ~1'b0 ;
  assign y11431 = ~n25375 ;
  assign y11432 = ~n25378 ;
  assign y11433 = n25380 ;
  assign y11434 = ~n25383 ;
  assign y11435 = n25390 ;
  assign y11436 = n25392 ;
  assign y11437 = ~n25393 ;
  assign y11438 = ~1'b0 ;
  assign y11439 = n25394 ;
  assign y11440 = n25403 ;
  assign y11441 = ~1'b0 ;
  assign y11442 = ~1'b0 ;
  assign y11443 = n25405 ;
  assign y11444 = n25410 ;
  assign y11445 = ~1'b0 ;
  assign y11446 = ~1'b0 ;
  assign y11447 = ~n25413 ;
  assign y11448 = n25416 ;
  assign y11449 = n25423 ;
  assign y11450 = n25425 ;
  assign y11451 = n25427 ;
  assign y11452 = n25428 ;
  assign y11453 = n2122 ;
  assign y11454 = ~n25432 ;
  assign y11455 = n25433 ;
  assign y11456 = ~1'b0 ;
  assign y11457 = ~n25435 ;
  assign y11458 = ~1'b0 ;
  assign y11459 = ~n25436 ;
  assign y11460 = n25441 ;
  assign y11461 = ~n13815 ;
  assign y11462 = n25442 ;
  assign y11463 = n25443 ;
  assign y11464 = ~1'b0 ;
  assign y11465 = ~1'b0 ;
  assign y11466 = ~1'b0 ;
  assign y11467 = n25444 ;
  assign y11468 = n25447 ;
  assign y11469 = ~1'b0 ;
  assign y11470 = ~n25449 ;
  assign y11471 = ~n25450 ;
  assign y11472 = n25451 ;
  assign y11473 = n25456 ;
  assign y11474 = ~1'b0 ;
  assign y11475 = ~1'b0 ;
  assign y11476 = n25457 ;
  assign y11477 = ~n25460 ;
  assign y11478 = ~n25466 ;
  assign y11479 = ~1'b0 ;
  assign y11480 = ~1'b0 ;
  assign y11481 = ~n8729 ;
  assign y11482 = 1'b0 ;
  assign y11483 = n25470 ;
  assign y11484 = ~n25473 ;
  assign y11485 = ~n25476 ;
  assign y11486 = ~1'b0 ;
  assign y11487 = ~1'b0 ;
  assign y11488 = ~n25478 ;
  assign y11489 = n25484 ;
  assign y11490 = ~1'b0 ;
  assign y11491 = n25487 ;
  assign y11492 = n25489 ;
  assign y11493 = ~1'b0 ;
  assign y11494 = 1'b0 ;
  assign y11495 = ~n25490 ;
  assign y11496 = n1279 ;
  assign y11497 = n25491 ;
  assign y11498 = ~n25492 ;
  assign y11499 = ~n25494 ;
  assign y11500 = ~n25496 ;
  assign y11501 = ~n25498 ;
  assign y11502 = n20971 ;
  assign y11503 = n25500 ;
  assign y11504 = ~1'b0 ;
  assign y11505 = ~n25501 ;
  assign y11506 = ~n25503 ;
  assign y11507 = ~n25505 ;
  assign y11508 = n2326 ;
  assign y11509 = n25506 ;
  assign y11510 = n25510 ;
  assign y11511 = ~n25513 ;
  assign y11512 = n25515 ;
  assign y11513 = n25517 ;
  assign y11514 = n25524 ;
  assign y11515 = ~1'b0 ;
  assign y11516 = n25525 ;
  assign y11517 = ~1'b0 ;
  assign y11518 = ~n23698 ;
  assign y11519 = ~n25528 ;
  assign y11520 = n25533 ;
  assign y11521 = ~n25534 ;
  assign y11522 = ~n25535 ;
  assign y11523 = ~1'b0 ;
  assign y11524 = n25537 ;
  assign y11525 = n25538 ;
  assign y11526 = ~n25542 ;
  assign y11527 = ~1'b0 ;
  assign y11528 = ~n25544 ;
  assign y11529 = ~1'b0 ;
  assign y11530 = ~1'b0 ;
  assign y11531 = n25546 ;
  assign y11532 = ~1'b0 ;
  assign y11533 = ~n25548 ;
  assign y11534 = n25552 ;
  assign y11535 = n25554 ;
  assign y11536 = n25556 ;
  assign y11537 = n25558 ;
  assign y11538 = n25563 ;
  assign y11539 = n25566 ;
  assign y11540 = ~1'b0 ;
  assign y11541 = ~n25569 ;
  assign y11542 = ~n25570 ;
  assign y11543 = ~1'b0 ;
  assign y11544 = n4422 ;
  assign y11545 = ~n25573 ;
  assign y11546 = n25575 ;
  assign y11547 = ~1'b0 ;
  assign y11548 = ~1'b0 ;
  assign y11549 = n25576 ;
  assign y11550 = ~1'b0 ;
  assign y11551 = ~n25579 ;
  assign y11552 = n25582 ;
  assign y11553 = ~n18702 ;
  assign y11554 = ~1'b0 ;
  assign y11555 = ~n25584 ;
  assign y11556 = ~n10269 ;
  assign y11557 = ~n25585 ;
  assign y11558 = ~n25586 ;
  assign y11559 = n25588 ;
  assign y11560 = ~1'b0 ;
  assign y11561 = ~n25595 ;
  assign y11562 = ~n25598 ;
  assign y11563 = ~1'b0 ;
  assign y11564 = ~n25600 ;
  assign y11565 = ~1'b0 ;
  assign y11566 = ~n25608 ;
  assign y11567 = ~1'b0 ;
  assign y11568 = n25609 ;
  assign y11569 = n25615 ;
  assign y11570 = ~1'b0 ;
  assign y11571 = ~1'b0 ;
  assign y11572 = n25618 ;
  assign y11573 = ~1'b0 ;
  assign y11574 = ~n25621 ;
  assign y11575 = n25629 ;
  assign y11576 = n25638 ;
  assign y11577 = n25639 ;
  assign y11578 = n25641 ;
  assign y11579 = n25646 ;
  assign y11580 = n25650 ;
  assign y11581 = n25651 ;
  assign y11582 = ~n25656 ;
  assign y11583 = n25659 ;
  assign y11584 = ~n25660 ;
  assign y11585 = 1'b0 ;
  assign y11586 = ~1'b0 ;
  assign y11587 = n25661 ;
  assign y11588 = n25666 ;
  assign y11589 = ~1'b0 ;
  assign y11590 = ~n25669 ;
  assign y11591 = ~n21395 ;
  assign y11592 = n25670 ;
  assign y11593 = ~1'b0 ;
  assign y11594 = ~n25672 ;
  assign y11595 = ~n24511 ;
  assign y11596 = ~n25673 ;
  assign y11597 = ~1'b0 ;
  assign y11598 = n25676 ;
  assign y11599 = ~n25677 ;
  assign y11600 = ~1'b0 ;
  assign y11601 = n25682 ;
  assign y11602 = n25684 ;
  assign y11603 = n25687 ;
  assign y11604 = ~n25691 ;
  assign y11605 = ~n25692 ;
  assign y11606 = n25694 ;
  assign y11607 = ~1'b0 ;
  assign y11608 = n1906 ;
  assign y11609 = ~n25696 ;
  assign y11610 = n25697 ;
  assign y11611 = ~1'b0 ;
  assign y11612 = n25700 ;
  assign y11613 = n25702 ;
  assign y11614 = n25709 ;
  assign y11615 = ~n25710 ;
  assign y11616 = ~n25711 ;
  assign y11617 = ~1'b0 ;
  assign y11618 = ~1'b0 ;
  assign y11619 = ~1'b0 ;
  assign y11620 = n25713 ;
  assign y11621 = n25714 ;
  assign y11622 = n25718 ;
  assign y11623 = n25720 ;
  assign y11624 = ~n25722 ;
  assign y11625 = ~n25726 ;
  assign y11626 = ~n25730 ;
  assign y11627 = n25733 ;
  assign y11628 = n25737 ;
  assign y11629 = ~n25738 ;
  assign y11630 = n25743 ;
  assign y11631 = ~n25744 ;
  assign y11632 = n25745 ;
  assign y11633 = ~n25751 ;
  assign y11634 = ~n25752 ;
  assign y11635 = ~n25754 ;
  assign y11636 = ~n25757 ;
  assign y11637 = ~1'b0 ;
  assign y11638 = 1'b0 ;
  assign y11639 = n25762 ;
  assign y11640 = n25764 ;
  assign y11641 = ~n25766 ;
  assign y11642 = n25772 ;
  assign y11643 = ~n11010 ;
  assign y11644 = ~1'b0 ;
  assign y11645 = ~n25773 ;
  assign y11646 = ~1'b0 ;
  assign y11647 = n25774 ;
  assign y11648 = ~n25778 ;
  assign y11649 = n21007 ;
  assign y11650 = n25781 ;
  assign y11651 = ~n25786 ;
  assign y11652 = ~n25793 ;
  assign y11653 = ~n25794 ;
  assign y11654 = ~n25797 ;
  assign y11655 = ~n25798 ;
  assign y11656 = ~n25803 ;
  assign y11657 = ~n25806 ;
  assign y11658 = ~n25808 ;
  assign y11659 = ~n25810 ;
  assign y11660 = n25815 ;
  assign y11661 = ~n25817 ;
  assign y11662 = n25820 ;
  assign y11663 = n25826 ;
  assign y11664 = ~n25831 ;
  assign y11665 = ~n25832 ;
  assign y11666 = ~n25834 ;
  assign y11667 = n25835 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = ~n25841 ;
  assign y11670 = n4908 ;
  assign y11671 = ~n3698 ;
  assign y11672 = n25842 ;
  assign y11673 = ~n25843 ;
  assign y11674 = n8566 ;
  assign y11675 = n25873 ;
  assign y11676 = n25876 ;
  assign y11677 = ~n25879 ;
  assign y11678 = n25880 ;
  assign y11679 = ~1'b0 ;
  assign y11680 = ~n25882 ;
  assign y11681 = ~n25891 ;
  assign y11682 = n25894 ;
  assign y11683 = n25896 ;
  assign y11684 = ~n25898 ;
  assign y11685 = n25902 ;
  assign y11686 = ~n25905 ;
  assign y11687 = ~1'b0 ;
  assign y11688 = ~n25909 ;
  assign y11689 = ~n25914 ;
  assign y11690 = n25918 ;
  assign y11691 = n25923 ;
  assign y11692 = 1'b0 ;
  assign y11693 = ~1'b0 ;
  assign y11694 = n25924 ;
  assign y11695 = ~n25926 ;
  assign y11696 = ~n25929 ;
  assign y11697 = ~1'b0 ;
  assign y11698 = n25930 ;
  assign y11699 = n25931 ;
  assign y11700 = ~n25933 ;
  assign y11701 = ~n25939 ;
  assign y11702 = ~n25940 ;
  assign y11703 = ~1'b0 ;
  assign y11704 = n25943 ;
  assign y11705 = ~n25947 ;
  assign y11706 = ~1'b0 ;
  assign y11707 = ~1'b0 ;
  assign y11708 = n25952 ;
  assign y11709 = n25953 ;
  assign y11710 = ~n25954 ;
  assign y11711 = ~n25957 ;
  assign y11712 = ~n25962 ;
  assign y11713 = n25965 ;
  assign y11714 = ~n25966 ;
  assign y11715 = n25967 ;
  assign y11716 = ~n25969 ;
  assign y11717 = ~n25972 ;
  assign y11718 = ~n25975 ;
  assign y11719 = n14876 ;
  assign y11720 = ~n25978 ;
  assign y11721 = n5053 ;
  assign y11722 = ~n25985 ;
  assign y11723 = ~1'b0 ;
  assign y11724 = ~n25988 ;
  assign y11725 = n25997 ;
  assign y11726 = ~n25999 ;
  assign y11727 = n1487 ;
  assign y11728 = n26002 ;
  assign y11729 = ~n26006 ;
  assign y11730 = n26009 ;
  assign y11731 = ~n26019 ;
  assign y11732 = ~1'b0 ;
  assign y11733 = ~n26021 ;
  assign y11734 = n26025 ;
  assign y11735 = ~1'b0 ;
  assign y11736 = ~n26027 ;
  assign y11737 = n24573 ;
  assign y11738 = ~1'b0 ;
  assign y11739 = ~n26029 ;
  assign y11740 = ~1'b0 ;
  assign y11741 = n26031 ;
  assign y11742 = ~n26032 ;
  assign y11743 = ~n26036 ;
  assign y11744 = ~n26039 ;
  assign y11745 = ~1'b0 ;
  assign y11746 = n26047 ;
  assign y11747 = ~n26050 ;
  assign y11748 = ~1'b0 ;
  assign y11749 = ~1'b0 ;
  assign y11750 = n26057 ;
  assign y11751 = n26059 ;
  assign y11752 = ~n26060 ;
  assign y11753 = n26061 ;
  assign y11754 = ~1'b0 ;
  assign y11755 = n26068 ;
  assign y11756 = ~1'b0 ;
  assign y11757 = n26069 ;
  assign y11758 = n26071 ;
  assign y11759 = ~1'b0 ;
  assign y11760 = ~1'b0 ;
  assign y11761 = ~1'b0 ;
  assign y11762 = n26074 ;
  assign y11763 = ~n26075 ;
  assign y11764 = n26078 ;
  assign y11765 = ~n5119 ;
  assign y11766 = ~n26081 ;
  assign y11767 = ~n26083 ;
  assign y11768 = n26086 ;
  assign y11769 = ~1'b0 ;
  assign y11770 = ~1'b0 ;
  assign y11771 = ~n26087 ;
  assign y11772 = ~n26091 ;
  assign y11773 = ~n26092 ;
  assign y11774 = n26098 ;
  assign y11775 = n26100 ;
  assign y11776 = n26101 ;
  assign y11777 = n26105 ;
  assign y11778 = n13359 ;
  assign y11779 = ~n26106 ;
  assign y11780 = ~1'b0 ;
  assign y11781 = ~n26111 ;
  assign y11782 = n26114 ;
  assign y11783 = ~n26115 ;
  assign y11784 = n1276 ;
  assign y11785 = n26116 ;
  assign y11786 = ~n26118 ;
  assign y11787 = ~n26120 ;
  assign y11788 = ~n26122 ;
  assign y11789 = n26123 ;
  assign y11790 = ~1'b0 ;
  assign y11791 = n26124 ;
  assign y11792 = ~n26125 ;
  assign y11793 = ~n26128 ;
  assign y11794 = n26129 ;
  assign y11795 = n26136 ;
  assign y11796 = ~1'b0 ;
  assign y11797 = ~1'b0 ;
  assign y11798 = ~n26138 ;
  assign y11799 = ~n26139 ;
  assign y11800 = ~n26143 ;
  assign y11801 = ~n25888 ;
  assign y11802 = ~n26146 ;
  assign y11803 = ~n26148 ;
  assign y11804 = ~n26155 ;
  assign y11805 = n26156 ;
  assign y11806 = ~1'b0 ;
  assign y11807 = n26157 ;
  assign y11808 = ~n26158 ;
  assign y11809 = n26161 ;
  assign y11810 = n26166 ;
  assign y11811 = ~n26167 ;
  assign y11812 = n26169 ;
  assign y11813 = ~1'b0 ;
  assign y11814 = n26170 ;
  assign y11815 = ~n26172 ;
  assign y11816 = n8882 ;
  assign y11817 = n26173 ;
  assign y11818 = ~n26178 ;
  assign y11819 = ~1'b0 ;
  assign y11820 = 1'b0 ;
  assign y11821 = ~n26180 ;
  assign y11822 = ~n26181 ;
  assign y11823 = n26184 ;
  assign y11824 = ~n26186 ;
  assign y11825 = ~1'b0 ;
  assign y11826 = n26188 ;
  assign y11827 = n26190 ;
  assign y11828 = ~1'b0 ;
  assign y11829 = n26193 ;
  assign y11830 = ~n26196 ;
  assign y11831 = ~n26198 ;
  assign y11832 = ~1'b0 ;
  assign y11833 = ~1'b0 ;
  assign y11834 = n26200 ;
  assign y11835 = n26201 ;
  assign y11836 = ~n6638 ;
  assign y11837 = ~n26208 ;
  assign y11838 = ~n26209 ;
  assign y11839 = ~1'b0 ;
  assign y11840 = ~n26212 ;
  assign y11841 = n23004 ;
  assign y11842 = ~n26213 ;
  assign y11843 = n26214 ;
  assign y11844 = n26217 ;
  assign y11845 = ~n26223 ;
  assign y11846 = ~n1746 ;
  assign y11847 = ~n26237 ;
  assign y11848 = n26239 ;
  assign y11849 = ~1'b0 ;
  assign y11850 = n26248 ;
  assign y11851 = ~n26250 ;
  assign y11852 = ~n26255 ;
  assign y11853 = ~1'b0 ;
  assign y11854 = ~1'b0 ;
  assign y11855 = ~n26258 ;
  assign y11856 = ~n26264 ;
  assign y11857 = n26269 ;
  assign y11858 = n26273 ;
  assign y11859 = ~n20638 ;
  assign y11860 = n26275 ;
  assign y11861 = n26281 ;
  assign y11862 = ~1'b0 ;
  assign y11863 = ~n26283 ;
  assign y11864 = n26285 ;
  assign y11865 = n26290 ;
  assign y11866 = n26292 ;
  assign y11867 = 1'b0 ;
  assign y11868 = ~n26293 ;
  assign y11869 = ~1'b0 ;
  assign y11870 = ~1'b0 ;
  assign y11871 = ~1'b0 ;
  assign y11872 = ~1'b0 ;
  assign y11873 = n26295 ;
  assign y11874 = n26301 ;
  assign y11875 = ~1'b0 ;
  assign y11876 = ~n26304 ;
  assign y11877 = ~n26308 ;
  assign y11878 = ~n26309 ;
  assign y11879 = ~n26315 ;
  assign y11880 = n26318 ;
  assign y11881 = ~1'b0 ;
  assign y11882 = ~n13003 ;
  assign y11883 = ~n26320 ;
  assign y11884 = n26322 ;
  assign y11885 = ~1'b0 ;
  assign y11886 = ~1'b0 ;
  assign y11887 = ~n26324 ;
  assign y11888 = n26325 ;
  assign y11889 = n26326 ;
  assign y11890 = n26330 ;
  assign y11891 = n26331 ;
  assign y11892 = ~n4060 ;
  assign y11893 = n26332 ;
  assign y11894 = ~1'b0 ;
  assign y11895 = n26333 ;
  assign y11896 = n26336 ;
  assign y11897 = ~n26338 ;
  assign y11898 = ~1'b0 ;
  assign y11899 = n26340 ;
  assign y11900 = ~n26055 ;
  assign y11901 = ~n26341 ;
  assign y11902 = 1'b0 ;
  assign y11903 = ~n26343 ;
  assign y11904 = ~1'b0 ;
  assign y11905 = n26348 ;
  assign y11906 = ~1'b0 ;
  assign y11907 = ~n26349 ;
  assign y11908 = ~n26351 ;
  assign y11909 = n26353 ;
  assign y11910 = n26355 ;
  assign y11911 = n26359 ;
  assign y11912 = ~n26362 ;
  assign y11913 = ~1'b0 ;
  assign y11914 = ~n26370 ;
  assign y11915 = ~n26377 ;
  assign y11916 = ~n26380 ;
  assign y11917 = ~1'b0 ;
  assign y11918 = ~n26381 ;
  assign y11919 = n26383 ;
  assign y11920 = ~1'b0 ;
  assign y11921 = n26385 ;
  assign y11922 = ~n26387 ;
  assign y11923 = ~1'b0 ;
  assign y11924 = n26388 ;
  assign y11925 = ~n26394 ;
  assign y11926 = ~n26396 ;
  assign y11927 = ~n26398 ;
  assign y11928 = ~n26399 ;
  assign y11929 = ~1'b0 ;
  assign y11930 = 1'b0 ;
  assign y11931 = ~n26401 ;
  assign y11932 = ~n26402 ;
  assign y11933 = ~n26405 ;
  assign y11934 = ~1'b0 ;
  assign y11935 = ~1'b0 ;
  assign y11936 = n26414 ;
  assign y11937 = ~n26415 ;
  assign y11938 = n26416 ;
  assign y11939 = ~n26418 ;
  assign y11940 = ~1'b0 ;
  assign y11941 = ~1'b0 ;
  assign y11942 = n26419 ;
  assign y11943 = ~n26420 ;
  assign y11944 = ~n26423 ;
  assign y11945 = n26430 ;
  assign y11946 = ~1'b0 ;
  assign y11947 = ~n26432 ;
  assign y11948 = n26436 ;
  assign y11949 = n26439 ;
  assign y11950 = n24380 ;
  assign y11951 = n26442 ;
  assign y11952 = n9995 ;
  assign y11953 = n26444 ;
  assign y11954 = n26445 ;
  assign y11955 = ~n26452 ;
  assign y11956 = ~n26455 ;
  assign y11957 = ~1'b0 ;
  assign y11958 = ~n26459 ;
  assign y11959 = n26460 ;
  assign y11960 = n26462 ;
  assign y11961 = n26464 ;
  assign y11962 = ~1'b0 ;
  assign y11963 = ~n26468 ;
  assign y11964 = n26470 ;
  assign y11965 = ~n26471 ;
  assign y11966 = n26478 ;
  assign y11967 = ~1'b0 ;
  assign y11968 = ~n26480 ;
  assign y11969 = ~1'b0 ;
  assign y11970 = n26481 ;
  assign y11971 = n26486 ;
  assign y11972 = ~n26488 ;
  assign y11973 = n26491 ;
  assign y11974 = n15046 ;
  assign y11975 = ~1'b0 ;
  assign y11976 = n26493 ;
  assign y11977 = ~n26498 ;
  assign y11978 = n26499 ;
  assign y11979 = ~n26500 ;
  assign y11980 = n26501 ;
  assign y11981 = ~1'b0 ;
  assign y11982 = ~n26502 ;
  assign y11983 = n26503 ;
  assign y11984 = ~n26507 ;
  assign y11985 = ~1'b0 ;
  assign y11986 = ~n26509 ;
  assign y11987 = n26511 ;
  assign y11988 = ~1'b0 ;
  assign y11989 = n26515 ;
  assign y11990 = ~n26516 ;
  assign y11991 = ~1'b0 ;
  assign y11992 = ~n26519 ;
  assign y11993 = n26521 ;
  assign y11994 = ~n26523 ;
  assign y11995 = n26529 ;
  assign y11996 = ~1'b0 ;
  assign y11997 = ~1'b0 ;
  assign y11998 = n26531 ;
  assign y11999 = ~1'b0 ;
  assign y12000 = n26534 ;
  assign y12001 = n26536 ;
  assign y12002 = n26539 ;
  assign y12003 = ~n26541 ;
  assign y12004 = ~n26543 ;
  assign y12005 = n26544 ;
  assign y12006 = ~n26546 ;
  assign y12007 = ~1'b0 ;
  assign y12008 = ~n26549 ;
  assign y12009 = ~n26550 ;
  assign y12010 = ~n26554 ;
  assign y12011 = n26556 ;
  assign y12012 = n26557 ;
  assign y12013 = ~1'b0 ;
  assign y12014 = ~n26559 ;
  assign y12015 = n26560 ;
  assign y12016 = ~n26562 ;
  assign y12017 = ~1'b0 ;
  assign y12018 = n26565 ;
  assign y12019 = ~1'b0 ;
  assign y12020 = ~1'b0 ;
  assign y12021 = n26567 ;
  assign y12022 = ~1'b0 ;
  assign y12023 = n26570 ;
  assign y12024 = n26572 ;
  assign y12025 = ~1'b0 ;
  assign y12026 = ~1'b0 ;
  assign y12027 = ~1'b0 ;
  assign y12028 = ~n4458 ;
  assign y12029 = ~n26574 ;
  assign y12030 = ~n26575 ;
  assign y12031 = ~1'b0 ;
  assign y12032 = ~n26587 ;
  assign y12033 = n2866 ;
  assign y12034 = ~1'b0 ;
  assign y12035 = ~n26590 ;
  assign y12036 = ~n26592 ;
  assign y12037 = n26593 ;
  assign y12038 = ~n26597 ;
  assign y12039 = ~n26602 ;
  assign y12040 = n26605 ;
  assign y12041 = ~1'b0 ;
  assign y12042 = n26607 ;
  assign y12043 = n26610 ;
  assign y12044 = ~n26616 ;
  assign y12045 = n19597 ;
  assign y12046 = ~n26623 ;
  assign y12047 = n26626 ;
  assign y12048 = ~1'b0 ;
  assign y12049 = ~1'b0 ;
  assign y12050 = n26627 ;
  assign y12051 = n26634 ;
  assign y12052 = ~1'b0 ;
  assign y12053 = ~n26636 ;
  assign y12054 = ~1'b0 ;
  assign y12055 = ~n26639 ;
  assign y12056 = ~n26640 ;
  assign y12057 = ~1'b0 ;
  assign y12058 = ~1'b0 ;
  assign y12059 = ~n26644 ;
  assign y12060 = 1'b0 ;
  assign y12061 = ~1'b0 ;
  assign y12062 = ~n26645 ;
  assign y12063 = ~1'b0 ;
  assign y12064 = ~1'b0 ;
  assign y12065 = ~1'b0 ;
  assign y12066 = ~1'b0 ;
  assign y12067 = n26649 ;
  assign y12068 = n26650 ;
  assign y12069 = n26653 ;
  assign y12070 = ~n26655 ;
  assign y12071 = n26656 ;
  assign y12072 = ~1'b0 ;
  assign y12073 = ~n26659 ;
  assign y12074 = ~n26660 ;
  assign y12075 = ~n26663 ;
  assign y12076 = ~n26675 ;
  assign y12077 = ~1'b0 ;
  assign y12078 = n26679 ;
  assign y12079 = ~1'b0 ;
  assign y12080 = ~n26681 ;
  assign y12081 = 1'b0 ;
  assign y12082 = ~n26687 ;
  assign y12083 = ~n26691 ;
  assign y12084 = n26692 ;
  assign y12085 = ~n26695 ;
  assign y12086 = n26697 ;
  assign y12087 = ~1'b0 ;
  assign y12088 = ~n26699 ;
  assign y12089 = n26700 ;
  assign y12090 = ~n3140 ;
  assign y12091 = ~n26702 ;
  assign y12092 = ~1'b0 ;
  assign y12093 = n26704 ;
  assign y12094 = ~n26707 ;
  assign y12095 = n26723 ;
  assign y12096 = ~n26728 ;
  assign y12097 = ~n26730 ;
  assign y12098 = n22534 ;
  assign y12099 = ~n26735 ;
  assign y12100 = ~n26736 ;
  assign y12101 = ~1'b0 ;
  assign y12102 = ~1'b0 ;
  assign y12103 = n26743 ;
  assign y12104 = n26745 ;
  assign y12105 = ~n26747 ;
  assign y12106 = ~1'b0 ;
  assign y12107 = ~n26752 ;
  assign y12108 = ~n26755 ;
  assign y12109 = n26757 ;
  assign y12110 = n26758 ;
  assign y12111 = ~n26761 ;
  assign y12112 = ~1'b0 ;
  assign y12113 = ~n18459 ;
  assign y12114 = n16828 ;
  assign y12115 = n26763 ;
  assign y12116 = ~1'b0 ;
  assign y12117 = n6546 ;
  assign y12118 = ~1'b0 ;
  assign y12119 = ~1'b0 ;
  assign y12120 = ~n26764 ;
  assign y12121 = n26765 ;
  assign y12122 = ~n26769 ;
  assign y12123 = n26770 ;
  assign y12124 = n26772 ;
  assign y12125 = n26774 ;
  assign y12126 = ~1'b0 ;
  assign y12127 = n26780 ;
  assign y12128 = n26784 ;
  assign y12129 = ~n26788 ;
  assign y12130 = ~1'b0 ;
  assign y12131 = n26791 ;
  assign y12132 = n26793 ;
  assign y12133 = n26794 ;
  assign y12134 = ~n26796 ;
  assign y12135 = ~n26799 ;
  assign y12136 = ~1'b0 ;
  assign y12137 = ~1'b0 ;
  assign y12138 = ~n26800 ;
  assign y12139 = ~n26803 ;
  assign y12140 = ~1'b0 ;
  assign y12141 = ~n26806 ;
  assign y12142 = ~n26807 ;
  assign y12143 = n26813 ;
  assign y12144 = ~n26817 ;
  assign y12145 = ~1'b0 ;
  assign y12146 = n26818 ;
  assign y12147 = ~1'b0 ;
  assign y12148 = ~n26824 ;
  assign y12149 = n26829 ;
  assign y12150 = ~n26832 ;
  assign y12151 = 1'b0 ;
  assign y12152 = ~n26834 ;
  assign y12153 = ~1'b0 ;
  assign y12154 = ~n26839 ;
  assign y12155 = ~n26843 ;
  assign y12156 = n26847 ;
  assign y12157 = n26855 ;
  assign y12158 = ~n26858 ;
  assign y12159 = ~n26862 ;
  assign y12160 = ~1'b0 ;
  assign y12161 = n26865 ;
  assign y12162 = ~n26866 ;
  assign y12163 = n13739 ;
  assign y12164 = ~n26870 ;
  assign y12165 = n9124 ;
  assign y12166 = n26871 ;
  assign y12167 = ~n26873 ;
  assign y12168 = ~1'b0 ;
  assign y12169 = ~1'b0 ;
  assign y12170 = n26874 ;
  assign y12171 = ~1'b0 ;
  assign y12172 = ~1'b0 ;
  assign y12173 = ~n26876 ;
  assign y12174 = ~n14227 ;
  assign y12175 = n26877 ;
  assign y12176 = ~n26883 ;
  assign y12177 = ~1'b0 ;
  assign y12178 = ~n98 ;
  assign y12179 = n11753 ;
  assign y12180 = ~n26885 ;
  assign y12181 = ~n26887 ;
  assign y12182 = ~n18014 ;
  assign y12183 = ~n26889 ;
  assign y12184 = n26907 ;
  assign y12185 = ~1'b0 ;
  assign y12186 = ~n26908 ;
  assign y12187 = n26915 ;
  assign y12188 = ~1'b0 ;
  assign y12189 = n26918 ;
  assign y12190 = n26919 ;
  assign y12191 = n26922 ;
  assign y12192 = ~n26925 ;
  assign y12193 = n26927 ;
  assign y12194 = n26928 ;
  assign y12195 = ~1'b0 ;
  assign y12196 = ~n26931 ;
  assign y12197 = ~1'b0 ;
  assign y12198 = ~1'b0 ;
  assign y12199 = n26933 ;
  assign y12200 = ~n26935 ;
  assign y12201 = n26936 ;
  assign y12202 = n26937 ;
  assign y12203 = 1'b0 ;
  assign y12204 = 1'b0 ;
  assign y12205 = ~1'b0 ;
  assign y12206 = ~1'b0 ;
  assign y12207 = n26926 ;
  assign y12208 = ~1'b0 ;
  assign y12209 = ~1'b0 ;
  assign y12210 = ~n26938 ;
  assign y12211 = n26939 ;
  assign y12212 = n26943 ;
  assign y12213 = ~n26948 ;
  assign y12214 = n26949 ;
  assign y12215 = n26952 ;
  assign y12216 = n26954 ;
  assign y12217 = ~n26955 ;
  assign y12218 = n26958 ;
  assign y12219 = n26960 ;
  assign y12220 = n26962 ;
  assign y12221 = ~1'b0 ;
  assign y12222 = n26964 ;
  assign y12223 = ~n26965 ;
  assign y12224 = ~n26968 ;
  assign y12225 = ~1'b0 ;
  assign y12226 = ~n26969 ;
  assign y12227 = n26970 ;
  assign y12228 = ~n26974 ;
  assign y12229 = ~1'b0 ;
  assign y12230 = ~n26985 ;
  assign y12231 = ~n26987 ;
  assign y12232 = n26988 ;
  assign y12233 = ~1'b0 ;
  assign y12234 = n26991 ;
  assign y12235 = ~n26993 ;
  assign y12236 = ~1'b0 ;
  assign y12237 = ~n27006 ;
  assign y12238 = ~1'b0 ;
  assign y12239 = ~1'b0 ;
  assign y12240 = ~1'b0 ;
  assign y12241 = n27009 ;
  assign y12242 = n27010 ;
  assign y12243 = ~n27012 ;
  assign y12244 = ~1'b0 ;
  assign y12245 = ~n27013 ;
  assign y12246 = ~1'b0 ;
  assign y12247 = ~n27015 ;
  assign y12248 = ~n19510 ;
  assign y12249 = n27026 ;
  assign y12250 = ~1'b0 ;
  assign y12251 = n27027 ;
  assign y12252 = ~1'b0 ;
  assign y12253 = n27028 ;
  assign y12254 = ~n27031 ;
  assign y12255 = ~n27032 ;
  assign y12256 = n27034 ;
  assign y12257 = 1'b0 ;
  assign y12258 = n27036 ;
  assign y12259 = n27038 ;
  assign y12260 = ~1'b0 ;
  assign y12261 = ~1'b0 ;
  assign y12262 = ~n23610 ;
  assign y12263 = ~n27051 ;
  assign y12264 = n4334 ;
  assign y12265 = n27053 ;
  assign y12266 = ~n27055 ;
  assign y12267 = n27057 ;
  assign y12268 = ~n27058 ;
  assign y12269 = ~1'b0 ;
  assign y12270 = ~1'b0 ;
  assign y12271 = ~n27070 ;
  assign y12272 = ~n27082 ;
  assign y12273 = n27084 ;
  assign y12274 = ~1'b0 ;
  assign y12275 = ~1'b0 ;
  assign y12276 = ~1'b0 ;
  assign y12277 = ~n27088 ;
  assign y12278 = n27089 ;
  assign y12279 = n3871 ;
  assign y12280 = ~1'b0 ;
  assign y12281 = ~1'b0 ;
  assign y12282 = ~n27090 ;
  assign y12283 = ~n27091 ;
  assign y12284 = ~n27094 ;
  assign y12285 = n27095 ;
  assign y12286 = ~n27099 ;
  assign y12287 = ~n27102 ;
  assign y12288 = ~1'b0 ;
  assign y12289 = n27113 ;
  assign y12290 = n27115 ;
  assign y12291 = n27126 ;
  assign y12292 = n27129 ;
  assign y12293 = n27131 ;
  assign y12294 = ~n27132 ;
  assign y12295 = ~1'b0 ;
  assign y12296 = ~1'b0 ;
  assign y12297 = n27133 ;
  assign y12298 = ~n27140 ;
  assign y12299 = ~1'b0 ;
  assign y12300 = ~1'b0 ;
  assign y12301 = ~1'b0 ;
  assign y12302 = ~n27144 ;
  assign y12303 = ~n27146 ;
  assign y12304 = ~1'b0 ;
  assign y12305 = ~n27148 ;
  assign y12306 = ~n27151 ;
  assign y12307 = n27152 ;
  assign y12308 = n27154 ;
  assign y12309 = ~n27158 ;
  assign y12310 = ~1'b0 ;
  assign y12311 = ~1'b0 ;
  assign y12312 = ~1'b0 ;
  assign y12313 = n27160 ;
  assign y12314 = n27162 ;
  assign y12315 = ~1'b0 ;
  assign y12316 = n27164 ;
  assign y12317 = ~1'b0 ;
  assign y12318 = ~1'b0 ;
  assign y12319 = ~n27169 ;
  assign y12320 = n27173 ;
  assign y12321 = ~1'b0 ;
  assign y12322 = ~1'b0 ;
  assign y12323 = ~n27175 ;
  assign y12324 = ~n20290 ;
  assign y12325 = ~n27184 ;
  assign y12326 = n27189 ;
  assign y12327 = n27192 ;
  assign y12328 = ~n27194 ;
  assign y12329 = ~1'b0 ;
  assign y12330 = ~n27196 ;
  assign y12331 = ~1'b0 ;
  assign y12332 = ~1'b0 ;
  assign y12333 = n27198 ;
  assign y12334 = ~n27201 ;
  assign y12335 = ~n27202 ;
  assign y12336 = n27206 ;
  assign y12337 = n27211 ;
  assign y12338 = ~1'b0 ;
  assign y12339 = ~n27213 ;
  assign y12340 = ~1'b0 ;
  assign y12341 = n27214 ;
  assign y12342 = n27219 ;
  assign y12343 = ~n27228 ;
  assign y12344 = ~n27231 ;
  assign y12345 = n27232 ;
  assign y12346 = ~n27235 ;
  assign y12347 = ~n27239 ;
  assign y12348 = ~n27242 ;
  assign y12349 = ~n27243 ;
  assign y12350 = ~1'b0 ;
  assign y12351 = ~n27244 ;
  assign y12352 = n27246 ;
  assign y12353 = ~1'b0 ;
  assign y12354 = n27249 ;
  assign y12355 = ~n27251 ;
  assign y12356 = ~n27252 ;
  assign y12357 = n27256 ;
  assign y12358 = ~n27257 ;
  assign y12359 = ~n27258 ;
  assign y12360 = ~1'b0 ;
  assign y12361 = ~1'b0 ;
  assign y12362 = n23483 ;
  assign y12363 = n27259 ;
  assign y12364 = ~1'b0 ;
  assign y12365 = ~1'b0 ;
  assign y12366 = n27264 ;
  assign y12367 = n24330 ;
  assign y12368 = ~n27269 ;
  assign y12369 = ~1'b0 ;
  assign y12370 = ~1'b0 ;
  assign y12371 = n27275 ;
  assign y12372 = ~n27279 ;
  assign y12373 = ~n27282 ;
  assign y12374 = ~1'b0 ;
  assign y12375 = n27283 ;
  assign y12376 = ~1'b0 ;
  assign y12377 = ~n27285 ;
  assign y12378 = n27286 ;
  assign y12379 = ~n27287 ;
  assign y12380 = ~1'b0 ;
  assign y12381 = ~n27290 ;
  assign y12382 = ~n27294 ;
  assign y12383 = n27298 ;
  assign y12384 = ~n27299 ;
  assign y12385 = ~n27301 ;
  assign y12386 = ~1'b0 ;
  assign y12387 = ~1'b0 ;
  assign y12388 = n27302 ;
  assign y12389 = n27308 ;
  assign y12390 = ~1'b0 ;
  assign y12391 = ~1'b0 ;
  assign y12392 = n27313 ;
  assign y12393 = ~1'b0 ;
  assign y12394 = n27314 ;
  assign y12395 = ~n27315 ;
  assign y12396 = n27316 ;
  assign y12397 = ~n27318 ;
  assign y12398 = ~1'b0 ;
  assign y12399 = ~n27319 ;
  assign y12400 = n27330 ;
  assign y12401 = ~1'b0 ;
  assign y12402 = ~n27337 ;
  assign y12403 = ~1'b0 ;
  assign y12404 = n27338 ;
  assign y12405 = ~1'b0 ;
  assign y12406 = n27345 ;
  assign y12407 = ~n27350 ;
  assign y12408 = n27354 ;
  assign y12409 = ~n27355 ;
  assign y12410 = ~n27357 ;
  assign y12411 = n27358 ;
  assign y12412 = ~n27361 ;
  assign y12413 = ~n27367 ;
  assign y12414 = ~n27369 ;
  assign y12415 = n27371 ;
  assign y12416 = n27381 ;
  assign y12417 = ~1'b0 ;
  assign y12418 = ~n27384 ;
  assign y12419 = n27392 ;
  assign y12420 = ~n27395 ;
  assign y12421 = n27397 ;
  assign y12422 = ~1'b0 ;
  assign y12423 = ~1'b0 ;
  assign y12424 = ~n27399 ;
  assign y12425 = ~n27400 ;
  assign y12426 = n27411 ;
  assign y12427 = ~1'b0 ;
  assign y12428 = n27413 ;
  assign y12429 = ~n27414 ;
  assign y12430 = n27417 ;
  assign y12431 = ~1'b0 ;
  assign y12432 = ~n27421 ;
  assign y12433 = ~n27423 ;
  assign y12434 = 1'b0 ;
  assign y12435 = ~1'b0 ;
  assign y12436 = ~1'b0 ;
  assign y12437 = ~1'b0 ;
  assign y12438 = n27424 ;
  assign y12439 = ~n27425 ;
  assign y12440 = n27426 ;
  assign y12441 = ~n27428 ;
  assign y12442 = ~n27431 ;
  assign y12443 = ~n27433 ;
  assign y12444 = ~n27435 ;
  assign y12445 = ~n27438 ;
  assign y12446 = ~n27441 ;
  assign y12447 = n27442 ;
  assign y12448 = ~1'b0 ;
  assign y12449 = ~n27443 ;
  assign y12450 = n27445 ;
  assign y12451 = ~n27447 ;
  assign y12452 = n27448 ;
  assign y12453 = ~1'b0 ;
  assign y12454 = 1'b0 ;
  assign y12455 = ~1'b0 ;
  assign y12456 = ~n27451 ;
  assign y12457 = n27456 ;
  assign y12458 = ~n3879 ;
  assign y12459 = n27458 ;
  assign y12460 = ~n27459 ;
  assign y12461 = n27460 ;
  assign y12462 = ~n27461 ;
  assign y12463 = ~1'b0 ;
  assign y12464 = ~n27463 ;
  assign y12465 = n27467 ;
  assign y12466 = n27478 ;
  assign y12467 = ~1'b0 ;
  assign y12468 = ~n27481 ;
  assign y12469 = n27484 ;
  assign y12470 = n27486 ;
  assign y12471 = ~n27488 ;
  assign y12472 = ~n26365 ;
  assign y12473 = n27489 ;
  assign y12474 = n27491 ;
  assign y12475 = ~n27496 ;
  assign y12476 = ~n27497 ;
  assign y12477 = n27498 ;
  assign y12478 = ~n27503 ;
  assign y12479 = ~n27508 ;
  assign y12480 = ~n27509 ;
  assign y12481 = ~1'b0 ;
  assign y12482 = ~1'b0 ;
  assign y12483 = ~n27512 ;
  assign y12484 = n27517 ;
  assign y12485 = n2695 ;
  assign y12486 = ~n27519 ;
  assign y12487 = ~1'b0 ;
  assign y12488 = ~1'b0 ;
  assign y12489 = ~n27523 ;
  assign y12490 = ~1'b0 ;
  assign y12491 = ~n27529 ;
  assign y12492 = n27530 ;
  assign y12493 = ~1'b0 ;
  assign y12494 = n27532 ;
  assign y12495 = n27534 ;
  assign y12496 = n12292 ;
  assign y12497 = ~n27538 ;
  assign y12498 = ~n27542 ;
  assign y12499 = ~n27547 ;
  assign y12500 = ~n27549 ;
  assign y12501 = ~1'b0 ;
  assign y12502 = ~1'b0 ;
  assign y12503 = ~n27550 ;
  assign y12504 = ~n27551 ;
  assign y12505 = ~n27555 ;
  assign y12506 = 1'b0 ;
  assign y12507 = n27556 ;
  assign y12508 = n27559 ;
  assign y12509 = ~1'b0 ;
  assign y12510 = ~n27568 ;
  assign y12511 = n27570 ;
  assign y12512 = n27572 ;
  assign y12513 = n27578 ;
  assign y12514 = ~n27580 ;
  assign y12515 = n27583 ;
  assign y12516 = ~1'b0 ;
  assign y12517 = n27586 ;
  assign y12518 = n27588 ;
  assign y12519 = ~1'b0 ;
  assign y12520 = ~1'b0 ;
  assign y12521 = ~1'b0 ;
  assign y12522 = ~1'b0 ;
  assign y12523 = n27590 ;
  assign y12524 = n27591 ;
  assign y12525 = ~n27593 ;
  assign y12526 = ~1'b0 ;
  assign y12527 = n27598 ;
  assign y12528 = ~n27600 ;
  assign y12529 = ~n27601 ;
  assign y12530 = ~1'b0 ;
  assign y12531 = ~n27602 ;
  assign y12532 = ~n27604 ;
  assign y12533 = n18928 ;
  assign y12534 = ~n27606 ;
  assign y12535 = ~n27610 ;
  assign y12536 = ~n27613 ;
  assign y12537 = ~n27615 ;
  assign y12538 = n27617 ;
  assign y12539 = n27618 ;
  assign y12540 = n27620 ;
  assign y12541 = n27623 ;
  assign y12542 = ~n16267 ;
  assign y12543 = ~1'b0 ;
  assign y12544 = ~n27625 ;
  assign y12545 = ~1'b0 ;
  assign y12546 = ~n27630 ;
  assign y12547 = ~n27632 ;
  assign y12548 = ~1'b0 ;
  assign y12549 = ~1'b0 ;
  assign y12550 = ~n27636 ;
  assign y12551 = ~1'b0 ;
  assign y12552 = n27637 ;
  assign y12553 = ~n27640 ;
  assign y12554 = ~1'b0 ;
  assign y12555 = ~1'b0 ;
  assign y12556 = ~n27644 ;
  assign y12557 = n27648 ;
  assign y12558 = n27653 ;
  assign y12559 = ~n27654 ;
  assign y12560 = ~1'b0 ;
  assign y12561 = n27655 ;
  assign y12562 = n27656 ;
  assign y12563 = ~1'b0 ;
  assign y12564 = ~n27657 ;
  assign y12565 = ~1'b0 ;
  assign y12566 = ~n27662 ;
  assign y12567 = ~n27664 ;
  assign y12568 = ~1'b0 ;
  assign y12569 = n27668 ;
  assign y12570 = ~n27677 ;
  assign y12571 = ~n27678 ;
  assign y12572 = ~n27679 ;
  assign y12573 = n27680 ;
  assign y12574 = n27681 ;
  assign y12575 = ~1'b0 ;
  assign y12576 = ~n27682 ;
  assign y12577 = ~1'b0 ;
  assign y12578 = ~n27683 ;
  assign y12579 = n27684 ;
  assign y12580 = n27695 ;
  assign y12581 = ~n27697 ;
  assign y12582 = ~n27701 ;
  assign y12583 = ~1'b0 ;
  assign y12584 = ~n27722 ;
  assign y12585 = n27724 ;
  assign y12586 = n27727 ;
  assign y12587 = ~n27730 ;
  assign y12588 = ~n27733 ;
  assign y12589 = n27735 ;
  assign y12590 = ~1'b0 ;
  assign y12591 = ~1'b0 ;
  assign y12592 = ~n27738 ;
  assign y12593 = n27740 ;
  assign y12594 = n27744 ;
  assign y12595 = n27745 ;
  assign y12596 = ~n27746 ;
  assign y12597 = ~n26845 ;
  assign y12598 = ~n27747 ;
  assign y12599 = ~1'b0 ;
  assign y12600 = 1'b0 ;
  assign y12601 = ~n27748 ;
  assign y12602 = ~n27751 ;
  assign y12603 = n27756 ;
  assign y12604 = ~1'b0 ;
  assign y12605 = ~n27761 ;
  assign y12606 = ~1'b0 ;
  assign y12607 = ~1'b0 ;
  assign y12608 = n27762 ;
  assign y12609 = ~n27764 ;
  assign y12610 = n27768 ;
  assign y12611 = ~n27772 ;
  assign y12612 = ~1'b0 ;
  assign y12613 = ~n27774 ;
  assign y12614 = n27775 ;
  assign y12615 = n27776 ;
  assign y12616 = n27777 ;
  assign y12617 = ~n27778 ;
  assign y12618 = n27780 ;
  assign y12619 = 1'b0 ;
  assign y12620 = n27785 ;
  assign y12621 = ~1'b0 ;
  assign y12622 = n37 ;
  assign y12623 = ~n27794 ;
  assign y12624 = ~1'b0 ;
  assign y12625 = ~n27798 ;
  assign y12626 = ~n5708 ;
  assign y12627 = ~n27801 ;
  assign y12628 = ~n7078 ;
  assign y12629 = ~1'b0 ;
  assign y12630 = n27803 ;
  assign y12631 = ~n27812 ;
  assign y12632 = n27813 ;
  assign y12633 = n27820 ;
  assign y12634 = ~n27821 ;
  assign y12635 = n27822 ;
  assign y12636 = ~1'b0 ;
  assign y12637 = ~1'b0 ;
  assign y12638 = n27828 ;
  assign y12639 = ~n27831 ;
  assign y12640 = ~n27833 ;
  assign y12641 = n27836 ;
  assign y12642 = ~n27843 ;
  assign y12643 = ~n27844 ;
  assign y12644 = ~1'b0 ;
  assign y12645 = ~n27847 ;
  assign y12646 = ~n27849 ;
  assign y12647 = ~n27854 ;
  assign y12648 = ~n27857 ;
  assign y12649 = ~1'b0 ;
  assign y12650 = ~1'b0 ;
  assign y12651 = ~1'b0 ;
  assign y12652 = n27858 ;
  assign y12653 = 1'b0 ;
  assign y12654 = ~1'b0 ;
  assign y12655 = ~n27859 ;
  assign y12656 = n27862 ;
  assign y12657 = n23987 ;
  assign y12658 = ~n27863 ;
  assign y12659 = n27866 ;
  assign y12660 = 1'b0 ;
  assign y12661 = ~1'b0 ;
  assign y12662 = n27869 ;
  assign y12663 = ~n27873 ;
  assign y12664 = ~n27876 ;
  assign y12665 = n21266 ;
  assign y12666 = ~1'b0 ;
  assign y12667 = ~n27882 ;
  assign y12668 = n27886 ;
  assign y12669 = ~1'b0 ;
  assign y12670 = n27890 ;
  assign y12671 = ~1'b0 ;
  assign y12672 = ~1'b0 ;
  assign y12673 = ~1'b0 ;
  assign y12674 = 1'b0 ;
  assign y12675 = ~n27891 ;
  assign y12676 = n27892 ;
  assign y12677 = n27893 ;
  assign y12678 = n27894 ;
  assign y12679 = ~1'b0 ;
  assign y12680 = ~1'b0 ;
  assign y12681 = n27900 ;
  assign y12682 = n27906 ;
  assign y12683 = ~n27907 ;
  assign y12684 = n27908 ;
  assign y12685 = n27909 ;
  assign y12686 = ~n27910 ;
  assign y12687 = n27914 ;
  assign y12688 = n27918 ;
  assign y12689 = ~n27921 ;
  assign y12690 = ~n27922 ;
  assign y12691 = ~n27925 ;
  assign y12692 = n27926 ;
  assign y12693 = n27928 ;
  assign y12694 = n27933 ;
  assign y12695 = ~n27938 ;
  assign y12696 = ~1'b0 ;
  assign y12697 = n27940 ;
  assign y12698 = ~1'b0 ;
  assign y12699 = ~1'b0 ;
  assign y12700 = ~1'b0 ;
  assign y12701 = ~n27948 ;
  assign y12702 = n27956 ;
  assign y12703 = ~1'b0 ;
  assign y12704 = ~n27958 ;
  assign y12705 = ~1'b0 ;
  assign y12706 = ~n27960 ;
  assign y12707 = n27962 ;
  assign y12708 = n27963 ;
  assign y12709 = ~1'b0 ;
  assign y12710 = n27966 ;
  assign y12711 = ~1'b0 ;
  assign y12712 = ~n27970 ;
  assign y12713 = ~n27974 ;
  assign y12714 = ~1'b0 ;
  assign y12715 = n12928 ;
  assign y12716 = n27977 ;
  assign y12717 = ~n27978 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = n27986 ;
  assign y12720 = ~1'b0 ;
  assign y12721 = ~n27987 ;
  assign y12722 = n5649 ;
  assign y12723 = ~n27995 ;
  assign y12724 = n27997 ;
  assign y12725 = n28004 ;
  assign y12726 = ~n25707 ;
  assign y12727 = n28007 ;
  assign y12728 = n28009 ;
  assign y12729 = ~n28010 ;
  assign y12730 = ~1'b0 ;
  assign y12731 = ~n28012 ;
  assign y12732 = n2644 ;
  assign y12733 = ~1'b0 ;
  assign y12734 = ~1'b0 ;
  assign y12735 = n28013 ;
  assign y12736 = n28016 ;
  assign y12737 = ~1'b0 ;
  assign y12738 = ~n1723 ;
  assign y12739 = ~n28018 ;
  assign y12740 = n11459 ;
  assign y12741 = n28028 ;
  assign y12742 = ~1'b0 ;
  assign y12743 = ~n28030 ;
  assign y12744 = n28034 ;
  assign y12745 = n28040 ;
  assign y12746 = n28046 ;
  assign y12747 = ~1'b0 ;
  assign y12748 = n28051 ;
  assign y12749 = ~1'b0 ;
  assign y12750 = n28053 ;
  assign y12751 = n28054 ;
  assign y12752 = ~1'b0 ;
  assign y12753 = 1'b0 ;
  assign y12754 = ~1'b0 ;
  assign y12755 = ~n28056 ;
  assign y12756 = ~1'b0 ;
  assign y12757 = ~n28059 ;
  assign y12758 = n28060 ;
  assign y12759 = n28064 ;
  assign y12760 = ~n16001 ;
  assign y12761 = n28065 ;
  assign y12762 = ~1'b0 ;
  assign y12763 = n28072 ;
  assign y12764 = ~n28073 ;
  assign y12765 = ~n28075 ;
  assign y12766 = ~1'b0 ;
  assign y12767 = ~1'b0 ;
  assign y12768 = ~n28080 ;
  assign y12769 = ~1'b0 ;
  assign y12770 = ~n28089 ;
  assign y12771 = ~n28095 ;
  assign y12772 = ~n28098 ;
  assign y12773 = n28099 ;
  assign y12774 = ~1'b0 ;
  assign y12775 = n28101 ;
  assign y12776 = ~n28103 ;
  assign y12777 = n28105 ;
  assign y12778 = n28109 ;
  assign y12779 = ~1'b0 ;
  assign y12780 = n28112 ;
  assign y12781 = n28116 ;
  assign y12782 = ~n28117 ;
  assign y12783 = ~n28119 ;
  assign y12784 = ~n28121 ;
  assign y12785 = n28122 ;
  assign y12786 = n28125 ;
  assign y12787 = n28126 ;
  assign y12788 = n28131 ;
  assign y12789 = ~n28133 ;
  assign y12790 = n28135 ;
  assign y12791 = n28136 ;
  assign y12792 = ~n28141 ;
  assign y12793 = n28145 ;
  assign y12794 = ~1'b0 ;
  assign y12795 = ~n28146 ;
  assign y12796 = n28150 ;
  assign y12797 = ~1'b0 ;
  assign y12798 = ~1'b0 ;
  assign y12799 = ~1'b0 ;
  assign y12800 = ~1'b0 ;
  assign y12801 = n28151 ;
  assign y12802 = ~n28154 ;
  assign y12803 = ~n28156 ;
  assign y12804 = ~n28157 ;
  assign y12805 = ~n28159 ;
  assign y12806 = n28165 ;
  assign y12807 = n28169 ;
  assign y12808 = n17692 ;
  assign y12809 = ~n28170 ;
  assign y12810 = ~n28171 ;
  assign y12811 = ~1'b0 ;
  assign y12812 = n28175 ;
  assign y12813 = ~1'b0 ;
  assign y12814 = ~1'b0 ;
  assign y12815 = ~n28176 ;
  assign y12816 = n28178 ;
  assign y12817 = ~n28180 ;
  assign y12818 = ~n28183 ;
  assign y12819 = ~n28187 ;
  assign y12820 = n28190 ;
  assign y12821 = n28193 ;
  assign y12822 = ~n28197 ;
  assign y12823 = ~n28202 ;
  assign y12824 = ~n28204 ;
  assign y12825 = ~1'b0 ;
  assign y12826 = n28208 ;
  assign y12827 = ~1'b0 ;
  assign y12828 = n28211 ;
  assign y12829 = ~1'b0 ;
  assign y12830 = n28216 ;
  assign y12831 = ~1'b0 ;
  assign y12832 = n28217 ;
  assign y12833 = n28219 ;
  assign y12834 = ~1'b0 ;
  assign y12835 = ~1'b0 ;
  assign y12836 = ~n28221 ;
  assign y12837 = ~n28225 ;
  assign y12838 = ~n10641 ;
  assign y12839 = ~1'b0 ;
  assign y12840 = ~1'b0 ;
  assign y12841 = ~n28227 ;
  assign y12842 = ~n28233 ;
  assign y12843 = ~n23227 ;
  assign y12844 = ~1'b0 ;
  assign y12845 = ~n28234 ;
  assign y12846 = n28238 ;
  assign y12847 = ~1'b0 ;
  assign y12848 = ~n28240 ;
  assign y12849 = ~1'b0 ;
  assign y12850 = ~1'b0 ;
  assign y12851 = n28241 ;
  assign y12852 = n11573 ;
  assign y12853 = ~n28244 ;
  assign y12854 = ~n28245 ;
  assign y12855 = n28246 ;
  assign y12856 = ~n28247 ;
  assign y12857 = ~n28248 ;
  assign y12858 = ~n28251 ;
  assign y12859 = ~n17245 ;
  assign y12860 = n28253 ;
  assign y12861 = ~1'b0 ;
  assign y12862 = ~n28259 ;
  assign y12863 = n28261 ;
  assign y12864 = n26596 ;
  assign y12865 = ~n28262 ;
  assign y12866 = ~1'b0 ;
  assign y12867 = ~n28265 ;
  assign y12868 = ~1'b0 ;
  assign y12869 = ~n16210 ;
  assign y12870 = ~1'b0 ;
  assign y12871 = ~n28267 ;
  assign y12872 = n28269 ;
  assign y12873 = ~n13449 ;
  assign y12874 = ~n28275 ;
  assign y12875 = ~n28277 ;
  assign y12876 = n28278 ;
  assign y12877 = n28285 ;
  assign y12878 = ~1'b0 ;
  assign y12879 = n28286 ;
  assign y12880 = ~n28288 ;
  assign y12881 = n28294 ;
  assign y12882 = n28295 ;
  assign y12883 = n28299 ;
  assign y12884 = ~n28302 ;
  assign y12885 = n28304 ;
  assign y12886 = ~n28312 ;
  assign y12887 = ~1'b0 ;
  assign y12888 = ~1'b0 ;
  assign y12889 = ~1'b0 ;
  assign y12890 = n28314 ;
  assign y12891 = ~1'b0 ;
  assign y12892 = n28318 ;
  assign y12893 = n28319 ;
  assign y12894 = n28320 ;
  assign y12895 = n28325 ;
  assign y12896 = ~n28326 ;
  assign y12897 = n28329 ;
  assign y12898 = ~1'b0 ;
  assign y12899 = n28332 ;
  assign y12900 = ~n28335 ;
  assign y12901 = ~n28336 ;
  assign y12902 = ~n28337 ;
  assign y12903 = ~n28341 ;
  assign y12904 = n28344 ;
  assign y12905 = ~n28348 ;
  assign y12906 = ~n28350 ;
  assign y12907 = ~1'b0 ;
  assign y12908 = n28354 ;
  assign y12909 = ~1'b0 ;
  assign y12910 = n28357 ;
  assign y12911 = n28358 ;
  assign y12912 = n28366 ;
  assign y12913 = ~1'b0 ;
  assign y12914 = ~1'b0 ;
  assign y12915 = ~n28370 ;
  assign y12916 = ~n28371 ;
  assign y12917 = n28374 ;
  assign y12918 = ~n28376 ;
  assign y12919 = ~n28378 ;
  assign y12920 = ~n28380 ;
  assign y12921 = n28381 ;
  assign y12922 = n28382 ;
  assign y12923 = ~n28385 ;
  assign y12924 = n28386 ;
  assign y12925 = n28388 ;
  assign y12926 = ~n28391 ;
  assign y12927 = ~1'b0 ;
  assign y12928 = n17306 ;
  assign y12929 = n28392 ;
  assign y12930 = ~1'b0 ;
  assign y12931 = ~1'b0 ;
  assign y12932 = ~n12530 ;
  assign y12933 = ~n28399 ;
  assign y12934 = ~1'b0 ;
  assign y12935 = ~n28402 ;
  assign y12936 = ~n28405 ;
  assign y12937 = ~1'b0 ;
  assign y12938 = n28407 ;
  assign y12939 = n28408 ;
  assign y12940 = ~n28410 ;
  assign y12941 = n28412 ;
  assign y12942 = ~1'b0 ;
  assign y12943 = ~n28417 ;
  assign y12944 = n28423 ;
  assign y12945 = ~n28424 ;
  assign y12946 = ~1'b0 ;
  assign y12947 = n28431 ;
  assign y12948 = ~n28433 ;
  assign y12949 = ~n28440 ;
  assign y12950 = n28441 ;
  assign y12951 = ~1'b0 ;
  assign y12952 = n28444 ;
  assign y12953 = ~1'b0 ;
  assign y12954 = n28447 ;
  assign y12955 = ~1'b0 ;
  assign y12956 = ~1'b0 ;
  assign y12957 = ~n28450 ;
  assign y12958 = ~n28451 ;
  assign y12959 = n28455 ;
  assign y12960 = ~1'b0 ;
  assign y12961 = n28458 ;
  assign y12962 = n28460 ;
  assign y12963 = ~n28462 ;
  assign y12964 = ~n28465 ;
  assign y12965 = ~1'b0 ;
  assign y12966 = ~n28467 ;
  assign y12967 = n28473 ;
  assign y12968 = ~1'b0 ;
  assign y12969 = ~1'b0 ;
  assign y12970 = ~n7471 ;
  assign y12971 = ~1'b0 ;
  assign y12972 = ~1'b0 ;
  assign y12973 = n28475 ;
  assign y12974 = n28476 ;
  assign y12975 = ~1'b0 ;
  assign y12976 = ~1'b0 ;
  assign y12977 = ~n28481 ;
  assign y12978 = ~n28482 ;
  assign y12979 = n28483 ;
  assign y12980 = n28487 ;
  assign y12981 = ~n28489 ;
  assign y12982 = n28491 ;
  assign y12983 = ~1'b0 ;
  assign y12984 = ~n1276 ;
  assign y12985 = n28494 ;
  assign y12986 = ~n13453 ;
  assign y12987 = n28496 ;
  assign y12988 = ~1'b0 ;
  assign y12989 = ~1'b0 ;
  assign y12990 = ~n28499 ;
  assign y12991 = ~1'b0 ;
  assign y12992 = n28505 ;
  assign y12993 = n28506 ;
  assign y12994 = ~n28508 ;
  assign y12995 = ~1'b0 ;
  assign y12996 = n28514 ;
  assign y12997 = n28515 ;
  assign y12998 = ~1'b0 ;
  assign y12999 = ~1'b0 ;
  assign y13000 = n28517 ;
  assign y13001 = ~n28518 ;
  assign y13002 = ~n28520 ;
  assign y13003 = ~n2060 ;
  assign y13004 = ~n28531 ;
  assign y13005 = n28533 ;
  assign y13006 = ~n16291 ;
  assign y13007 = n28535 ;
  assign y13008 = n28539 ;
  assign y13009 = n28540 ;
  assign y13010 = ~1'b0 ;
  assign y13011 = ~1'b0 ;
  assign y13012 = ~n3569 ;
  assign y13013 = ~n7096 ;
  assign y13014 = ~n25604 ;
  assign y13015 = 1'b0 ;
  assign y13016 = ~1'b0 ;
  assign y13017 = ~n28541 ;
  assign y13018 = n28547 ;
  assign y13019 = ~1'b0 ;
  assign y13020 = ~1'b0 ;
  assign y13021 = n28550 ;
  assign y13022 = ~n28559 ;
  assign y13023 = ~n28560 ;
  assign y13024 = n28561 ;
  assign y13025 = ~n28563 ;
  assign y13026 = ~n28565 ;
  assign y13027 = ~1'b0 ;
  assign y13028 = ~n28568 ;
  assign y13029 = ~n28570 ;
  assign y13030 = ~n28571 ;
  assign y13031 = ~n28574 ;
  assign y13032 = n28578 ;
  assign y13033 = ~n28580 ;
  assign y13034 = n28583 ;
  assign y13035 = ~n9653 ;
  assign y13036 = n28586 ;
  assign y13037 = ~n28590 ;
  assign y13038 = n10950 ;
  assign y13039 = n28593 ;
  assign y13040 = n28594 ;
  assign y13041 = n28598 ;
  assign y13042 = ~n28601 ;
  assign y13043 = ~n28602 ;
  assign y13044 = ~1'b0 ;
  assign y13045 = ~1'b0 ;
  assign y13046 = ~n28609 ;
  assign y13047 = ~1'b0 ;
  assign y13048 = 1'b0 ;
  assign y13049 = ~n28610 ;
  assign y13050 = ~n28612 ;
  assign y13051 = ~n28615 ;
  assign y13052 = n28616 ;
  assign y13053 = ~1'b0 ;
  assign y13054 = ~n28617 ;
  assign y13055 = n28623 ;
  assign y13056 = n28624 ;
  assign y13057 = ~n28625 ;
  assign y13058 = ~n28629 ;
  assign y13059 = ~n3310 ;
  assign y13060 = ~n28633 ;
  assign y13061 = n28638 ;
  assign y13062 = ~n28642 ;
  assign y13063 = ~1'b0 ;
  assign y13064 = ~n28644 ;
  assign y13065 = ~1'b0 ;
  assign y13066 = ~n28648 ;
  assign y13067 = ~n28650 ;
  assign y13068 = ~1'b0 ;
  assign y13069 = ~1'b0 ;
  assign y13070 = ~n28653 ;
  assign y13071 = ~1'b0 ;
  assign y13072 = ~n28657 ;
  assign y13073 = ~1'b0 ;
  assign y13074 = ~1'b0 ;
  assign y13075 = n28658 ;
  assign y13076 = n28660 ;
  assign y13077 = n28662 ;
  assign y13078 = ~n28666 ;
  assign y13079 = ~n28672 ;
  assign y13080 = ~1'b0 ;
  assign y13081 = n28682 ;
  assign y13082 = n28684 ;
  assign y13083 = ~1'b0 ;
  assign y13084 = ~n28685 ;
  assign y13085 = ~1'b0 ;
  assign y13086 = n28689 ;
  assign y13087 = ~n28692 ;
  assign y13088 = ~1'b0 ;
  assign y13089 = ~n28695 ;
  assign y13090 = n28696 ;
  assign y13091 = ~1'b0 ;
  assign y13092 = ~n28698 ;
  assign y13093 = n28701 ;
  assign y13094 = ~n28702 ;
  assign y13095 = n28704 ;
  assign y13096 = n15730 ;
  assign y13097 = n28705 ;
  assign y13098 = ~n28706 ;
  assign y13099 = n28707 ;
  assign y13100 = ~n28708 ;
  assign y13101 = n28711 ;
  assign y13102 = n6426 ;
  assign y13103 = ~n28712 ;
  assign y13104 = ~n28713 ;
  assign y13105 = ~1'b0 ;
  assign y13106 = ~1'b0 ;
  assign y13107 = n28715 ;
  assign y13108 = ~n28719 ;
  assign y13109 = n1166 ;
  assign y13110 = ~n28722 ;
  assign y13111 = n28723 ;
  assign y13112 = ~n28724 ;
  assign y13113 = ~n28731 ;
  assign y13114 = ~1'b0 ;
  assign y13115 = ~1'b0 ;
  assign y13116 = n28733 ;
  assign y13117 = n4620 ;
  assign y13118 = ~n28736 ;
  assign y13119 = ~n28737 ;
  assign y13120 = ~n28738 ;
  assign y13121 = n28740 ;
  assign y13122 = ~1'b0 ;
  assign y13123 = ~1'b0 ;
  assign y13124 = ~1'b0 ;
  assign y13125 = n28744 ;
  assign y13126 = ~1'b0 ;
  assign y13127 = n28745 ;
  assign y13128 = n28748 ;
  assign y13129 = ~n28751 ;
  assign y13130 = n28752 ;
  assign y13131 = ~n28753 ;
  assign y13132 = ~n28755 ;
  assign y13133 = ~n28758 ;
  assign y13134 = n28764 ;
  assign y13135 = n28765 ;
  assign y13136 = ~1'b0 ;
  assign y13137 = n28768 ;
  assign y13138 = 1'b0 ;
  assign y13139 = ~n28771 ;
  assign y13140 = ~n28774 ;
  assign y13141 = ~1'b0 ;
  assign y13142 = n28775 ;
  assign y13143 = ~n2596 ;
  assign y13144 = n28777 ;
  assign y13145 = n12126 ;
  assign y13146 = ~n4602 ;
  assign y13147 = n28779 ;
  assign y13148 = n28787 ;
  assign y13149 = n28788 ;
  assign y13150 = ~1'b0 ;
  assign y13151 = n28789 ;
  assign y13152 = n28792 ;
  assign y13153 = ~n28796 ;
  assign y13154 = ~1'b0 ;
  assign y13155 = n28799 ;
  assign y13156 = n7862 ;
  assign y13157 = n28800 ;
  assign y13158 = n28803 ;
  assign y13159 = ~1'b0 ;
  assign y13160 = ~1'b0 ;
  assign y13161 = ~n28806 ;
  assign y13162 = n21052 ;
  assign y13163 = ~n28814 ;
  assign y13164 = ~n28816 ;
  assign y13165 = n28817 ;
  assign y13166 = 1'b0 ;
  assign y13167 = n28818 ;
  assign y13168 = ~n28821 ;
  assign y13169 = ~n28829 ;
  assign y13170 = ~n28830 ;
  assign y13171 = ~n25103 ;
  assign y13172 = n5337 ;
  assign y13173 = ~1'b0 ;
  assign y13174 = ~n28831 ;
  assign y13175 = ~n28838 ;
  assign y13176 = ~n28839 ;
  assign y13177 = n28840 ;
  assign y13178 = 1'b0 ;
  assign y13179 = ~n5874 ;
  assign y13180 = n28848 ;
  assign y13181 = ~n1370 ;
  assign y13182 = ~n28849 ;
  assign y13183 = ~1'b0 ;
  assign y13184 = ~1'b0 ;
  assign y13185 = ~1'b0 ;
  assign y13186 = ~n28853 ;
  assign y13187 = ~n18780 ;
  assign y13188 = ~n15989 ;
  assign y13189 = n22985 ;
  assign y13190 = n28858 ;
  assign y13191 = n28860 ;
  assign y13192 = ~n28864 ;
  assign y13193 = ~1'b0 ;
  assign y13194 = n7468 ;
  assign y13195 = n28870 ;
  assign y13196 = ~1'b0 ;
  assign y13197 = n28874 ;
  assign y13198 = ~1'b0 ;
  assign y13199 = n28879 ;
  assign y13200 = ~n28880 ;
  assign y13201 = ~1'b0 ;
  assign y13202 = n16232 ;
  assign y13203 = ~n27000 ;
  assign y13204 = n28887 ;
  assign y13205 = ~n28889 ;
  assign y13206 = n28890 ;
  assign y13207 = ~1'b0 ;
  assign y13208 = n28897 ;
  assign y13209 = ~1'b0 ;
  assign y13210 = n28899 ;
  assign y13211 = ~n28902 ;
  assign y13212 = ~n28906 ;
  assign y13213 = n28908 ;
  assign y13214 = ~n28913 ;
  assign y13215 = n28915 ;
  assign y13216 = ~n28917 ;
  assign y13217 = ~n28919 ;
  assign y13218 = n28920 ;
  assign y13219 = n28923 ;
  assign y13220 = ~1'b0 ;
  assign y13221 = n28932 ;
  assign y13222 = 1'b0 ;
  assign y13223 = n28934 ;
  assign y13224 = ~1'b0 ;
  assign y13225 = ~n28936 ;
  assign y13226 = n28937 ;
  assign y13227 = n28938 ;
  assign y13228 = ~n28941 ;
  assign y13229 = ~1'b0 ;
  assign y13230 = ~n28943 ;
  assign y13231 = n10316 ;
  assign y13232 = ~n28945 ;
  assign y13233 = ~n12887 ;
  assign y13234 = ~1'b0 ;
  assign y13235 = ~n28949 ;
  assign y13236 = ~n28953 ;
  assign y13237 = ~n28954 ;
  assign y13238 = n28958 ;
  assign y13239 = ~n28960 ;
  assign y13240 = ~n28962 ;
  assign y13241 = ~n28966 ;
  assign y13242 = ~n28968 ;
  assign y13243 = ~n28969 ;
  assign y13244 = ~1'b0 ;
  assign y13245 = ~1'b0 ;
  assign y13246 = n28973 ;
  assign y13247 = n28567 ;
  assign y13248 = n28975 ;
  assign y13249 = n28976 ;
  assign y13250 = n28980 ;
  assign y13251 = n28981 ;
  assign y13252 = n28982 ;
  assign y13253 = n28989 ;
  assign y13254 = 1'b0 ;
  assign y13255 = ~n28990 ;
  assign y13256 = ~n28992 ;
  assign y13257 = ~1'b0 ;
  assign y13258 = n28995 ;
  assign y13259 = ~1'b0 ;
  assign y13260 = n28996 ;
  assign y13261 = ~n28997 ;
  assign y13262 = ~n28999 ;
  assign y13263 = n29002 ;
  assign y13264 = n29005 ;
  assign y13265 = ~1'b0 ;
  assign y13266 = n29008 ;
  assign y13267 = ~n29012 ;
  assign y13268 = ~n29015 ;
  assign y13269 = n24235 ;
  assign y13270 = n29019 ;
  assign y13271 = n29020 ;
  assign y13272 = ~1'b0 ;
  assign y13273 = ~n19642 ;
  assign y13274 = ~n29021 ;
  assign y13275 = ~n29026 ;
  assign y13276 = ~n29030 ;
  assign y13277 = ~n29031 ;
  assign y13278 = ~n29032 ;
  assign y13279 = ~1'b0 ;
  assign y13280 = ~1'b0 ;
  assign y13281 = n29033 ;
  assign y13282 = ~1'b0 ;
  assign y13283 = ~n29035 ;
  assign y13284 = n29037 ;
  assign y13285 = ~1'b0 ;
  assign y13286 = ~1'b0 ;
  assign y13287 = ~n29042 ;
  assign y13288 = n29045 ;
  assign y13289 = n29046 ;
  assign y13290 = n29049 ;
  assign y13291 = n29050 ;
  assign y13292 = n29052 ;
  assign y13293 = ~n29058 ;
  assign y13294 = n29062 ;
  assign y13295 = ~1'b0 ;
  assign y13296 = ~n29065 ;
  assign y13297 = ~n29070 ;
  assign y13298 = ~n29071 ;
  assign y13299 = n29076 ;
  assign y13300 = n29081 ;
  assign y13301 = ~1'b0 ;
  assign y13302 = ~n29082 ;
  assign y13303 = ~n29085 ;
  assign y13304 = ~n29087 ;
  assign y13305 = ~n29093 ;
  assign y13306 = ~n2088 ;
  assign y13307 = n16407 ;
  assign y13308 = ~n29095 ;
  assign y13309 = ~n29099 ;
  assign y13310 = ~1'b0 ;
  assign y13311 = n7684 ;
  assign y13312 = n29100 ;
  assign y13313 = ~1'b0 ;
  assign y13314 = ~1'b0 ;
  assign y13315 = ~1'b0 ;
  assign y13316 = ~1'b0 ;
  assign y13317 = n29102 ;
  assign y13318 = ~n29104 ;
  assign y13319 = ~n29110 ;
  assign y13320 = ~1'b0 ;
  assign y13321 = n29113 ;
  assign y13322 = ~n29118 ;
  assign y13323 = n29119 ;
  assign y13324 = n29123 ;
  assign y13325 = ~n29125 ;
  assign y13326 = n29130 ;
  assign y13327 = ~n29132 ;
  assign y13328 = n29137 ;
  assign y13329 = ~n29138 ;
  assign y13330 = ~n29140 ;
  assign y13331 = ~n29144 ;
  assign y13332 = n29148 ;
  assign y13333 = n29150 ;
  assign y13334 = n29151 ;
  assign y13335 = ~n29157 ;
  assign y13336 = ~n29158 ;
  assign y13337 = ~1'b0 ;
  assign y13338 = ~n29162 ;
  assign y13339 = ~n29165 ;
  assign y13340 = ~n29167 ;
  assign y13341 = n29168 ;
  assign y13342 = ~1'b0 ;
  assign y13343 = ~n29170 ;
  assign y13344 = ~n29172 ;
  assign y13345 = ~n29179 ;
  assign y13346 = ~1'b0 ;
  assign y13347 = ~1'b0 ;
  assign y13348 = n29181 ;
  assign y13349 = n29186 ;
  assign y13350 = ~n29190 ;
  assign y13351 = ~1'b0 ;
  assign y13352 = ~n29191 ;
  assign y13353 = ~1'b0 ;
  assign y13354 = n29195 ;
  assign y13355 = ~n29196 ;
  assign y13356 = ~n29197 ;
  assign y13357 = ~n29199 ;
  assign y13358 = ~1'b0 ;
  assign y13359 = ~n29202 ;
  assign y13360 = ~n29209 ;
  assign y13361 = ~n7530 ;
  assign y13362 = ~n29211 ;
  assign y13363 = ~n29221 ;
  assign y13364 = ~1'b0 ;
  assign y13365 = ~n29223 ;
  assign y13366 = ~n29231 ;
  assign y13367 = n29233 ;
  assign y13368 = ~n12058 ;
  assign y13369 = n29236 ;
  assign y13370 = ~n29239 ;
  assign y13371 = n29242 ;
  assign y13372 = n29245 ;
  assign y13373 = ~1'b0 ;
  assign y13374 = n29248 ;
  assign y13375 = ~n29249 ;
  assign y13376 = ~1'b0 ;
  assign y13377 = n29250 ;
  assign y13378 = ~n29254 ;
  assign y13379 = ~n26982 ;
  assign y13380 = ~n29259 ;
  assign y13381 = ~1'b0 ;
  assign y13382 = ~n29263 ;
  assign y13383 = ~n29264 ;
  assign y13384 = ~n29270 ;
  assign y13385 = n29272 ;
  assign y13386 = ~x0 ;
  assign y13387 = n29273 ;
  assign y13388 = n29275 ;
  assign y13389 = ~1'b0 ;
  assign y13390 = ~n5212 ;
  assign y13391 = n29278 ;
  assign y13392 = ~n29280 ;
  assign y13393 = n29282 ;
  assign y13394 = ~n29283 ;
  assign y13395 = ~1'b0 ;
  assign y13396 = ~n29286 ;
  assign y13397 = n29291 ;
  assign y13398 = ~n29292 ;
  assign y13399 = ~1'b0 ;
  assign y13400 = ~n29296 ;
  assign y13401 = n29300 ;
  assign y13402 = ~1'b0 ;
  assign y13403 = ~1'b0 ;
  assign y13404 = ~n29304 ;
  assign y13405 = ~n29306 ;
  assign y13406 = n29308 ;
  assign y13407 = n29309 ;
  assign y13408 = ~1'b0 ;
  assign y13409 = ~n29316 ;
  assign y13410 = n29321 ;
  assign y13411 = ~n29322 ;
  assign y13412 = n29324 ;
  assign y13413 = n29325 ;
  assign y13414 = ~n29326 ;
  assign y13415 = ~n29333 ;
  assign y13416 = n29334 ;
  assign y13417 = ~n29339 ;
  assign y13418 = n29344 ;
  assign y13419 = ~n29346 ;
  assign y13420 = ~1'b0 ;
  assign y13421 = ~1'b0 ;
  assign y13422 = n29347 ;
  assign y13423 = n29348 ;
  assign y13424 = n29349 ;
  assign y13425 = ~1'b0 ;
  assign y13426 = ~n29351 ;
  assign y13427 = ~1'b0 ;
  assign y13428 = n29352 ;
  assign y13429 = n29353 ;
  assign y13430 = n29354 ;
  assign y13431 = n29357 ;
  assign y13432 = ~1'b0 ;
  assign y13433 = ~n29360 ;
  assign y13434 = ~1'b0 ;
  assign y13435 = ~n29362 ;
  assign y13436 = ~n29363 ;
  assign y13437 = ~n29364 ;
  assign y13438 = n29366 ;
  assign y13439 = ~1'b0 ;
  assign y13440 = n29369 ;
  assign y13441 = ~n29371 ;
  assign y13442 = ~n29378 ;
  assign y13443 = ~1'b0 ;
  assign y13444 = ~n29380 ;
  assign y13445 = n29381 ;
  assign y13446 = ~1'b0 ;
  assign y13447 = ~1'b0 ;
  assign y13448 = n29383 ;
  assign y13449 = ~n12578 ;
  assign y13450 = n29386 ;
  assign y13451 = ~n29388 ;
  assign y13452 = ~1'b0 ;
  assign y13453 = n29389 ;
  assign y13454 = ~n29390 ;
  assign y13455 = n29391 ;
  assign y13456 = ~1'b0 ;
  assign y13457 = ~1'b0 ;
  assign y13458 = n29396 ;
  assign y13459 = n29398 ;
  assign y13460 = n29400 ;
  assign y13461 = n29404 ;
  assign y13462 = n29405 ;
  assign y13463 = n29406 ;
  assign y13464 = n29407 ;
  assign y13465 = ~n29411 ;
  assign y13466 = ~n29415 ;
  assign y13467 = n29416 ;
  assign y13468 = n10549 ;
  assign y13469 = n29418 ;
  assign y13470 = n29420 ;
  assign y13471 = n29421 ;
  assign y13472 = ~n29424 ;
  assign y13473 = n29426 ;
  assign y13474 = n29427 ;
  assign y13475 = n29430 ;
  assign y13476 = n29431 ;
  assign y13477 = ~1'b0 ;
  assign y13478 = ~n29435 ;
  assign y13479 = ~n29439 ;
  assign y13480 = ~n29443 ;
  assign y13481 = ~n29445 ;
  assign y13482 = n29453 ;
  assign y13483 = ~n29456 ;
  assign y13484 = n29464 ;
  assign y13485 = n29465 ;
  assign y13486 = n29468 ;
  assign y13487 = n29469 ;
  assign y13488 = ~n29471 ;
  assign y13489 = ~1'b0 ;
  assign y13490 = n29472 ;
  assign y13491 = n29473 ;
  assign y13492 = n29475 ;
  assign y13493 = ~1'b0 ;
  assign y13494 = ~n29481 ;
  assign y13495 = ~n29487 ;
  assign y13496 = ~n29488 ;
  assign y13497 = ~n29490 ;
  assign y13498 = ~n29491 ;
  assign y13499 = ~n29494 ;
  assign y13500 = n29495 ;
  assign y13501 = n29496 ;
  assign y13502 = n29499 ;
  assign y13503 = ~1'b0 ;
  assign y13504 = ~n29501 ;
  assign y13505 = n29502 ;
  assign y13506 = ~n29504 ;
  assign y13507 = n26917 ;
  assign y13508 = n29506 ;
  assign y13509 = n29513 ;
  assign y13510 = ~1'b0 ;
  assign y13511 = ~1'b0 ;
  assign y13512 = ~n29518 ;
  assign y13513 = n29519 ;
  assign y13514 = n29521 ;
  assign y13515 = n29522 ;
  assign y13516 = n29525 ;
  assign y13517 = n29529 ;
  assign y13518 = ~1'b0 ;
  assign y13519 = n29532 ;
  assign y13520 = n29534 ;
  assign y13521 = ~n29535 ;
  assign y13522 = n29536 ;
  assign y13523 = n29540 ;
  assign y13524 = n29545 ;
  assign y13525 = ~1'b0 ;
  assign y13526 = ~1'b0 ;
  assign y13527 = ~n29546 ;
  assign y13528 = ~1'b0 ;
  assign y13529 = ~n29550 ;
  assign y13530 = ~n29556 ;
  assign y13531 = ~n29558 ;
  assign y13532 = n29561 ;
  assign y13533 = ~n29564 ;
  assign y13534 = ~n29569 ;
  assign y13535 = ~n29577 ;
  assign y13536 = n29579 ;
  assign y13537 = ~n29581 ;
  assign y13538 = ~n29583 ;
  assign y13539 = ~n29589 ;
  assign y13540 = n4507 ;
  assign y13541 = ~1'b0 ;
  assign y13542 = ~n29590 ;
  assign y13543 = ~n29591 ;
  assign y13544 = ~n29597 ;
  assign y13545 = ~n29602 ;
  assign y13546 = ~n29603 ;
  assign y13547 = ~1'b0 ;
  assign y13548 = ~1'b0 ;
  assign y13549 = ~n29607 ;
  assign y13550 = ~1'b0 ;
  assign y13551 = ~1'b0 ;
  assign y13552 = ~n29608 ;
  assign y13553 = n29615 ;
  assign y13554 = ~n29619 ;
  assign y13555 = ~n29623 ;
  assign y13556 = ~n29627 ;
  assign y13557 = n29631 ;
  assign y13558 = n29636 ;
  assign y13559 = ~n10044 ;
  assign y13560 = n29637 ;
  assign y13561 = ~n29641 ;
  assign y13562 = ~n29647 ;
  assign y13563 = ~n29648 ;
  assign y13564 = n5511 ;
  assign y13565 = ~n29649 ;
  assign y13566 = 1'b0 ;
  assign y13567 = n29651 ;
  assign y13568 = n29656 ;
  assign y13569 = ~n29663 ;
  assign y13570 = ~1'b0 ;
  assign y13571 = ~1'b0 ;
  assign y13572 = ~1'b0 ;
  assign y13573 = ~n29665 ;
  assign y13574 = ~n29667 ;
  assign y13575 = ~n29669 ;
  assign y13576 = ~1'b0 ;
  assign y13577 = ~n29670 ;
  assign y13578 = ~n29671 ;
  assign y13579 = n29673 ;
  assign y13580 = ~1'b0 ;
  assign y13581 = ~1'b0 ;
  assign y13582 = ~n20589 ;
  assign y13583 = ~n29674 ;
  assign y13584 = ~n29677 ;
  assign y13585 = 1'b0 ;
  assign y13586 = n29681 ;
  assign y13587 = ~1'b0 ;
  assign y13588 = ~n29682 ;
  assign y13589 = n29689 ;
  assign y13590 = n29691 ;
  assign y13591 = n29694 ;
  assign y13592 = ~n29696 ;
  assign y13593 = ~n29699 ;
  assign y13594 = ~n29712 ;
  assign y13595 = ~n29715 ;
  assign y13596 = ~1'b0 ;
  assign y13597 = n29718 ;
  assign y13598 = ~n29720 ;
  assign y13599 = n29722 ;
  assign y13600 = ~n29724 ;
  assign y13601 = ~1'b0 ;
  assign y13602 = ~n29733 ;
  assign y13603 = ~n29734 ;
  assign y13604 = n29736 ;
  assign y13605 = n29738 ;
  assign y13606 = ~1'b0 ;
  assign y13607 = n29739 ;
  assign y13608 = n29742 ;
  assign y13609 = ~n29745 ;
  assign y13610 = n29746 ;
  assign y13611 = ~n29748 ;
  assign y13612 = ~n29749 ;
  assign y13613 = n29750 ;
  assign y13614 = ~1'b0 ;
  assign y13615 = ~n29756 ;
  assign y13616 = ~n29757 ;
  assign y13617 = ~n29762 ;
  assign y13618 = ~1'b0 ;
  assign y13619 = n29764 ;
  assign y13620 = ~1'b0 ;
  assign y13621 = ~n29766 ;
  assign y13622 = ~n29773 ;
  assign y13623 = ~1'b0 ;
  assign y13624 = ~1'b0 ;
  assign y13625 = n29777 ;
  assign y13626 = ~n29781 ;
  assign y13627 = n29782 ;
  assign y13628 = n29785 ;
  assign y13629 = ~n29786 ;
  assign y13630 = n29787 ;
  assign y13631 = n29790 ;
  assign y13632 = ~1'b0 ;
  assign y13633 = n519 ;
  assign y13634 = n29796 ;
  assign y13635 = ~n29797 ;
  assign y13636 = 1'b0 ;
  assign y13637 = ~n29800 ;
  assign y13638 = ~n29804 ;
  assign y13639 = ~1'b0 ;
  assign y13640 = ~n29806 ;
  assign y13641 = n29807 ;
  assign y13642 = ~1'b0 ;
  assign y13643 = ~1'b0 ;
  assign y13644 = n29810 ;
  assign y13645 = n1777 ;
  assign y13646 = n29811 ;
  assign y13647 = ~n29812 ;
  assign y13648 = n29813 ;
  assign y13649 = n29814 ;
  assign y13650 = n29816 ;
  assign y13651 = n29817 ;
  assign y13652 = n29822 ;
  assign y13653 = ~n29828 ;
  assign y13654 = ~n29832 ;
  assign y13655 = ~1'b0 ;
  assign y13656 = n29834 ;
  assign y13657 = ~1'b0 ;
  assign y13658 = ~n29836 ;
  assign y13659 = n29840 ;
  assign y13660 = n29844 ;
  assign y13661 = ~1'b0 ;
  assign y13662 = ~1'b0 ;
  assign y13663 = 1'b0 ;
  assign y13664 = n29852 ;
  assign y13665 = n29853 ;
  assign y13666 = ~n29858 ;
  assign y13667 = n29859 ;
  assign y13668 = ~n29862 ;
  assign y13669 = ~1'b0 ;
  assign y13670 = ~1'b0 ;
  assign y13671 = n29865 ;
  assign y13672 = ~n29868 ;
  assign y13673 = ~n29870 ;
  assign y13674 = ~1'b0 ;
  assign y13675 = n29873 ;
  assign y13676 = ~1'b0 ;
  assign y13677 = ~1'b0 ;
  assign y13678 = n29874 ;
  assign y13679 = ~n29880 ;
  assign y13680 = ~n29887 ;
  assign y13681 = n29892 ;
  assign y13682 = n29903 ;
  assign y13683 = n29906 ;
  assign y13684 = n29907 ;
  assign y13685 = n29908 ;
  assign y13686 = ~n29916 ;
  assign y13687 = n29917 ;
  assign y13688 = n29919 ;
  assign y13689 = ~n29920 ;
  assign y13690 = ~n29921 ;
  assign y13691 = ~n29924 ;
  assign y13692 = n29927 ;
  assign y13693 = ~1'b0 ;
  assign y13694 = ~n14972 ;
  assign y13695 = ~1'b0 ;
  assign y13696 = ~n29928 ;
  assign y13697 = n29929 ;
  assign y13698 = ~1'b0 ;
  assign y13699 = ~n29931 ;
  assign y13700 = n29937 ;
  assign y13701 = ~1'b0 ;
  assign y13702 = ~1'b0 ;
  assign y13703 = n29943 ;
  assign y13704 = ~n29944 ;
  assign y13705 = n29945 ;
  assign y13706 = ~n29946 ;
  assign y13707 = n29949 ;
  assign y13708 = ~n29950 ;
  assign y13709 = n29953 ;
  assign y13710 = n29955 ;
  assign y13711 = ~1'b0 ;
  assign y13712 = ~1'b0 ;
  assign y13713 = ~n29957 ;
  assign y13714 = ~n29958 ;
  assign y13715 = ~n29962 ;
  assign y13716 = ~1'b0 ;
  assign y13717 = ~n29964 ;
  assign y13718 = ~1'b0 ;
  assign y13719 = ~1'b0 ;
  assign y13720 = ~1'b0 ;
  assign y13721 = ~n29968 ;
  assign y13722 = n29969 ;
  assign y13723 = n29972 ;
  assign y13724 = n29973 ;
  assign y13725 = n29976 ;
  assign y13726 = n5225 ;
  assign y13727 = n29977 ;
  assign y13728 = ~1'b0 ;
  assign y13729 = n29978 ;
  assign y13730 = 1'b0 ;
  assign y13731 = n29979 ;
  assign y13732 = ~n29980 ;
  assign y13733 = n29985 ;
  assign y13734 = n29990 ;
  assign y13735 = n29992 ;
  assign y13736 = n29994 ;
  assign y13737 = n29995 ;
  assign y13738 = n29999 ;
  assign y13739 = ~1'b0 ;
  assign y13740 = ~1'b0 ;
  assign y13741 = n30000 ;
  assign y13742 = ~n30003 ;
  assign y13743 = ~1'b0 ;
  assign y13744 = ~n30004 ;
  assign y13745 = n30005 ;
  assign y13746 = ~1'b0 ;
  assign y13747 = n30008 ;
  assign y13748 = ~1'b0 ;
  assign y13749 = ~n30011 ;
  assign y13750 = ~1'b0 ;
  assign y13751 = ~1'b0 ;
  assign y13752 = n30018 ;
  assign y13753 = n30019 ;
  assign y13754 = ~n30020 ;
  assign y13755 = ~n30021 ;
  assign y13756 = ~n30022 ;
  assign y13757 = ~1'b0 ;
  assign y13758 = n30023 ;
  assign y13759 = ~n30027 ;
  assign y13760 = ~n30033 ;
  assign y13761 = ~1'b0 ;
  assign y13762 = ~1'b0 ;
  assign y13763 = ~1'b0 ;
  assign y13764 = ~n30034 ;
  assign y13765 = n30038 ;
  assign y13766 = ~1'b0 ;
  assign y13767 = n30039 ;
  assign y13768 = n30040 ;
  assign y13769 = ~1'b0 ;
  assign y13770 = ~n30042 ;
  assign y13771 = ~n30044 ;
  assign y13772 = ~n13164 ;
  assign y13773 = n30054 ;
  assign y13774 = n30061 ;
  assign y13775 = n30065 ;
  assign y13776 = n30067 ;
  assign y13777 = ~n3430 ;
  assign y13778 = ~1'b0 ;
  assign y13779 = ~1'b0 ;
  assign y13780 = n30072 ;
  assign y13781 = n30082 ;
  assign y13782 = ~n30085 ;
  assign y13783 = n30087 ;
  assign y13784 = n17861 ;
  assign y13785 = n30092 ;
  assign y13786 = ~n30093 ;
  assign y13787 = ~n30098 ;
  assign y13788 = ~1'b0 ;
  assign y13789 = ~n30100 ;
  assign y13790 = ~n30102 ;
  assign y13791 = ~n30104 ;
  assign y13792 = ~n30112 ;
  assign y13793 = n30119 ;
  assign y13794 = n30121 ;
  assign y13795 = ~n30126 ;
  assign y13796 = ~1'b0 ;
  assign y13797 = ~n30129 ;
  assign y13798 = ~n852 ;
  assign y13799 = ~1'b0 ;
  assign y13800 = n30130 ;
  assign y13801 = ~n30133 ;
  assign y13802 = n17783 ;
  assign y13803 = ~n30134 ;
  assign y13804 = ~n30136 ;
  assign y13805 = n30137 ;
  assign y13806 = ~n30140 ;
  assign y13807 = ~n30141 ;
  assign y13808 = ~n30145 ;
  assign y13809 = ~n30146 ;
  assign y13810 = ~n30148 ;
  assign y13811 = ~n30150 ;
  assign y13812 = ~n30152 ;
  assign y13813 = ~n30159 ;
  assign y13814 = ~n30165 ;
  assign y13815 = n30166 ;
  assign y13816 = ~n30172 ;
  assign y13817 = ~1'b0 ;
  assign y13818 = ~1'b0 ;
  assign y13819 = ~n30173 ;
  assign y13820 = n30174 ;
  assign y13821 = ~n30178 ;
  assign y13822 = ~1'b0 ;
  assign y13823 = ~1'b0 ;
  assign y13824 = ~1'b0 ;
  assign y13825 = ~n30180 ;
  assign y13826 = n30181 ;
  assign y13827 = ~n12784 ;
  assign y13828 = n30183 ;
  assign y13829 = n30184 ;
  assign y13830 = ~n30186 ;
  assign y13831 = ~n30188 ;
  assign y13832 = n30189 ;
  assign y13833 = ~n16321 ;
  assign y13834 = ~1'b0 ;
  assign y13835 = ~1'b0 ;
  assign y13836 = n30192 ;
  assign y13837 = ~1'b0 ;
  assign y13838 = n30193 ;
  assign y13839 = n30194 ;
  assign y13840 = ~n30199 ;
  assign y13841 = 1'b0 ;
  assign y13842 = ~n30206 ;
  assign y13843 = ~n30207 ;
  assign y13844 = ~n30208 ;
  assign y13845 = ~1'b0 ;
  assign y13846 = n6605 ;
  assign y13847 = ~1'b0 ;
  assign y13848 = ~n5329 ;
  assign y13849 = n30210 ;
  assign y13850 = n30211 ;
  assign y13851 = ~1'b0 ;
  assign y13852 = n30215 ;
  assign y13853 = ~n30222 ;
  assign y13854 = n30225 ;
  assign y13855 = ~1'b0 ;
  assign y13856 = ~n30233 ;
  assign y13857 = ~1'b0 ;
  assign y13858 = ~n30237 ;
  assign y13859 = ~n30238 ;
  assign y13860 = ~n30240 ;
  assign y13861 = n30244 ;
  assign y13862 = 1'b0 ;
  assign y13863 = ~n30246 ;
  assign y13864 = n30248 ;
  assign y13865 = ~n30252 ;
  assign y13866 = n30254 ;
  assign y13867 = ~1'b0 ;
  assign y13868 = n30257 ;
  assign y13869 = ~n30258 ;
  assign y13870 = n30263 ;
  assign y13871 = ~n30265 ;
  assign y13872 = ~n30269 ;
  assign y13873 = ~n30271 ;
  assign y13874 = ~n30272 ;
  assign y13875 = ~n30277 ;
  assign y13876 = ~n30279 ;
  assign y13877 = ~1'b0 ;
  assign y13878 = n30282 ;
  assign y13879 = ~n30283 ;
  assign y13880 = ~n30284 ;
  assign y13881 = ~n30286 ;
  assign y13882 = ~n30287 ;
  assign y13883 = ~n10995 ;
  assign y13884 = n30290 ;
  assign y13885 = ~1'b0 ;
  assign y13886 = ~n30293 ;
  assign y13887 = n8374 ;
  assign y13888 = n30302 ;
  assign y13889 = ~1'b0 ;
  assign y13890 = ~n30304 ;
  assign y13891 = ~1'b0 ;
  assign y13892 = ~n30305 ;
  assign y13893 = n30309 ;
  assign y13894 = n30312 ;
  assign y13895 = ~n30313 ;
  assign y13896 = ~n30315 ;
  assign y13897 = n30328 ;
  assign y13898 = ~n30330 ;
  assign y13899 = ~n20405 ;
  assign y13900 = ~n30340 ;
  assign y13901 = n30342 ;
  assign y13902 = n30344 ;
  assign y13903 = n30346 ;
  assign y13904 = ~1'b0 ;
  assign y13905 = n30348 ;
  assign y13906 = n30349 ;
  assign y13907 = ~n30352 ;
  assign y13908 = n30354 ;
  assign y13909 = ~n30357 ;
  assign y13910 = ~1'b0 ;
  assign y13911 = ~1'b0 ;
  assign y13912 = ~1'b0 ;
  assign y13913 = ~n30359 ;
  assign y13914 = ~n30363 ;
  assign y13915 = n30375 ;
  assign y13916 = ~1'b0 ;
  assign y13917 = ~n3260 ;
  assign y13918 = ~n11736 ;
  assign y13919 = n30378 ;
  assign y13920 = n30383 ;
  assign y13921 = ~n24891 ;
  assign y13922 = ~n30388 ;
  assign y13923 = n30389 ;
  assign y13924 = n30390 ;
  assign y13925 = ~1'b0 ;
  assign y13926 = n30396 ;
  assign y13927 = n30397 ;
  assign y13928 = n30403 ;
  assign y13929 = ~n30409 ;
  assign y13930 = ~n30410 ;
  assign y13931 = n30412 ;
  assign y13932 = ~n30413 ;
  assign y13933 = n30414 ;
  assign y13934 = ~n30417 ;
  assign y13935 = n30421 ;
  assign y13936 = ~n30423 ;
  assign y13937 = ~n30426 ;
  assign y13938 = n30429 ;
  assign y13939 = ~1'b0 ;
  assign y13940 = ~1'b0 ;
  assign y13941 = ~n30436 ;
  assign y13942 = ~n30440 ;
  assign y13943 = ~n30447 ;
  assign y13944 = n30458 ;
  assign y13945 = ~1'b0 ;
  assign y13946 = n30462 ;
  assign y13947 = ~n30464 ;
  assign y13948 = n30468 ;
  assign y13949 = ~n30469 ;
  assign y13950 = n30470 ;
  assign y13951 = ~n30471 ;
  assign y13952 = ~n30472 ;
  assign y13953 = ~n30473 ;
  assign y13954 = ~n30477 ;
  assign y13955 = ~n30478 ;
  assign y13956 = ~n30479 ;
  assign y13957 = ~n692 ;
  assign y13958 = n30480 ;
  assign y13959 = n30484 ;
  assign y13960 = ~n30486 ;
  assign y13961 = ~n30487 ;
  assign y13962 = n30490 ;
  assign y13963 = ~1'b0 ;
  assign y13964 = n30491 ;
  assign y13965 = ~1'b0 ;
  assign y13966 = n30493 ;
  assign y13967 = ~1'b0 ;
  assign y13968 = ~1'b0 ;
  assign y13969 = ~n30494 ;
  assign y13970 = n30495 ;
  assign y13971 = ~n30497 ;
  assign y13972 = ~1'b0 ;
  assign y13973 = ~1'b0 ;
  assign y13974 = n30501 ;
  assign y13975 = ~1'b0 ;
  assign y13976 = ~n30502 ;
  assign y13977 = ~1'b0 ;
  assign y13978 = ~n30504 ;
  assign y13979 = ~n30505 ;
  assign y13980 = ~n30510 ;
  assign y13981 = n30511 ;
  assign y13982 = n30516 ;
  assign y13983 = ~n30517 ;
  assign y13984 = ~1'b0 ;
  assign y13985 = 1'b0 ;
  assign y13986 = ~n30519 ;
  assign y13987 = n30521 ;
  assign y13988 = n30522 ;
  assign y13989 = n30523 ;
  assign y13990 = n30525 ;
  assign y13991 = n30527 ;
  assign y13992 = n30528 ;
  assign y13993 = ~n30531 ;
  assign y13994 = ~n30532 ;
  assign y13995 = n30535 ;
  assign y13996 = n30536 ;
  assign y13997 = ~n30539 ;
  assign y13998 = ~n30541 ;
  assign y13999 = n30542 ;
  assign y14000 = ~n30544 ;
  assign y14001 = n30547 ;
  assign y14002 = n30548 ;
  assign y14003 = ~n30549 ;
  assign y14004 = n30551 ;
  assign y14005 = ~1'b0 ;
  assign y14006 = n30556 ;
  assign y14007 = ~n30557 ;
  assign y14008 = n30562 ;
  assign y14009 = ~n30564 ;
  assign y14010 = n30565 ;
  assign y14011 = ~1'b0 ;
  assign y14012 = ~1'b0 ;
  assign y14013 = n30567 ;
  assign y14014 = ~1'b0 ;
  assign y14015 = ~n30570 ;
  assign y14016 = ~1'b0 ;
  assign y14017 = ~n30572 ;
  assign y14018 = n9416 ;
  assign y14019 = n30575 ;
  assign y14020 = ~n30576 ;
  assign y14021 = n30578 ;
  assign y14022 = ~1'b0 ;
  assign y14023 = ~1'b0 ;
  assign y14024 = n30582 ;
  assign y14025 = n30583 ;
  assign y14026 = n30587 ;
  assign y14027 = ~n30591 ;
  assign y14028 = ~n30594 ;
  assign y14029 = ~n30595 ;
  assign y14030 = ~1'b0 ;
  assign y14031 = ~1'b0 ;
  assign y14032 = ~1'b0 ;
  assign y14033 = ~n30597 ;
  assign y14034 = n30598 ;
  assign y14035 = n30600 ;
  assign y14036 = ~n30605 ;
  assign y14037 = ~n30606 ;
  assign y14038 = n30612 ;
  assign y14039 = ~1'b0 ;
  assign y14040 = ~n30618 ;
  assign y14041 = ~1'b0 ;
  assign y14042 = ~n30623 ;
  assign y14043 = n30625 ;
  assign y14044 = n30629 ;
  assign y14045 = n30632 ;
  assign y14046 = n30637 ;
  assign y14047 = n30659 ;
  assign y14048 = ~n30677 ;
  assign y14049 = ~n30683 ;
  assign y14050 = ~n30684 ;
  assign y14051 = ~n30686 ;
  assign y14052 = ~n30688 ;
  assign y14053 = n30690 ;
  assign y14054 = ~n30694 ;
  assign y14055 = ~n17490 ;
  assign y14056 = ~n30695 ;
  assign y14057 = ~1'b0 ;
  assign y14058 = ~n30696 ;
  assign y14059 = n30697 ;
  assign y14060 = ~n30699 ;
  assign y14061 = ~n30701 ;
  assign y14062 = ~1'b0 ;
  assign y14063 = ~n30703 ;
  assign y14064 = ~n30704 ;
  assign y14065 = ~n30709 ;
  assign y14066 = ~n30711 ;
  assign y14067 = n30716 ;
  assign y14068 = n30720 ;
  assign y14069 = ~n30721 ;
  assign y14070 = ~n30722 ;
  assign y14071 = n30726 ;
  assign y14072 = ~n30731 ;
  assign y14073 = ~n30733 ;
  assign y14074 = ~n30741 ;
  assign y14075 = n30744 ;
  assign y14076 = ~1'b0 ;
  assign y14077 = n30747 ;
  assign y14078 = n30750 ;
  assign y14079 = ~1'b0 ;
  assign y14080 = ~n30751 ;
  assign y14081 = ~n2546 ;
  assign y14082 = ~n25242 ;
  assign y14083 = n30755 ;
  assign y14084 = ~1'b0 ;
  assign y14085 = ~1'b0 ;
  assign y14086 = ~n30757 ;
  assign y14087 = ~n30762 ;
  assign y14088 = ~n30765 ;
  assign y14089 = n30768 ;
  assign y14090 = ~1'b0 ;
  assign y14091 = ~1'b0 ;
  assign y14092 = ~1'b0 ;
  assign y14093 = ~n30770 ;
  assign y14094 = n30774 ;
  assign y14095 = n30777 ;
  assign y14096 = ~n30779 ;
  assign y14097 = ~1'b0 ;
  assign y14098 = n30783 ;
  assign y14099 = ~n2281 ;
  assign y14100 = ~1'b0 ;
  assign y14101 = ~n30786 ;
  assign y14102 = n30789 ;
  assign y14103 = ~n30792 ;
  assign y14104 = ~1'b0 ;
  assign y14105 = ~n30794 ;
  assign y14106 = ~n30795 ;
  assign y14107 = ~n30804 ;
  assign y14108 = n30808 ;
  assign y14109 = n30811 ;
  assign y14110 = ~1'b0 ;
  assign y14111 = n30814 ;
  assign y14112 = ~1'b0 ;
  assign y14113 = ~n30816 ;
  assign y14114 = ~n30819 ;
  assign y14115 = ~1'b0 ;
  assign y14116 = ~n30820 ;
  assign y14117 = ~1'b0 ;
  assign y14118 = ~1'b0 ;
  assign y14119 = ~1'b0 ;
  assign y14120 = n30830 ;
  assign y14121 = ~1'b0 ;
  assign y14122 = ~n2425 ;
  assign y14123 = n30835 ;
  assign y14124 = ~n30838 ;
  assign y14125 = n30839 ;
  assign y14126 = ~n30843 ;
  assign y14127 = ~n30844 ;
  assign y14128 = n30848 ;
  assign y14129 = ~n30850 ;
  assign y14130 = ~1'b0 ;
  assign y14131 = ~1'b0 ;
  assign y14132 = n30853 ;
  assign y14133 = ~1'b0 ;
  assign y14134 = ~n30855 ;
  assign y14135 = ~n30859 ;
  assign y14136 = n30865 ;
  assign y14137 = ~1'b0 ;
  assign y14138 = n30868 ;
  assign y14139 = ~n30869 ;
  assign y14140 = ~n30871 ;
  assign y14141 = ~n30873 ;
  assign y14142 = ~n30875 ;
  assign y14143 = ~n30878 ;
  assign y14144 = ~n30879 ;
  assign y14145 = n10721 ;
  assign y14146 = ~n30880 ;
  assign y14147 = n30884 ;
  assign y14148 = ~1'b0 ;
  assign y14149 = ~n30890 ;
  assign y14150 = ~1'b0 ;
  assign y14151 = n30892 ;
  assign y14152 = ~n4892 ;
  assign y14153 = ~n18048 ;
  assign y14154 = ~n1461 ;
  assign y14155 = n30896 ;
  assign y14156 = ~n30900 ;
  assign y14157 = ~n30903 ;
  assign y14158 = n30910 ;
  assign y14159 = n30911 ;
  assign y14160 = ~n30913 ;
  assign y14161 = n30915 ;
  assign y14162 = ~1'b0 ;
  assign y14163 = n30917 ;
  assign y14164 = ~1'b0 ;
  assign y14165 = ~n30920 ;
  assign y14166 = ~n30923 ;
  assign y14167 = n30926 ;
  assign y14168 = ~n30929 ;
  assign y14169 = n30931 ;
  assign y14170 = ~1'b0 ;
  assign y14171 = ~n30932 ;
  assign y14172 = n30933 ;
  assign y14173 = ~n30937 ;
  assign y14174 = n30938 ;
  assign y14175 = n30946 ;
  assign y14176 = ~n30952 ;
  assign y14177 = ~1'b0 ;
  assign y14178 = n30954 ;
  assign y14179 = ~n30956 ;
  assign y14180 = ~n30958 ;
  assign y14181 = n30961 ;
  assign y14182 = ~1'b0 ;
  assign y14183 = ~1'b0 ;
  assign y14184 = ~1'b0 ;
  assign y14185 = ~1'b0 ;
  assign y14186 = ~n30963 ;
  assign y14187 = ~n30964 ;
  assign y14188 = ~n30969 ;
  assign y14189 = n30975 ;
  assign y14190 = ~n30976 ;
  assign y14191 = ~1'b0 ;
  assign y14192 = ~1'b0 ;
  assign y14193 = n30977 ;
  assign y14194 = n11969 ;
  assign y14195 = ~n30978 ;
  assign y14196 = ~1'b0 ;
  assign y14197 = ~n30981 ;
  assign y14198 = ~n30984 ;
  assign y14199 = ~n30987 ;
  assign y14200 = n30994 ;
  assign y14201 = ~1'b0 ;
  assign y14202 = ~1'b0 ;
  assign y14203 = ~1'b0 ;
  assign y14204 = n30995 ;
  assign y14205 = n30998 ;
  assign y14206 = n8767 ;
  assign y14207 = n31004 ;
  assign y14208 = n31009 ;
  assign y14209 = n31012 ;
  assign y14210 = ~n31014 ;
  assign y14211 = ~1'b0 ;
  assign y14212 = ~1'b0 ;
  assign y14213 = n5224 ;
  assign y14214 = ~n31017 ;
  assign y14215 = ~n31018 ;
  assign y14216 = 1'b0 ;
  assign y14217 = ~1'b0 ;
  assign y14218 = ~n31028 ;
  assign y14219 = ~1'b0 ;
  assign y14220 = n31033 ;
  assign y14221 = n31034 ;
  assign y14222 = ~n31038 ;
  assign y14223 = ~n31040 ;
  assign y14224 = ~1'b0 ;
  assign y14225 = ~n31042 ;
  assign y14226 = n31043 ;
  assign y14227 = ~1'b0 ;
  assign y14228 = ~1'b0 ;
  assign y14229 = ~n31045 ;
  assign y14230 = ~n31049 ;
  assign y14231 = 1'b0 ;
  assign y14232 = n31051 ;
  assign y14233 = ~1'b0 ;
  assign y14234 = ~n31054 ;
  assign y14235 = n31056 ;
  assign y14236 = n31059 ;
  assign y14237 = n31064 ;
  assign y14238 = n31065 ;
  assign y14239 = ~n31067 ;
  assign y14240 = ~1'b0 ;
  assign y14241 = ~n4826 ;
  assign y14242 = ~1'b0 ;
  assign y14243 = ~1'b0 ;
  assign y14244 = n31069 ;
  assign y14245 = ~n31073 ;
  assign y14246 = ~n31075 ;
  assign y14247 = n31081 ;
  assign y14248 = n31083 ;
  assign y14249 = ~1'b0 ;
  assign y14250 = ~n31091 ;
  assign y14251 = ~n31095 ;
  assign y14252 = ~1'b0 ;
  assign y14253 = ~n31101 ;
  assign y14254 = ~n31104 ;
  assign y14255 = ~1'b0 ;
  assign y14256 = ~1'b0 ;
  assign y14257 = n31106 ;
  assign y14258 = 1'b0 ;
  assign y14259 = n31107 ;
  assign y14260 = ~1'b0 ;
  assign y14261 = ~n31110 ;
  assign y14262 = ~1'b0 ;
  assign y14263 = ~1'b0 ;
  assign y14264 = ~n31112 ;
  assign y14265 = ~1'b0 ;
  assign y14266 = n31117 ;
  assign y14267 = ~1'b0 ;
  assign y14268 = ~n31118 ;
  assign y14269 = ~1'b0 ;
  assign y14270 = ~n14758 ;
  assign y14271 = ~n31120 ;
  assign y14272 = n612 ;
  assign y14273 = n31122 ;
  assign y14274 = ~n31123 ;
  assign y14275 = ~1'b0 ;
  assign y14276 = n31127 ;
  assign y14277 = ~1'b0 ;
  assign y14278 = n31128 ;
  assign y14279 = n4914 ;
  assign y14280 = ~n31131 ;
  assign y14281 = 1'b0 ;
  assign y14282 = n31134 ;
  assign y14283 = n31136 ;
  assign y14284 = n31138 ;
  assign y14285 = ~1'b0 ;
  assign y14286 = ~n31141 ;
  assign y14287 = n31144 ;
  assign y14288 = n31147 ;
  assign y14289 = ~n31151 ;
  assign y14290 = ~n31154 ;
  assign y14291 = n31156 ;
  assign y14292 = ~n31157 ;
  assign y14293 = n31159 ;
  assign y14294 = ~1'b0 ;
  assign y14295 = ~n31160 ;
  assign y14296 = ~n31162 ;
  assign y14297 = n31165 ;
  assign y14298 = n31167 ;
  assign y14299 = ~1'b0 ;
  assign y14300 = ~1'b0 ;
  assign y14301 = n31168 ;
  assign y14302 = ~n31172 ;
  assign y14303 = n31173 ;
  assign y14304 = ~1'b0 ;
  assign y14305 = ~1'b0 ;
  assign y14306 = n31176 ;
  assign y14307 = ~n31178 ;
  assign y14308 = n31184 ;
  assign y14309 = ~n5781 ;
  assign y14310 = ~1'b0 ;
  assign y14311 = ~1'b0 ;
  assign y14312 = ~n31186 ;
  assign y14313 = n31188 ;
  assign y14314 = ~n31189 ;
  assign y14315 = n31190 ;
  assign y14316 = ~1'b0 ;
  assign y14317 = ~n31191 ;
  assign y14318 = n31193 ;
  assign y14319 = n12249 ;
  assign y14320 = ~1'b0 ;
  assign y14321 = ~n31195 ;
  assign y14322 = ~1'b0 ;
  assign y14323 = n31198 ;
  assign y14324 = ~n31204 ;
  assign y14325 = ~1'b0 ;
  assign y14326 = ~n31207 ;
  assign y14327 = ~1'b0 ;
  assign y14328 = ~1'b0 ;
  assign y14329 = ~1'b0 ;
  assign y14330 = ~n31209 ;
  assign y14331 = n31212 ;
  assign y14332 = n31215 ;
  assign y14333 = ~1'b0 ;
  assign y14334 = ~1'b0 ;
  assign y14335 = ~n31217 ;
  assign y14336 = ~1'b0 ;
  assign y14337 = ~1'b0 ;
  assign y14338 = ~n31218 ;
  assign y14339 = ~n31219 ;
  assign y14340 = ~n31221 ;
  assign y14341 = n31223 ;
  assign y14342 = ~1'b0 ;
  assign y14343 = ~n31224 ;
  assign y14344 = ~n10649 ;
  assign y14345 = n31225 ;
  assign y14346 = ~n31231 ;
  assign y14347 = ~1'b0 ;
  assign y14348 = n31232 ;
  assign y14349 = n31236 ;
  assign y14350 = ~n31237 ;
  assign y14351 = n31238 ;
  assign y14352 = ~n31242 ;
  assign y14353 = n31243 ;
  assign y14354 = ~n31247 ;
  assign y14355 = ~1'b0 ;
  assign y14356 = ~n31251 ;
  assign y14357 = ~1'b0 ;
  assign y14358 = ~1'b0 ;
  assign y14359 = ~1'b0 ;
  assign y14360 = ~n31252 ;
  assign y14361 = ~n31253 ;
  assign y14362 = n31255 ;
  assign y14363 = ~1'b0 ;
  assign y14364 = ~1'b0 ;
  assign y14365 = n31257 ;
  assign y14366 = ~n31261 ;
  assign y14367 = n31262 ;
  assign y14368 = ~1'b0 ;
  assign y14369 = ~n31265 ;
  assign y14370 = ~n31270 ;
  assign y14371 = ~n31273 ;
  assign y14372 = ~n31274 ;
  assign y14373 = n31277 ;
  assign y14374 = ~1'b0 ;
  assign y14375 = ~n31279 ;
  assign y14376 = n31282 ;
  assign y14377 = ~1'b0 ;
  assign y14378 = ~1'b0 ;
  assign y14379 = ~n31283 ;
  assign y14380 = ~n31288 ;
  assign y14381 = 1'b0 ;
  assign y14382 = n31292 ;
  assign y14383 = n31293 ;
  assign y14384 = n31295 ;
  assign y14385 = ~1'b0 ;
  assign y14386 = ~n31297 ;
  assign y14387 = ~n31303 ;
  assign y14388 = ~n31306 ;
  assign y14389 = n31308 ;
  assign y14390 = ~1'b0 ;
  assign y14391 = ~n31310 ;
  assign y14392 = ~n31311 ;
  assign y14393 = ~1'b0 ;
  assign y14394 = ~1'b0 ;
  assign y14395 = ~n31314 ;
  assign y14396 = n31318 ;
  assign y14397 = ~1'b0 ;
  assign y14398 = n31322 ;
  assign y14399 = n31323 ;
  assign y14400 = n31326 ;
  assign y14401 = ~1'b0 ;
  assign y14402 = ~n31329 ;
  assign y14403 = ~n31339 ;
  assign y14404 = ~n31340 ;
  assign y14405 = ~1'b0 ;
  assign y14406 = ~1'b0 ;
  assign y14407 = ~n31341 ;
  assign y14408 = ~n31344 ;
  assign y14409 = ~n31346 ;
  assign y14410 = ~n31349 ;
  assign y14411 = ~n31350 ;
  assign y14412 = n31353 ;
  assign y14413 = ~n31355 ;
  assign y14414 = n31356 ;
  assign y14415 = ~1'b0 ;
  assign y14416 = ~1'b0 ;
  assign y14417 = n31357 ;
  assign y14418 = n31360 ;
  assign y14419 = n31364 ;
  assign y14420 = n31372 ;
  assign y14421 = ~1'b0 ;
  assign y14422 = n31373 ;
  assign y14423 = n31375 ;
  assign y14424 = ~1'b0 ;
  assign y14425 = n31376 ;
  assign y14426 = ~1'b0 ;
  assign y14427 = ~n31379 ;
  assign y14428 = n31380 ;
  assign y14429 = n31383 ;
  assign y14430 = ~1'b0 ;
  assign y14431 = n31384 ;
  assign y14432 = ~n31391 ;
  assign y14433 = ~n31395 ;
  assign y14434 = ~1'b0 ;
  assign y14435 = ~1'b0 ;
  assign y14436 = ~n31398 ;
  assign y14437 = ~n15677 ;
  assign y14438 = n31404 ;
  assign y14439 = n31406 ;
  assign y14440 = n31408 ;
  assign y14441 = n31409 ;
  assign y14442 = n31414 ;
  assign y14443 = ~n31418 ;
  assign y14444 = n31422 ;
  assign y14445 = n31424 ;
  assign y14446 = n31425 ;
  assign y14447 = ~n31426 ;
  assign y14448 = n31427 ;
  assign y14449 = n31428 ;
  assign y14450 = ~n31429 ;
  assign y14451 = ~n31433 ;
  assign y14452 = n31435 ;
  assign y14453 = ~1'b0 ;
  assign y14454 = n31436 ;
  assign y14455 = n31437 ;
  assign y14456 = n31440 ;
  assign y14457 = ~n31446 ;
  assign y14458 = n31448 ;
  assign y14459 = n31452 ;
  assign y14460 = ~n31453 ;
  assign y14461 = n31454 ;
  assign y14462 = n31456 ;
  assign y14463 = ~n31458 ;
  assign y14464 = ~1'b0 ;
  assign y14465 = n31469 ;
  assign y14466 = ~n31471 ;
  assign y14467 = n31476 ;
  assign y14468 = ~n31477 ;
  assign y14469 = ~n31481 ;
  assign y14470 = 1'b0 ;
  assign y14471 = n31485 ;
  assign y14472 = ~n31488 ;
  assign y14473 = ~1'b0 ;
  assign y14474 = ~n31491 ;
  assign y14475 = ~n31492 ;
  assign y14476 = ~1'b0 ;
  assign y14477 = ~1'b0 ;
  assign y14478 = 1'b0 ;
  assign y14479 = n31496 ;
  assign y14480 = ~n31498 ;
  assign y14481 = ~1'b0 ;
  assign y14482 = n31503 ;
  assign y14483 = ~n31507 ;
  assign y14484 = ~1'b0 ;
  assign y14485 = n31508 ;
  assign y14486 = ~n935 ;
  assign y14487 = ~n31509 ;
  assign y14488 = n31510 ;
  assign y14489 = n31511 ;
  assign y14490 = ~n31515 ;
  assign y14491 = ~n31516 ;
  assign y14492 = ~n31517 ;
  assign y14493 = ~1'b0 ;
  assign y14494 = ~n31518 ;
  assign y14495 = n31519 ;
  assign y14496 = ~1'b0 ;
  assign y14497 = n31522 ;
  assign y14498 = ~n31526 ;
  assign y14499 = n31528 ;
  assign y14500 = n10321 ;
  assign y14501 = n31532 ;
  assign y14502 = ~n31538 ;
  assign y14503 = ~n31540 ;
  assign y14504 = n9686 ;
  assign y14505 = ~1'b0 ;
  assign y14506 = ~n31541 ;
  assign y14507 = ~1'b0 ;
  assign y14508 = ~1'b0 ;
  assign y14509 = n31546 ;
  assign y14510 = n31552 ;
  assign y14511 = n31553 ;
  assign y14512 = ~n31554 ;
  assign y14513 = n31560 ;
  assign y14514 = ~n31561 ;
  assign y14515 = n24908 ;
  assign y14516 = ~n31562 ;
  assign y14517 = n31564 ;
  assign y14518 = ~1'b0 ;
  assign y14519 = ~n31566 ;
  assign y14520 = ~n31567 ;
  assign y14521 = n31568 ;
  assign y14522 = ~n31574 ;
  assign y14523 = ~n32 ;
  assign y14524 = ~n31578 ;
  assign y14525 = ~n31579 ;
  assign y14526 = ~1'b0 ;
  assign y14527 = ~n31581 ;
  assign y14528 = n23548 ;
  assign y14529 = ~n31585 ;
  assign y14530 = n31587 ;
  assign y14531 = ~n31589 ;
  assign y14532 = ~1'b0 ;
  assign y14533 = ~1'b0 ;
  assign y14534 = ~n31595 ;
  assign y14535 = ~n31597 ;
  assign y14536 = ~n31601 ;
  assign y14537 = n31606 ;
  assign y14538 = n31608 ;
  assign y14539 = n31609 ;
  assign y14540 = n31610 ;
  assign y14541 = n31611 ;
  assign y14542 = n31624 ;
  assign y14543 = ~n31626 ;
  assign y14544 = ~n31627 ;
  assign y14545 = ~1'b0 ;
  assign y14546 = ~1'b0 ;
  assign y14547 = ~n31630 ;
  assign y14548 = n31631 ;
  assign y14549 = ~n31632 ;
  assign y14550 = ~1'b0 ;
  assign y14551 = ~n31633 ;
  assign y14552 = n31635 ;
  assign y14553 = ~1'b0 ;
  assign y14554 = ~n31637 ;
  assign y14555 = ~n31639 ;
  assign y14556 = ~1'b0 ;
  assign y14557 = n31641 ;
  assign y14558 = ~n31643 ;
  assign y14559 = n31645 ;
  assign y14560 = ~n31649 ;
  assign y14561 = ~n31651 ;
  assign y14562 = n31654 ;
  assign y14563 = ~n24647 ;
  assign y14564 = ~1'b0 ;
  assign y14565 = ~1'b0 ;
  assign y14566 = ~1'b0 ;
  assign y14567 = n31656 ;
  assign y14568 = ~n31659 ;
  assign y14569 = ~1'b0 ;
  assign y14570 = ~n31662 ;
  assign y14571 = ~1'b0 ;
  assign y14572 = n31664 ;
  assign y14573 = ~1'b0 ;
  assign y14574 = ~n31667 ;
  assign y14575 = ~1'b0 ;
  assign y14576 = ~n31669 ;
  assign y14577 = ~n31672 ;
  assign y14578 = ~n31675 ;
  assign y14579 = ~1'b0 ;
  assign y14580 = ~n2995 ;
  assign y14581 = n31676 ;
  assign y14582 = ~n31680 ;
  assign y14583 = n31684 ;
  assign y14584 = n31685 ;
  assign y14585 = ~1'b0 ;
  assign y14586 = n31692 ;
  assign y14587 = n12198 ;
  assign y14588 = ~1'b0 ;
  assign y14589 = ~n31693 ;
  assign y14590 = n31697 ;
  assign y14591 = n31700 ;
  assign y14592 = ~n31702 ;
  assign y14593 = ~1'b0 ;
  assign y14594 = ~1'b0 ;
  assign y14595 = ~n31703 ;
  assign y14596 = ~n31704 ;
  assign y14597 = ~n31710 ;
  assign y14598 = 1'b0 ;
  assign y14599 = ~n12612 ;
  assign y14600 = n31712 ;
  assign y14601 = n29095 ;
  assign y14602 = ~n31714 ;
  assign y14603 = n31718 ;
  assign y14604 = ~1'b0 ;
  assign y14605 = ~n31728 ;
  assign y14606 = n31730 ;
  assign y14607 = ~1'b0 ;
  assign y14608 = ~1'b0 ;
  assign y14609 = n31733 ;
  assign y14610 = n31735 ;
  assign y14611 = ~1'b0 ;
  assign y14612 = ~1'b0 ;
  assign y14613 = n31738 ;
  assign y14614 = ~1'b0 ;
  assign y14615 = ~n16328 ;
  assign y14616 = ~n31739 ;
  assign y14617 = n31740 ;
  assign y14618 = n31742 ;
  assign y14619 = ~1'b0 ;
  assign y14620 = ~n31745 ;
  assign y14621 = ~1'b0 ;
  assign y14622 = ~n31746 ;
  assign y14623 = ~1'b0 ;
  assign y14624 = n31747 ;
  assign y14625 = ~n31748 ;
  assign y14626 = ~n31749 ;
  assign y14627 = ~n31750 ;
  assign y14628 = ~n31752 ;
  assign y14629 = ~1'b0 ;
  assign y14630 = ~1'b0 ;
  assign y14631 = ~1'b0 ;
  assign y14632 = ~n31754 ;
  assign y14633 = ~n26373 ;
  assign y14634 = ~n31759 ;
  assign y14635 = ~1'b0 ;
  assign y14636 = n31760 ;
  assign y14637 = n31762 ;
  assign y14638 = n31767 ;
  assign y14639 = n30117 ;
  assign y14640 = n31768 ;
  assign y14641 = n31771 ;
  assign y14642 = ~1'b0 ;
  assign y14643 = ~n31775 ;
  assign y14644 = n31778 ;
  assign y14645 = ~n24304 ;
  assign y14646 = n31780 ;
  assign y14647 = n31781 ;
  assign y14648 = ~1'b0 ;
  assign y14649 = n31783 ;
  assign y14650 = n31784 ;
  assign y14651 = n31790 ;
  assign y14652 = ~1'b0 ;
  assign y14653 = ~n31793 ;
  assign y14654 = n31798 ;
  assign y14655 = n31800 ;
  assign y14656 = ~1'b0 ;
  assign y14657 = ~n31804 ;
  assign y14658 = n31805 ;
  assign y14659 = n31810 ;
  assign y14660 = n31811 ;
  assign y14661 = ~n26809 ;
  assign y14662 = ~n18875 ;
  assign y14663 = ~1'b0 ;
  assign y14664 = ~n31815 ;
  assign y14665 = n25164 ;
  assign y14666 = ~n31818 ;
  assign y14667 = ~1'b0 ;
  assign y14668 = ~n31821 ;
  assign y14669 = n31825 ;
  assign y14670 = ~n31827 ;
  assign y14671 = n31828 ;
  assign y14672 = ~n31831 ;
  assign y14673 = n31837 ;
  assign y14674 = ~1'b0 ;
  assign y14675 = n31839 ;
  assign y14676 = ~1'b0 ;
  assign y14677 = ~1'b0 ;
  assign y14678 = n22893 ;
  assign y14679 = n31844 ;
  assign y14680 = ~n31846 ;
  assign y14681 = ~n31849 ;
  assign y14682 = n31850 ;
  assign y14683 = ~1'b0 ;
  assign y14684 = ~n31855 ;
  assign y14685 = ~1'b0 ;
  assign y14686 = n31860 ;
  assign y14687 = ~1'b0 ;
  assign y14688 = n31862 ;
  assign y14689 = ~n31873 ;
  assign y14690 = ~1'b0 ;
  assign y14691 = ~n31876 ;
  assign y14692 = ~1'b0 ;
  assign y14693 = ~n31877 ;
  assign y14694 = ~n31882 ;
  assign y14695 = n31883 ;
  assign y14696 = n31887 ;
  assign y14697 = ~n31891 ;
  assign y14698 = ~1'b0 ;
  assign y14699 = ~1'b0 ;
  assign y14700 = ~1'b0 ;
  assign y14701 = n31899 ;
  assign y14702 = ~n31900 ;
  assign y14703 = ~n31902 ;
  assign y14704 = ~n31907 ;
  assign y14705 = n31912 ;
  assign y14706 = ~n31919 ;
  assign y14707 = ~1'b0 ;
  assign y14708 = ~n31920 ;
  assign y14709 = ~n31921 ;
  assign y14710 = n31923 ;
  assign y14711 = n31927 ;
  assign y14712 = ~1'b0 ;
  assign y14713 = ~n31934 ;
  assign y14714 = ~n31936 ;
  assign y14715 = n31938 ;
  assign y14716 = ~n31940 ;
  assign y14717 = ~n31941 ;
  assign y14718 = 1'b0 ;
  assign y14719 = n31943 ;
  assign y14720 = n31947 ;
  assign y14721 = n31949 ;
  assign y14722 = ~n31951 ;
  assign y14723 = ~n31952 ;
  assign y14724 = ~1'b0 ;
  assign y14725 = ~n31959 ;
  assign y14726 = ~1'b0 ;
  assign y14727 = n31960 ;
  assign y14728 = ~1'b0 ;
  assign y14729 = n31966 ;
  assign y14730 = ~n31967 ;
  assign y14731 = ~1'b0 ;
  assign y14732 = ~n31969 ;
  assign y14733 = n31970 ;
  assign y14734 = ~1'b0 ;
  assign y14735 = n27793 ;
  assign y14736 = ~1'b0 ;
  assign y14737 = ~n31972 ;
  assign y14738 = n31977 ;
  assign y14739 = ~n31981 ;
  assign y14740 = n31982 ;
  assign y14741 = n31986 ;
  assign y14742 = 1'b0 ;
  assign y14743 = ~1'b0 ;
  assign y14744 = ~1'b0 ;
  assign y14745 = ~n31987 ;
  assign y14746 = ~n31988 ;
  assign y14747 = ~1'b0 ;
  assign y14748 = ~1'b0 ;
  assign y14749 = ~1'b0 ;
  assign y14750 = ~n15958 ;
  assign y14751 = ~n31993 ;
  assign y14752 = ~n32000 ;
  assign y14753 = ~n32002 ;
  assign y14754 = ~1'b0 ;
  assign y14755 = ~n5711 ;
  assign y14756 = n32011 ;
  assign y14757 = n32012 ;
  assign y14758 = ~1'b0 ;
  assign y14759 = ~n32014 ;
  assign y14760 = ~n32019 ;
  assign y14761 = ~1'b0 ;
  assign y14762 = ~n32020 ;
  assign y14763 = ~n32024 ;
  assign y14764 = ~n22483 ;
  assign y14765 = ~n32026 ;
  assign y14766 = n32032 ;
  assign y14767 = ~1'b0 ;
  assign y14768 = n32036 ;
  assign y14769 = ~n32038 ;
  assign y14770 = ~1'b0 ;
  assign y14771 = ~n26197 ;
  assign y14772 = ~n32041 ;
  assign y14773 = ~1'b0 ;
  assign y14774 = n32043 ;
  assign y14775 = ~n32044 ;
  assign y14776 = ~1'b0 ;
  assign y14777 = n32048 ;
  assign y14778 = n32053 ;
  assign y14779 = ~n32057 ;
  assign y14780 = ~n6126 ;
  assign y14781 = ~1'b0 ;
  assign y14782 = ~n32059 ;
  assign y14783 = n32061 ;
  assign y14784 = ~n32063 ;
  assign y14785 = ~n32065 ;
  assign y14786 = ~1'b0 ;
  assign y14787 = ~n32066 ;
  assign y14788 = n32067 ;
  assign y14789 = n32068 ;
  assign y14790 = ~n32071 ;
  assign y14791 = ~1'b0 ;
  assign y14792 = ~1'b0 ;
  assign y14793 = ~1'b0 ;
  assign y14794 = n32073 ;
  assign y14795 = n32074 ;
  assign y14796 = ~n32076 ;
  assign y14797 = n32079 ;
  assign y14798 = ~n32092 ;
  assign y14799 = n32093 ;
  assign y14800 = n32094 ;
  assign y14801 = ~n32095 ;
  assign y14802 = n32098 ;
  assign y14803 = ~n7617 ;
  assign y14804 = n32100 ;
  assign y14805 = ~n32101 ;
  assign y14806 = ~n32102 ;
  assign y14807 = ~n32103 ;
  assign y14808 = ~1'b0 ;
  assign y14809 = ~1'b0 ;
  assign y14810 = ~n32105 ;
  assign y14811 = n32108 ;
  assign y14812 = n32111 ;
  assign y14813 = n32115 ;
  assign y14814 = ~1'b0 ;
  assign y14815 = ~n8822 ;
  assign y14816 = ~1'b0 ;
  assign y14817 = n32118 ;
  assign y14818 = ~n32119 ;
  assign y14819 = ~1'b0 ;
  assign y14820 = ~n32121 ;
  assign y14821 = ~n32122 ;
  assign y14822 = ~1'b0 ;
  assign y14823 = ~1'b0 ;
  assign y14824 = n32123 ;
  assign y14825 = ~n32124 ;
  assign y14826 = ~n32125 ;
  assign y14827 = n32126 ;
  assign y14828 = ~n32130 ;
  assign y14829 = n32138 ;
  assign y14830 = ~n32140 ;
  assign y14831 = ~1'b0 ;
  assign y14832 = ~n32142 ;
  assign y14833 = n7493 ;
  assign y14834 = ~n32143 ;
  assign y14835 = n32145 ;
  assign y14836 = ~1'b0 ;
  assign y14837 = n32147 ;
  assign y14838 = n32151 ;
  assign y14839 = n32152 ;
  assign y14840 = ~1'b0 ;
  assign y14841 = ~n32154 ;
  assign y14842 = ~n32157 ;
  assign y14843 = n32159 ;
  assign y14844 = n7917 ;
  assign y14845 = ~n32162 ;
  assign y14846 = ~1'b0 ;
  assign y14847 = ~n32163 ;
  assign y14848 = n32165 ;
  assign y14849 = n32168 ;
  assign y14850 = ~n32176 ;
  assign y14851 = n11874 ;
  assign y14852 = n32178 ;
  assign y14853 = ~n32181 ;
  assign y14854 = n32184 ;
  assign y14855 = n32185 ;
  assign y14856 = ~1'b0 ;
  assign y14857 = n32187 ;
  assign y14858 = n32194 ;
  assign y14859 = n32196 ;
  assign y14860 = n32197 ;
  assign y14861 = n32198 ;
  assign y14862 = ~1'b0 ;
  assign y14863 = n32204 ;
  assign y14864 = ~n32209 ;
  assign y14865 = ~1'b0 ;
  assign y14866 = ~1'b0 ;
  assign y14867 = ~n32213 ;
  assign y14868 = ~n32214 ;
  assign y14869 = n10854 ;
  assign y14870 = n32216 ;
  assign y14871 = ~n32218 ;
  assign y14872 = n32220 ;
  assign y14873 = ~1'b0 ;
  assign y14874 = ~n32221 ;
  assign y14875 = n18100 ;
  assign y14876 = ~1'b0 ;
  assign y14877 = ~1'b0 ;
  assign y14878 = ~1'b0 ;
  assign y14879 = ~1'b0 ;
  assign y14880 = ~n32223 ;
  assign y14881 = ~1'b0 ;
  assign y14882 = ~n32225 ;
  assign y14883 = n32231 ;
  assign y14884 = n32233 ;
  assign y14885 = n32235 ;
  assign y14886 = 1'b0 ;
  assign y14887 = ~1'b0 ;
  assign y14888 = ~1'b0 ;
  assign y14889 = ~n32236 ;
  assign y14890 = ~1'b0 ;
  assign y14891 = 1'b0 ;
  assign y14892 = ~1'b0 ;
  assign y14893 = ~n32238 ;
  assign y14894 = ~n1487 ;
  assign y14895 = ~1'b0 ;
  assign y14896 = ~n32242 ;
  assign y14897 = n32245 ;
  assign y14898 = ~n32247 ;
  assign y14899 = ~1'b0 ;
  assign y14900 = ~n32249 ;
  assign y14901 = ~1'b0 ;
  assign y14902 = ~1'b0 ;
  assign y14903 = n32251 ;
  assign y14904 = ~n32252 ;
  assign y14905 = ~n32254 ;
  assign y14906 = ~n32255 ;
  assign y14907 = n32269 ;
  assign y14908 = ~1'b0 ;
  assign y14909 = ~1'b0 ;
  assign y14910 = n32271 ;
  assign y14911 = n32274 ;
  assign y14912 = n32275 ;
  assign y14913 = ~n32280 ;
  assign y14914 = ~n6634 ;
  assign y14915 = ~n32282 ;
  assign y14916 = n32286 ;
  assign y14917 = ~n32287 ;
  assign y14918 = ~n2180 ;
  assign y14919 = ~n32291 ;
  assign y14920 = ~n32297 ;
  assign y14921 = ~n32298 ;
  assign y14922 = ~n32299 ;
  assign y14923 = n1387 ;
  assign y14924 = ~1'b0 ;
  assign y14925 = n20057 ;
  assign y14926 = ~n32300 ;
  assign y14927 = ~1'b0 ;
  assign y14928 = ~1'b0 ;
  assign y14929 = ~n32302 ;
  assign y14930 = ~n32304 ;
  assign y14931 = ~n32305 ;
  assign y14932 = ~1'b0 ;
  assign y14933 = ~n32313 ;
  assign y14934 = ~n32315 ;
  assign y14935 = n32316 ;
  assign y14936 = ~n32320 ;
  assign y14937 = ~1'b0 ;
  assign y14938 = ~n32321 ;
  assign y14939 = ~1'b0 ;
  assign y14940 = ~n32326 ;
  assign y14941 = ~1'b0 ;
  assign y14942 = ~n32329 ;
  assign y14943 = ~n32337 ;
  assign y14944 = ~n32342 ;
  assign y14945 = ~1'b0 ;
  assign y14946 = n32345 ;
  assign y14947 = n32347 ;
  assign y14948 = n32350 ;
  assign y14949 = ~1'b0 ;
  assign y14950 = n32354 ;
  assign y14951 = ~n2635 ;
  assign y14952 = ~1'b0 ;
  assign y14953 = n32361 ;
  assign y14954 = ~1'b0 ;
  assign y14955 = n32362 ;
  assign y14956 = ~1'b0 ;
  assign y14957 = n32365 ;
  assign y14958 = n32366 ;
  assign y14959 = n32372 ;
  assign y14960 = n32373 ;
  assign y14961 = n32374 ;
  assign y14962 = n32378 ;
  assign y14963 = n32384 ;
  assign y14964 = ~1'b0 ;
  assign y14965 = ~1'b0 ;
  assign y14966 = n16068 ;
  assign y14967 = ~1'b0 ;
  assign y14968 = ~n32385 ;
  assign y14969 = ~n9277 ;
  assign y14970 = ~n32386 ;
  assign y14971 = ~1'b0 ;
  assign y14972 = ~n26138 ;
  assign y14973 = ~1'b0 ;
  assign y14974 = ~n32389 ;
  assign y14975 = ~n32392 ;
  assign y14976 = ~n32395 ;
  assign y14977 = ~n24202 ;
  assign y14978 = n32399 ;
  assign y14979 = ~n13111 ;
  assign y14980 = 1'b0 ;
  assign y14981 = ~n32402 ;
  assign y14982 = ~1'b0 ;
  assign y14983 = 1'b0 ;
  assign y14984 = n32404 ;
  assign y14985 = n32405 ;
  assign y14986 = n32411 ;
  assign y14987 = n32416 ;
  assign y14988 = n32421 ;
  assign y14989 = ~1'b0 ;
  assign y14990 = ~1'b0 ;
  assign y14991 = ~1'b0 ;
  assign y14992 = 1'b0 ;
  assign y14993 = n32422 ;
  assign y14994 = n2262 ;
  assign y14995 = ~n32423 ;
  assign y14996 = n32425 ;
  assign y14997 = ~n20443 ;
  assign y14998 = ~1'b0 ;
  assign y14999 = ~n32427 ;
  assign y15000 = ~n32436 ;
  assign y15001 = ~1'b0 ;
  assign y15002 = ~n32437 ;
  assign y15003 = ~1'b0 ;
  assign y15004 = ~1'b0 ;
  assign y15005 = n32439 ;
  assign y15006 = n32441 ;
  assign y15007 = ~n32446 ;
  assign y15008 = ~1'b0 ;
  assign y15009 = ~n32448 ;
  assign y15010 = n32449 ;
  assign y15011 = n32451 ;
  assign y15012 = ~n32452 ;
  assign y15013 = ~n32453 ;
  assign y15014 = ~1'b0 ;
  assign y15015 = n32454 ;
  assign y15016 = n32458 ;
  assign y15017 = n32459 ;
  assign y15018 = ~n32461 ;
  assign y15019 = n32466 ;
  assign y15020 = ~n32474 ;
  assign y15021 = ~n32476 ;
  assign y15022 = 1'b0 ;
  assign y15023 = ~n32478 ;
  assign y15024 = n32479 ;
  assign y15025 = ~1'b0 ;
  assign y15026 = n32481 ;
  assign y15027 = ~n32488 ;
  assign y15028 = ~n32489 ;
  assign y15029 = 1'b0 ;
  assign y15030 = ~n32494 ;
  assign y15031 = ~n32496 ;
  assign y15032 = n32500 ;
  assign y15033 = n32502 ;
  assign y15034 = ~1'b0 ;
  assign y15035 = ~n32505 ;
  assign y15036 = n32506 ;
  assign y15037 = ~1'b0 ;
  assign y15038 = ~1'b0 ;
  assign y15039 = ~1'b0 ;
  assign y15040 = n32510 ;
  assign y15041 = ~n32511 ;
  assign y15042 = n32513 ;
  assign y15043 = ~1'b0 ;
  assign y15044 = ~n32514 ;
  assign y15045 = n32515 ;
  assign y15046 = n32516 ;
  assign y15047 = ~n32520 ;
  assign y15048 = ~n32528 ;
  assign y15049 = ~n32535 ;
  assign y15050 = ~n32536 ;
  assign y15051 = ~n9274 ;
  assign y15052 = ~n32538 ;
  assign y15053 = ~1'b0 ;
  assign y15054 = n32539 ;
  assign y15055 = n32540 ;
  assign y15056 = n32546 ;
  assign y15057 = ~1'b0 ;
  assign y15058 = ~n32547 ;
  assign y15059 = ~n32549 ;
  assign y15060 = ~1'b0 ;
  assign y15061 = n32551 ;
  assign y15062 = ~n32556 ;
  assign y15063 = ~n32557 ;
  assign y15064 = n32558 ;
  assign y15065 = ~1'b0 ;
  assign y15066 = ~1'b0 ;
  assign y15067 = ~n32559 ;
  assign y15068 = ~n32560 ;
  assign y15069 = ~n32561 ;
  assign y15070 = ~1'b0 ;
  assign y15071 = n32562 ;
  assign y15072 = ~n32564 ;
  assign y15073 = ~n32568 ;
  assign y15074 = n32571 ;
  assign y15075 = ~1'b0 ;
  assign y15076 = ~n32578 ;
  assign y15077 = ~n32588 ;
  assign y15078 = n32589 ;
  assign y15079 = ~1'b0 ;
  assign y15080 = ~n32590 ;
  assign y15081 = n32592 ;
  assign y15082 = ~n32593 ;
  assign y15083 = ~n32594 ;
  assign y15084 = n32596 ;
  assign y15085 = n32599 ;
  assign y15086 = n16794 ;
  assign y15087 = ~1'b0 ;
  assign y15088 = ~n32601 ;
  assign y15089 = ~1'b0 ;
  assign y15090 = n32604 ;
  assign y15091 = ~n32607 ;
  assign y15092 = ~n32609 ;
  assign y15093 = ~n32611 ;
  assign y15094 = 1'b0 ;
  assign y15095 = ~n32612 ;
  assign y15096 = ~n32617 ;
  assign y15097 = n32620 ;
  assign y15098 = ~1'b0 ;
  assign y15099 = n32622 ;
  assign y15100 = ~n32627 ;
  assign y15101 = n32628 ;
  assign y15102 = ~n18100 ;
  assign y15103 = n32630 ;
  assign y15104 = n32634 ;
  assign y15105 = ~1'b0 ;
  assign y15106 = ~n32636 ;
  assign y15107 = n32637 ;
  assign y15108 = ~1'b0 ;
  assign y15109 = ~n1862 ;
  assign y15110 = ~1'b0 ;
  assign y15111 = n32641 ;
  assign y15112 = ~n32644 ;
  assign y15113 = ~n32646 ;
  assign y15114 = ~n32647 ;
  assign y15115 = ~n32649 ;
  assign y15116 = n32653 ;
  assign y15117 = ~1'b0 ;
  assign y15118 = ~n32655 ;
  assign y15119 = n32658 ;
  assign y15120 = n17020 ;
  assign y15121 = ~1'b0 ;
  assign y15122 = ~1'b0 ;
  assign y15123 = ~1'b0 ;
  assign y15124 = n32663 ;
  assign y15125 = ~1'b0 ;
  assign y15126 = n32664 ;
  assign y15127 = ~n32670 ;
  assign y15128 = ~1'b0 ;
  assign y15129 = n32672 ;
  assign y15130 = ~n32674 ;
  assign y15131 = n32677 ;
  assign y15132 = n32679 ;
  assign y15133 = ~1'b0 ;
  assign y15134 = n32690 ;
  assign y15135 = ~n32691 ;
  assign y15136 = ~n32697 ;
  assign y15137 = ~1'b0 ;
  assign y15138 = ~n32705 ;
  assign y15139 = ~n32708 ;
  assign y15140 = n32709 ;
  assign y15141 = ~n32713 ;
  assign y15142 = n32714 ;
  assign y15143 = ~n32719 ;
  assign y15144 = ~n32722 ;
  assign y15145 = ~1'b0 ;
  assign y15146 = ~1'b0 ;
  assign y15147 = ~1'b0 ;
  assign y15148 = ~n32724 ;
  assign y15149 = ~1'b0 ;
  assign y15150 = n32725 ;
  assign y15151 = ~n32726 ;
  assign y15152 = n392 ;
  assign y15153 = ~n32729 ;
  assign y15154 = n32734 ;
  assign y15155 = n32735 ;
  assign y15156 = n32737 ;
  assign y15157 = ~1'b0 ;
  assign y15158 = ~n32738 ;
  assign y15159 = ~1'b0 ;
  assign y15160 = ~1'b0 ;
  assign y15161 = n32740 ;
  assign y15162 = ~n32745 ;
  assign y15163 = ~n32748 ;
  assign y15164 = n32749 ;
  assign y15165 = ~1'b0 ;
  assign y15166 = ~n32752 ;
  assign y15167 = n7049 ;
  assign y15168 = ~1'b0 ;
  assign y15169 = ~1'b0 ;
  assign y15170 = ~1'b0 ;
  assign y15171 = n32753 ;
  assign y15172 = ~1'b0 ;
  assign y15173 = ~1'b0 ;
  assign y15174 = ~n32756 ;
  assign y15175 = n32758 ;
  assign y15176 = ~n32763 ;
  assign y15177 = n32764 ;
  assign y15178 = n32766 ;
  assign y15179 = ~n32767 ;
  assign y15180 = ~1'b0 ;
  assign y15181 = ~1'b0 ;
  assign y15182 = n32768 ;
  assign y15183 = ~n32770 ;
  assign y15184 = n32772 ;
  assign y15185 = ~n32775 ;
  assign y15186 = ~1'b0 ;
  assign y15187 = ~n32492 ;
  assign y15188 = ~n32783 ;
  assign y15189 = n32784 ;
  assign y15190 = ~1'b0 ;
  assign y15191 = n32785 ;
  assign y15192 = ~1'b0 ;
  assign y15193 = ~1'b0 ;
  assign y15194 = ~n32787 ;
  assign y15195 = ~1'b0 ;
  assign y15196 = n700 ;
  assign y15197 = ~1'b0 ;
  assign y15198 = ~1'b0 ;
  assign y15199 = ~1'b0 ;
  assign y15200 = ~n11973 ;
  assign y15201 = ~n32789 ;
  assign y15202 = ~n32797 ;
  assign y15203 = ~n21787 ;
  assign y15204 = ~1'b0 ;
  assign y15205 = ~1'b0 ;
  assign y15206 = ~1'b0 ;
  assign y15207 = n32798 ;
  assign y15208 = n32799 ;
  assign y15209 = ~1'b0 ;
  assign y15210 = ~n32805 ;
  assign y15211 = ~1'b0 ;
  assign y15212 = n32806 ;
  assign y15213 = ~n32809 ;
  assign y15214 = ~n32810 ;
  assign y15215 = ~1'b0 ;
  assign y15216 = ~n32811 ;
  assign y15217 = ~1'b0 ;
  assign y15218 = ~n32816 ;
  assign y15219 = ~1'b0 ;
  assign y15220 = ~1'b0 ;
  assign y15221 = ~n32819 ;
  assign y15222 = ~n32834 ;
  assign y15223 = ~1'b0 ;
  assign y15224 = ~n11372 ;
  assign y15225 = ~n32835 ;
  assign y15226 = ~n32839 ;
  assign y15227 = n32841 ;
  assign y15228 = ~n32842 ;
  assign y15229 = ~1'b0 ;
  assign y15230 = ~1'b0 ;
  assign y15231 = ~n32844 ;
  assign y15232 = ~n32846 ;
  assign y15233 = n32849 ;
  assign y15234 = ~1'b0 ;
  assign y15235 = ~1'b0 ;
  assign y15236 = n32853 ;
  assign y15237 = n32859 ;
  assign y15238 = 1'b0 ;
  assign y15239 = ~1'b0 ;
  assign y15240 = ~n32864 ;
  assign y15241 = ~n32865 ;
  assign y15242 = ~n32868 ;
  assign y15243 = ~n32870 ;
  assign y15244 = ~1'b0 ;
  assign y15245 = ~n32876 ;
  assign y15246 = ~n32879 ;
  assign y15247 = ~1'b0 ;
  assign y15248 = ~n32884 ;
  assign y15249 = n32889 ;
  assign y15250 = ~n32893 ;
  assign y15251 = n32899 ;
  assign y15252 = n32906 ;
  assign y15253 = n32907 ;
  assign y15254 = ~1'b0 ;
  assign y15255 = ~1'b0 ;
  assign y15256 = ~n32909 ;
  assign y15257 = ~n32911 ;
  assign y15258 = ~1'b0 ;
  assign y15259 = n32912 ;
  assign y15260 = ~1'b0 ;
  assign y15261 = ~n32920 ;
  assign y15262 = n32926 ;
  assign y15263 = ~1'b0 ;
  assign y15264 = ~1'b0 ;
  assign y15265 = ~1'b0 ;
  assign y15266 = ~1'b0 ;
  assign y15267 = ~n14781 ;
  assign y15268 = ~1'b0 ;
  assign y15269 = n32929 ;
  assign y15270 = 1'b0 ;
  assign y15271 = ~n32934 ;
  assign y15272 = n32935 ;
  assign y15273 = ~n32940 ;
  assign y15274 = ~1'b0 ;
  assign y15275 = n32941 ;
  assign y15276 = ~1'b0 ;
  assign y15277 = n32942 ;
  assign y15278 = ~n32945 ;
  assign y15279 = ~n32948 ;
  assign y15280 = ~n32949 ;
  assign y15281 = n32951 ;
  assign y15282 = ~1'b0 ;
  assign y15283 = n32954 ;
  assign y15284 = ~n16372 ;
  assign y15285 = ~n32956 ;
  assign y15286 = n32958 ;
  assign y15287 = n32960 ;
  assign y15288 = ~1'b0 ;
  assign y15289 = ~n24663 ;
  assign y15290 = ~n32961 ;
  assign y15291 = ~1'b0 ;
  assign y15292 = ~n32965 ;
  assign y15293 = ~n32968 ;
  assign y15294 = n21807 ;
  assign y15295 = ~n32969 ;
  assign y15296 = ~n32970 ;
  assign y15297 = ~n32973 ;
  assign y15298 = n32974 ;
  assign y15299 = ~n32977 ;
  assign y15300 = n32986 ;
  assign y15301 = n20448 ;
  assign y15302 = ~n32987 ;
  assign y15303 = ~1'b0 ;
  assign y15304 = n32990 ;
  assign y15305 = ~n32991 ;
  assign y15306 = ~1'b0 ;
  assign y15307 = n32994 ;
  assign y15308 = n32997 ;
  assign y15309 = ~n33002 ;
  assign y15310 = ~n33004 ;
  assign y15311 = n33005 ;
  assign y15312 = ~1'b0 ;
  assign y15313 = ~1'b0 ;
  assign y15314 = ~n33008 ;
  assign y15315 = n33009 ;
  assign y15316 = ~n33010 ;
  assign y15317 = n33012 ;
  assign y15318 = ~1'b0 ;
  assign y15319 = ~1'b0 ;
  assign y15320 = ~n33019 ;
  assign y15321 = ~n33020 ;
  assign y15322 = ~1'b0 ;
  assign y15323 = n33026 ;
  assign y15324 = ~1'b0 ;
  assign y15325 = ~n33028 ;
  assign y15326 = n33030 ;
  assign y15327 = n33034 ;
  assign y15328 = ~n33035 ;
  assign y15329 = n33036 ;
  assign y15330 = ~n33040 ;
  assign y15331 = ~n33041 ;
  assign y15332 = ~1'b0 ;
  assign y15333 = ~n6570 ;
  assign y15334 = ~n33042 ;
  assign y15335 = ~n33044 ;
  assign y15336 = ~n33049 ;
  assign y15337 = ~n33051 ;
  assign y15338 = 1'b0 ;
  assign y15339 = ~1'b0 ;
  assign y15340 = ~n33060 ;
  assign y15341 = n33062 ;
  assign y15342 = ~n29198 ;
  assign y15343 = ~n33068 ;
  assign y15344 = ~1'b0 ;
  assign y15345 = n33074 ;
  assign y15346 = ~1'b0 ;
  assign y15347 = ~n33075 ;
  assign y15348 = n33081 ;
  assign y15349 = ~1'b0 ;
  assign y15350 = n33082 ;
  assign y15351 = ~1'b0 ;
  assign y15352 = ~n33084 ;
  assign y15353 = n33085 ;
  assign y15354 = n33087 ;
  assign y15355 = ~1'b0 ;
  assign y15356 = ~1'b0 ;
  assign y15357 = n33088 ;
  assign y15358 = ~n33092 ;
  assign y15359 = ~n33095 ;
  assign y15360 = ~n33098 ;
  assign y15361 = n33106 ;
  assign y15362 = n33111 ;
  assign y15363 = ~1'b0 ;
  assign y15364 = ~1'b0 ;
  assign y15365 = n33114 ;
  assign y15366 = n33116 ;
  assign y15367 = ~n33119 ;
  assign y15368 = ~1'b0 ;
  assign y15369 = ~n33121 ;
  assign y15370 = n33123 ;
  assign y15371 = ~1'b0 ;
  assign y15372 = ~1'b0 ;
  assign y15373 = n33126 ;
  assign y15374 = ~1'b0 ;
  assign y15375 = n11292 ;
  assign y15376 = ~1'b0 ;
  assign y15377 = n13947 ;
  assign y15378 = ~n33127 ;
  assign y15379 = ~n33134 ;
  assign y15380 = ~1'b0 ;
  assign y15381 = n33139 ;
  assign y15382 = n33140 ;
  assign y15383 = ~1'b0 ;
  assign y15384 = ~n33143 ;
  assign y15385 = ~n33144 ;
  assign y15386 = n33148 ;
  assign y15387 = ~n33149 ;
  assign y15388 = ~n33150 ;
  assign y15389 = n33152 ;
  assign y15390 = ~1'b0 ;
  assign y15391 = ~n33156 ;
  assign y15392 = ~1'b0 ;
  assign y15393 = n33166 ;
  assign y15394 = n33171 ;
  assign y15395 = ~n33173 ;
  assign y15396 = n33175 ;
  assign y15397 = ~n33177 ;
  assign y15398 = ~n33178 ;
  assign y15399 = n33181 ;
  assign y15400 = ~n33183 ;
  assign y15401 = n33185 ;
  assign y15402 = ~n33187 ;
  assign y15403 = n33190 ;
  assign y15404 = n33197 ;
  assign y15405 = ~n33200 ;
  assign y15406 = n33201 ;
  assign y15407 = n33202 ;
  assign y15408 = n33205 ;
  assign y15409 = ~1'b0 ;
  assign y15410 = ~n33206 ;
  assign y15411 = ~1'b0 ;
  assign y15412 = n33211 ;
  assign y15413 = n33213 ;
  assign y15414 = ~n33215 ;
  assign y15415 = n33217 ;
  assign y15416 = ~1'b0 ;
  assign y15417 = ~n33219 ;
  assign y15418 = ~n33222 ;
  assign y15419 = ~n33224 ;
  assign y15420 = ~n33226 ;
  assign y15421 = n33230 ;
  assign y15422 = ~n33233 ;
  assign y15423 = n33235 ;
  assign y15424 = ~n33238 ;
  assign y15425 = n33240 ;
  assign y15426 = n33243 ;
  assign y15427 = ~n33251 ;
  assign y15428 = n33256 ;
  assign y15429 = n33257 ;
  assign y15430 = ~n33259 ;
  assign y15431 = n33261 ;
  assign y15432 = 1'b0 ;
  assign y15433 = ~1'b0 ;
  assign y15434 = n33264 ;
  assign y15435 = ~n33265 ;
  assign y15436 = ~n33266 ;
  assign y15437 = ~n33271 ;
  assign y15438 = ~n33272 ;
  assign y15439 = n20277 ;
  assign y15440 = n30379 ;
  assign y15441 = 1'b0 ;
  assign y15442 = ~n9452 ;
  assign y15443 = ~n33281 ;
  assign y15444 = ~n33282 ;
  assign y15445 = ~1'b0 ;
  assign y15446 = ~1'b0 ;
  assign y15447 = ~1'b0 ;
  assign y15448 = ~n33284 ;
  assign y15449 = ~n25392 ;
  assign y15450 = ~n33285 ;
  assign y15451 = ~n33287 ;
  assign y15452 = ~1'b0 ;
  assign y15453 = ~1'b0 ;
  assign y15454 = n33292 ;
  assign y15455 = n33294 ;
  assign y15456 = n33296 ;
  assign y15457 = ~1'b0 ;
  assign y15458 = ~n33297 ;
  assign y15459 = ~n33302 ;
  assign y15460 = ~n33306 ;
  assign y15461 = n33310 ;
  assign y15462 = ~1'b0 ;
  assign y15463 = ~n33311 ;
  assign y15464 = ~n33313 ;
  assign y15465 = n29531 ;
  assign y15466 = n33314 ;
  assign y15467 = ~n33315 ;
  assign y15468 = ~n33317 ;
  assign y15469 = ~n33319 ;
  assign y15470 = n33323 ;
  assign y15471 = ~n33324 ;
  assign y15472 = n33327 ;
  assign y15473 = ~1'b0 ;
  assign y15474 = ~n33331 ;
  assign y15475 = n33336 ;
  assign y15476 = n33338 ;
  assign y15477 = ~n33341 ;
  assign y15478 = n33342 ;
  assign y15479 = n33345 ;
  assign y15480 = n33352 ;
  assign y15481 = ~n33354 ;
  assign y15482 = ~n33355 ;
  assign y15483 = ~n30123 ;
  assign y15484 = ~n33358 ;
  assign y15485 = n33360 ;
  assign y15486 = ~1'b0 ;
  assign y15487 = ~n33362 ;
  assign y15488 = ~1'b0 ;
  assign y15489 = ~n33364 ;
  assign y15490 = ~1'b0 ;
  assign y15491 = n33371 ;
  assign y15492 = ~n33373 ;
  assign y15493 = ~1'b0 ;
  assign y15494 = ~1'b0 ;
  assign y15495 = ~n33376 ;
  assign y15496 = ~n33379 ;
  assign y15497 = ~n33380 ;
  assign y15498 = ~n33383 ;
  assign y15499 = n33385 ;
  assign y15500 = ~1'b0 ;
  assign y15501 = ~n33386 ;
  assign y15502 = ~n33387 ;
  assign y15503 = ~n33389 ;
  assign y15504 = n33392 ;
  assign y15505 = n33396 ;
  assign y15506 = ~n33404 ;
  assign y15507 = ~n33407 ;
  assign y15508 = ~n33408 ;
  assign y15509 = ~n33409 ;
  assign y15510 = n33412 ;
  assign y15511 = n29521 ;
  assign y15512 = n33414 ;
  assign y15513 = ~1'b0 ;
  assign y15514 = ~1'b0 ;
  assign y15515 = ~1'b0 ;
  assign y15516 = n33416 ;
  assign y15517 = n33417 ;
  assign y15518 = ~n33419 ;
  assign y15519 = ~1'b0 ;
  assign y15520 = ~1'b0 ;
  assign y15521 = 1'b0 ;
  assign y15522 = ~n7221 ;
  assign y15523 = n33426 ;
  assign y15524 = ~n33433 ;
  assign y15525 = n33434 ;
  assign y15526 = ~n29434 ;
  assign y15527 = ~n33440 ;
  assign y15528 = ~1'b0 ;
  assign y15529 = ~n33446 ;
  assign y15530 = ~n33450 ;
  assign y15531 = ~1'b0 ;
  assign y15532 = n33454 ;
  assign y15533 = ~1'b0 ;
  assign y15534 = ~1'b0 ;
  assign y15535 = n33456 ;
  assign y15536 = ~n33459 ;
  assign y15537 = n33460 ;
  assign y15538 = ~1'b0 ;
  assign y15539 = n33461 ;
  assign y15540 = ~n33463 ;
  assign y15541 = ~1'b0 ;
  assign y15542 = ~1'b0 ;
  assign y15543 = ~n791 ;
  assign y15544 = ~n33467 ;
  assign y15545 = 1'b0 ;
  assign y15546 = ~n33471 ;
  assign y15547 = ~n33473 ;
  assign y15548 = n33474 ;
  assign y15549 = ~n33476 ;
  assign y15550 = ~1'b0 ;
  assign y15551 = ~1'b0 ;
  assign y15552 = n33477 ;
  assign y15553 = ~n33478 ;
  assign y15554 = ~1'b0 ;
  assign y15555 = ~1'b0 ;
  assign y15556 = ~n33479 ;
  assign y15557 = ~n33485 ;
  assign y15558 = ~1'b0 ;
  assign y15559 = ~n33486 ;
  assign y15560 = ~n17005 ;
  assign y15561 = ~1'b0 ;
  assign y15562 = ~n33488 ;
  assign y15563 = n33491 ;
  assign y15564 = ~n33492 ;
  assign y15565 = ~n33493 ;
  assign y15566 = n33499 ;
  assign y15567 = ~1'b0 ;
  assign y15568 = ~1'b0 ;
  assign y15569 = ~n33503 ;
  assign y15570 = 1'b0 ;
  assign y15571 = ~1'b0 ;
  assign y15572 = ~n33505 ;
  assign y15573 = n33509 ;
  assign y15574 = n33512 ;
  assign y15575 = n33517 ;
  assign y15576 = ~1'b0 ;
  assign y15577 = ~1'b0 ;
  assign y15578 = n33518 ;
  assign y15579 = n33521 ;
  assign y15580 = n33524 ;
  assign y15581 = ~n33527 ;
  assign y15582 = ~n33528 ;
  assign y15583 = ~n33531 ;
  assign y15584 = n33532 ;
  assign y15585 = ~n33536 ;
  assign y15586 = 1'b0 ;
  assign y15587 = ~1'b0 ;
  assign y15588 = n33539 ;
  assign y15589 = ~n33540 ;
  assign y15590 = ~n7868 ;
  assign y15591 = n33542 ;
  assign y15592 = ~n33543 ;
  assign y15593 = ~n33545 ;
  assign y15594 = n33546 ;
  assign y15595 = ~1'b0 ;
  assign y15596 = ~n33547 ;
  assign y15597 = ~n33548 ;
  assign y15598 = n33552 ;
  assign y15599 = ~1'b0 ;
  assign y15600 = ~1'b0 ;
  assign y15601 = ~n33555 ;
  assign y15602 = ~1'b0 ;
  assign y15603 = n33556 ;
  assign y15604 = ~n33559 ;
  assign y15605 = ~n33560 ;
  assign y15606 = ~n33562 ;
  assign y15607 = ~1'b0 ;
  assign y15608 = ~n21664 ;
  assign y15609 = ~1'b0 ;
  assign y15610 = n4834 ;
  assign y15611 = ~n33564 ;
  assign y15612 = ~n33566 ;
  assign y15613 = n13077 ;
  assign y15614 = ~n6487 ;
  assign y15615 = n33568 ;
  assign y15616 = ~n33576 ;
  assign y15617 = n33577 ;
  assign y15618 = ~1'b0 ;
  assign y15619 = ~n33587 ;
  assign y15620 = ~n33588 ;
  assign y15621 = ~1'b0 ;
  assign y15622 = ~1'b0 ;
  assign y15623 = ~n33591 ;
  assign y15624 = n33593 ;
  assign y15625 = n33594 ;
  assign y15626 = ~n33600 ;
  assign y15627 = ~n33602 ;
  assign y15628 = ~n33604 ;
  assign y15629 = ~n33606 ;
  assign y15630 = n11290 ;
  assign y15631 = ~n33607 ;
  assign y15632 = ~n33608 ;
  assign y15633 = ~n33610 ;
  assign y15634 = n33611 ;
  assign y15635 = ~1'b0 ;
  assign y15636 = ~n33612 ;
  assign y15637 = ~n33615 ;
  assign y15638 = ~n8418 ;
  assign y15639 = n33616 ;
  assign y15640 = n33618 ;
  assign y15641 = ~1'b0 ;
  assign y15642 = n4729 ;
  assign y15643 = n33619 ;
  assign y15644 = n33621 ;
  assign y15645 = n33626 ;
  assign y15646 = n33627 ;
  assign y15647 = ~n33628 ;
  assign y15648 = ~1'b0 ;
  assign y15649 = ~1'b0 ;
  assign y15650 = ~1'b0 ;
  assign y15651 = ~n33629 ;
  assign y15652 = ~1'b0 ;
  assign y15653 = n33632 ;
  assign y15654 = ~n33634 ;
  assign y15655 = ~n33636 ;
  assign y15656 = ~1'b0 ;
  assign y15657 = ~1'b0 ;
  assign y15658 = n33638 ;
  assign y15659 = ~n33639 ;
  assign y15660 = 1'b0 ;
  assign y15661 = ~n33649 ;
  assign y15662 = n33654 ;
  assign y15663 = ~n33656 ;
  assign y15664 = n33658 ;
  assign y15665 = n33659 ;
  assign y15666 = ~n33661 ;
  assign y15667 = ~n33663 ;
  assign y15668 = n33666 ;
  assign y15669 = ~n33669 ;
  assign y15670 = n33670 ;
  assign y15671 = n33673 ;
  assign y15672 = n33675 ;
  assign y15673 = n33676 ;
  assign y15674 = ~n7183 ;
  assign y15675 = ~1'b0 ;
  assign y15676 = ~1'b0 ;
  assign y15677 = ~1'b0 ;
  assign y15678 = n33680 ;
  assign y15679 = n33682 ;
  assign y15680 = ~n33684 ;
  assign y15681 = n33685 ;
  assign y15682 = n13561 ;
  assign y15683 = 1'b0 ;
  assign y15684 = ~n33687 ;
  assign y15685 = n33691 ;
  assign y15686 = n33692 ;
  assign y15687 = n33693 ;
  assign y15688 = n33694 ;
  assign y15689 = ~1'b0 ;
  assign y15690 = n33700 ;
  assign y15691 = ~1'b0 ;
  assign y15692 = ~n33703 ;
  assign y15693 = ~n33704 ;
  assign y15694 = n33705 ;
  assign y15695 = ~n33707 ;
  assign y15696 = ~n33709 ;
  assign y15697 = ~n33714 ;
  assign y15698 = ~n33717 ;
  assign y15699 = ~n22580 ;
  assign y15700 = n12197 ;
  assign y15701 = ~1'b0 ;
  assign y15702 = n23265 ;
  assign y15703 = n33718 ;
  assign y15704 = ~n33723 ;
  assign y15705 = ~n33730 ;
  assign y15706 = ~1'b0 ;
  assign y15707 = n33735 ;
  assign y15708 = 1'b0 ;
  assign y15709 = ~n33738 ;
  assign y15710 = n33746 ;
  assign y15711 = n33753 ;
  assign y15712 = ~n33762 ;
  assign y15713 = ~n33763 ;
  assign y15714 = ~n33767 ;
  assign y15715 = ~n33773 ;
  assign y15716 = n33782 ;
  assign y15717 = ~1'b0 ;
  assign y15718 = ~n33789 ;
  assign y15719 = ~n33792 ;
  assign y15720 = n33793 ;
  assign y15721 = ~n33796 ;
  assign y15722 = ~n33798 ;
  assign y15723 = ~n33800 ;
  assign y15724 = ~1'b0 ;
  assign y15725 = ~1'b0 ;
  assign y15726 = ~n33801 ;
  assign y15727 = n33804 ;
  assign y15728 = ~1'b0 ;
  assign y15729 = ~1'b0 ;
  assign y15730 = ~n33805 ;
  assign y15731 = ~1'b0 ;
  assign y15732 = 1'b0 ;
  assign y15733 = ~n33806 ;
  assign y15734 = ~n33808 ;
  assign y15735 = ~n33812 ;
  assign y15736 = ~1'b0 ;
  assign y15737 = ~n33814 ;
  assign y15738 = n33815 ;
  assign y15739 = ~1'b0 ;
  assign y15740 = ~1'b0 ;
  assign y15741 = n33816 ;
  assign y15742 = n33817 ;
  assign y15743 = ~n33819 ;
  assign y15744 = ~n33820 ;
  assign y15745 = n33824 ;
  assign y15746 = n33826 ;
  assign y15747 = n33827 ;
  assign y15748 = ~n8319 ;
  assign y15749 = n33828 ;
  assign y15750 = n33830 ;
  assign y15751 = ~n33833 ;
  assign y15752 = ~n33837 ;
  assign y15753 = ~1'b0 ;
  assign y15754 = ~1'b0 ;
  assign y15755 = n33838 ;
  assign y15756 = n33845 ;
  assign y15757 = ~n33851 ;
  assign y15758 = ~1'b0 ;
  assign y15759 = ~n33854 ;
  assign y15760 = ~n33857 ;
  assign y15761 = n33864 ;
  assign y15762 = ~n33868 ;
  assign y15763 = ~1'b0 ;
  assign y15764 = n33871 ;
  assign y15765 = ~1'b0 ;
  assign y15766 = n33874 ;
  assign y15767 = ~1'b0 ;
  assign y15768 = ~1'b0 ;
  assign y15769 = ~n33876 ;
  assign y15770 = ~n33878 ;
  assign y15771 = ~1'b0 ;
  assign y15772 = ~1'b0 ;
  assign y15773 = n33884 ;
  assign y15774 = ~1'b0 ;
  assign y15775 = ~n33886 ;
  assign y15776 = ~n33887 ;
  assign y15777 = ~1'b0 ;
  assign y15778 = n33889 ;
  assign y15779 = ~n33892 ;
  assign y15780 = ~1'b0 ;
  assign y15781 = n33895 ;
  assign y15782 = ~n33902 ;
  assign y15783 = ~n33903 ;
  assign y15784 = n15815 ;
  assign y15785 = ~1'b0 ;
  assign y15786 = ~1'b0 ;
  assign y15787 = ~n33907 ;
  assign y15788 = ~n33908 ;
  assign y15789 = n33911 ;
  assign y15790 = ~n33914 ;
  assign y15791 = ~n33915 ;
  assign y15792 = n33921 ;
  assign y15793 = n33925 ;
  assign y15794 = n33926 ;
  assign y15795 = ~n9357 ;
  assign y15796 = n33935 ;
  assign y15797 = n33937 ;
  assign y15798 = n33940 ;
  assign y15799 = n10217 ;
  assign y15800 = ~1'b0 ;
  assign y15801 = n33943 ;
  assign y15802 = n33944 ;
  assign y15803 = ~n33945 ;
  assign y15804 = ~n33946 ;
  assign y15805 = ~n33952 ;
  assign y15806 = n33954 ;
  assign y15807 = n33959 ;
  assign y15808 = n23 ;
  assign y15809 = n33964 ;
  assign y15810 = n33966 ;
  assign y15811 = ~1'b0 ;
  assign y15812 = ~n33967 ;
  assign y15813 = ~n33969 ;
  assign y15814 = ~n33971 ;
  assign y15815 = ~n33972 ;
  assign y15816 = n33974 ;
  assign y15817 = ~n33975 ;
  assign y15818 = ~n33976 ;
  assign y15819 = ~1'b0 ;
  assign y15820 = ~n33978 ;
  assign y15821 = n33981 ;
  assign y15822 = ~n6844 ;
  assign y15823 = n33982 ;
  assign y15824 = n33983 ;
  assign y15825 = ~1'b0 ;
  assign y15826 = ~1'b0 ;
  assign y15827 = n33985 ;
  assign y15828 = n33987 ;
  assign y15829 = n33989 ;
  assign y15830 = ~n33990 ;
  assign y15831 = ~n33992 ;
  assign y15832 = n33995 ;
  assign y15833 = n33997 ;
  assign y15834 = ~1'b0 ;
  assign y15835 = n33999 ;
  assign y15836 = 1'b0 ;
  assign y15837 = ~n23036 ;
  assign y15838 = ~n34003 ;
  assign y15839 = n34006 ;
  assign y15840 = n34009 ;
  assign y15841 = ~1'b0 ;
  assign y15842 = ~1'b0 ;
  assign y15843 = ~1'b0 ;
  assign y15844 = ~n34012 ;
  assign y15845 = n34014 ;
  assign y15846 = ~1'b0 ;
  assign y15847 = n34017 ;
  assign y15848 = ~n34020 ;
  assign y15849 = n34023 ;
  assign y15850 = n3307 ;
  assign y15851 = ~n34025 ;
  assign y15852 = ~n34026 ;
  assign y15853 = n34030 ;
  assign y15854 = n34031 ;
  assign y15855 = ~n34033 ;
  assign y15856 = ~n34034 ;
  assign y15857 = n34038 ;
  assign y15858 = ~1'b0 ;
  assign y15859 = ~1'b0 ;
  assign y15860 = ~1'b0 ;
  assign y15861 = ~1'b0 ;
  assign y15862 = ~n34039 ;
  assign y15863 = 1'b0 ;
  assign y15864 = ~n34044 ;
  assign y15865 = n34047 ;
  assign y15866 = ~1'b0 ;
  assign y15867 = ~1'b0 ;
  assign y15868 = ~n34048 ;
  assign y15869 = n34049 ;
  assign y15870 = ~1'b0 ;
  assign y15871 = ~1'b0 ;
  assign y15872 = n34052 ;
  assign y15873 = n34053 ;
  assign y15874 = n34055 ;
  assign y15875 = ~n34057 ;
  assign y15876 = n34060 ;
  assign y15877 = ~n34062 ;
  assign y15878 = ~1'b0 ;
  assign y15879 = ~1'b0 ;
  assign y15880 = ~1'b0 ;
  assign y15881 = ~1'b0 ;
  assign y15882 = n34063 ;
  assign y15883 = n34064 ;
  assign y15884 = ~n34065 ;
  assign y15885 = ~n17042 ;
  assign y15886 = n34071 ;
  assign y15887 = 1'b0 ;
  assign y15888 = ~1'b0 ;
  assign y15889 = ~n34074 ;
  assign y15890 = ~1'b0 ;
  assign y15891 = ~1'b0 ;
  assign y15892 = ~n34075 ;
  assign y15893 = ~n34081 ;
  assign y15894 = ~1'b0 ;
  assign y15895 = ~1'b0 ;
  assign y15896 = ~n34083 ;
  assign y15897 = ~n34086 ;
  assign y15898 = n34090 ;
  assign y15899 = n34091 ;
  assign y15900 = ~1'b0 ;
  assign y15901 = n34092 ;
  assign y15902 = n34094 ;
  assign y15903 = ~n34099 ;
  assign y15904 = ~1'b0 ;
  assign y15905 = ~n34102 ;
  assign y15906 = n34103 ;
  assign y15907 = ~n34104 ;
  assign y15908 = n10587 ;
  assign y15909 = n34105 ;
  assign y15910 = ~n34106 ;
  assign y15911 = ~1'b0 ;
  assign y15912 = n34107 ;
  assign y15913 = ~n34109 ;
  assign y15914 = ~1'b0 ;
  assign y15915 = n34113 ;
  assign y15916 = n34116 ;
  assign y15917 = ~n34117 ;
  assign y15918 = ~1'b0 ;
  assign y15919 = n34118 ;
  assign y15920 = ~n34124 ;
  assign y15921 = ~n34133 ;
  assign y15922 = n34134 ;
  assign y15923 = n34138 ;
  assign y15924 = n34139 ;
  assign y15925 = n34141 ;
  assign y15926 = n34142 ;
  assign y15927 = ~1'b0 ;
  assign y15928 = ~n34147 ;
  assign y15929 = n34149 ;
  assign y15930 = n34151 ;
  assign y15931 = ~n34153 ;
  assign y15932 = ~n34154 ;
  assign y15933 = ~n34155 ;
  assign y15934 = ~1'b0 ;
  assign y15935 = ~1'b0 ;
  assign y15936 = n34159 ;
  assign y15937 = n34161 ;
  assign y15938 = ~1'b0 ;
  assign y15939 = ~1'b0 ;
  assign y15940 = n34165 ;
  assign y15941 = ~n3762 ;
  assign y15942 = n34167 ;
  assign y15943 = n34169 ;
  assign y15944 = ~n34171 ;
  assign y15945 = ~1'b0 ;
  assign y15946 = n34172 ;
  assign y15947 = ~n34176 ;
  assign y15948 = n11871 ;
  assign y15949 = ~1'b0 ;
  assign y15950 = ~1'b0 ;
  assign y15951 = ~1'b0 ;
  assign y15952 = n34177 ;
  assign y15953 = ~1'b0 ;
  assign y15954 = ~n34179 ;
  assign y15955 = n34183 ;
  assign y15956 = ~1'b0 ;
  assign y15957 = ~1'b0 ;
  assign y15958 = ~1'b0 ;
  assign y15959 = ~1'b0 ;
  assign y15960 = ~1'b0 ;
  assign y15961 = n34185 ;
  assign y15962 = ~1'b0 ;
  assign y15963 = ~1'b0 ;
  assign y15964 = ~n34187 ;
  assign y15965 = ~n34189 ;
  assign y15966 = ~n34190 ;
  assign y15967 = ~n34191 ;
  assign y15968 = ~n34193 ;
  assign y15969 = n34195 ;
  assign y15970 = ~1'b0 ;
  assign y15971 = n3552 ;
  assign y15972 = n25603 ;
  assign y15973 = ~n34196 ;
  assign y15974 = n34198 ;
  assign y15975 = n34202 ;
  assign y15976 = n34204 ;
  assign y15977 = ~n34209 ;
  assign y15978 = ~n34211 ;
  assign y15979 = ~1'b0 ;
  assign y15980 = n34214 ;
  assign y15981 = n34216 ;
  assign y15982 = n34220 ;
  assign y15983 = n34222 ;
  assign y15984 = ~1'b0 ;
  assign y15985 = ~n34224 ;
  assign y15986 = ~n34225 ;
  assign y15987 = n34227 ;
  assign y15988 = ~n6618 ;
  assign y15989 = ~n34228 ;
  assign y15990 = ~1'b0 ;
  assign y15991 = ~n34234 ;
  assign y15992 = n34237 ;
  assign y15993 = ~n34239 ;
  assign y15994 = ~n34241 ;
  assign y15995 = ~1'b0 ;
  assign y15996 = ~n34242 ;
  assign y15997 = ~n34244 ;
  assign y15998 = ~1'b0 ;
  assign y15999 = ~1'b0 ;
  assign y16000 = 1'b0 ;
  assign y16001 = ~1'b0 ;
  assign y16002 = ~1'b0 ;
  assign y16003 = ~n34247 ;
  assign y16004 = ~n34253 ;
  assign y16005 = ~n34255 ;
  assign y16006 = ~n34256 ;
  assign y16007 = ~n34258 ;
  assign y16008 = ~1'b0 ;
  assign y16009 = ~n18679 ;
  assign y16010 = ~n34269 ;
  assign y16011 = n34270 ;
  assign y16012 = n34276 ;
  assign y16013 = 1'b0 ;
  assign y16014 = ~n34280 ;
  assign y16015 = ~n34285 ;
  assign y16016 = n34287 ;
  assign y16017 = n34289 ;
  assign y16018 = ~1'b0 ;
  assign y16019 = ~n34294 ;
  assign y16020 = n22330 ;
  assign y16021 = ~1'b0 ;
  assign y16022 = n22427 ;
  assign y16023 = ~n34296 ;
  assign y16024 = ~n34300 ;
  assign y16025 = ~1'b0 ;
  assign y16026 = ~n34301 ;
  assign y16027 = ~n34309 ;
  assign y16028 = n34310 ;
  assign y16029 = ~n34313 ;
  assign y16030 = ~1'b0 ;
  assign y16031 = ~n34316 ;
  assign y16032 = ~1'b0 ;
  assign y16033 = ~n34322 ;
  assign y16034 = ~n34324 ;
  assign y16035 = ~n34328 ;
  assign y16036 = ~n34330 ;
  assign y16037 = ~n34333 ;
  assign y16038 = n34336 ;
  assign y16039 = ~n34340 ;
  assign y16040 = ~n34342 ;
  assign y16041 = ~n34350 ;
  assign y16042 = ~n34354 ;
  assign y16043 = n34359 ;
  assign y16044 = n34360 ;
  assign y16045 = n34362 ;
  assign y16046 = ~n34365 ;
  assign y16047 = ~n34368 ;
  assign y16048 = ~1'b0 ;
  assign y16049 = n34370 ;
  assign y16050 = n34371 ;
  assign y16051 = ~1'b0 ;
  assign y16052 = n34375 ;
  assign y16053 = ~1'b0 ;
  assign y16054 = n34380 ;
  assign y16055 = n34381 ;
  assign y16056 = n34382 ;
  assign y16057 = ~n34384 ;
  assign y16058 = ~n34385 ;
  assign y16059 = ~1'b0 ;
  assign y16060 = n34386 ;
  assign y16061 = n34388 ;
  assign y16062 = n34392 ;
  assign y16063 = ~n34394 ;
  assign y16064 = ~n34396 ;
  assign y16065 = ~1'b0 ;
  assign y16066 = n34400 ;
  assign y16067 = ~n16197 ;
  assign y16068 = ~n34401 ;
  assign y16069 = ~n34402 ;
  assign y16070 = n34404 ;
  assign y16071 = n34409 ;
  assign y16072 = ~1'b0 ;
  assign y16073 = ~n34415 ;
  assign y16074 = ~n34420 ;
  assign y16075 = n34421 ;
  assign y16076 = n34422 ;
  assign y16077 = ~1'b0 ;
  assign y16078 = ~n34428 ;
  assign y16079 = n34430 ;
  assign y16080 = ~n34433 ;
  assign y16081 = ~n34434 ;
  assign y16082 = ~n34436 ;
  assign y16083 = ~1'b0 ;
  assign y16084 = ~1'b0 ;
  assign y16085 = ~n34437 ;
  assign y16086 = ~1'b0 ;
  assign y16087 = ~1'b0 ;
  assign y16088 = ~n34439 ;
  assign y16089 = ~n23610 ;
  assign y16090 = ~1'b0 ;
  assign y16091 = ~n34441 ;
  assign y16092 = n34446 ;
  assign y16093 = ~n34451 ;
  assign y16094 = ~n34452 ;
  assign y16095 = ~1'b0 ;
  assign y16096 = ~n34457 ;
  assign y16097 = n34458 ;
  assign y16098 = ~n34459 ;
  assign y16099 = ~1'b0 ;
  assign y16100 = n34465 ;
  assign y16101 = ~1'b0 ;
  assign y16102 = n34467 ;
  assign y16103 = ~n34475 ;
  assign y16104 = n34476 ;
  assign y16105 = n34477 ;
  assign y16106 = ~n34478 ;
  assign y16107 = ~n34480 ;
  assign y16108 = ~1'b0 ;
  assign y16109 = n34484 ;
  assign y16110 = ~1'b0 ;
  assign y16111 = n34485 ;
  assign y16112 = ~n34491 ;
  assign y16113 = n34492 ;
  assign y16114 = ~n34495 ;
  assign y16115 = ~1'b0 ;
  assign y16116 = n13426 ;
  assign y16117 = n34497 ;
  assign y16118 = ~n34498 ;
  assign y16119 = ~1'b0 ;
  assign y16120 = ~n34501 ;
  assign y16121 = ~1'b0 ;
  assign y16122 = n34502 ;
  assign y16123 = ~1'b0 ;
  assign y16124 = ~1'b0 ;
  assign y16125 = ~n34505 ;
  assign y16126 = ~1'b0 ;
  assign y16127 = n34514 ;
  assign y16128 = ~1'b0 ;
  assign y16129 = n34517 ;
  assign y16130 = n34520 ;
  assign y16131 = n34526 ;
  assign y16132 = n34531 ;
  assign y16133 = ~1'b0 ;
  assign y16134 = n34532 ;
  assign y16135 = n34533 ;
  assign y16136 = ~n34534 ;
  assign y16137 = ~n34538 ;
  assign y16138 = n34539 ;
  assign y16139 = ~1'b0 ;
  assign y16140 = ~n34543 ;
  assign y16141 = ~n34549 ;
  assign y16142 = n34553 ;
  assign y16143 = ~1'b0 ;
  assign y16144 = ~n34557 ;
  assign y16145 = ~n34559 ;
  assign y16146 = ~1'b0 ;
  assign y16147 = ~1'b0 ;
  assign y16148 = n34565 ;
  assign y16149 = ~n34568 ;
  assign y16150 = ~n34570 ;
  assign y16151 = ~n34573 ;
  assign y16152 = ~1'b0 ;
  assign y16153 = ~n34575 ;
  assign y16154 = ~1'b0 ;
  assign y16155 = ~n34579 ;
  assign y16156 = n34580 ;
  assign y16157 = ~n34583 ;
  assign y16158 = ~n34584 ;
  assign y16159 = ~1'b0 ;
  assign y16160 = ~n34585 ;
  assign y16161 = ~n34587 ;
  assign y16162 = n34592 ;
  assign y16163 = ~1'b0 ;
  assign y16164 = ~n34594 ;
  assign y16165 = ~1'b0 ;
  assign y16166 = ~1'b0 ;
  assign y16167 = n34597 ;
  assign y16168 = n34599 ;
  assign y16169 = n34602 ;
  assign y16170 = ~n34604 ;
  assign y16171 = n34608 ;
  assign y16172 = ~n34610 ;
  assign y16173 = n34616 ;
  assign y16174 = ~n34618 ;
  assign y16175 = n34623 ;
  assign y16176 = ~n34626 ;
  assign y16177 = ~n34628 ;
  assign y16178 = ~n34632 ;
  assign y16179 = n34636 ;
  assign y16180 = n34637 ;
  assign y16181 = ~1'b0 ;
  assign y16182 = n27319 ;
  assign y16183 = ~n34639 ;
  assign y16184 = ~n34641 ;
  assign y16185 = ~n25068 ;
  assign y16186 = ~1'b0 ;
  assign y16187 = ~1'b0 ;
  assign y16188 = ~1'b0 ;
  assign y16189 = ~1'b0 ;
  assign y16190 = n14590 ;
  assign y16191 = ~n34644 ;
  assign y16192 = n34648 ;
  assign y16193 = n18688 ;
  assign y16194 = ~n34650 ;
  assign y16195 = ~n34651 ;
  assign y16196 = n34653 ;
  assign y16197 = 1'b0 ;
  assign y16198 = n34654 ;
  assign y16199 = ~n34661 ;
  assign y16200 = ~1'b0 ;
  assign y16201 = ~n34668 ;
  assign y16202 = ~1'b0 ;
  assign y16203 = n34670 ;
  assign y16204 = n34671 ;
  assign y16205 = ~n34675 ;
  assign y16206 = ~n34682 ;
  assign y16207 = ~n34683 ;
  assign y16208 = n34691 ;
  assign y16209 = ~1'b0 ;
  assign y16210 = ~n34694 ;
  assign y16211 = n34699 ;
  assign y16212 = ~n34701 ;
  assign y16213 = ~n9197 ;
  assign y16214 = n34703 ;
  assign y16215 = n34711 ;
  assign y16216 = ~n34715 ;
  assign y16217 = ~n34716 ;
  assign y16218 = n34719 ;
  assign y16219 = ~1'b0 ;
  assign y16220 = ~n34722 ;
  assign y16221 = n34726 ;
  assign y16222 = ~1'b0 ;
  assign y16223 = n34731 ;
  assign y16224 = ~n4983 ;
  assign y16225 = ~n34736 ;
  assign y16226 = ~n34737 ;
  assign y16227 = n34739 ;
  assign y16228 = ~1'b0 ;
  assign y16229 = n34740 ;
  assign y16230 = ~n34742 ;
  assign y16231 = ~n34744 ;
  assign y16232 = ~n34747 ;
  assign y16233 = ~n34749 ;
  assign y16234 = ~n34750 ;
  assign y16235 = ~n34752 ;
  assign y16236 = 1'b0 ;
  assign y16237 = 1'b0 ;
  assign y16238 = n34754 ;
  assign y16239 = n34759 ;
  assign y16240 = ~1'b0 ;
  assign y16241 = n34762 ;
  assign y16242 = ~1'b0 ;
  assign y16243 = ~1'b0 ;
  assign y16244 = n34763 ;
  assign y16245 = ~n34765 ;
  assign y16246 = n34769 ;
  assign y16247 = n34773 ;
  assign y16248 = ~n34774 ;
  assign y16249 = ~1'b0 ;
  assign y16250 = n34778 ;
  assign y16251 = n34780 ;
  assign y16252 = ~n34784 ;
  assign y16253 = n34786 ;
  assign y16254 = n34787 ;
  assign y16255 = n34797 ;
  assign y16256 = ~n34799 ;
  assign y16257 = ~n34800 ;
  assign y16258 = ~n34808 ;
  assign y16259 = ~1'b0 ;
  assign y16260 = ~n34810 ;
  assign y16261 = ~1'b0 ;
  assign y16262 = n34815 ;
  assign y16263 = ~n34816 ;
  assign y16264 = n34817 ;
  assign y16265 = n34818 ;
  assign y16266 = ~n34821 ;
  assign y16267 = ~1'b0 ;
  assign y16268 = ~n34822 ;
  assign y16269 = n34826 ;
  assign y16270 = 1'b0 ;
  assign y16271 = 1'b0 ;
  assign y16272 = ~n34829 ;
  assign y16273 = ~n34831 ;
  assign y16274 = n34832 ;
  assign y16275 = ~1'b0 ;
  assign y16276 = n34833 ;
  assign y16277 = ~1'b0 ;
  assign y16278 = ~n34834 ;
  assign y16279 = ~n34838 ;
  assign y16280 = n34840 ;
  assign y16281 = n10617 ;
  assign y16282 = ~1'b0 ;
  assign y16283 = ~n34841 ;
  assign y16284 = ~1'b0 ;
  assign y16285 = ~1'b0 ;
  assign y16286 = ~1'b0 ;
  assign y16287 = ~1'b0 ;
  assign y16288 = ~1'b0 ;
  assign y16289 = ~n34845 ;
  assign y16290 = n34848 ;
  assign y16291 = n8592 ;
  assign y16292 = ~1'b0 ;
  assign y16293 = ~n34851 ;
  assign y16294 = ~n34852 ;
  assign y16295 = ~n34858 ;
  assign y16296 = n34864 ;
  assign y16297 = ~n34866 ;
  assign y16298 = ~n34869 ;
  assign y16299 = ~1'b0 ;
  assign y16300 = ~n34871 ;
  assign y16301 = n18357 ;
  assign y16302 = n34875 ;
  assign y16303 = ~1'b0 ;
  assign y16304 = n34876 ;
  assign y16305 = ~n34878 ;
  assign y16306 = n34879 ;
  assign y16307 = ~n34882 ;
  assign y16308 = ~n34883 ;
  assign y16309 = n34886 ;
  assign y16310 = ~n34888 ;
  assign y16311 = ~n17384 ;
  assign y16312 = ~n34890 ;
  assign y16313 = n34893 ;
  assign y16314 = n34898 ;
  assign y16315 = n34899 ;
  assign y16316 = ~n34900 ;
  assign y16317 = ~n30297 ;
  assign y16318 = n34904 ;
  assign y16319 = n34907 ;
  assign y16320 = ~n34909 ;
  assign y16321 = n34914 ;
  assign y16322 = ~n34918 ;
  assign y16323 = n28307 ;
  assign y16324 = ~n34921 ;
  assign y16325 = n34924 ;
  assign y16326 = n34928 ;
  assign y16327 = 1'b0 ;
  assign y16328 = n10218 ;
  assign y16329 = n34932 ;
  assign y16330 = ~n15870 ;
  assign y16331 = ~1'b0 ;
  assign y16332 = ~1'b0 ;
  assign y16333 = ~n34933 ;
  assign y16334 = ~n34939 ;
  assign y16335 = n34944 ;
  assign y16336 = n34945 ;
  assign y16337 = ~n34946 ;
  assign y16338 = n34950 ;
  assign y16339 = 1'b0 ;
  assign y16340 = n34952 ;
  assign y16341 = ~1'b0 ;
  assign y16342 = 1'b0 ;
  assign y16343 = n25560 ;
  assign y16344 = n34957 ;
  assign y16345 = ~n34961 ;
  assign y16346 = 1'b0 ;
  assign y16347 = ~1'b0 ;
  assign y16348 = ~1'b0 ;
  assign y16349 = ~n34964 ;
  assign y16350 = ~n15627 ;
  assign y16351 = n34967 ;
  assign y16352 = n26363 ;
  assign y16353 = ~n34971 ;
  assign y16354 = ~n34976 ;
  assign y16355 = ~n34979 ;
  assign y16356 = ~n34980 ;
  assign y16357 = ~1'b0 ;
  assign y16358 = n34983 ;
  assign y16359 = n34984 ;
  assign y16360 = ~1'b0 ;
  assign y16361 = n34986 ;
  assign y16362 = ~n34988 ;
  assign y16363 = ~n34992 ;
  assign y16364 = ~1'b0 ;
  assign y16365 = n34999 ;
  assign y16366 = n35002 ;
  assign y16367 = ~n35003 ;
  assign y16368 = n17737 ;
  assign y16369 = n35012 ;
  assign y16370 = n35014 ;
  assign y16371 = n35017 ;
  assign y16372 = ~n35020 ;
  assign y16373 = n35024 ;
  assign y16374 = ~n35025 ;
  assign y16375 = ~1'b0 ;
  assign y16376 = n35027 ;
  assign y16377 = ~n35031 ;
  assign y16378 = n35032 ;
  assign y16379 = ~n35033 ;
  assign y16380 = ~n35037 ;
  assign y16381 = n35038 ;
  assign y16382 = n29746 ;
  assign y16383 = n35043 ;
  assign y16384 = ~n35044 ;
  assign y16385 = n6286 ;
  assign y16386 = ~1'b0 ;
  assign y16387 = ~n35047 ;
  assign y16388 = n35050 ;
  assign y16389 = n35051 ;
  assign y16390 = ~n2785 ;
  assign y16391 = ~1'b0 ;
  assign y16392 = ~n35053 ;
  assign y16393 = ~n35055 ;
  assign y16394 = n35056 ;
  assign y16395 = n35058 ;
  assign y16396 = 1'b0 ;
  assign y16397 = ~1'b0 ;
  assign y16398 = n35061 ;
  assign y16399 = ~1'b0 ;
  assign y16400 = ~1'b0 ;
  assign y16401 = n35065 ;
  assign y16402 = ~n35068 ;
  assign y16403 = n35070 ;
  assign y16404 = n35071 ;
  assign y16405 = ~1'b0 ;
  assign y16406 = ~n35076 ;
  assign y16407 = n35077 ;
  assign y16408 = ~1'b0 ;
  assign y16409 = ~1'b0 ;
  assign y16410 = ~n35078 ;
  assign y16411 = ~1'b0 ;
  assign y16412 = n35081 ;
  assign y16413 = ~1'b0 ;
  assign y16414 = n35083 ;
  assign y16415 = ~n35086 ;
  assign y16416 = ~n8478 ;
  assign y16417 = ~n35090 ;
  assign y16418 = ~n35092 ;
  assign y16419 = n35095 ;
  assign y16420 = n35099 ;
  assign y16421 = n5167 ;
  assign y16422 = ~1'b0 ;
  assign y16423 = n35100 ;
  assign y16424 = n35103 ;
  assign y16425 = ~1'b0 ;
  assign y16426 = ~1'b0 ;
  assign y16427 = n35104 ;
  assign y16428 = ~n35108 ;
  assign y16429 = ~1'b0 ;
  assign y16430 = 1'b0 ;
  assign y16431 = n35115 ;
  assign y16432 = n35119 ;
  assign y16433 = ~n35123 ;
  assign y16434 = ~1'b0 ;
  assign y16435 = ~n35127 ;
  assign y16436 = n35135 ;
  assign y16437 = ~n35140 ;
  assign y16438 = n35141 ;
  assign y16439 = ~1'b0 ;
  assign y16440 = n35148 ;
  assign y16441 = ~n35150 ;
  assign y16442 = ~n35152 ;
  assign y16443 = ~1'b0 ;
  assign y16444 = ~n35154 ;
  assign y16445 = ~n35155 ;
  assign y16446 = n6908 ;
  assign y16447 = n35156 ;
  assign y16448 = ~1'b0 ;
  assign y16449 = n35157 ;
  assign y16450 = ~1'b0 ;
  assign y16451 = n35158 ;
  assign y16452 = n35160 ;
  assign y16453 = ~n25503 ;
  assign y16454 = ~n35165 ;
  assign y16455 = ~n35166 ;
  assign y16456 = n35167 ;
  assign y16457 = ~n10772 ;
  assign y16458 = n35170 ;
  assign y16459 = n35171 ;
  assign y16460 = ~n35179 ;
  assign y16461 = 1'b0 ;
  assign y16462 = ~1'b0 ;
  assign y16463 = ~n35181 ;
  assign y16464 = ~1'b0 ;
  assign y16465 = 1'b0 ;
  assign y16466 = ~n35182 ;
  assign y16467 = n35186 ;
  assign y16468 = ~n35201 ;
  assign y16469 = ~n35206 ;
  assign y16470 = n35208 ;
  assign y16471 = ~1'b0 ;
  assign y16472 = ~n35209 ;
  assign y16473 = ~n35212 ;
  assign y16474 = ~n35217 ;
  assign y16475 = ~n35219 ;
  assign y16476 = n35222 ;
  assign y16477 = n35224 ;
  assign y16478 = ~1'b0 ;
  assign y16479 = n35225 ;
  assign y16480 = ~1'b0 ;
  assign y16481 = ~n35226 ;
  assign y16482 = n35227 ;
  assign y16483 = ~1'b0 ;
  assign y16484 = ~n35233 ;
  assign y16485 = ~1'b0 ;
  assign y16486 = ~n35235 ;
  assign y16487 = n35240 ;
  assign y16488 = n35241 ;
  assign y16489 = n35244 ;
  assign y16490 = n35248 ;
  assign y16491 = ~1'b0 ;
  assign y16492 = n28763 ;
  assign y16493 = n12032 ;
  assign y16494 = ~n13057 ;
  assign y16495 = n35250 ;
  assign y16496 = ~1'b0 ;
  assign y16497 = n35253 ;
  assign y16498 = n35259 ;
  assign y16499 = ~1'b0 ;
  assign y16500 = n35263 ;
  assign y16501 = ~n35268 ;
  assign y16502 = ~n35271 ;
  assign y16503 = n35272 ;
  assign y16504 = ~n35273 ;
  assign y16505 = n35274 ;
  assign y16506 = ~1'b0 ;
  assign y16507 = ~n35276 ;
  assign y16508 = ~1'b0 ;
  assign y16509 = ~n35277 ;
  assign y16510 = n35281 ;
  assign y16511 = n35283 ;
  assign y16512 = ~1'b0 ;
  assign y16513 = n35287 ;
  assign y16514 = n35289 ;
  assign y16515 = n35290 ;
  assign y16516 = ~n35296 ;
  assign y16517 = ~n35299 ;
  assign y16518 = n35303 ;
  assign y16519 = n35304 ;
  assign y16520 = ~1'b0 ;
  assign y16521 = ~n35310 ;
  assign y16522 = ~n35311 ;
  assign y16523 = ~n35317 ;
  assign y16524 = ~1'b0 ;
  assign y16525 = n35319 ;
  assign y16526 = ~n35327 ;
  assign y16527 = n35331 ;
  assign y16528 = ~1'b0 ;
  assign y16529 = ~1'b0 ;
  assign y16530 = ~n35332 ;
  assign y16531 = n35333 ;
  assign y16532 = ~1'b0 ;
  assign y16533 = ~n35337 ;
  assign y16534 = n35338 ;
  assign y16535 = n35342 ;
  assign y16536 = ~n35345 ;
  assign y16537 = ~n35347 ;
  assign y16538 = n35350 ;
  assign y16539 = ~1'b0 ;
  assign y16540 = n35351 ;
  assign y16541 = 1'b0 ;
  assign y16542 = ~1'b0 ;
  assign y16543 = n35352 ;
  assign y16544 = n35353 ;
  assign y16545 = ~1'b0 ;
  assign y16546 = ~1'b0 ;
  assign y16547 = ~1'b0 ;
  assign y16548 = ~1'b0 ;
  assign y16549 = n35354 ;
  assign y16550 = ~n35355 ;
  assign y16551 = ~n35357 ;
  assign y16552 = ~n35361 ;
  assign y16553 = ~1'b0 ;
  assign y16554 = n35362 ;
  assign y16555 = n35363 ;
  assign y16556 = 1'b0 ;
  assign y16557 = n7968 ;
  assign y16558 = n35366 ;
  assign y16559 = ~n35368 ;
  assign y16560 = ~n35369 ;
  assign y16561 = ~n35372 ;
  assign y16562 = ~n16369 ;
  assign y16563 = ~n35373 ;
  assign y16564 = n35381 ;
  assign y16565 = ~n35382 ;
  assign y16566 = n18866 ;
  assign y16567 = ~n35386 ;
  assign y16568 = ~1'b0 ;
  assign y16569 = n35388 ;
  assign y16570 = ~n35389 ;
  assign y16571 = n35391 ;
  assign y16572 = n35393 ;
  assign y16573 = n35398 ;
  assign y16574 = ~n35400 ;
  assign y16575 = ~1'b0 ;
  assign y16576 = n35402 ;
  assign y16577 = ~n35408 ;
  assign y16578 = n35411 ;
  assign y16579 = ~n35412 ;
  assign y16580 = ~n35416 ;
  assign y16581 = ~n35419 ;
  assign y16582 = ~n7343 ;
  assign y16583 = ~n35420 ;
  assign y16584 = n35425 ;
  assign y16585 = ~n35434 ;
  assign y16586 = 1'b0 ;
  assign y16587 = ~n35440 ;
  assign y16588 = n29987 ;
  assign y16589 = n35448 ;
  assign y16590 = n35452 ;
  assign y16591 = ~n35455 ;
  assign y16592 = ~n35456 ;
  assign y16593 = ~1'b0 ;
  assign y16594 = n35461 ;
  assign y16595 = ~n35462 ;
  assign y16596 = ~n35464 ;
  assign y16597 = n35466 ;
  assign y16598 = ~1'b0 ;
  assign y16599 = ~n35468 ;
  assign y16600 = ~1'b0 ;
  assign y16601 = n35469 ;
  assign y16602 = ~n35470 ;
  assign y16603 = ~n35471 ;
  assign y16604 = ~n35473 ;
  assign y16605 = ~1'b0 ;
  assign y16606 = n35474 ;
  assign y16607 = n35477 ;
  assign y16608 = 1'b0 ;
  assign y16609 = ~1'b0 ;
  assign y16610 = ~n35489 ;
  assign y16611 = ~1'b0 ;
  assign y16612 = n35493 ;
  assign y16613 = ~n35494 ;
  assign y16614 = 1'b0 ;
  assign y16615 = ~1'b0 ;
  assign y16616 = ~1'b0 ;
  assign y16617 = ~1'b0 ;
  assign y16618 = ~n35498 ;
  assign y16619 = ~1'b0 ;
  assign y16620 = ~n35502 ;
  assign y16621 = ~n35504 ;
  assign y16622 = n35505 ;
  assign y16623 = ~n35508 ;
  assign y16624 = ~n35510 ;
  assign y16625 = ~n35512 ;
  assign y16626 = ~n35517 ;
  assign y16627 = ~n35518 ;
  assign y16628 = ~n35519 ;
  assign y16629 = ~1'b0 ;
  assign y16630 = ~1'b0 ;
  assign y16631 = n35520 ;
  assign y16632 = ~1'b0 ;
  assign y16633 = ~n35523 ;
  assign y16634 = ~n35524 ;
  assign y16635 = n35526 ;
  assign y16636 = 1'b0 ;
  assign y16637 = ~1'b0 ;
  assign y16638 = ~n2271 ;
  assign y16639 = ~n35528 ;
  assign y16640 = n35529 ;
  assign y16641 = ~n35530 ;
  assign y16642 = n35533 ;
  assign y16643 = n35539 ;
  assign y16644 = ~n35541 ;
  assign y16645 = ~n29685 ;
  assign y16646 = ~n35545 ;
  assign y16647 = n35547 ;
  assign y16648 = n35550 ;
  assign y16649 = ~n35554 ;
  assign y16650 = ~1'b0 ;
  assign y16651 = n5749 ;
  assign y16652 = ~1'b0 ;
  assign y16653 = ~n35561 ;
  assign y16654 = ~n35566 ;
  assign y16655 = ~n24766 ;
  assign y16656 = ~1'b0 ;
  assign y16657 = ~1'b0 ;
  assign y16658 = ~n35568 ;
  assign y16659 = n35570 ;
  assign y16660 = ~n35575 ;
  assign y16661 = ~n35577 ;
  assign y16662 = 1'b0 ;
  assign y16663 = ~1'b0 ;
  assign y16664 = ~n35582 ;
  assign y16665 = ~n35586 ;
  assign y16666 = ~n35587 ;
  assign y16667 = n12123 ;
  assign y16668 = ~n35589 ;
  assign y16669 = ~1'b0 ;
  assign y16670 = ~n35590 ;
  assign y16671 = ~1'b0 ;
  assign y16672 = ~n35596 ;
  assign y16673 = ~n35597 ;
  assign y16674 = ~1'b0 ;
  assign y16675 = ~n35599 ;
  assign y16676 = ~1'b0 ;
  assign y16677 = ~n35604 ;
  assign y16678 = n15838 ;
  assign y16679 = n35606 ;
  assign y16680 = n35607 ;
  assign y16681 = ~n8158 ;
  assign y16682 = n35608 ;
  assign y16683 = n35612 ;
  assign y16684 = n17493 ;
  assign y16685 = n35613 ;
  assign y16686 = n35617 ;
  assign y16687 = n35619 ;
  assign y16688 = ~1'b0 ;
  assign y16689 = n35627 ;
  assign y16690 = ~1'b0 ;
  assign y16691 = ~n35628 ;
  assign y16692 = ~n35629 ;
  assign y16693 = n35634 ;
  assign y16694 = ~n35638 ;
  assign y16695 = ~n35642 ;
  assign y16696 = ~1'b0 ;
  assign y16697 = ~n35643 ;
  assign y16698 = n35644 ;
  assign y16699 = ~n35648 ;
  assign y16700 = ~1'b0 ;
  assign y16701 = n35655 ;
  assign y16702 = n35657 ;
  assign y16703 = n19344 ;
  assign y16704 = n35658 ;
  assign y16705 = ~n6653 ;
  assign y16706 = ~n35662 ;
  assign y16707 = ~n35667 ;
  assign y16708 = ~n6068 ;
  assign y16709 = ~1'b0 ;
  assign y16710 = ~1'b0 ;
  assign y16711 = ~n35668 ;
  assign y16712 = n35670 ;
  assign y16713 = n35673 ;
  assign y16714 = ~n35680 ;
  assign y16715 = n35686 ;
  assign y16716 = ~n15807 ;
  assign y16717 = ~1'b0 ;
  assign y16718 = n35688 ;
  assign y16719 = n35718 ;
  assign y16720 = ~1'b0 ;
  assign y16721 = n35720 ;
  assign y16722 = n35723 ;
  assign y16723 = n35724 ;
  assign y16724 = ~n35725 ;
  assign y16725 = ~1'b0 ;
  assign y16726 = ~n15461 ;
  assign y16727 = ~1'b0 ;
  assign y16728 = n35726 ;
  assign y16729 = n35728 ;
  assign y16730 = n35729 ;
  assign y16731 = ~1'b0 ;
  assign y16732 = ~n35731 ;
  assign y16733 = ~1'b0 ;
  assign y16734 = n35733 ;
  assign y16735 = ~n35735 ;
  assign y16736 = n35736 ;
  assign y16737 = n35738 ;
  assign y16738 = ~1'b0 ;
  assign y16739 = ~1'b0 ;
  assign y16740 = n35744 ;
  assign y16741 = ~1'b0 ;
  assign y16742 = n35749 ;
  assign y16743 = ~n35750 ;
  assign y16744 = n35755 ;
  assign y16745 = ~n35756 ;
  assign y16746 = ~1'b0 ;
  assign y16747 = ~1'b0 ;
  assign y16748 = ~1'b0 ;
  assign y16749 = ~1'b0 ;
  assign y16750 = ~n35758 ;
  assign y16751 = ~n35761 ;
  assign y16752 = ~n35763 ;
  assign y16753 = ~n35765 ;
  assign y16754 = ~n35766 ;
  assign y16755 = n35767 ;
  assign y16756 = ~n35768 ;
  assign y16757 = ~n35769 ;
  assign y16758 = ~n35770 ;
  assign y16759 = ~n35772 ;
  assign y16760 = ~1'b0 ;
  assign y16761 = ~1'b0 ;
  assign y16762 = ~1'b0 ;
  assign y16763 = ~1'b0 ;
  assign y16764 = ~n35773 ;
  assign y16765 = ~1'b0 ;
  assign y16766 = ~n35774 ;
  assign y16767 = ~n35776 ;
  assign y16768 = ~1'b0 ;
  assign y16769 = ~1'b0 ;
  assign y16770 = ~1'b0 ;
  assign y16771 = ~n35777 ;
  assign y16772 = n35779 ;
  assign y16773 = n35781 ;
  assign y16774 = ~n35782 ;
  assign y16775 = ~n35784 ;
  assign y16776 = n35805 ;
  assign y16777 = ~n35808 ;
  assign y16778 = n35810 ;
  assign y16779 = ~1'b0 ;
  assign y16780 = ~n35811 ;
  assign y16781 = ~n35814 ;
  assign y16782 = n35816 ;
  assign y16783 = n35819 ;
  assign y16784 = ~n35821 ;
  assign y16785 = ~n35823 ;
  assign y16786 = n35826 ;
  assign y16787 = ~1'b0 ;
  assign y16788 = ~1'b0 ;
  assign y16789 = ~1'b0 ;
  assign y16790 = ~n35827 ;
  assign y16791 = ~1'b0 ;
  assign y16792 = n35830 ;
  assign y16793 = n35835 ;
  assign y16794 = ~n35837 ;
  assign y16795 = ~1'b0 ;
  assign y16796 = n35839 ;
  assign y16797 = ~n35843 ;
  assign y16798 = ~n35845 ;
  assign y16799 = ~n35849 ;
  assign y16800 = ~n35851 ;
  assign y16801 = n35853 ;
  assign y16802 = 1'b0 ;
  assign y16803 = ~1'b0 ;
  assign y16804 = ~n35856 ;
  assign y16805 = ~n35857 ;
  assign y16806 = ~1'b0 ;
  assign y16807 = ~n35859 ;
  assign y16808 = 1'b0 ;
  assign y16809 = n35862 ;
  assign y16810 = ~n35863 ;
  assign y16811 = n35864 ;
  assign y16812 = n963 ;
  assign y16813 = ~n35867 ;
  assign y16814 = ~1'b0 ;
  assign y16815 = ~1'b0 ;
  assign y16816 = ~n35868 ;
  assign y16817 = ~1'b0 ;
  assign y16818 = n35870 ;
  assign y16819 = ~1'b0 ;
  assign y16820 = ~n35871 ;
  assign y16821 = ~n35874 ;
  assign y16822 = ~1'b0 ;
  assign y16823 = ~n35875 ;
  assign y16824 = ~n35876 ;
  assign y16825 = ~n35879 ;
  assign y16826 = ~n35884 ;
  assign y16827 = ~n35885 ;
  assign y16828 = ~n35889 ;
  assign y16829 = ~1'b0 ;
  assign y16830 = ~1'b0 ;
  assign y16831 = n35890 ;
  assign y16832 = ~1'b0 ;
  assign y16833 = n35891 ;
  assign y16834 = 1'b0 ;
  assign y16835 = n35896 ;
  assign y16836 = ~n35899 ;
  assign y16837 = ~n35900 ;
  assign y16838 = n35901 ;
  assign y16839 = n35902 ;
  assign y16840 = n35905 ;
  assign y16841 = n35908 ;
  assign y16842 = ~n35912 ;
  assign y16843 = ~1'b0 ;
  assign y16844 = n35914 ;
  assign y16845 = n35916 ;
  assign y16846 = ~1'b0 ;
  assign y16847 = ~n35918 ;
  assign y16848 = ~n35921 ;
  assign y16849 = ~1'b0 ;
  assign y16850 = ~1'b0 ;
  assign y16851 = n35922 ;
  assign y16852 = n15024 ;
  assign y16853 = ~n35923 ;
  assign y16854 = n32538 ;
  assign y16855 = ~1'b0 ;
  assign y16856 = ~1'b0 ;
  assign y16857 = ~1'b0 ;
  assign y16858 = n35925 ;
  assign y16859 = 1'b0 ;
  assign y16860 = n35927 ;
  assign y16861 = n16259 ;
  assign y16862 = n35929 ;
  assign y16863 = n35931 ;
  assign y16864 = 1'b0 ;
  assign y16865 = ~n35932 ;
  assign y16866 = ~n35939 ;
  assign y16867 = ~n9036 ;
  assign y16868 = n35943 ;
  assign y16869 = n35948 ;
  assign y16870 = ~1'b0 ;
  assign y16871 = ~1'b0 ;
  assign y16872 = ~n35949 ;
  assign y16873 = ~n35954 ;
  assign y16874 = n35956 ;
  assign y16875 = ~1'b0 ;
  assign y16876 = ~1'b0 ;
  assign y16877 = ~n33273 ;
  assign y16878 = n35957 ;
  assign y16879 = n35962 ;
  assign y16880 = ~n1182 ;
  assign y16881 = ~n35965 ;
  assign y16882 = ~n35966 ;
  assign y16883 = ~n35971 ;
  assign y16884 = n35973 ;
  assign y16885 = n35975 ;
  assign y16886 = n35977 ;
  assign y16887 = ~n35979 ;
  assign y16888 = ~n35980 ;
  assign y16889 = n8304 ;
  assign y16890 = ~n35981 ;
  assign y16891 = n35986 ;
  assign y16892 = ~n35988 ;
  assign y16893 = ~n17623 ;
  assign y16894 = n35991 ;
  assign y16895 = ~n35993 ;
  assign y16896 = n35994 ;
  assign y16897 = ~1'b0 ;
  assign y16898 = n35996 ;
  assign y16899 = ~1'b0 ;
  assign y16900 = n36003 ;
  assign y16901 = n36006 ;
  assign y16902 = ~n36014 ;
  assign y16903 = ~1'b0 ;
  assign y16904 = ~1'b0 ;
  assign y16905 = n36015 ;
  assign y16906 = ~n36020 ;
  assign y16907 = n36023 ;
  assign y16908 = ~1'b0 ;
  assign y16909 = n36025 ;
  assign y16910 = n36027 ;
  assign y16911 = ~n36028 ;
  assign y16912 = ~1'b0 ;
  assign y16913 = ~n36031 ;
  assign y16914 = ~n36033 ;
  assign y16915 = n36040 ;
  assign y16916 = n31130 ;
  assign y16917 = n36044 ;
  assign y16918 = ~n36049 ;
  assign y16919 = n29845 ;
  assign y16920 = n36056 ;
  assign y16921 = ~n1689 ;
  assign y16922 = ~n20385 ;
  assign y16923 = ~n36057 ;
  assign y16924 = ~n36060 ;
  assign y16925 = ~1'b0 ;
  assign y16926 = ~n1713 ;
  assign y16927 = ~n36061 ;
  assign y16928 = ~n34152 ;
  assign y16929 = ~1'b0 ;
  assign y16930 = n36062 ;
  assign y16931 = n36066 ;
  assign y16932 = ~1'b0 ;
  assign y16933 = ~1'b0 ;
  assign y16934 = ~n36068 ;
  assign y16935 = n36070 ;
  assign y16936 = ~n36072 ;
  assign y16937 = ~n16245 ;
  assign y16938 = ~1'b0 ;
  assign y16939 = ~n36073 ;
  assign y16940 = ~n36074 ;
  assign y16941 = ~1'b0 ;
  assign y16942 = n36075 ;
  assign y16943 = ~n36076 ;
  assign y16944 = n36078 ;
  assign y16945 = ~1'b0 ;
  assign y16946 = n36079 ;
  assign y16947 = n36080 ;
  assign y16948 = ~n36082 ;
  assign y16949 = ~1'b0 ;
  assign y16950 = ~1'b0 ;
  assign y16951 = ~n36088 ;
  assign y16952 = n36092 ;
  assign y16953 = ~1'b0 ;
  assign y16954 = n36099 ;
  assign y16955 = n36100 ;
  assign y16956 = n36101 ;
  assign y16957 = n36102 ;
  assign y16958 = ~1'b0 ;
  assign y16959 = ~n36103 ;
  assign y16960 = ~1'b0 ;
  assign y16961 = n36104 ;
  assign y16962 = n36105 ;
  assign y16963 = ~n23946 ;
  assign y16964 = ~n13133 ;
  assign y16965 = ~1'b0 ;
  assign y16966 = ~1'b0 ;
  assign y16967 = ~n36111 ;
  assign y16968 = n36115 ;
  assign y16969 = n36116 ;
  assign y16970 = n26514 ;
  assign y16971 = n36117 ;
  assign y16972 = ~1'b0 ;
  assign y16973 = ~n36119 ;
  assign y16974 = n36121 ;
  assign y16975 = n36124 ;
  assign y16976 = n10274 ;
  assign y16977 = n36127 ;
  assign y16978 = ~n36129 ;
  assign y16979 = ~n36131 ;
  assign y16980 = ~1'b0 ;
  assign y16981 = ~n9528 ;
  assign y16982 = n36132 ;
  assign y16983 = 1'b0 ;
  assign y16984 = ~1'b0 ;
  assign y16985 = n36134 ;
  assign y16986 = ~1'b0 ;
  assign y16987 = ~1'b0 ;
  assign y16988 = n36135 ;
  assign y16989 = ~1'b0 ;
  assign y16990 = ~n36137 ;
  assign y16991 = ~n13567 ;
  assign y16992 = n36139 ;
  assign y16993 = n36142 ;
  assign y16994 = ~n36145 ;
  assign y16995 = ~1'b0 ;
  assign y16996 = ~1'b0 ;
  assign y16997 = ~1'b0 ;
  assign y16998 = ~n36147 ;
  assign y16999 = ~1'b0 ;
  assign y17000 = ~n36148 ;
  assign y17001 = ~n36150 ;
  assign y17002 = n36154 ;
  assign y17003 = n36157 ;
  assign y17004 = ~n36159 ;
  assign y17005 = ~1'b0 ;
  assign y17006 = n36160 ;
  assign y17007 = ~n36161 ;
  assign y17008 = ~1'b0 ;
  assign y17009 = n36167 ;
  assign y17010 = n36168 ;
  assign y17011 = ~n36170 ;
  assign y17012 = ~n36175 ;
  assign y17013 = ~n36177 ;
  assign y17014 = ~n36179 ;
  assign y17015 = ~n32667 ;
  assign y17016 = ~n36181 ;
  assign y17017 = n36183 ;
  assign y17018 = n36184 ;
  assign y17019 = ~n36187 ;
  assign y17020 = ~1'b0 ;
  assign y17021 = 1'b0 ;
  assign y17022 = n36189 ;
  assign y17023 = ~n36190 ;
  assign y17024 = ~n36192 ;
  assign y17025 = ~n36196 ;
  assign y17026 = ~n36197 ;
  assign y17027 = ~n36199 ;
  assign y17028 = n17949 ;
  assign y17029 = ~n36203 ;
  assign y17030 = ~n36204 ;
  assign y17031 = ~n36205 ;
  assign y17032 = ~1'b0 ;
  assign y17033 = n36208 ;
  assign y17034 = ~n36211 ;
  assign y17035 = n36212 ;
  assign y17036 = ~n36214 ;
  assign y17037 = ~n7864 ;
  assign y17038 = ~1'b0 ;
  assign y17039 = n36215 ;
  assign y17040 = ~1'b0 ;
  assign y17041 = ~n36217 ;
  assign y17042 = ~n36220 ;
  assign y17043 = ~1'b0 ;
  assign y17044 = n36223 ;
  assign y17045 = 1'b0 ;
  assign y17046 = ~n36226 ;
  assign y17047 = ~1'b0 ;
  assign y17048 = ~1'b0 ;
  assign y17049 = ~1'b0 ;
  assign y17050 = ~n36236 ;
  assign y17051 = ~n36239 ;
  assign y17052 = n36240 ;
  assign y17053 = n36246 ;
  assign y17054 = n36248 ;
  assign y17055 = n36253 ;
  assign y17056 = ~1'b0 ;
  assign y17057 = ~n36258 ;
  assign y17058 = n36262 ;
  assign y17059 = n36263 ;
  assign y17060 = ~1'b0 ;
  assign y17061 = ~1'b0 ;
  assign y17062 = n36265 ;
  assign y17063 = ~n36270 ;
  assign y17064 = ~n36271 ;
  assign y17065 = ~n36272 ;
  assign y17066 = n772 ;
  assign y17067 = ~n19332 ;
  assign y17068 = ~n36273 ;
  assign y17069 = ~n36275 ;
  assign y17070 = ~n36277 ;
  assign y17071 = ~1'b0 ;
  assign y17072 = ~n36278 ;
  assign y17073 = n36289 ;
  assign y17074 = ~n36290 ;
  assign y17075 = ~1'b0 ;
  assign y17076 = ~1'b0 ;
  assign y17077 = ~n36292 ;
  assign y17078 = n36294 ;
  assign y17079 = ~n36295 ;
  assign y17080 = ~n36297 ;
  assign y17081 = n36298 ;
  assign y17082 = ~n36306 ;
  assign y17083 = ~1'b0 ;
  assign y17084 = ~n22899 ;
  assign y17085 = ~1'b0 ;
  assign y17086 = ~n36307 ;
  assign y17087 = ~n36308 ;
  assign y17088 = ~1'b0 ;
  assign y17089 = ~1'b0 ;
  assign y17090 = ~1'b0 ;
  assign y17091 = ~n36310 ;
  assign y17092 = n36312 ;
  assign y17093 = ~n36315 ;
  assign y17094 = n36319 ;
  assign y17095 = ~n36320 ;
  assign y17096 = ~n36324 ;
  assign y17097 = ~1'b0 ;
  assign y17098 = ~1'b0 ;
  assign y17099 = n36325 ;
  assign y17100 = ~n36330 ;
  assign y17101 = ~n36333 ;
  assign y17102 = ~n36335 ;
  assign y17103 = n36336 ;
  assign y17104 = ~1'b0 ;
  assign y17105 = ~n36341 ;
  assign y17106 = ~1'b0 ;
  assign y17107 = ~n36342 ;
  assign y17108 = ~n36343 ;
  assign y17109 = n36345 ;
  assign y17110 = ~1'b0 ;
  assign y17111 = ~n36350 ;
  assign y17112 = n36353 ;
  assign y17113 = ~1'b0 ;
  assign y17114 = n36355 ;
  assign y17115 = ~n36358 ;
  assign y17116 = ~n36359 ;
  assign y17117 = ~n36365 ;
  assign y17118 = ~n36371 ;
  assign y17119 = n36372 ;
  assign y17120 = ~1'b0 ;
  assign y17121 = n36374 ;
  assign y17122 = ~1'b0 ;
  assign y17123 = ~n36380 ;
  assign y17124 = n36390 ;
  assign y17125 = ~1'b0 ;
  assign y17126 = n36391 ;
  assign y17127 = ~n36394 ;
  assign y17128 = n36396 ;
  assign y17129 = ~n36398 ;
  assign y17130 = ~n36400 ;
  assign y17131 = n36401 ;
  assign y17132 = ~n36402 ;
  assign y17133 = ~n36404 ;
  assign y17134 = ~1'b0 ;
  assign y17135 = ~1'b0 ;
  assign y17136 = n36405 ;
  assign y17137 = n36406 ;
  assign y17138 = ~n36409 ;
  assign y17139 = ~n36410 ;
  assign y17140 = n21628 ;
  assign y17141 = ~n36415 ;
  assign y17142 = ~1'b0 ;
  assign y17143 = ~1'b0 ;
  assign y17144 = n36417 ;
  assign y17145 = ~n36421 ;
  assign y17146 = n36423 ;
  assign y17147 = ~1'b0 ;
  assign y17148 = ~1'b0 ;
  assign y17149 = n36424 ;
  assign y17150 = ~n36431 ;
  assign y17151 = n36439 ;
  assign y17152 = ~1'b0 ;
  assign y17153 = ~n36443 ;
  assign y17154 = ~n36448 ;
  assign y17155 = ~1'b0 ;
  assign y17156 = ~1'b0 ;
  assign y17157 = n36451 ;
  assign y17158 = ~n36452 ;
  assign y17159 = ~n36455 ;
  assign y17160 = n36457 ;
  assign y17161 = ~1'b0 ;
  assign y17162 = ~1'b0 ;
  assign y17163 = ~n36462 ;
  assign y17164 = n36464 ;
  assign y17165 = ~n36465 ;
  assign y17166 = ~1'b0 ;
  assign y17167 = 1'b0 ;
  assign y17168 = n36466 ;
  assign y17169 = ~1'b0 ;
  assign y17170 = ~n36467 ;
  assign y17171 = n36468 ;
  assign y17172 = n36483 ;
  assign y17173 = n36485 ;
  assign y17174 = 1'b0 ;
  assign y17175 = ~1'b0 ;
  assign y17176 = n6825 ;
  assign y17177 = ~n36486 ;
  assign y17178 = ~n36492 ;
  assign y17179 = ~n36496 ;
  assign y17180 = ~n34973 ;
  assign y17181 = ~1'b0 ;
  assign y17182 = n36500 ;
  assign y17183 = ~1'b0 ;
  assign y17184 = ~n36505 ;
  assign y17185 = ~n7238 ;
  assign y17186 = n36506 ;
  assign y17187 = n36508 ;
  assign y17188 = ~n36510 ;
  assign y17189 = ~1'b0 ;
  assign y17190 = ~n36513 ;
  assign y17191 = n36515 ;
  assign y17192 = ~1'b0 ;
  assign y17193 = ~1'b0 ;
  assign y17194 = n36516 ;
  assign y17195 = n36517 ;
  assign y17196 = ~n36520 ;
  assign y17197 = ~1'b0 ;
  assign y17198 = ~1'b0 ;
  assign y17199 = n36521 ;
  assign y17200 = n36523 ;
  assign y17201 = n36524 ;
  assign y17202 = ~1'b0 ;
  assign y17203 = ~1'b0 ;
  assign y17204 = n36525 ;
  assign y17205 = ~1'b0 ;
  assign y17206 = ~1'b0 ;
  assign y17207 = ~1'b0 ;
  assign y17208 = ~n36527 ;
  assign y17209 = n2723 ;
  assign y17210 = ~n36528 ;
  assign y17211 = ~1'b0 ;
  assign y17212 = n36536 ;
  assign y17213 = ~1'b0 ;
  assign y17214 = ~1'b0 ;
  assign y17215 = ~1'b0 ;
  assign y17216 = ~1'b0 ;
  assign y17217 = ~n36539 ;
  assign y17218 = n36540 ;
  assign y17219 = ~n36542 ;
  assign y17220 = ~n36547 ;
  assign y17221 = n36549 ;
  assign y17222 = ~n36553 ;
  assign y17223 = ~n36554 ;
  assign y17224 = 1'b0 ;
  assign y17225 = ~n36555 ;
  assign y17226 = n36556 ;
  assign y17227 = n7237 ;
  assign y17228 = ~n36557 ;
  assign y17229 = n36558 ;
  assign y17230 = n36559 ;
  assign y17231 = n36561 ;
  assign y17232 = 1'b0 ;
  assign y17233 = ~n36562 ;
  assign y17234 = ~n36563 ;
  assign y17235 = ~n36564 ;
  assign y17236 = n36567 ;
  assign y17237 = ~n36569 ;
  assign y17238 = n36572 ;
  assign y17239 = 1'b0 ;
  assign y17240 = ~n36574 ;
  assign y17241 = n36577 ;
  assign y17242 = 1'b0 ;
  assign y17243 = ~n36578 ;
  assign y17244 = n36581 ;
  assign y17245 = n36583 ;
  assign y17246 = n36589 ;
  assign y17247 = n36590 ;
  assign y17248 = n36593 ;
  assign y17249 = ~1'b0 ;
  assign y17250 = ~1'b0 ;
  assign y17251 = n36598 ;
  assign y17252 = n36602 ;
  assign y17253 = n36603 ;
  assign y17254 = ~n36606 ;
  assign y17255 = ~1'b0 ;
  assign y17256 = ~n36611 ;
  assign y17257 = n36613 ;
  assign y17258 = n36617 ;
  assign y17259 = ~n36618 ;
  assign y17260 = n143 ;
  assign y17261 = n36623 ;
  assign y17262 = ~n36630 ;
  assign y17263 = ~n36633 ;
  assign y17264 = n36634 ;
  assign y17265 = ~1'b0 ;
  assign y17266 = n36636 ;
  assign y17267 = ~n36639 ;
  assign y17268 = n36640 ;
  assign y17269 = n36643 ;
  assign y17270 = ~1'b0 ;
  assign y17271 = ~1'b0 ;
  assign y17272 = ~1'b0 ;
  assign y17273 = ~1'b0 ;
  assign y17274 = ~n36648 ;
  assign y17275 = ~n36649 ;
  assign y17276 = n36653 ;
  assign y17277 = ~1'b0 ;
  assign y17278 = n36654 ;
  assign y17279 = ~n36658 ;
  assign y17280 = ~n36660 ;
  assign y17281 = n32823 ;
  assign y17282 = n36669 ;
  assign y17283 = 1'b0 ;
  assign y17284 = ~n36670 ;
  assign y17285 = ~n36672 ;
  assign y17286 = ~n36673 ;
  assign y17287 = ~1'b0 ;
  assign y17288 = ~n36674 ;
  assign y17289 = ~n36676 ;
  assign y17290 = ~1'b0 ;
  assign y17291 = ~n26 ;
  assign y17292 = n36679 ;
  assign y17293 = ~n36682 ;
  assign y17294 = n36687 ;
  assign y17295 = n36688 ;
  assign y17296 = ~n36697 ;
  assign y17297 = n36702 ;
  assign y17298 = n36704 ;
  assign y17299 = ~n36705 ;
  assign y17300 = ~n36708 ;
  assign y17301 = n36711 ;
  assign y17302 = n36715 ;
  assign y17303 = ~n36717 ;
  assign y17304 = ~1'b0 ;
  assign y17305 = ~n36721 ;
  assign y17306 = ~n36722 ;
  assign y17307 = ~n36726 ;
  assign y17308 = ~1'b0 ;
  assign y17309 = ~n36728 ;
  assign y17310 = n36731 ;
  assign y17311 = n3745 ;
  assign y17312 = n36732 ;
  assign y17313 = ~n36733 ;
  assign y17314 = ~n36736 ;
  assign y17315 = ~n36739 ;
  assign y17316 = n36748 ;
  assign y17317 = ~1'b0 ;
  assign y17318 = ~n36749 ;
  assign y17319 = ~n36751 ;
  assign y17320 = ~1'b0 ;
  assign y17321 = ~n36754 ;
  assign y17322 = n36755 ;
  assign y17323 = ~1'b0 ;
  assign y17324 = ~1'b0 ;
  assign y17325 = ~n24205 ;
  assign y17326 = n36759 ;
  assign y17327 = ~n36760 ;
  assign y17328 = n36761 ;
  assign y17329 = ~n31177 ;
  assign y17330 = ~n36762 ;
  assign y17331 = ~n36763 ;
  assign y17332 = ~n36765 ;
  assign y17333 = ~n36766 ;
  assign y17334 = n36769 ;
  assign y17335 = ~n3567 ;
  assign y17336 = n36774 ;
  assign y17337 = ~1'b0 ;
  assign y17338 = n36778 ;
  assign y17339 = ~n36780 ;
  assign y17340 = n36782 ;
  assign y17341 = n36787 ;
  assign y17342 = ~1'b0 ;
  assign y17343 = n36788 ;
  assign y17344 = ~n36793 ;
  assign y17345 = ~1'b0 ;
  assign y17346 = ~n36794 ;
  assign y17347 = ~n36796 ;
  assign y17348 = n36797 ;
  assign y17349 = ~n36798 ;
  assign y17350 = n36799 ;
  assign y17351 = n36802 ;
  assign y17352 = n36804 ;
  assign y17353 = ~1'b0 ;
  assign y17354 = ~n36806 ;
  assign y17355 = n36807 ;
  assign y17356 = n36813 ;
  assign y17357 = n36816 ;
  assign y17358 = n36817 ;
  assign y17359 = ~1'b0 ;
  assign y17360 = ~1'b0 ;
  assign y17361 = ~n36820 ;
  assign y17362 = n1840 ;
  assign y17363 = ~1'b0 ;
  assign y17364 = n36821 ;
  assign y17365 = n36826 ;
  assign y17366 = ~n36827 ;
  assign y17367 = n36831 ;
  assign y17368 = ~n36836 ;
  assign y17369 = n36838 ;
  assign y17370 = n36840 ;
  assign y17371 = ~1'b0 ;
  assign y17372 = n36842 ;
  assign y17373 = ~1'b0 ;
  assign y17374 = ~1'b0 ;
  assign y17375 = ~n36844 ;
  assign y17376 = ~1'b0 ;
  assign y17377 = ~1'b0 ;
  assign y17378 = ~1'b0 ;
  assign y17379 = ~n36845 ;
  assign y17380 = n36849 ;
  assign y17381 = n36851 ;
  assign y17382 = ~n36853 ;
  assign y17383 = ~1'b0 ;
  assign y17384 = ~1'b0 ;
  assign y17385 = ~n36855 ;
  assign y17386 = n36862 ;
  assign y17387 = ~n36865 ;
  assign y17388 = ~n36868 ;
  assign y17389 = n36870 ;
  assign y17390 = n36871 ;
  assign y17391 = ~1'b0 ;
  assign y17392 = ~n36878 ;
  assign y17393 = ~n36879 ;
  assign y17394 = ~1'b0 ;
  assign y17395 = ~n36882 ;
  assign y17396 = n36892 ;
  assign y17397 = ~n36895 ;
  assign y17398 = ~n36900 ;
  assign y17399 = ~n36904 ;
  assign y17400 = 1'b0 ;
  assign y17401 = ~1'b0 ;
  assign y17402 = ~1'b0 ;
  assign y17403 = ~n36910 ;
  assign y17404 = n36912 ;
  assign y17405 = ~1'b0 ;
  assign y17406 = ~n36913 ;
  assign y17407 = n36917 ;
  assign y17408 = n36919 ;
  assign y17409 = ~n11736 ;
  assign y17410 = n36920 ;
  assign y17411 = ~n36925 ;
  assign y17412 = n36927 ;
  assign y17413 = n36931 ;
  assign y17414 = ~1'b0 ;
  assign y17415 = ~1'b0 ;
  assign y17416 = ~n36932 ;
  assign y17417 = n36934 ;
  assign y17418 = ~n36935 ;
  assign y17419 = n36937 ;
  assign y17420 = ~n36939 ;
  assign y17421 = ~n36940 ;
  assign y17422 = n36941 ;
  assign y17423 = ~1'b0 ;
  assign y17424 = n36942 ;
  assign y17425 = ~n36944 ;
  assign y17426 = n36948 ;
  assign y17427 = 1'b0 ;
  assign y17428 = ~n36951 ;
  assign y17429 = n36955 ;
  assign y17430 = ~n36956 ;
  assign y17431 = n36961 ;
  assign y17432 = ~1'b0 ;
  assign y17433 = n36964 ;
  assign y17434 = n36965 ;
  assign y17435 = ~n36966 ;
  assign y17436 = n36967 ;
  assign y17437 = n36974 ;
  assign y17438 = ~n36977 ;
  assign y17439 = ~1'b0 ;
  assign y17440 = n36978 ;
  assign y17441 = ~1'b0 ;
  assign y17442 = n36980 ;
  assign y17443 = ~n36988 ;
  assign y17444 = n36990 ;
  assign y17445 = ~n36993 ;
  assign y17446 = n36994 ;
  assign y17447 = ~n36997 ;
  assign y17448 = ~n37001 ;
  assign y17449 = n37003 ;
  assign y17450 = n37006 ;
  assign y17451 = n37007 ;
  assign y17452 = ~n37011 ;
  assign y17453 = n37012 ;
  assign y17454 = n37014 ;
  assign y17455 = ~n37017 ;
  assign y17456 = ~n37020 ;
  assign y17457 = ~1'b0 ;
  assign y17458 = ~1'b0 ;
  assign y17459 = ~n37023 ;
  assign y17460 = ~n18583 ;
  assign y17461 = n37025 ;
  assign y17462 = ~n37027 ;
  assign y17463 = ~1'b0 ;
  assign y17464 = n37030 ;
  assign y17465 = n5872 ;
  assign y17466 = n37031 ;
  assign y17467 = n37032 ;
  assign y17468 = ~n37041 ;
  assign y17469 = n37042 ;
  assign y17470 = ~1'b0 ;
  assign y17471 = ~1'b0 ;
  assign y17472 = ~n37043 ;
  assign y17473 = ~n37044 ;
  assign y17474 = ~1'b0 ;
  assign y17475 = ~1'b0 ;
  assign y17476 = n37048 ;
  assign y17477 = 1'b0 ;
  assign y17478 = n37049 ;
  assign y17479 = ~1'b0 ;
  assign y17480 = ~1'b0 ;
  assign y17481 = ~n37051 ;
  assign y17482 = ~n37055 ;
  assign y17483 = ~1'b0 ;
  assign y17484 = ~n37057 ;
  assign y17485 = n1894 ;
  assign y17486 = ~n37058 ;
  assign y17487 = ~n37066 ;
  assign y17488 = n37068 ;
  assign y17489 = ~n37070 ;
  assign y17490 = ~n37076 ;
  assign y17491 = ~1'b0 ;
  assign y17492 = ~n37079 ;
  assign y17493 = ~n37082 ;
  assign y17494 = n37083 ;
  assign y17495 = n37084 ;
  assign y17496 = ~n37085 ;
  assign y17497 = ~1'b0 ;
  assign y17498 = ~n37088 ;
  assign y17499 = ~1'b0 ;
  assign y17500 = ~1'b0 ;
  assign y17501 = ~1'b0 ;
  assign y17502 = ~n37091 ;
  assign y17503 = ~n37096 ;
  assign y17504 = ~n37105 ;
  assign y17505 = n37108 ;
  assign y17506 = ~1'b0 ;
  assign y17507 = 1'b0 ;
  assign y17508 = ~n37109 ;
  assign y17509 = ~n37115 ;
  assign y17510 = ~n37116 ;
  assign y17511 = ~1'b0 ;
  assign y17512 = ~1'b0 ;
  assign y17513 = ~1'b0 ;
  assign y17514 = ~1'b0 ;
  assign y17515 = 1'b0 ;
  assign y17516 = ~1'b0 ;
  assign y17517 = n37117 ;
  assign y17518 = n24585 ;
  assign y17519 = n37119 ;
  assign y17520 = ~n37120 ;
  assign y17521 = ~1'b0 ;
  assign y17522 = n37121 ;
  assign y17523 = ~n37123 ;
  assign y17524 = ~n37127 ;
  assign y17525 = ~1'b0 ;
  assign y17526 = n37134 ;
  assign y17527 = n37136 ;
  assign y17528 = n37138 ;
  assign y17529 = ~1'b0 ;
  assign y17530 = ~1'b0 ;
  assign y17531 = ~1'b0 ;
  assign y17532 = ~n37142 ;
  assign y17533 = ~1'b0 ;
  assign y17534 = ~1'b0 ;
  assign y17535 = ~1'b0 ;
  assign y17536 = n37144 ;
  assign y17537 = ~n37147 ;
  assign y17538 = ~n37148 ;
  assign y17539 = ~n37154 ;
  assign y17540 = ~n18748 ;
  assign y17541 = ~n37157 ;
  assign y17542 = ~n37160 ;
  assign y17543 = ~n37166 ;
  assign y17544 = n37171 ;
  assign y17545 = ~n37177 ;
  assign y17546 = n37178 ;
  assign y17547 = n37186 ;
  assign y17548 = ~n37187 ;
  assign y17549 = n37192 ;
  assign y17550 = ~n37194 ;
  assign y17551 = ~n37195 ;
  assign y17552 = n37198 ;
  assign y17553 = ~n37200 ;
  assign y17554 = ~1'b0 ;
  assign y17555 = n37203 ;
  assign y17556 = ~n37205 ;
  assign y17557 = ~1'b0 ;
  assign y17558 = ~n37206 ;
  assign y17559 = ~1'b0 ;
  assign y17560 = n37207 ;
  assign y17561 = ~1'b0 ;
  assign y17562 = ~1'b0 ;
  assign y17563 = n37209 ;
  assign y17564 = n37211 ;
  assign y17565 = ~n37215 ;
  assign y17566 = n37218 ;
  assign y17567 = n25152 ;
  assign y17568 = ~n37219 ;
  assign y17569 = ~n37220 ;
  assign y17570 = n37225 ;
  assign y17571 = ~n12678 ;
  assign y17572 = n24400 ;
  assign y17573 = ~n37226 ;
  assign y17574 = ~1'b0 ;
  assign y17575 = 1'b0 ;
  assign y17576 = ~n37228 ;
  assign y17577 = ~1'b0 ;
  assign y17578 = ~1'b0 ;
  assign y17579 = n37229 ;
  assign y17580 = ~1'b0 ;
  assign y17581 = n37230 ;
  assign y17582 = ~n37232 ;
  assign y17583 = ~n37240 ;
  assign y17584 = n37241 ;
  assign y17585 = n37244 ;
  assign y17586 = n37245 ;
  assign y17587 = n37246 ;
  assign y17588 = n37247 ;
  assign y17589 = ~n37254 ;
  assign y17590 = ~1'b0 ;
  assign y17591 = ~1'b0 ;
  assign y17592 = n37256 ;
  assign y17593 = ~n37260 ;
  assign y17594 = n37261 ;
  assign y17595 = n37264 ;
  assign y17596 = ~n37268 ;
  assign y17597 = n37269 ;
  assign y17598 = ~n37271 ;
  assign y17599 = ~n37276 ;
  assign y17600 = ~n37277 ;
  assign y17601 = ~n37283 ;
  assign y17602 = n37284 ;
  assign y17603 = n4263 ;
  assign y17604 = n24864 ;
  assign y17605 = n37286 ;
  assign y17606 = n37288 ;
  assign y17607 = ~1'b0 ;
  assign y17608 = ~1'b0 ;
  assign y17609 = ~n37290 ;
  assign y17610 = ~1'b0 ;
  assign y17611 = ~1'b0 ;
  assign y17612 = ~n37294 ;
  assign y17613 = ~1'b0 ;
  assign y17614 = ~1'b0 ;
  assign y17615 = n37296 ;
  assign y17616 = n37297 ;
  assign y17617 = ~n37299 ;
  assign y17618 = n37300 ;
  assign y17619 = ~n37302 ;
  assign y17620 = n37304 ;
  assign y17621 = n37306 ;
  assign y17622 = n37308 ;
  assign y17623 = n37315 ;
  assign y17624 = ~n37316 ;
  assign y17625 = ~n37319 ;
  assign y17626 = ~1'b0 ;
  assign y17627 = n37322 ;
  assign y17628 = ~n37323 ;
  assign y17629 = ~1'b0 ;
  assign y17630 = n37326 ;
  assign y17631 = ~n2621 ;
  assign y17632 = ~1'b0 ;
  assign y17633 = 1'b0 ;
  assign y17634 = ~1'b0 ;
  assign y17635 = ~n37330 ;
  assign y17636 = n37334 ;
  assign y17637 = ~n37336 ;
  assign y17638 = ~1'b0 ;
  assign y17639 = ~n37337 ;
  assign y17640 = n2566 ;
  assign y17641 = ~n37344 ;
  assign y17642 = n37346 ;
  assign y17643 = n37353 ;
  assign y17644 = ~n37356 ;
  assign y17645 = n37357 ;
  assign y17646 = ~n37362 ;
  assign y17647 = ~1'b0 ;
  assign y17648 = n37363 ;
  assign y17649 = ~n37364 ;
  assign y17650 = ~n37373 ;
  assign y17651 = n25072 ;
  assign y17652 = n37376 ;
  assign y17653 = ~1'b0 ;
  assign y17654 = ~n37378 ;
  assign y17655 = ~1'b0 ;
  assign y17656 = n37379 ;
  assign y17657 = n37381 ;
  assign y17658 = n37382 ;
  assign y17659 = ~1'b0 ;
  assign y17660 = ~n37385 ;
  assign y17661 = ~1'b0 ;
  assign y17662 = ~n37386 ;
  assign y17663 = n37390 ;
  assign y17664 = ~n29828 ;
  assign y17665 = n37392 ;
  assign y17666 = ~1'b0 ;
  assign y17667 = ~n37397 ;
  assign y17668 = ~n37400 ;
  assign y17669 = ~1'b0 ;
  assign y17670 = ~1'b0 ;
  assign y17671 = ~n37406 ;
  assign y17672 = ~n37410 ;
  assign y17673 = n37412 ;
  assign y17674 = ~n37413 ;
  assign y17675 = ~n37414 ;
  assign y17676 = n37417 ;
  assign y17677 = ~n37418 ;
  assign y17678 = ~n37420 ;
  assign y17679 = n37422 ;
  assign y17680 = ~n6133 ;
  assign y17681 = ~n37424 ;
  assign y17682 = n37425 ;
  assign y17683 = n28086 ;
  assign y17684 = ~n37426 ;
  assign y17685 = ~1'b0 ;
  assign y17686 = ~n37427 ;
  assign y17687 = n37429 ;
  assign y17688 = ~n37432 ;
  assign y17689 = n37437 ;
  assign y17690 = ~n37439 ;
  assign y17691 = n37441 ;
  assign y17692 = ~1'b0 ;
  assign y17693 = n37444 ;
  assign y17694 = ~1'b0 ;
  assign y17695 = n37447 ;
  assign y17696 = ~n37448 ;
  assign y17697 = ~n37451 ;
  assign y17698 = n37455 ;
  assign y17699 = n37456 ;
  assign y17700 = n37460 ;
  assign y17701 = ~n33412 ;
  assign y17702 = ~n37461 ;
  assign y17703 = ~n37463 ;
  assign y17704 = n37465 ;
  assign y17705 = n37468 ;
  assign y17706 = n37469 ;
  assign y17707 = n37470 ;
  assign y17708 = ~n37472 ;
  assign y17709 = n37473 ;
  assign y17710 = ~n37475 ;
  assign y17711 = ~n37476 ;
  assign y17712 = ~1'b0 ;
  assign y17713 = n37477 ;
  assign y17714 = ~n37478 ;
  assign y17715 = ~1'b0 ;
  assign y17716 = ~n37480 ;
  assign y17717 = ~n22286 ;
  assign y17718 = n37482 ;
  assign y17719 = ~n37487 ;
  assign y17720 = n37488 ;
  assign y17721 = n37489 ;
  assign y17722 = n37490 ;
  assign y17723 = ~n37498 ;
  assign y17724 = ~1'b0 ;
  assign y17725 = n37500 ;
  assign y17726 = ~1'b0 ;
  assign y17727 = ~n37505 ;
  assign y17728 = ~n37506 ;
  assign y17729 = n37507 ;
  assign y17730 = n37513 ;
  assign y17731 = ~n37515 ;
  assign y17732 = ~1'b0 ;
  assign y17733 = ~1'b0 ;
  assign y17734 = n37517 ;
  assign y17735 = ~n37518 ;
  assign y17736 = ~n37522 ;
  assign y17737 = ~n37525 ;
  assign y17738 = n37530 ;
  assign y17739 = ~n37533 ;
  assign y17740 = ~1'b0 ;
  assign y17741 = n37535 ;
  assign y17742 = ~n37539 ;
  assign y17743 = ~n37542 ;
  assign y17744 = ~n37543 ;
  assign y17745 = ~1'b0 ;
  assign y17746 = ~1'b0 ;
  assign y17747 = ~1'b0 ;
  assign y17748 = n37545 ;
  assign y17749 = ~1'b0 ;
  assign y17750 = ~1'b0 ;
  assign y17751 = ~n16778 ;
  assign y17752 = ~n37549 ;
  assign y17753 = n260 ;
  assign y17754 = n37550 ;
  assign y17755 = n37552 ;
  assign y17756 = ~n2612 ;
  assign y17757 = ~1'b0 ;
  assign y17758 = ~n37555 ;
  assign y17759 = ~n37558 ;
  assign y17760 = n18778 ;
  assign y17761 = ~n3644 ;
  assign y17762 = ~1'b0 ;
  assign y17763 = ~n37561 ;
  assign y17764 = ~1'b0 ;
  assign y17765 = ~n37564 ;
  assign y17766 = ~n37566 ;
  assign y17767 = n37568 ;
  assign y17768 = n37569 ;
  assign y17769 = ~n37573 ;
  assign y17770 = n37574 ;
  assign y17771 = n37579 ;
  assign y17772 = ~1'b0 ;
  assign y17773 = ~n37580 ;
  assign y17774 = 1'b0 ;
  assign y17775 = n37582 ;
  assign y17776 = n37583 ;
  assign y17777 = n37584 ;
  assign y17778 = ~1'b0 ;
  assign y17779 = ~n34324 ;
  assign y17780 = ~n37586 ;
  assign y17781 = ~1'b0 ;
  assign y17782 = ~n37594 ;
  assign y17783 = ~n37597 ;
  assign y17784 = n37599 ;
  assign y17785 = ~n37603 ;
  assign y17786 = ~n1766 ;
  assign y17787 = ~1'b0 ;
  assign y17788 = n37606 ;
  assign y17789 = ~n37609 ;
  assign y17790 = ~n37612 ;
  assign y17791 = ~1'b0 ;
  assign y17792 = ~n37614 ;
  assign y17793 = n37618 ;
  assign y17794 = n37619 ;
  assign y17795 = ~n37620 ;
  assign y17796 = ~1'b0 ;
  assign y17797 = ~n37624 ;
  assign y17798 = ~n37627 ;
  assign y17799 = ~1'b0 ;
  assign y17800 = ~n37628 ;
  assign y17801 = ~1'b0 ;
  assign y17802 = ~n37631 ;
  assign y17803 = n8159 ;
  assign y17804 = n37634 ;
  assign y17805 = n37637 ;
  assign y17806 = ~1'b0 ;
  assign y17807 = ~1'b0 ;
  assign y17808 = n37641 ;
  assign y17809 = n37642 ;
  assign y17810 = n37643 ;
  assign y17811 = n37644 ;
  assign y17812 = 1'b0 ;
  assign y17813 = ~n37649 ;
  assign y17814 = n37650 ;
  assign y17815 = n37651 ;
  assign y17816 = ~n37653 ;
  assign y17817 = ~n37658 ;
  assign y17818 = n37659 ;
  assign y17819 = n37666 ;
  assign y17820 = ~n37667 ;
  assign y17821 = ~1'b0 ;
  assign y17822 = ~n37673 ;
  assign y17823 = ~n37674 ;
  assign y17824 = n37675 ;
  assign y17825 = n37679 ;
  assign y17826 = n37680 ;
  assign y17827 = n37681 ;
  assign y17828 = n37682 ;
  assign y17829 = ~1'b0 ;
  assign y17830 = ~1'b0 ;
  assign y17831 = ~1'b0 ;
  assign y17832 = ~1'b0 ;
  assign y17833 = ~n20364 ;
  assign y17834 = ~n37686 ;
  assign y17835 = ~n37687 ;
  assign y17836 = ~n37690 ;
  assign y17837 = ~1'b0 ;
  assign y17838 = ~n37692 ;
  assign y17839 = ~1'b0 ;
  assign y17840 = n37693 ;
  assign y17841 = n37695 ;
  assign y17842 = ~n37696 ;
  assign y17843 = ~n37708 ;
  assign y17844 = n37711 ;
  assign y17845 = n37714 ;
  assign y17846 = n37719 ;
  assign y17847 = ~n37720 ;
  assign y17848 = n37722 ;
  assign y17849 = ~n37723 ;
  assign y17850 = n37724 ;
  assign y17851 = n37725 ;
  assign y17852 = ~n37726 ;
  assign y17853 = ~1'b0 ;
  assign y17854 = n37729 ;
  assign y17855 = ~n37735 ;
  assign y17856 = ~n37737 ;
  assign y17857 = ~1'b0 ;
  assign y17858 = ~n37739 ;
  assign y17859 = ~n37740 ;
  assign y17860 = n37741 ;
  assign y17861 = n37747 ;
  assign y17862 = n37750 ;
  assign y17863 = ~n37751 ;
  assign y17864 = ~n37752 ;
  assign y17865 = ~1'b0 ;
  assign y17866 = n32343 ;
  assign y17867 = ~n37754 ;
  assign y17868 = ~1'b0 ;
  assign y17869 = n37756 ;
  assign y17870 = ~n37759 ;
  assign y17871 = ~n37760 ;
  assign y17872 = ~n37765 ;
  assign y17873 = n37767 ;
  assign y17874 = ~1'b0 ;
  assign y17875 = n37769 ;
  assign y17876 = n37770 ;
  assign y17877 = ~1'b0 ;
  assign y17878 = ~n37779 ;
  assign y17879 = 1'b0 ;
  assign y17880 = n7701 ;
  assign y17881 = 1'b0 ;
  assign y17882 = ~1'b0 ;
  assign y17883 = n29942 ;
  assign y17884 = ~n37780 ;
  assign y17885 = ~n37784 ;
  assign y17886 = ~1'b0 ;
  assign y17887 = ~1'b0 ;
  assign y17888 = ~1'b0 ;
  assign y17889 = ~n37788 ;
  assign y17890 = n37789 ;
  assign y17891 = n37790 ;
  assign y17892 = ~n37791 ;
  assign y17893 = n37795 ;
  assign y17894 = ~n37796 ;
  assign y17895 = ~1'b0 ;
  assign y17896 = n37797 ;
  assign y17897 = n37800 ;
  assign y17898 = n9196 ;
  assign y17899 = ~n37804 ;
  assign y17900 = n37805 ;
  assign y17901 = n37807 ;
  assign y17902 = ~1'b0 ;
  assign y17903 = 1'b0 ;
  assign y17904 = ~n37808 ;
  assign y17905 = n3447 ;
  assign y17906 = ~n37810 ;
  assign y17907 = n37812 ;
  assign y17908 = n37814 ;
  assign y17909 = ~1'b0 ;
  assign y17910 = ~n37815 ;
  assign y17911 = ~n37819 ;
  assign y17912 = ~n37820 ;
  assign y17913 = n37821 ;
  assign y17914 = ~n37825 ;
  assign y17915 = n37826 ;
  assign y17916 = 1'b0 ;
  assign y17917 = n37830 ;
  assign y17918 = n37834 ;
  assign y17919 = ~n37837 ;
  assign y17920 = ~n37838 ;
  assign y17921 = ~n37841 ;
  assign y17922 = ~1'b0 ;
  assign y17923 = 1'b0 ;
  assign y17924 = n37842 ;
  assign y17925 = n37844 ;
  assign y17926 = n37846 ;
  assign y17927 = n37848 ;
  assign y17928 = ~n37850 ;
  assign y17929 = n37854 ;
  assign y17930 = ~n37856 ;
  assign y17931 = ~n37858 ;
  assign y17932 = n37860 ;
  assign y17933 = n37865 ;
  assign y17934 = ~n23953 ;
  assign y17935 = ~n37867 ;
  assign y17936 = ~1'b0 ;
  assign y17937 = ~1'b0 ;
  assign y17938 = n37868 ;
  assign y17939 = n37871 ;
  assign y17940 = n37873 ;
  assign y17941 = ~n37874 ;
  assign y17942 = ~1'b0 ;
  assign y17943 = n37878 ;
  assign y17944 = ~1'b0 ;
  assign y17945 = ~1'b0 ;
  assign y17946 = n37882 ;
  assign y17947 = ~n37885 ;
  assign y17948 = ~n37887 ;
  assign y17949 = ~n37888 ;
  assign y17950 = ~n37890 ;
  assign y17951 = ~1'b0 ;
  assign y17952 = ~1'b0 ;
  assign y17953 = ~1'b0 ;
  assign y17954 = ~n37892 ;
  assign y17955 = ~1'b0 ;
  assign y17956 = ~n37893 ;
  assign y17957 = ~1'b0 ;
  assign y17958 = ~1'b0 ;
  assign y17959 = n37894 ;
  assign y17960 = ~n37898 ;
  assign y17961 = ~n37900 ;
  assign y17962 = n556 ;
  assign y17963 = n37905 ;
  assign y17964 = ~1'b0 ;
  assign y17965 = ~n37908 ;
  assign y17966 = n37909 ;
  assign y17967 = ~1'b0 ;
  assign y17968 = n37912 ;
  assign y17969 = ~n37919 ;
  assign y17970 = n37920 ;
  assign y17971 = ~n37923 ;
  assign y17972 = ~n37928 ;
  assign y17973 = ~n37932 ;
  assign y17974 = ~1'b0 ;
  assign y17975 = n37934 ;
  assign y17976 = ~n37935 ;
  assign y17977 = ~n37937 ;
  assign y17978 = ~1'b0 ;
  assign y17979 = n37940 ;
  assign y17980 = n37941 ;
  assign y17981 = ~n37942 ;
  assign y17982 = ~1'b0 ;
  assign y17983 = n37947 ;
  assign y17984 = ~n37949 ;
  assign y17985 = ~1'b0 ;
  assign y17986 = ~n37955 ;
  assign y17987 = ~1'b0 ;
  assign y17988 = n37959 ;
  assign y17989 = n37964 ;
  assign y17990 = n37966 ;
  assign y17991 = ~n37968 ;
  assign y17992 = ~1'b0 ;
  assign y17993 = n37970 ;
  assign y17994 = ~1'b0 ;
  assign y17995 = ~1'b0 ;
  assign y17996 = ~n37974 ;
  assign y17997 = n37976 ;
  assign y17998 = ~n37983 ;
  assign y17999 = ~n37984 ;
  assign y18000 = ~1'b0 ;
  assign y18001 = ~n37986 ;
  assign y18002 = n37990 ;
  assign y18003 = ~1'b0 ;
  assign y18004 = n37991 ;
  assign y18005 = ~1'b0 ;
  assign y18006 = ~n37993 ;
  assign y18007 = n37994 ;
  assign y18008 = ~n37996 ;
  assign y18009 = n38002 ;
  assign y18010 = ~n8242 ;
  assign y18011 = ~n38005 ;
  assign y18012 = ~1'b0 ;
  assign y18013 = n38009 ;
  assign y18014 = ~n38011 ;
  assign y18015 = ~1'b0 ;
  assign y18016 = ~1'b0 ;
  assign y18017 = ~1'b0 ;
  assign y18018 = ~n38013 ;
  assign y18019 = ~n38015 ;
  assign y18020 = n38022 ;
  assign y18021 = ~1'b0 ;
  assign y18022 = ~1'b0 ;
  assign y18023 = ~1'b0 ;
  assign y18024 = n38024 ;
  assign y18025 = ~n38027 ;
  assign y18026 = ~n38032 ;
  assign y18027 = n38034 ;
  assign y18028 = n28760 ;
  assign y18029 = ~n38036 ;
  assign y18030 = ~1'b0 ;
  assign y18031 = ~n38039 ;
  assign y18032 = n38040 ;
  assign y18033 = ~n36899 ;
  assign y18034 = n38041 ;
  assign y18035 = ~n38043 ;
  assign y18036 = ~1'b0 ;
  assign y18037 = ~n38044 ;
  assign y18038 = ~n38047 ;
  assign y18039 = n38049 ;
  assign y18040 = n38055 ;
  assign y18041 = ~1'b0 ;
  assign y18042 = ~1'b0 ;
  assign y18043 = ~1'b0 ;
  assign y18044 = ~n38059 ;
  assign y18045 = ~n38064 ;
  assign y18046 = ~n38066 ;
  assign y18047 = n38068 ;
  assign y18048 = ~1'b0 ;
  assign y18049 = ~n38070 ;
  assign y18050 = n38071 ;
  assign y18051 = n38081 ;
  assign y18052 = ~n1545 ;
  assign y18053 = n38083 ;
  assign y18054 = ~1'b0 ;
  assign y18055 = ~n38087 ;
  assign y18056 = ~n38088 ;
  assign y18057 = ~1'b0 ;
  assign y18058 = ~n38092 ;
  assign y18059 = ~n38096 ;
  assign y18060 = n38098 ;
  assign y18061 = n38099 ;
  assign y18062 = n38101 ;
  assign y18063 = ~n38103 ;
  assign y18064 = ~n11594 ;
  assign y18065 = ~n38107 ;
  assign y18066 = ~n38108 ;
  assign y18067 = n38109 ;
  assign y18068 = n38111 ;
  assign y18069 = ~1'b0 ;
  assign y18070 = ~1'b0 ;
  assign y18071 = ~n38112 ;
  assign y18072 = ~n38113 ;
  assign y18073 = ~n38118 ;
  assign y18074 = n38119 ;
  assign y18075 = ~n11691 ;
  assign y18076 = ~n7631 ;
  assign y18077 = n38120 ;
  assign y18078 = ~1'b0 ;
  assign y18079 = ~n38122 ;
  assign y18080 = n38127 ;
  assign y18081 = ~n38129 ;
  assign y18082 = n38131 ;
  assign y18083 = ~1'b0 ;
  assign y18084 = n38135 ;
  assign y18085 = n38137 ;
  assign y18086 = ~n38138 ;
  assign y18087 = ~n38145 ;
  assign y18088 = ~1'b0 ;
  assign y18089 = ~n38146 ;
  assign y18090 = ~n18720 ;
  assign y18091 = ~1'b0 ;
  assign y18092 = n38149 ;
  assign y18093 = n38150 ;
  assign y18094 = ~1'b0 ;
  assign y18095 = ~n38153 ;
  assign y18096 = ~1'b0 ;
  assign y18097 = ~1'b0 ;
  assign y18098 = ~n38157 ;
  assign y18099 = n38158 ;
  assign y18100 = n38159 ;
  assign y18101 = n38161 ;
  assign y18102 = ~1'b0 ;
  assign y18103 = n38164 ;
  assign y18104 = ~n38165 ;
  assign y18105 = n38169 ;
  assign y18106 = ~n38176 ;
  assign y18107 = ~1'b0 ;
  assign y18108 = n38177 ;
  assign y18109 = 1'b0 ;
  assign y18110 = ~n38179 ;
  assign y18111 = ~1'b0 ;
  assign y18112 = n38180 ;
  assign y18113 = n6105 ;
  assign y18114 = 1'b0 ;
  assign y18115 = n38182 ;
  assign y18116 = ~1'b0 ;
  assign y18117 = ~1'b0 ;
  assign y18118 = n38184 ;
  assign y18119 = ~n38186 ;
  assign y18120 = ~1'b0 ;
  assign y18121 = n38192 ;
  assign y18122 = n38193 ;
  assign y18123 = ~1'b0 ;
  assign y18124 = ~n38196 ;
  assign y18125 = ~1'b0 ;
  assign y18126 = ~1'b0 ;
  assign y18127 = ~n38198 ;
  assign y18128 = n38207 ;
  assign y18129 = ~n38208 ;
  assign y18130 = ~n38212 ;
  assign y18131 = ~n38214 ;
  assign y18132 = ~1'b0 ;
  assign y18133 = 1'b0 ;
  assign y18134 = n38220 ;
  assign y18135 = ~n38222 ;
  assign y18136 = ~n37150 ;
  assign y18137 = ~n38223 ;
  assign y18138 = n38226 ;
  assign y18139 = ~1'b0 ;
  assign y18140 = ~n38229 ;
  assign y18141 = n37788 ;
  assign y18142 = n1853 ;
  assign y18143 = 1'b0 ;
  assign y18144 = ~1'b0 ;
  assign y18145 = ~1'b0 ;
  assign y18146 = ~1'b0 ;
  assign y18147 = ~1'b0 ;
  assign y18148 = ~n38232 ;
  assign y18149 = 1'b0 ;
  assign y18150 = ~n38235 ;
  assign y18151 = ~1'b0 ;
  assign y18152 = n38237 ;
  assign y18153 = ~n38238 ;
  assign y18154 = n38241 ;
  assign y18155 = ~1'b0 ;
  assign y18156 = ~n38243 ;
  assign y18157 = ~1'b0 ;
  assign y18158 = ~n38246 ;
  assign y18159 = ~n38248 ;
  assign y18160 = ~n38252 ;
  assign y18161 = ~1'b0 ;
  assign y18162 = n38255 ;
  assign y18163 = n38256 ;
  assign y18164 = ~1'b0 ;
  assign y18165 = ~1'b0 ;
  assign y18166 = ~1'b0 ;
  assign y18167 = ~n38259 ;
  assign y18168 = n38267 ;
  assign y18169 = ~n38268 ;
  assign y18170 = n38269 ;
  assign y18171 = ~1'b0 ;
  assign y18172 = ~n38272 ;
  assign y18173 = ~n38282 ;
  assign y18174 = ~1'b0 ;
  assign y18175 = n38283 ;
  assign y18176 = n38294 ;
  assign y18177 = ~n38297 ;
  assign y18178 = ~1'b0 ;
  assign y18179 = n38299 ;
  assign y18180 = ~n38302 ;
  assign y18181 = n38306 ;
  assign y18182 = n38313 ;
  assign y18183 = ~n38321 ;
  assign y18184 = ~1'b0 ;
  assign y18185 = ~n38325 ;
  assign y18186 = ~n11558 ;
  assign y18187 = ~1'b0 ;
  assign y18188 = n38329 ;
  assign y18189 = ~n30598 ;
  assign y18190 = ~1'b0 ;
  assign y18191 = n38330 ;
  assign y18192 = ~1'b0 ;
  assign y18193 = n38331 ;
  assign y18194 = ~n38335 ;
  assign y18195 = n38338 ;
  assign y18196 = ~1'b0 ;
  assign y18197 = n38340 ;
  assign y18198 = n38342 ;
  assign y18199 = n38345 ;
  assign y18200 = ~n38349 ;
  assign y18201 = n38350 ;
  assign y18202 = n38358 ;
  assign y18203 = ~1'b0 ;
  assign y18204 = ~n38360 ;
  assign y18205 = ~n38361 ;
  assign y18206 = ~1'b0 ;
  assign y18207 = ~n38363 ;
  assign y18208 = n38364 ;
  assign y18209 = ~n38365 ;
  assign y18210 = n38368 ;
  assign y18211 = ~n32334 ;
  assign y18212 = ~n38370 ;
  assign y18213 = ~1'b0 ;
  assign y18214 = n38373 ;
  assign y18215 = n38375 ;
  assign y18216 = ~n38377 ;
  assign y18217 = n38381 ;
  assign y18218 = n38384 ;
  assign y18219 = ~n38387 ;
  assign y18220 = ~n38391 ;
  assign y18221 = n38395 ;
  assign y18222 = n38396 ;
  assign y18223 = ~1'b0 ;
  assign y18224 = ~n38402 ;
  assign y18225 = n38403 ;
  assign y18226 = ~n38404 ;
  assign y18227 = ~1'b0 ;
  assign y18228 = ~n38407 ;
  assign y18229 = ~n38410 ;
  assign y18230 = n22951 ;
  assign y18231 = ~n38411 ;
  assign y18232 = n38412 ;
  assign y18233 = ~n31401 ;
  assign y18234 = n38416 ;
  assign y18235 = ~n38417 ;
  assign y18236 = n38418 ;
  assign y18237 = ~n38420 ;
  assign y18238 = ~1'b0 ;
  assign y18239 = n4216 ;
  assign y18240 = ~n38423 ;
  assign y18241 = ~n38425 ;
  assign y18242 = ~n38429 ;
  assign y18243 = ~n38430 ;
  assign y18244 = n38433 ;
  assign y18245 = ~n38438 ;
  assign y18246 = n38440 ;
  assign y18247 = ~n38441 ;
  assign y18248 = ~1'b0 ;
  assign y18249 = ~n38443 ;
  assign y18250 = ~1'b0 ;
  assign y18251 = ~1'b0 ;
  assign y18252 = ~n38449 ;
  assign y18253 = ~n38450 ;
  assign y18254 = ~n38452 ;
  assign y18255 = n38453 ;
  assign y18256 = ~n38454 ;
  assign y18257 = n38456 ;
  assign y18258 = ~n38463 ;
  assign y18259 = ~n38465 ;
  assign y18260 = ~1'b0 ;
  assign y18261 = n8536 ;
  assign y18262 = ~1'b0 ;
  assign y18263 = n38466 ;
  assign y18264 = ~1'b0 ;
  assign y18265 = n38467 ;
  assign y18266 = ~n38468 ;
  assign y18267 = n38469 ;
  assign y18268 = ~n38471 ;
  assign y18269 = ~n38473 ;
  assign y18270 = ~n38476 ;
  assign y18271 = ~n38478 ;
  assign y18272 = ~1'b0 ;
  assign y18273 = n38481 ;
  assign y18274 = ~1'b0 ;
  assign y18275 = ~n38483 ;
  assign y18276 = ~n38485 ;
  assign y18277 = ~1'b0 ;
  assign y18278 = ~1'b0 ;
  assign y18279 = ~1'b0 ;
  assign y18280 = n38486 ;
  assign y18281 = n38487 ;
  assign y18282 = ~n38499 ;
  assign y18283 = n11695 ;
  assign y18284 = ~n38507 ;
  assign y18285 = ~n38510 ;
  assign y18286 = 1'b0 ;
  assign y18287 = ~n38511 ;
  assign y18288 = n38515 ;
  assign y18289 = n38518 ;
  assign y18290 = ~n38520 ;
  assign y18291 = ~n38522 ;
  assign y18292 = ~n38523 ;
  assign y18293 = ~n38527 ;
  assign y18294 = n38529 ;
  assign y18295 = ~1'b0 ;
  assign y18296 = n38531 ;
  assign y18297 = n29476 ;
  assign y18298 = ~n38533 ;
  assign y18299 = n38534 ;
  assign y18300 = ~1'b0 ;
  assign y18301 = ~1'b0 ;
  assign y18302 = n38535 ;
  assign y18303 = n38537 ;
  assign y18304 = ~1'b0 ;
  assign y18305 = ~n38540 ;
  assign y18306 = n38542 ;
  assign y18307 = n38545 ;
  assign y18308 = ~n38547 ;
  assign y18309 = n38550 ;
  assign y18310 = ~1'b0 ;
  assign y18311 = ~1'b0 ;
  assign y18312 = n38553 ;
  assign y18313 = ~n38558 ;
  assign y18314 = n38559 ;
  assign y18315 = n38560 ;
  assign y18316 = ~n38565 ;
  assign y18317 = n38571 ;
  assign y18318 = n38573 ;
  assign y18319 = n38575 ;
  assign y18320 = ~1'b0 ;
  assign y18321 = ~n38577 ;
  assign y18322 = ~n38579 ;
  assign y18323 = ~n38583 ;
  assign y18324 = ~n8651 ;
  assign y18325 = ~n38590 ;
  assign y18326 = n38591 ;
  assign y18327 = ~n38594 ;
  assign y18328 = ~n38602 ;
  assign y18329 = ~n38604 ;
  assign y18330 = n38605 ;
  assign y18331 = n38609 ;
  assign y18332 = ~n38611 ;
  assign y18333 = ~n22900 ;
  assign y18334 = ~1'b0 ;
  assign y18335 = ~1'b0 ;
  assign y18336 = ~1'b0 ;
  assign y18337 = n38618 ;
  assign y18338 = ~n11032 ;
  assign y18339 = ~n38620 ;
  assign y18340 = ~n38622 ;
  assign y18341 = n38626 ;
  assign y18342 = ~1'b0 ;
  assign y18343 = n38628 ;
  assign y18344 = ~n38629 ;
  assign y18345 = 1'b0 ;
  assign y18346 = ~n31904 ;
  assign y18347 = ~1'b0 ;
  assign y18348 = ~1'b0 ;
  assign y18349 = ~n38630 ;
  assign y18350 = ~n38633 ;
  assign y18351 = ~1'b0 ;
  assign y18352 = n11078 ;
  assign y18353 = ~1'b0 ;
  assign y18354 = ~1'b0 ;
  assign y18355 = n38635 ;
  assign y18356 = ~n38640 ;
  assign y18357 = ~1'b0 ;
  assign y18358 = ~n9698 ;
  assign y18359 = ~n38644 ;
  assign y18360 = ~1'b0 ;
  assign y18361 = 1'b0 ;
  assign y18362 = n38647 ;
  assign y18363 = ~1'b0 ;
  assign y18364 = n38650 ;
  assign y18365 = ~1'b0 ;
  assign y18366 = n38652 ;
  assign y18367 = n38656 ;
  assign y18368 = ~1'b0 ;
  assign y18369 = ~n38658 ;
  assign y18370 = ~1'b0 ;
  assign y18371 = n38659 ;
  assign y18372 = ~n9012 ;
  assign y18373 = ~1'b0 ;
  assign y18374 = ~1'b0 ;
  assign y18375 = ~1'b0 ;
  assign y18376 = ~n38661 ;
  assign y18377 = n38663 ;
  assign y18378 = ~n38664 ;
  assign y18379 = ~n38670 ;
  assign y18380 = ~1'b0 ;
  assign y18381 = n38673 ;
  assign y18382 = ~1'b0 ;
  assign y18383 = n38675 ;
  assign y18384 = ~1'b0 ;
  assign y18385 = ~1'b0 ;
  assign y18386 = ~1'b0 ;
  assign y18387 = n38678 ;
  assign y18388 = ~1'b0 ;
  assign y18389 = ~1'b0 ;
  assign y18390 = n38680 ;
  assign y18391 = n26214 ;
  assign y18392 = n38681 ;
  assign y18393 = ~1'b0 ;
  assign y18394 = n38685 ;
  assign y18395 = ~n38694 ;
  assign y18396 = ~1'b0 ;
  assign y18397 = ~1'b0 ;
  assign y18398 = n22119 ;
  assign y18399 = ~1'b0 ;
  assign y18400 = n38696 ;
  assign y18401 = n38698 ;
  assign y18402 = ~n38700 ;
  assign y18403 = ~1'b0 ;
  assign y18404 = ~n38702 ;
  assign y18405 = ~1'b0 ;
  assign y18406 = ~n38705 ;
  assign y18407 = ~n38706 ;
  assign y18408 = ~n38707 ;
  assign y18409 = n17310 ;
  assign y18410 = ~1'b0 ;
  assign y18411 = ~n38708 ;
  assign y18412 = ~n38716 ;
  assign y18413 = ~n38718 ;
  assign y18414 = n38722 ;
  assign y18415 = ~1'b0 ;
  assign y18416 = n38729 ;
  assign y18417 = ~n38730 ;
  assign y18418 = n38733 ;
  assign y18419 = ~1'b0 ;
  assign y18420 = ~1'b0 ;
  assign y18421 = ~n38736 ;
  assign y18422 = ~1'b0 ;
  assign y18423 = ~1'b0 ;
  assign y18424 = ~n38737 ;
  assign y18425 = ~n38740 ;
  assign y18426 = ~n38741 ;
  assign y18427 = ~1'b0 ;
  assign y18428 = n38745 ;
  assign y18429 = n954 ;
  assign y18430 = n38746 ;
  assign y18431 = n38747 ;
  assign y18432 = n38748 ;
  assign y18433 = ~n38749 ;
  assign y18434 = n38754 ;
  assign y18435 = ~1'b0 ;
  assign y18436 = ~n38758 ;
  assign y18437 = ~n38759 ;
  assign y18438 = 1'b0 ;
  assign y18439 = ~n38761 ;
  assign y18440 = n38765 ;
  assign y18441 = ~n38773 ;
  assign y18442 = ~1'b0 ;
  assign y18443 = ~n38777 ;
  assign y18444 = ~n33102 ;
  assign y18445 = ~n38778 ;
  assign y18446 = ~n38779 ;
  assign y18447 = ~1'b0 ;
  assign y18448 = ~1'b0 ;
  assign y18449 = ~1'b0 ;
  assign y18450 = n7717 ;
  assign y18451 = ~n38780 ;
  assign y18452 = n14891 ;
  assign y18453 = ~n29747 ;
  assign y18454 = n38782 ;
  assign y18455 = n38783 ;
  assign y18456 = ~n38788 ;
  assign y18457 = ~n38790 ;
  assign y18458 = n38794 ;
  assign y18459 = ~1'b0 ;
  assign y18460 = ~1'b0 ;
  assign y18461 = ~n38798 ;
  assign y18462 = n38800 ;
  assign y18463 = n38807 ;
  assign y18464 = ~n38809 ;
  assign y18465 = ~1'b0 ;
  assign y18466 = ~n38811 ;
  assign y18467 = n38814 ;
  assign y18468 = n38818 ;
  assign y18469 = n38820 ;
  assign y18470 = ~n38822 ;
  assign y18471 = ~n38824 ;
  assign y18472 = ~n6278 ;
  assign y18473 = n38829 ;
  assign y18474 = n38830 ;
  assign y18475 = ~n18069 ;
  assign y18476 = ~n38832 ;
  assign y18477 = n38834 ;
  assign y18478 = ~1'b0 ;
  assign y18479 = ~1'b0 ;
  assign y18480 = n38836 ;
  assign y18481 = n38843 ;
  assign y18482 = ~n38844 ;
  assign y18483 = ~1'b0 ;
  assign y18484 = ~1'b0 ;
  assign y18485 = n38845 ;
  assign y18486 = n38847 ;
  assign y18487 = ~n38851 ;
  assign y18488 = n38857 ;
  assign y18489 = n38861 ;
  assign y18490 = ~1'b0 ;
  assign y18491 = ~1'b0 ;
  assign y18492 = ~n38864 ;
  assign y18493 = ~1'b0 ;
  assign y18494 = n38869 ;
  assign y18495 = ~n38873 ;
  assign y18496 = n38876 ;
  assign y18497 = ~n38878 ;
  assign y18498 = ~n38880 ;
  assign y18499 = ~n38882 ;
  assign y18500 = ~n38885 ;
  assign y18501 = ~1'b0 ;
  assign y18502 = ~1'b0 ;
  assign y18503 = ~1'b0 ;
  assign y18504 = n38887 ;
  assign y18505 = n38892 ;
  assign y18506 = n38897 ;
  assign y18507 = ~n38899 ;
  assign y18508 = ~n38904 ;
  assign y18509 = n38905 ;
  assign y18510 = n38907 ;
  assign y18511 = ~1'b0 ;
  assign y18512 = ~1'b0 ;
  assign y18513 = ~n38909 ;
  assign y18514 = ~n38912 ;
  assign y18515 = ~n38913 ;
  assign y18516 = ~1'b0 ;
  assign y18517 = ~n38914 ;
  assign y18518 = ~1'b0 ;
  assign y18519 = ~n38920 ;
  assign y18520 = ~1'b0 ;
  assign y18521 = ~n38922 ;
  assign y18522 = ~n38925 ;
  assign y18523 = n38926 ;
  assign y18524 = ~n38927 ;
  assign y18525 = n38928 ;
  assign y18526 = ~1'b0 ;
  assign y18527 = ~n38929 ;
  assign y18528 = n22278 ;
  assign y18529 = ~n38931 ;
  assign y18530 = n38932 ;
  assign y18531 = n38934 ;
  assign y18532 = ~n38937 ;
  assign y18533 = n38941 ;
  assign y18534 = ~n38945 ;
  assign y18535 = ~n38946 ;
  assign y18536 = ~n38948 ;
  assign y18537 = ~n38951 ;
  assign y18538 = n38958 ;
  assign y18539 = ~1'b0 ;
  assign y18540 = n38963 ;
  assign y18541 = ~1'b0 ;
  assign y18542 = ~n38972 ;
  assign y18543 = n38974 ;
  assign y18544 = ~1'b0 ;
  assign y18545 = ~1'b0 ;
  assign y18546 = n38976 ;
  assign y18547 = n38978 ;
  assign y18548 = n38979 ;
  assign y18549 = n38980 ;
  assign y18550 = ~n22267 ;
  assign y18551 = ~n38981 ;
  assign y18552 = n20280 ;
  assign y18553 = ~1'b0 ;
  assign y18554 = ~n38982 ;
  assign y18555 = n38989 ;
  assign y18556 = ~n38991 ;
  assign y18557 = 1'b0 ;
  assign y18558 = n38992 ;
  assign y18559 = ~1'b0 ;
  assign y18560 = ~n19411 ;
  assign y18561 = ~n38993 ;
  assign y18562 = ~n38997 ;
  assign y18563 = ~n38998 ;
  assign y18564 = n38999 ;
  assign y18565 = n39007 ;
  assign y18566 = ~1'b0 ;
  assign y18567 = ~n39009 ;
  assign y18568 = ~n39011 ;
  assign y18569 = n39012 ;
  assign y18570 = ~1'b0 ;
  assign y18571 = ~n39016 ;
  assign y18572 = ~n39021 ;
  assign y18573 = n39022 ;
  assign y18574 = ~n39023 ;
  assign y18575 = n39024 ;
  assign y18576 = ~n39026 ;
  assign y18577 = ~n39028 ;
  assign y18578 = n39031 ;
  assign y18579 = n39032 ;
  assign y18580 = n39034 ;
  assign y18581 = n39036 ;
  assign y18582 = ~n39043 ;
  assign y18583 = ~1'b0 ;
  assign y18584 = n39044 ;
  assign y18585 = n39047 ;
  assign y18586 = ~1'b0 ;
  assign y18587 = n39048 ;
  assign y18588 = n39054 ;
  assign y18589 = n39057 ;
  assign y18590 = ~1'b0 ;
  assign y18591 = ~1'b0 ;
  assign y18592 = ~n39059 ;
  assign y18593 = ~1'b0 ;
  assign y18594 = ~n39061 ;
  assign y18595 = n39062 ;
  assign y18596 = ~1'b0 ;
  assign y18597 = n39063 ;
  assign y18598 = n39069 ;
  assign y18599 = ~1'b0 ;
  assign y18600 = ~1'b0 ;
  assign y18601 = ~n39072 ;
  assign y18602 = ~1'b0 ;
  assign y18603 = 1'b0 ;
  assign y18604 = ~n39074 ;
  assign y18605 = n39076 ;
  assign y18606 = ~n39081 ;
  assign y18607 = n39082 ;
  assign y18608 = ~n39083 ;
  assign y18609 = ~1'b0 ;
  assign y18610 = n39085 ;
  assign y18611 = ~1'b0 ;
  assign y18612 = ~1'b0 ;
  assign y18613 = ~1'b0 ;
  assign y18614 = ~1'b0 ;
  assign y18615 = ~n39088 ;
  assign y18616 = n39092 ;
  assign y18617 = ~n39098 ;
  assign y18618 = n39103 ;
  assign y18619 = ~n39108 ;
  assign y18620 = ~1'b0 ;
  assign y18621 = 1'b0 ;
  assign y18622 = ~n39110 ;
  assign y18623 = n39112 ;
  assign y18624 = n39115 ;
  assign y18625 = n39118 ;
  assign y18626 = ~n39120 ;
  assign y18627 = n39124 ;
  assign y18628 = n39129 ;
  assign y18629 = ~n39133 ;
  assign y18630 = ~n39136 ;
  assign y18631 = ~1'b0 ;
  assign y18632 = ~n39139 ;
  assign y18633 = n39142 ;
  assign y18634 = n39143 ;
  assign y18635 = ~1'b0 ;
  assign y18636 = n39146 ;
  assign y18637 = ~1'b0 ;
  assign y18638 = n39147 ;
  assign y18639 = n39148 ;
  assign y18640 = n39152 ;
  assign y18641 = n39153 ;
  assign y18642 = ~1'b0 ;
  assign y18643 = ~1'b0 ;
  assign y18644 = ~1'b0 ;
  assign y18645 = ~1'b0 ;
  assign y18646 = n39154 ;
  assign y18647 = ~n39156 ;
  assign y18648 = n39157 ;
  assign y18649 = ~n39159 ;
  assign y18650 = ~n12105 ;
  assign y18651 = ~1'b0 ;
  assign y18652 = ~1'b0 ;
  assign y18653 = n39162 ;
  assign y18654 = n39169 ;
  assign y18655 = ~n39173 ;
  assign y18656 = ~n9995 ;
  assign y18657 = ~n39179 ;
  assign y18658 = ~n39187 ;
  assign y18659 = ~1'b0 ;
  assign y18660 = ~1'b0 ;
  assign y18661 = ~n39188 ;
  assign y18662 = n39189 ;
  assign y18663 = ~n29944 ;
  assign y18664 = ~n39193 ;
  assign y18665 = ~1'b0 ;
  assign y18666 = n39197 ;
  assign y18667 = n39198 ;
  assign y18668 = n39199 ;
  assign y18669 = n39210 ;
  assign y18670 = ~n39213 ;
  assign y18671 = ~n39215 ;
  assign y18672 = ~n39218 ;
  assign y18673 = ~n39220 ;
  assign y18674 = ~n39223 ;
  assign y18675 = n39224 ;
  assign y18676 = ~1'b0 ;
  assign y18677 = ~n39229 ;
  assign y18678 = n39232 ;
  assign y18679 = n39235 ;
  assign y18680 = ~1'b0 ;
  assign y18681 = ~n29944 ;
  assign y18682 = ~1'b0 ;
  assign y18683 = ~1'b0 ;
  assign y18684 = 1'b0 ;
  assign y18685 = n39236 ;
  assign y18686 = n39240 ;
  assign y18687 = ~n39245 ;
  assign y18688 = n39257 ;
  assign y18689 = n39264 ;
  assign y18690 = ~n39266 ;
  assign y18691 = ~1'b0 ;
  assign y18692 = ~1'b0 ;
  assign y18693 = n39268 ;
  assign y18694 = ~n39269 ;
  assign y18695 = n39272 ;
  assign y18696 = n39275 ;
  assign y18697 = ~n39276 ;
  assign y18698 = ~n39283 ;
  assign y18699 = ~1'b0 ;
  assign y18700 = n39284 ;
  assign y18701 = n39285 ;
  assign y18702 = ~n39289 ;
  assign y18703 = n39291 ;
  assign y18704 = ~n39293 ;
  assign y18705 = n39295 ;
  assign y18706 = ~n39297 ;
  assign y18707 = ~n13438 ;
  assign y18708 = ~n39301 ;
  assign y18709 = n39305 ;
  assign y18710 = n39311 ;
  assign y18711 = ~n39317 ;
  assign y18712 = ~1'b0 ;
  assign y18713 = ~n39318 ;
  assign y18714 = ~n39319 ;
  assign y18715 = ~1'b0 ;
  assign y18716 = ~n39321 ;
  assign y18717 = ~1'b0 ;
  assign y18718 = ~n9979 ;
  assign y18719 = n39322 ;
  assign y18720 = ~n39326 ;
  assign y18721 = n39328 ;
  assign y18722 = ~n39331 ;
  assign y18723 = ~1'b0 ;
  assign y18724 = ~n39335 ;
  assign y18725 = n13006 ;
  assign y18726 = ~1'b0 ;
  assign y18727 = ~n39339 ;
  assign y18728 = ~n39343 ;
  assign y18729 = 1'b0 ;
  assign y18730 = n39344 ;
  assign y18731 = ~1'b0 ;
  assign y18732 = ~n39345 ;
  assign y18733 = n39349 ;
  assign y18734 = ~n39355 ;
  assign y18735 = n39360 ;
  assign y18736 = ~n39361 ;
  assign y18737 = ~n39362 ;
  assign y18738 = n39364 ;
  assign y18739 = n39366 ;
  assign y18740 = ~1'b0 ;
  assign y18741 = ~1'b0 ;
  assign y18742 = ~1'b0 ;
  assign y18743 = n39369 ;
  assign y18744 = ~1'b0 ;
  assign y18745 = ~n39370 ;
  assign y18746 = ~n39372 ;
  assign y18747 = n39374 ;
  assign y18748 = ~n39376 ;
  assign y18749 = ~1'b0 ;
  assign y18750 = n39379 ;
  assign y18751 = n39381 ;
  assign y18752 = n39385 ;
  assign y18753 = n39386 ;
  assign y18754 = ~n39393 ;
  assign y18755 = ~1'b0 ;
  assign y18756 = ~n39395 ;
  assign y18757 = ~n39398 ;
  assign y18758 = ~n39400 ;
  assign y18759 = 1'b0 ;
  assign y18760 = ~n39402 ;
  assign y18761 = ~n39404 ;
  assign y18762 = n39406 ;
  assign y18763 = n39409 ;
  assign y18764 = ~1'b0 ;
  assign y18765 = n39414 ;
  assign y18766 = n39415 ;
  assign y18767 = ~n39419 ;
  assign y18768 = n39426 ;
  assign y18769 = n38835 ;
  assign y18770 = ~n39427 ;
  assign y18771 = ~n19923 ;
  assign y18772 = ~n39429 ;
  assign y18773 = ~1'b0 ;
  assign y18774 = n39431 ;
  assign y18775 = n39432 ;
  assign y18776 = ~n39434 ;
  assign y18777 = ~n39435 ;
  assign y18778 = ~1'b0 ;
  assign y18779 = ~1'b0 ;
  assign y18780 = ~1'b0 ;
  assign y18781 = ~1'b0 ;
  assign y18782 = ~n39437 ;
  assign y18783 = ~n39440 ;
  assign y18784 = ~1'b0 ;
  assign y18785 = n39442 ;
  assign y18786 = n39444 ;
  assign y18787 = n39451 ;
  assign y18788 = ~n39454 ;
  assign y18789 = ~1'b0 ;
  assign y18790 = ~n39457 ;
  assign y18791 = n39460 ;
  assign y18792 = n39461 ;
  assign y18793 = n39463 ;
  assign y18794 = ~n39468 ;
  assign y18795 = ~n39476 ;
  assign y18796 = ~n39482 ;
  assign y18797 = ~n39487 ;
  assign y18798 = n39491 ;
  assign y18799 = n39493 ;
  assign y18800 = ~1'b0 ;
  assign y18801 = ~n39494 ;
  assign y18802 = n39497 ;
  assign y18803 = n16403 ;
  assign y18804 = ~1'b0 ;
  assign y18805 = n39498 ;
  assign y18806 = ~n39503 ;
  assign y18807 = ~1'b0 ;
  assign y18808 = n39504 ;
  assign y18809 = n20740 ;
  assign y18810 = n39506 ;
  assign y18811 = ~n39512 ;
  assign y18812 = ~1'b0 ;
  assign y18813 = ~n39513 ;
  assign y18814 = n39514 ;
  assign y18815 = ~1'b0 ;
  assign y18816 = n7147 ;
  assign y18817 = ~1'b0 ;
  assign y18818 = ~1'b0 ;
  assign y18819 = ~n39515 ;
  assign y18820 = ~n39517 ;
  assign y18821 = n39518 ;
  assign y18822 = n23264 ;
  assign y18823 = ~n39524 ;
  assign y18824 = ~1'b0 ;
  assign y18825 = ~n39531 ;
  assign y18826 = ~1'b0 ;
  assign y18827 = ~n39533 ;
  assign y18828 = n39535 ;
  assign y18829 = ~1'b0 ;
  assign y18830 = n39536 ;
  assign y18831 = n39540 ;
  assign y18832 = ~n39548 ;
  assign y18833 = n39549 ;
  assign y18834 = ~1'b0 ;
  assign y18835 = ~n39552 ;
  assign y18836 = ~n12058 ;
  assign y18837 = ~1'b0 ;
  assign y18838 = ~n39554 ;
  assign y18839 = 1'b0 ;
  assign y18840 = ~1'b0 ;
  assign y18841 = n34320 ;
  assign y18842 = n39557 ;
  assign y18843 = n39559 ;
  assign y18844 = ~1'b0 ;
  assign y18845 = n39561 ;
  assign y18846 = ~n39563 ;
  assign y18847 = ~1'b0 ;
  assign y18848 = ~n39565 ;
  assign y18849 = n39569 ;
  assign y18850 = ~n39571 ;
  assign y18851 = ~n39574 ;
  assign y18852 = ~1'b0 ;
  assign y18853 = n39575 ;
  assign y18854 = ~n1661 ;
  assign y18855 = ~1'b0 ;
  assign y18856 = ~1'b0 ;
  assign y18857 = n39583 ;
  assign y18858 = ~1'b0 ;
  assign y18859 = ~n39588 ;
  assign y18860 = ~1'b0 ;
  assign y18861 = ~n39591 ;
  assign y18862 = ~n39601 ;
  assign y18863 = ~n39603 ;
  assign y18864 = ~1'b0 ;
  assign y18865 = ~1'b0 ;
  assign y18866 = n39610 ;
  assign y18867 = n39614 ;
  assign y18868 = n39615 ;
  assign y18869 = ~n39619 ;
  assign y18870 = n39624 ;
  assign y18871 = n39625 ;
  assign y18872 = ~1'b0 ;
  assign y18873 = ~1'b0 ;
  assign y18874 = n39626 ;
  assign y18875 = ~n39629 ;
  assign y18876 = n39630 ;
  assign y18877 = ~n39632 ;
  assign y18878 = n39634 ;
  assign y18879 = ~1'b0 ;
  assign y18880 = n39635 ;
  assign y18881 = ~n39637 ;
  assign y18882 = ~1'b0 ;
  assign y18883 = n39639 ;
  assign y18884 = n39649 ;
  assign y18885 = n39651 ;
  assign y18886 = n39652 ;
  assign y18887 = ~n39657 ;
  assign y18888 = ~n39659 ;
  assign y18889 = n39661 ;
  assign y18890 = ~n39665 ;
  assign y18891 = ~n39666 ;
  assign y18892 = ~n39668 ;
  assign y18893 = 1'b0 ;
  assign y18894 = n39672 ;
  assign y18895 = ~n39674 ;
  assign y18896 = n39677 ;
  assign y18897 = ~n39679 ;
  assign y18898 = ~n39683 ;
  assign y18899 = ~n39687 ;
  assign y18900 = n39692 ;
  assign y18901 = n39693 ;
  assign y18902 = n39697 ;
  assign y18903 = 1'b0 ;
  assign y18904 = ~n39699 ;
  assign y18905 = ~n39700 ;
  assign y18906 = ~1'b0 ;
  assign y18907 = ~n39704 ;
  assign y18908 = ~n39707 ;
  assign y18909 = ~1'b0 ;
  assign y18910 = ~n39708 ;
  assign y18911 = n39716 ;
  assign y18912 = n39717 ;
  assign y18913 = ~n39721 ;
  assign y18914 = n39726 ;
  assign y18915 = ~n39728 ;
  assign y18916 = n39732 ;
  assign y18917 = n39737 ;
  assign y18918 = ~1'b0 ;
  assign y18919 = n39739 ;
  assign y18920 = ~n39742 ;
  assign y18921 = ~n39745 ;
  assign y18922 = ~n39746 ;
  assign y18923 = n39748 ;
  assign y18924 = ~n39750 ;
  assign y18925 = n39754 ;
  assign y18926 = ~1'b0 ;
  assign y18927 = ~n39756 ;
  assign y18928 = 1'b0 ;
  assign y18929 = n39762 ;
  assign y18930 = ~n39763 ;
  assign y18931 = n39765 ;
  assign y18932 = ~n39775 ;
  assign y18933 = ~n39776 ;
  assign y18934 = ~1'b0 ;
  assign y18935 = ~1'b0 ;
  assign y18936 = n39778 ;
  assign y18937 = n36657 ;
  assign y18938 = ~1'b0 ;
  assign y18939 = n39779 ;
  assign y18940 = ~1'b0 ;
  assign y18941 = ~1'b0 ;
  assign y18942 = n39780 ;
  assign y18943 = n39783 ;
  assign y18944 = ~n39784 ;
  assign y18945 = ~1'b0 ;
  assign y18946 = n39785 ;
  assign y18947 = ~n39786 ;
  assign y18948 = ~1'b0 ;
  assign y18949 = n39788 ;
  assign y18950 = ~n39789 ;
  assign y18951 = ~n39790 ;
  assign y18952 = n39791 ;
  assign y18953 = ~1'b0 ;
  assign y18954 = ~1'b0 ;
  assign y18955 = n39793 ;
  assign y18956 = ~n39795 ;
  assign y18957 = ~n39800 ;
  assign y18958 = ~1'b0 ;
  assign y18959 = n23 ;
  assign y18960 = ~n39802 ;
  assign y18961 = n39803 ;
  assign y18962 = ~n22052 ;
  assign y18963 = ~n39804 ;
  assign y18964 = n39806 ;
  assign y18965 = ~n3581 ;
  assign y18966 = n39811 ;
  assign y18967 = 1'b0 ;
  assign y18968 = n39813 ;
  assign y18969 = n39815 ;
  assign y18970 = 1'b0 ;
  assign y18971 = ~n39816 ;
  assign y18972 = n39817 ;
  assign y18973 = ~1'b0 ;
  assign y18974 = ~n39819 ;
  assign y18975 = ~1'b0 ;
  assign y18976 = ~n39827 ;
  assign y18977 = ~n39828 ;
  assign y18978 = n39830 ;
  assign y18979 = ~1'b0 ;
  assign y18980 = ~n21751 ;
  assign y18981 = ~1'b0 ;
  assign y18982 = n39835 ;
  assign y18983 = ~1'b0 ;
  assign y18984 = ~1'b0 ;
  assign y18985 = n39837 ;
  assign y18986 = ~1'b0 ;
  assign y18987 = n39840 ;
  assign y18988 = ~1'b0 ;
  assign y18989 = ~n39847 ;
  assign y18990 = ~n39849 ;
  assign y18991 = n39850 ;
  assign y18992 = ~1'b0 ;
  assign y18993 = ~n39854 ;
  assign y18994 = ~1'b0 ;
  assign y18995 = ~n39855 ;
  assign y18996 = ~n691 ;
  assign y18997 = ~n39859 ;
  assign y18998 = ~n39861 ;
  assign y18999 = n39863 ;
  assign y19000 = n39866 ;
  assign y19001 = ~1'b0 ;
  assign y19002 = n39867 ;
  assign y19003 = ~n39868 ;
  assign y19004 = ~n39871 ;
  assign y19005 = ~1'b0 ;
  assign y19006 = ~1'b0 ;
  assign y19007 = ~n39872 ;
  assign y19008 = 1'b0 ;
  assign y19009 = ~n39875 ;
  assign y19010 = n39877 ;
  assign y19011 = n39880 ;
  assign y19012 = ~1'b0 ;
  assign y19013 = n39885 ;
  assign y19014 = ~n13509 ;
  assign y19015 = n39886 ;
  assign y19016 = ~1'b0 ;
  assign y19017 = n39888 ;
  assign y19018 = n39890 ;
  assign y19019 = ~n39891 ;
  assign y19020 = ~n39893 ;
  assign y19021 = ~n39901 ;
  assign y19022 = ~n39903 ;
  assign y19023 = n39904 ;
  assign y19024 = n39182 ;
  assign y19025 = 1'b0 ;
  assign y19026 = ~n39906 ;
  assign y19027 = n39907 ;
  assign y19028 = ~n39909 ;
  assign y19029 = ~n39914 ;
  assign y19030 = n39916 ;
  assign y19031 = ~1'b0 ;
  assign y19032 = ~1'b0 ;
  assign y19033 = ~1'b0 ;
  assign y19034 = ~n39918 ;
  assign y19035 = n39919 ;
  assign y19036 = n39921 ;
  assign y19037 = ~n39923 ;
  assign y19038 = ~n39924 ;
  assign y19039 = ~1'b0 ;
  assign y19040 = n39926 ;
  assign y19041 = ~1'b0 ;
  assign y19042 = n39928 ;
  assign y19043 = ~n39930 ;
  assign y19044 = ~1'b0 ;
  assign y19045 = n39932 ;
  assign y19046 = ~n39934 ;
  assign y19047 = ~n25543 ;
  assign y19048 = ~1'b0 ;
  assign y19049 = n39943 ;
  assign y19050 = 1'b0 ;
  assign y19051 = ~n39944 ;
  assign y19052 = n39945 ;
  assign y19053 = ~n39947 ;
  assign y19054 = ~n39954 ;
  assign y19055 = n1235 ;
  assign y19056 = ~1'b0 ;
  assign y19057 = ~n39955 ;
  assign y19058 = n39958 ;
  assign y19059 = ~n39960 ;
  assign y19060 = n39963 ;
  assign y19061 = ~n16192 ;
  assign y19062 = ~n4226 ;
  assign y19063 = ~1'b0 ;
  assign y19064 = ~1'b0 ;
  assign y19065 = ~n3656 ;
  assign y19066 = ~n3694 ;
  assign y19067 = ~n39964 ;
  assign y19068 = ~1'b0 ;
  assign y19069 = n39965 ;
  assign y19070 = ~1'b0 ;
  assign y19071 = n39967 ;
  assign y19072 = n39971 ;
  assign y19073 = n2628 ;
  assign y19074 = ~n39974 ;
  assign y19075 = ~1'b0 ;
  assign y19076 = ~n6229 ;
  assign y19077 = n34643 ;
  assign y19078 = n3606 ;
  assign y19079 = ~1'b0 ;
  assign y19080 = n39978 ;
  assign y19081 = n39981 ;
  assign y19082 = ~n39982 ;
  assign y19083 = n39983 ;
  assign y19084 = n39985 ;
  assign y19085 = n39992 ;
  assign y19086 = ~1'b0 ;
  assign y19087 = ~n39996 ;
  assign y19088 = ~n40000 ;
  assign y19089 = n40001 ;
  assign y19090 = n40002 ;
  assign y19091 = n1442 ;
  assign y19092 = n40005 ;
  assign y19093 = ~1'b0 ;
  assign y19094 = ~n40011 ;
  assign y19095 = ~n40015 ;
  assign y19096 = ~n40019 ;
  assign y19097 = n40024 ;
  assign y19098 = n40032 ;
  assign y19099 = 1'b0 ;
  assign y19100 = ~n40035 ;
  assign y19101 = ~1'b0 ;
  assign y19102 = ~n40038 ;
  assign y19103 = ~n40043 ;
  assign y19104 = n40045 ;
  assign y19105 = ~1'b0 ;
  assign y19106 = ~n40049 ;
  assign y19107 = 1'b0 ;
  assign y19108 = ~n40051 ;
  assign y19109 = ~1'b0 ;
  assign y19110 = n40052 ;
  assign y19111 = ~n40053 ;
  assign y19112 = ~n3192 ;
  assign y19113 = ~n40056 ;
  assign y19114 = ~n40058 ;
  assign y19115 = n40060 ;
  assign y19116 = ~n40061 ;
  assign y19117 = ~1'b0 ;
  assign y19118 = n40062 ;
  assign y19119 = n40070 ;
  assign y19120 = n40071 ;
  assign y19121 = ~n40072 ;
  assign y19122 = ~n40075 ;
  assign y19123 = ~1'b0 ;
  assign y19124 = n32692 ;
  assign y19125 = n40078 ;
  assign y19126 = ~1'b0 ;
  assign y19127 = ~1'b0 ;
  assign y19128 = n40079 ;
  assign y19129 = ~n40080 ;
  assign y19130 = ~n40082 ;
  assign y19131 = ~n8684 ;
  assign y19132 = ~n40084 ;
  assign y19133 = ~n40086 ;
  assign y19134 = n40087 ;
  assign y19135 = ~n40089 ;
  assign y19136 = ~1'b0 ;
  assign y19137 = ~1'b0 ;
  assign y19138 = ~1'b0 ;
  assign y19139 = ~1'b0 ;
  assign y19140 = n40092 ;
  assign y19141 = ~n40107 ;
  assign y19142 = n40109 ;
  assign y19143 = ~n40110 ;
  assign y19144 = ~n40114 ;
  assign y19145 = n40117 ;
  assign y19146 = ~n40123 ;
  assign y19147 = n40124 ;
  assign y19148 = ~n40126 ;
  assign y19149 = ~n40127 ;
  assign y19150 = ~n40132 ;
  assign y19151 = ~n40133 ;
  assign y19152 = ~n40134 ;
  assign y19153 = ~1'b0 ;
  assign y19154 = ~n40136 ;
  assign y19155 = n40139 ;
  assign y19156 = n6047 ;
  assign y19157 = n40140 ;
  assign y19158 = ~1'b0 ;
  assign y19159 = n40145 ;
  assign y19160 = ~n40151 ;
  assign y19161 = ~n40158 ;
  assign y19162 = ~1'b0 ;
  assign y19163 = n40161 ;
  assign y19164 = ~n17765 ;
  assign y19165 = ~n40164 ;
  assign y19166 = ~1'b0 ;
  assign y19167 = n40167 ;
  assign y19168 = ~n40168 ;
  assign y19169 = ~n40170 ;
  assign y19170 = n40173 ;
  assign y19171 = ~n40175 ;
  assign y19172 = ~n40177 ;
  assign y19173 = ~n20505 ;
  assign y19174 = ~n40179 ;
  assign y19175 = n40181 ;
  assign y19176 = ~1'b0 ;
  assign y19177 = ~1'b0 ;
  assign y19178 = ~n40184 ;
  assign y19179 = ~n40187 ;
  assign y19180 = ~n40188 ;
  assign y19181 = n40189 ;
  assign y19182 = ~1'b0 ;
  assign y19183 = ~1'b0 ;
  assign y19184 = 1'b0 ;
  assign y19185 = n40194 ;
  assign y19186 = n40196 ;
  assign y19187 = n40198 ;
  assign y19188 = n40199 ;
  assign y19189 = n40202 ;
  assign y19190 = ~1'b0 ;
  assign y19191 = ~n40204 ;
  assign y19192 = ~1'b0 ;
  assign y19193 = n40206 ;
  assign y19194 = ~1'b0 ;
  assign y19195 = n40207 ;
  assign y19196 = ~1'b0 ;
  assign y19197 = ~1'b0 ;
  assign y19198 = ~n40214 ;
  assign y19199 = n40221 ;
  assign y19200 = 1'b0 ;
  assign y19201 = ~n40223 ;
  assign y19202 = n40224 ;
  assign y19203 = n40232 ;
  assign y19204 = n40234 ;
  assign y19205 = ~n40235 ;
  assign y19206 = ~1'b0 ;
  assign y19207 = ~1'b0 ;
  assign y19208 = ~n40236 ;
  assign y19209 = ~n40240 ;
  assign y19210 = ~n40241 ;
  assign y19211 = ~n8829 ;
  assign y19212 = n40245 ;
  assign y19213 = n40246 ;
  assign y19214 = ~1'b0 ;
  assign y19215 = n40249 ;
  assign y19216 = n40252 ;
  assign y19217 = n40254 ;
  assign y19218 = ~1'b0 ;
  assign y19219 = n40256 ;
  assign y19220 = ~n40257 ;
  assign y19221 = n40260 ;
  assign y19222 = ~1'b0 ;
  assign y19223 = n40269 ;
  assign y19224 = ~1'b0 ;
  assign y19225 = ~n17102 ;
  assign y19226 = ~1'b0 ;
  assign y19227 = ~n40272 ;
  assign y19228 = ~n40273 ;
  assign y19229 = ~n39970 ;
  assign y19230 = n40277 ;
  assign y19231 = n40278 ;
  assign y19232 = ~1'b0 ;
  assign y19233 = n40302 ;
  assign y19234 = ~n40305 ;
  assign y19235 = ~n40310 ;
  assign y19236 = n40311 ;
  assign y19237 = n40316 ;
  assign y19238 = ~1'b0 ;
  assign y19239 = n40318 ;
  assign y19240 = ~1'b0 ;
  assign y19241 = n22900 ;
  assign y19242 = ~n40319 ;
  assign y19243 = n40323 ;
  assign y19244 = ~1'b0 ;
  assign y19245 = ~n40324 ;
  assign y19246 = ~1'b0 ;
  assign y19247 = ~1'b0 ;
  assign y19248 = ~n40327 ;
  assign y19249 = n40331 ;
  assign y19250 = n40334 ;
  assign y19251 = ~n40340 ;
  assign y19252 = ~n40342 ;
  assign y19253 = ~1'b0 ;
  assign y19254 = n40343 ;
  assign y19255 = n40346 ;
  assign y19256 = ~n40348 ;
  assign y19257 = ~1'b0 ;
  assign y19258 = ~n19371 ;
  assign y19259 = n40355 ;
  assign y19260 = ~1'b0 ;
  assign y19261 = n40358 ;
  assign y19262 = ~n40360 ;
  assign y19263 = n40362 ;
  assign y19264 = ~n40365 ;
  assign y19265 = ~1'b0 ;
  assign y19266 = ~n40370 ;
  assign y19267 = n40373 ;
  assign y19268 = n40377 ;
  assign y19269 = ~1'b0 ;
  assign y19270 = ~n40381 ;
  assign y19271 = ~1'b0 ;
  assign y19272 = ~n40382 ;
  assign y19273 = ~n14671 ;
  assign y19274 = n40383 ;
  assign y19275 = ~n40384 ;
  assign y19276 = ~n40385 ;
  assign y19277 = n4204 ;
  assign y19278 = ~1'b0 ;
  assign y19279 = n40387 ;
  assign y19280 = n20679 ;
  assign y19281 = ~1'b0 ;
  assign y19282 = ~1'b0 ;
  assign y19283 = ~1'b0 ;
  assign y19284 = ~n40389 ;
  assign y19285 = ~n40392 ;
  assign y19286 = n32276 ;
  assign y19287 = ~n40395 ;
  assign y19288 = ~1'b0 ;
  assign y19289 = n16082 ;
  assign y19290 = ~1'b0 ;
  assign y19291 = n40396 ;
  assign y19292 = ~1'b0 ;
  assign y19293 = n40398 ;
  assign y19294 = ~n40401 ;
  assign y19295 = ~1'b0 ;
  assign y19296 = ~1'b0 ;
  assign y19297 = ~n40402 ;
  assign y19298 = ~n40404 ;
  assign y19299 = ~n40405 ;
  assign y19300 = n40406 ;
  assign y19301 = ~n21571 ;
  assign y19302 = ~n40408 ;
  assign y19303 = ~1'b0 ;
  assign y19304 = ~n40413 ;
  assign y19305 = n40414 ;
  assign y19306 = ~n10221 ;
  assign y19307 = n40418 ;
  assign y19308 = ~1'b0 ;
  assign y19309 = n40419 ;
  assign y19310 = n40420 ;
  assign y19311 = ~1'b0 ;
  assign y19312 = ~1'b0 ;
  assign y19313 = n40421 ;
  assign y19314 = ~1'b0 ;
  assign y19315 = n2620 ;
  assign y19316 = n40422 ;
  assign y19317 = ~n40424 ;
  assign y19318 = ~1'b0 ;
  assign y19319 = ~n40425 ;
  assign y19320 = ~n40426 ;
  assign y19321 = ~n40429 ;
  assign y19322 = ~n40431 ;
  assign y19323 = n40432 ;
  assign y19324 = ~1'b0 ;
  assign y19325 = n40434 ;
  assign y19326 = ~1'b0 ;
  assign y19327 = ~n40441 ;
  assign y19328 = n40442 ;
  assign y19329 = n40444 ;
  assign y19330 = ~1'b0 ;
  assign y19331 = n40447 ;
  assign y19332 = ~n40449 ;
  assign y19333 = n40450 ;
  assign y19334 = ~1'b0 ;
  assign y19335 = ~n40453 ;
  assign y19336 = n40457 ;
  assign y19337 = ~n40460 ;
  assign y19338 = n17042 ;
  assign y19339 = ~n40464 ;
  assign y19340 = ~n40469 ;
  assign y19341 = ~n40473 ;
  assign y19342 = n40478 ;
  assign y19343 = n40480 ;
  assign y19344 = n40483 ;
  assign y19345 = ~1'b0 ;
  assign y19346 = ~1'b0 ;
  assign y19347 = ~1'b0 ;
  assign y19348 = ~1'b0 ;
  assign y19349 = n40485 ;
  assign y19350 = ~n40487 ;
  assign y19351 = n40488 ;
  assign y19352 = ~n40491 ;
  assign y19353 = ~n40493 ;
  assign y19354 = ~1'b0 ;
  assign y19355 = n40495 ;
  assign y19356 = ~n39112 ;
  assign y19357 = n40498 ;
  assign y19358 = n40499 ;
  assign y19359 = n15730 ;
  assign y19360 = ~1'b0 ;
  assign y19361 = ~1'b0 ;
  assign y19362 = n40501 ;
  assign y19363 = ~n40502 ;
  assign y19364 = ~n40503 ;
  assign y19365 = n40508 ;
  assign y19366 = ~1'b0 ;
  assign y19367 = ~1'b0 ;
  assign y19368 = n40510 ;
  assign y19369 = ~n40511 ;
  assign y19370 = ~n3607 ;
  assign y19371 = ~n40512 ;
  assign y19372 = ~1'b0 ;
  assign y19373 = n40514 ;
  assign y19374 = n40515 ;
  assign y19375 = ~n1768 ;
  assign y19376 = ~n40520 ;
  assign y19377 = ~n40521 ;
  assign y19378 = ~n40527 ;
  assign y19379 = ~1'b0 ;
  assign y19380 = ~n16488 ;
  assign y19381 = ~n7516 ;
  assign y19382 = n40529 ;
  assign y19383 = ~n40531 ;
  assign y19384 = ~n40533 ;
  assign y19385 = ~n40536 ;
  assign y19386 = ~n40538 ;
  assign y19387 = ~n40539 ;
  assign y19388 = 1'b0 ;
  assign y19389 = ~1'b0 ;
  assign y19390 = n40542 ;
  assign y19391 = ~n40543 ;
  assign y19392 = n40545 ;
  assign y19393 = ~n40546 ;
  assign y19394 = n40547 ;
  assign y19395 = n40549 ;
  assign y19396 = ~n40550 ;
  assign y19397 = n40552 ;
  assign y19398 = n40554 ;
  assign y19399 = ~n40558 ;
  assign y19400 = ~1'b0 ;
  assign y19401 = ~n40563 ;
  assign y19402 = ~n1846 ;
  assign y19403 = ~n40565 ;
  assign y19404 = ~n40567 ;
  assign y19405 = 1'b0 ;
  assign y19406 = ~n40569 ;
  assign y19407 = n40574 ;
  assign y19408 = ~1'b0 ;
  assign y19409 = n40577 ;
  assign y19410 = ~n40584 ;
  assign y19411 = ~n40585 ;
  assign y19412 = 1'b0 ;
  assign y19413 = ~n40588 ;
  assign y19414 = ~n40589 ;
  assign y19415 = ~1'b0 ;
  assign y19416 = n40591 ;
  assign y19417 = ~1'b0 ;
  assign y19418 = n40592 ;
  assign y19419 = n40595 ;
  assign y19420 = ~n40596 ;
  assign y19421 = n35057 ;
  assign y19422 = ~n40603 ;
  assign y19423 = ~1'b0 ;
  assign y19424 = ~n40606 ;
  assign y19425 = ~1'b0 ;
  assign y19426 = ~1'b0 ;
  assign y19427 = ~1'b0 ;
  assign y19428 = n3196 ;
  assign y19429 = ~n32808 ;
  assign y19430 = n40611 ;
  assign y19431 = n40612 ;
  assign y19432 = ~n40613 ;
  assign y19433 = 1'b0 ;
  assign y19434 = ~n1308 ;
  assign y19435 = ~1'b0 ;
  assign y19436 = n40617 ;
  assign y19437 = ~n40620 ;
  assign y19438 = ~1'b0 ;
  assign y19439 = n40626 ;
  assign y19440 = n40630 ;
  assign y19441 = ~n40633 ;
  assign y19442 = ~1'b0 ;
  assign y19443 = ~1'b0 ;
  assign y19444 = ~1'b0 ;
  assign y19445 = ~n40634 ;
  assign y19446 = n40635 ;
  assign y19447 = ~n19450 ;
  assign y19448 = n40637 ;
  assign y19449 = ~n40638 ;
  assign y19450 = ~n40044 ;
  assign y19451 = ~n40640 ;
  assign y19452 = ~n40642 ;
  assign y19453 = n40643 ;
  assign y19454 = n40645 ;
  assign y19455 = ~1'b0 ;
  assign y19456 = n40647 ;
  assign y19457 = ~1'b0 ;
  assign y19458 = ~n40648 ;
  assign y19459 = ~n40655 ;
  assign y19460 = n40657 ;
  assign y19461 = n40659 ;
  assign y19462 = ~n40660 ;
  assign y19463 = ~1'b0 ;
  assign y19464 = n40663 ;
  assign y19465 = ~1'b0 ;
  assign y19466 = ~n4639 ;
  assign y19467 = n29643 ;
  assign y19468 = ~n40666 ;
  assign y19469 = ~1'b0 ;
  assign y19470 = ~n40668 ;
  assign y19471 = ~n40677 ;
  assign y19472 = ~1'b0 ;
  assign y19473 = n40681 ;
  assign y19474 = ~n40682 ;
  assign y19475 = ~1'b0 ;
  assign y19476 = ~1'b0 ;
  assign y19477 = ~1'b0 ;
  assign y19478 = n40687 ;
  assign y19479 = n40688 ;
  assign y19480 = ~n40692 ;
  assign y19481 = ~n40693 ;
  assign y19482 = ~1'b0 ;
  assign y19483 = n40699 ;
  assign y19484 = n40700 ;
  assign y19485 = n40701 ;
  assign y19486 = ~1'b0 ;
  assign y19487 = n40704 ;
  assign y19488 = ~n40705 ;
  assign y19489 = ~n40706 ;
  assign y19490 = ~n40707 ;
  assign y19491 = n40709 ;
  assign y19492 = n40715 ;
  assign y19493 = n40718 ;
  assign y19494 = ~n40719 ;
  assign y19495 = ~n40722 ;
  assign y19496 = ~1'b0 ;
  assign y19497 = ~n40726 ;
  assign y19498 = ~1'b0 ;
  assign y19499 = n40730 ;
  assign y19500 = ~n40732 ;
  assign y19501 = ~n40733 ;
  assign y19502 = n40734 ;
  assign y19503 = 1'b0 ;
  assign y19504 = n40737 ;
  assign y19505 = n40740 ;
  assign y19506 = n40746 ;
  assign y19507 = n40750 ;
  assign y19508 = ~1'b0 ;
  assign y19509 = ~n40754 ;
  assign y19510 = n40760 ;
  assign y19511 = ~1'b0 ;
  assign y19512 = ~1'b0 ;
  assign y19513 = ~1'b0 ;
  assign y19514 = ~1'b0 ;
  assign y19515 = ~1'b0 ;
  assign y19516 = n40761 ;
  assign y19517 = ~1'b0 ;
  assign y19518 = ~n40767 ;
  assign y19519 = ~n40769 ;
  assign y19520 = ~n24462 ;
  assign y19521 = ~n16291 ;
  assign y19522 = n40772 ;
  assign y19523 = ~n40773 ;
  assign y19524 = ~1'b0 ;
  assign y19525 = ~1'b0 ;
  assign y19526 = ~n40779 ;
  assign y19527 = ~n40783 ;
  assign y19528 = ~1'b0 ;
  assign y19529 = n40785 ;
  assign y19530 = ~n40789 ;
  assign y19531 = n8355 ;
  assign y19532 = ~1'b0 ;
  assign y19533 = ~1'b0 ;
  assign y19534 = ~n40791 ;
  assign y19535 = ~1'b0 ;
  assign y19536 = ~1'b0 ;
  assign y19537 = n40793 ;
  assign y19538 = n40796 ;
  assign y19539 = ~n14671 ;
  assign y19540 = n40797 ;
  assign y19541 = n40798 ;
  assign y19542 = n40799 ;
  assign y19543 = ~n40802 ;
  assign y19544 = n40803 ;
  assign y19545 = ~1'b0 ;
  assign y19546 = ~n40813 ;
  assign y19547 = n19623 ;
  assign y19548 = n40814 ;
  assign y19549 = n40817 ;
  assign y19550 = n40818 ;
  assign y19551 = 1'b0 ;
  assign y19552 = ~1'b0 ;
  assign y19553 = ~n40821 ;
  assign y19554 = ~n40825 ;
  assign y19555 = ~n40827 ;
  assign y19556 = 1'b0 ;
  assign y19557 = ~n40830 ;
  assign y19558 = ~n40833 ;
  assign y19559 = ~1'b0 ;
  assign y19560 = ~1'b0 ;
  assign y19561 = ~n40835 ;
  assign y19562 = n40836 ;
  assign y19563 = ~n40838 ;
  assign y19564 = n40840 ;
  assign y19565 = n40841 ;
  assign y19566 = n40844 ;
  assign y19567 = n40845 ;
  assign y19568 = n40847 ;
  assign y19569 = ~n40848 ;
  assign y19570 = ~n40850 ;
  assign y19571 = n960 ;
  assign y19572 = n40852 ;
  assign y19573 = n40856 ;
  assign y19574 = ~1'b0 ;
  assign y19575 = ~n40858 ;
  assign y19576 = n40860 ;
  assign y19577 = n40861 ;
  assign y19578 = ~n26928 ;
  assign y19579 = ~n40864 ;
  assign y19580 = ~1'b0 ;
  assign y19581 = ~n40870 ;
  assign y19582 = ~1'b0 ;
  assign y19583 = ~n40871 ;
  assign y19584 = ~n40878 ;
  assign y19585 = ~1'b0 ;
  assign y19586 = ~n40880 ;
  assign y19587 = ~n40884 ;
  assign y19588 = ~n40885 ;
  assign y19589 = n40887 ;
  assign y19590 = ~1'b0 ;
  assign y19591 = ~n40888 ;
  assign y19592 = ~n40889 ;
  assign y19593 = ~n40895 ;
  assign y19594 = ~n40896 ;
  assign y19595 = ~n40897 ;
  assign y19596 = ~1'b0 ;
  assign y19597 = ~1'b0 ;
  assign y19598 = ~1'b0 ;
  assign y19599 = ~n22103 ;
  assign y19600 = n40898 ;
  assign y19601 = ~n40900 ;
  assign y19602 = 1'b0 ;
  assign y19603 = 1'b0 ;
  assign y19604 = n20487 ;
  assign y19605 = n40905 ;
  assign y19606 = ~1'b0 ;
  assign y19607 = n40907 ;
  assign y19608 = n40915 ;
  assign y19609 = ~1'b0 ;
  assign y19610 = ~1'b0 ;
  assign y19611 = ~n40916 ;
  assign y19612 = ~1'b0 ;
  assign y19613 = ~1'b0 ;
  assign y19614 = ~n40918 ;
  assign y19615 = ~n40920 ;
  assign y19616 = ~n40923 ;
  assign y19617 = n40926 ;
  assign y19618 = ~n40927 ;
  assign y19619 = ~1'b0 ;
  assign y19620 = ~n40931 ;
  assign y19621 = ~n40937 ;
  assign y19622 = n40939 ;
  assign y19623 = ~n40942 ;
  assign y19624 = ~n40945 ;
  assign y19625 = n5501 ;
  assign y19626 = ~1'b0 ;
  assign y19627 = ~n40950 ;
  assign y19628 = ~1'b0 ;
  assign y19629 = ~n40952 ;
  assign y19630 = ~n40956 ;
  assign y19631 = n40959 ;
  assign y19632 = ~1'b0 ;
  assign y19633 = n40961 ;
  assign y19634 = ~n40963 ;
  assign y19635 = ~n40964 ;
  assign y19636 = ~1'b0 ;
  assign y19637 = n40968 ;
  assign y19638 = ~n40970 ;
  assign y19639 = n40971 ;
  assign y19640 = ~n40972 ;
  assign y19641 = n40974 ;
  assign y19642 = ~1'b0 ;
  assign y19643 = ~1'b0 ;
  assign y19644 = n40975 ;
  assign y19645 = ~n40976 ;
  assign y19646 = n40979 ;
  assign y19647 = 1'b0 ;
  assign y19648 = ~n40980 ;
  assign y19649 = n40981 ;
  assign y19650 = ~1'b0 ;
  assign y19651 = ~1'b0 ;
  assign y19652 = n40983 ;
  assign y19653 = ~n40985 ;
  assign y19654 = n40986 ;
  assign y19655 = ~1'b0 ;
  assign y19656 = n19714 ;
  assign y19657 = n40992 ;
  assign y19658 = n40995 ;
  assign y19659 = ~1'b0 ;
  assign y19660 = 1'b0 ;
  assign y19661 = ~1'b0 ;
  assign y19662 = n40999 ;
  assign y19663 = n41001 ;
  assign y19664 = ~1'b0 ;
  assign y19665 = n9286 ;
  assign y19666 = ~n41006 ;
  assign y19667 = n41008 ;
  assign y19668 = n41009 ;
  assign y19669 = ~n41011 ;
  assign y19670 = n5128 ;
  assign y19671 = ~1'b0 ;
  assign y19672 = n41012 ;
  assign y19673 = ~n41014 ;
  assign y19674 = n41015 ;
  assign y19675 = ~n41018 ;
  assign y19676 = ~n13730 ;
  assign y19677 = ~n41024 ;
  assign y19678 = ~1'b0 ;
  assign y19679 = ~n41026 ;
  assign y19680 = n41027 ;
  assign y19681 = n41028 ;
  assign y19682 = ~n41031 ;
  assign y19683 = n41034 ;
  assign y19684 = n62 ;
  assign y19685 = n41035 ;
  assign y19686 = n41036 ;
  assign y19687 = ~1'b0 ;
  assign y19688 = ~1'b0 ;
  assign y19689 = ~1'b0 ;
  assign y19690 = ~n41038 ;
  assign y19691 = ~n41040 ;
  assign y19692 = ~n41045 ;
  assign y19693 = ~1'b0 ;
  assign y19694 = n41050 ;
  assign y19695 = ~n41053 ;
  assign y19696 = n41054 ;
  assign y19697 = ~n41057 ;
  assign y19698 = ~1'b0 ;
  assign y19699 = ~n41061 ;
  assign y19700 = ~1'b0 ;
  assign y19701 = n41064 ;
  assign y19702 = ~n41066 ;
  assign y19703 = ~n41069 ;
  assign y19704 = n41073 ;
  assign y19705 = n41075 ;
  assign y19706 = ~n41076 ;
  assign y19707 = ~1'b0 ;
  assign y19708 = ~1'b0 ;
  assign y19709 = ~n41078 ;
  assign y19710 = ~n41081 ;
  assign y19711 = ~n41086 ;
  assign y19712 = ~1'b0 ;
  assign y19713 = n41091 ;
  assign y19714 = ~n41092 ;
  assign y19715 = ~1'b0 ;
  assign y19716 = ~1'b0 ;
  assign y19717 = ~1'b0 ;
  assign y19718 = n41094 ;
  assign y19719 = n41095 ;
  assign y19720 = n41102 ;
  assign y19721 = ~n41103 ;
  assign y19722 = n41104 ;
  assign y19723 = ~1'b0 ;
  assign y19724 = ~n41108 ;
  assign y19725 = ~1'b0 ;
  assign y19726 = n41109 ;
  assign y19727 = ~n1359 ;
  assign y19728 = n41112 ;
  assign y19729 = ~n41117 ;
  assign y19730 = ~1'b0 ;
  assign y19731 = n41119 ;
  assign y19732 = ~n41121 ;
  assign y19733 = ~n41123 ;
  assign y19734 = n41124 ;
  assign y19735 = ~1'b0 ;
  assign y19736 = n41125 ;
  assign y19737 = ~n41129 ;
  assign y19738 = n41131 ;
  assign y19739 = ~n41132 ;
  assign y19740 = ~n41136 ;
  assign y19741 = ~n41138 ;
  assign y19742 = ~n41140 ;
  assign y19743 = n41144 ;
  assign y19744 = ~n24212 ;
  assign y19745 = ~1'b0 ;
  assign y19746 = n41146 ;
  assign y19747 = ~1'b0 ;
  assign y19748 = ~n41148 ;
  assign y19749 = ~n41152 ;
  assign y19750 = n41154 ;
  assign y19751 = n41159 ;
  assign y19752 = ~n41160 ;
  assign y19753 = ~1'b0 ;
  assign y19754 = ~n5831 ;
  assign y19755 = ~n41162 ;
  assign y19756 = ~1'b0 ;
  assign y19757 = ~n41164 ;
  assign y19758 = n41165 ;
  assign y19759 = ~1'b0 ;
  assign y19760 = n41166 ;
  assign y19761 = n18950 ;
  assign y19762 = n41167 ;
  assign y19763 = n41170 ;
  assign y19764 = n41173 ;
  assign y19765 = ~1'b0 ;
  assign y19766 = ~n2776 ;
  assign y19767 = ~1'b0 ;
  assign y19768 = n41176 ;
  assign y19769 = n41180 ;
  assign y19770 = ~n41184 ;
  assign y19771 = ~1'b0 ;
  assign y19772 = ~1'b0 ;
  assign y19773 = ~n41185 ;
  assign y19774 = ~n41188 ;
  assign y19775 = n41190 ;
  assign y19776 = ~n41191 ;
  assign y19777 = ~n41192 ;
  assign y19778 = n41193 ;
  assign y19779 = ~1'b0 ;
  assign y19780 = n41198 ;
  assign y19781 = ~n41200 ;
  assign y19782 = ~n41201 ;
  assign y19783 = ~n41202 ;
  assign y19784 = n41208 ;
  assign y19785 = ~n41212 ;
  assign y19786 = n41215 ;
  assign y19787 = ~n41217 ;
  assign y19788 = n41219 ;
  assign y19789 = ~1'b0 ;
  assign y19790 = ~1'b0 ;
  assign y19791 = ~1'b0 ;
  assign y19792 = ~n41220 ;
  assign y19793 = ~1'b0 ;
  assign y19794 = ~1'b0 ;
  assign y19795 = n41221 ;
  assign y19796 = n41222 ;
  assign y19797 = ~n41224 ;
  assign y19798 = ~1'b0 ;
  assign y19799 = n41227 ;
  assign y19800 = ~n304 ;
  assign y19801 = n41228 ;
  assign y19802 = n41232 ;
  assign y19803 = n41236 ;
  assign y19804 = ~n41237 ;
  assign y19805 = n41243 ;
  assign y19806 = n41244 ;
  assign y19807 = ~n41245 ;
  assign y19808 = n41247 ;
  assign y19809 = ~n41251 ;
  assign y19810 = n41257 ;
  assign y19811 = ~1'b0 ;
  assign y19812 = ~n41260 ;
  assign y19813 = n41264 ;
  assign y19814 = n41266 ;
  assign y19815 = ~1'b0 ;
  assign y19816 = n22888 ;
  assign y19817 = ~n41267 ;
  assign y19818 = n41274 ;
  assign y19819 = ~n41275 ;
  assign y19820 = ~1'b0 ;
  assign y19821 = ~n41277 ;
  assign y19822 = ~1'b0 ;
  assign y19823 = ~1'b0 ;
  assign y19824 = ~n41279 ;
  assign y19825 = ~n41280 ;
  assign y19826 = n41282 ;
  assign y19827 = n27916 ;
  assign y19828 = ~1'b0 ;
  assign y19829 = n41284 ;
  assign y19830 = ~1'b0 ;
  assign y19831 = ~n41289 ;
  assign y19832 = ~n41290 ;
  assign y19833 = n41294 ;
  assign y19834 = ~n41299 ;
  assign y19835 = ~1'b0 ;
  assign y19836 = n41301 ;
  assign y19837 = ~n41306 ;
  assign y19838 = n41310 ;
  assign y19839 = ~n41314 ;
  assign y19840 = ~n41322 ;
  assign y19841 = ~n41324 ;
  assign y19842 = ~n41326 ;
  assign y19843 = ~1'b0 ;
  assign y19844 = ~1'b0 ;
  assign y19845 = ~n41329 ;
  assign y19846 = n41334 ;
  assign y19847 = ~n41336 ;
  assign y19848 = ~n41338 ;
  assign y19849 = n41342 ;
  assign y19850 = ~1'b0 ;
  assign y19851 = n36265 ;
  assign y19852 = ~n41343 ;
  assign y19853 = ~n41349 ;
  assign y19854 = n41352 ;
  assign y19855 = ~1'b0 ;
  assign y19856 = n41355 ;
  assign y19857 = ~n41370 ;
  assign y19858 = n41371 ;
  assign y19859 = ~1'b0 ;
  assign y19860 = ~n28442 ;
  assign y19861 = ~n41372 ;
  assign y19862 = ~n41376 ;
  assign y19863 = ~n40675 ;
  assign y19864 = ~1'b0 ;
  assign y19865 = n41377 ;
  assign y19866 = ~n41378 ;
  assign y19867 = ~1'b0 ;
  assign y19868 = n41379 ;
  assign y19869 = n41382 ;
  assign y19870 = ~1'b0 ;
  assign y19871 = ~1'b0 ;
  assign y19872 = n41386 ;
  assign y19873 = ~n41388 ;
  assign y19874 = ~n41389 ;
  assign y19875 = ~1'b0 ;
  assign y19876 = ~1'b0 ;
  assign y19877 = ~n41399 ;
  assign y19878 = n41402 ;
  assign y19879 = ~n41403 ;
  assign y19880 = n41405 ;
  assign y19881 = ~1'b0 ;
  assign y19882 = ~1'b0 ;
  assign y19883 = ~1'b0 ;
  assign y19884 = ~n41406 ;
  assign y19885 = ~n41408 ;
  assign y19886 = ~n36296 ;
  assign y19887 = ~n41409 ;
  assign y19888 = n41412 ;
  assign y19889 = ~n41416 ;
  assign y19890 = ~n41418 ;
  assign y19891 = 1'b0 ;
  assign y19892 = n41420 ;
  assign y19893 = ~n41422 ;
  assign y19894 = ~n41423 ;
  assign y19895 = n41427 ;
  assign y19896 = ~n34320 ;
  assign y19897 = n41429 ;
  assign y19898 = ~1'b0 ;
  assign y19899 = ~1'b0 ;
  assign y19900 = n41431 ;
  assign y19901 = n41436 ;
  assign y19902 = ~n41437 ;
  assign y19903 = ~n41440 ;
  assign y19904 = n41442 ;
  assign y19905 = ~1'b0 ;
  assign y19906 = ~n7363 ;
  assign y19907 = n41443 ;
  assign y19908 = n41445 ;
  assign y19909 = ~n41446 ;
  assign y19910 = ~1'b0 ;
  assign y19911 = n41449 ;
  assign y19912 = ~1'b0 ;
  assign y19913 = n41453 ;
  assign y19914 = ~n41456 ;
  assign y19915 = n41467 ;
  assign y19916 = n41468 ;
  assign y19917 = n41469 ;
  assign y19918 = ~1'b0 ;
  assign y19919 = n41473 ;
  assign y19920 = ~n41474 ;
  assign y19921 = n41478 ;
  assign y19922 = ~1'b0 ;
  assign y19923 = ~1'b0 ;
  assign y19924 = ~n41479 ;
  assign y19925 = ~n41480 ;
  assign y19926 = ~1'b0 ;
  assign y19927 = 1'b0 ;
  assign y19928 = ~1'b0 ;
  assign y19929 = ~1'b0 ;
  assign y19930 = n11660 ;
  assign y19931 = n41485 ;
  assign y19932 = n41489 ;
  assign y19933 = ~1'b0 ;
  assign y19934 = ~1'b0 ;
  assign y19935 = ~n41492 ;
  assign y19936 = ~1'b0 ;
  assign y19937 = n41498 ;
  assign y19938 = n41500 ;
  assign y19939 = n41503 ;
  assign y19940 = ~n41504 ;
  assign y19941 = 1'b0 ;
  assign y19942 = ~1'b0 ;
  assign y19943 = ~1'b0 ;
  assign y19944 = ~n41505 ;
  assign y19945 = n41507 ;
  assign y19946 = n41508 ;
  assign y19947 = ~n41509 ;
  assign y19948 = ~n41510 ;
  assign y19949 = ~1'b0 ;
  assign y19950 = n41511 ;
  assign y19951 = 1'b0 ;
  assign y19952 = ~n41514 ;
  assign y19953 = ~n41521 ;
  assign y19954 = ~n41523 ;
  assign y19955 = ~1'b0 ;
  assign y19956 = ~1'b0 ;
  assign y19957 = ~1'b0 ;
  assign y19958 = ~n41531 ;
  assign y19959 = ~1'b0 ;
  assign y19960 = ~n41533 ;
  assign y19961 = n41534 ;
  assign y19962 = ~n41535 ;
  assign y19963 = n22847 ;
  assign y19964 = n41537 ;
  assign y19965 = n7713 ;
  assign y19966 = n41539 ;
  assign y19967 = n41540 ;
  assign y19968 = ~n41542 ;
  assign y19969 = n41546 ;
  assign y19970 = ~n17203 ;
  assign y19971 = ~1'b0 ;
  assign y19972 = ~n41548 ;
  assign y19973 = ~n41550 ;
  assign y19974 = n41551 ;
  assign y19975 = ~n41554 ;
  assign y19976 = n41559 ;
  assign y19977 = ~n41560 ;
  assign y19978 = ~1'b0 ;
  assign y19979 = ~1'b0 ;
  assign y19980 = ~n41561 ;
  assign y19981 = ~n41565 ;
  assign y19982 = ~1'b0 ;
  assign y19983 = ~1'b0 ;
  assign y19984 = n41566 ;
  assign y19985 = n41568 ;
  assign y19986 = ~n41571 ;
  assign y19987 = ~n41572 ;
  assign y19988 = ~n41573 ;
  assign y19989 = ~n41576 ;
  assign y19990 = ~n41578 ;
  assign y19991 = ~1'b0 ;
  assign y19992 = ~n41579 ;
  assign y19993 = ~n41582 ;
  assign y19994 = n41583 ;
  assign y19995 = n41584 ;
  assign y19996 = n41587 ;
  assign y19997 = ~n41590 ;
  assign y19998 = ~1'b0 ;
  assign y19999 = ~1'b0 ;
  assign y20000 = n41592 ;
  assign y20001 = ~1'b0 ;
  assign y20002 = ~n41593 ;
  assign y20003 = n41594 ;
  assign y20004 = ~n41595 ;
  assign y20005 = ~n41596 ;
  assign y20006 = ~n41603 ;
  assign y20007 = ~n41604 ;
  assign y20008 = ~1'b0 ;
  assign y20009 = ~n41606 ;
  assign y20010 = n41607 ;
  assign y20011 = ~n41608 ;
  assign y20012 = n41612 ;
  assign y20013 = ~n41616 ;
  assign y20014 = ~n41620 ;
  assign y20015 = n41623 ;
  assign y20016 = ~n41626 ;
  assign y20017 = ~n41627 ;
  assign y20018 = n41629 ;
  assign y20019 = ~n41635 ;
  assign y20020 = ~n41638 ;
  assign y20021 = ~n41645 ;
  assign y20022 = ~n41647 ;
  assign y20023 = n41650 ;
  assign y20024 = n41654 ;
  assign y20025 = ~n41656 ;
  assign y20026 = n41658 ;
  assign y20027 = n25164 ;
  assign y20028 = ~1'b0 ;
  assign y20029 = n41660 ;
  assign y20030 = n41662 ;
  assign y20031 = n41667 ;
  assign y20032 = ~n41668 ;
  assign y20033 = n41672 ;
  assign y20034 = n41674 ;
  assign y20035 = n41678 ;
  assign y20036 = ~n41679 ;
  assign y20037 = n41682 ;
  assign y20038 = n41684 ;
  assign y20039 = ~n41686 ;
  assign y20040 = ~n22844 ;
  assign y20041 = ~1'b0 ;
  assign y20042 = ~n41688 ;
  assign y20043 = n41696 ;
  assign y20044 = 1'b0 ;
  assign y20045 = ~1'b0 ;
  assign y20046 = ~1'b0 ;
  assign y20047 = ~n41697 ;
  assign y20048 = n41702 ;
  assign y20049 = n41705 ;
  assign y20050 = n41706 ;
  assign y20051 = n41707 ;
  assign y20052 = n41710 ;
  assign y20053 = ~n41712 ;
  assign y20054 = ~1'b0 ;
  assign y20055 = n17296 ;
  assign y20056 = ~n41716 ;
  assign y20057 = ~1'b0 ;
  assign y20058 = ~n41718 ;
  assign y20059 = n41719 ;
  assign y20060 = ~n41721 ;
  assign y20061 = ~1'b0 ;
  assign y20062 = ~1'b0 ;
  assign y20063 = n41725 ;
  assign y20064 = ~n41727 ;
  assign y20065 = ~n41728 ;
  assign y20066 = n41729 ;
  assign y20067 = n41731 ;
  assign y20068 = n41733 ;
  assign y20069 = ~1'b0 ;
  assign y20070 = ~1'b0 ;
  assign y20071 = ~1'b0 ;
  assign y20072 = n18492 ;
  assign y20073 = n41736 ;
  assign y20074 = n41737 ;
  assign y20075 = ~n8346 ;
  assign y20076 = ~n41738 ;
  assign y20077 = ~n41739 ;
  assign y20078 = n41742 ;
  assign y20079 = n41744 ;
  assign y20080 = ~n41752 ;
  assign y20081 = n41753 ;
  assign y20082 = ~n41755 ;
  assign y20083 = n41756 ;
  assign y20084 = n41757 ;
  assign y20085 = ~1'b0 ;
  assign y20086 = ~1'b0 ;
  assign y20087 = n21339 ;
  assign y20088 = ~n41760 ;
  assign y20089 = 1'b0 ;
  assign y20090 = ~n41763 ;
  assign y20091 = n41766 ;
  assign y20092 = n41767 ;
  assign y20093 = ~n41773 ;
  assign y20094 = ~n41778 ;
  assign y20095 = ~n41780 ;
  assign y20096 = n41782 ;
  assign y20097 = 1'b0 ;
  assign y20098 = n41786 ;
  assign y20099 = ~n41788 ;
  assign y20100 = n41790 ;
  assign y20101 = n41793 ;
  assign y20102 = n41799 ;
  assign y20103 = ~n41802 ;
  assign y20104 = ~n34753 ;
  assign y20105 = ~n41804 ;
  assign y20106 = ~n41805 ;
  assign y20107 = ~1'b0 ;
  assign y20108 = ~n41806 ;
  assign y20109 = n41807 ;
  assign y20110 = ~1'b0 ;
  assign y20111 = ~1'b0 ;
  assign y20112 = n41811 ;
  assign y20113 = n41814 ;
  assign y20114 = ~1'b0 ;
  assign y20115 = ~n38422 ;
  assign y20116 = ~n41817 ;
  assign y20117 = ~n41822 ;
  assign y20118 = n41823 ;
  assign y20119 = n41828 ;
  assign y20120 = n41830 ;
  assign y20121 = ~n41831 ;
  assign y20122 = n41834 ;
  assign y20123 = ~n621 ;
  assign y20124 = n41835 ;
  assign y20125 = n41837 ;
  assign y20126 = n41839 ;
  assign y20127 = ~1'b0 ;
  assign y20128 = ~1'b0 ;
  assign y20129 = n41841 ;
  assign y20130 = n41842 ;
  assign y20131 = ~n41843 ;
  assign y20132 = ~n30299 ;
  assign y20133 = ~n41845 ;
  assign y20134 = n41847 ;
  assign y20135 = ~1'b0 ;
  assign y20136 = ~n41848 ;
  assign y20137 = n41850 ;
  assign y20138 = ~n41853 ;
  assign y20139 = n3337 ;
  assign y20140 = ~n41859 ;
  assign y20141 = ~n41861 ;
  assign y20142 = n41863 ;
  assign y20143 = ~1'b0 ;
  assign y20144 = ~1'b0 ;
  assign y20145 = n41864 ;
  assign y20146 = ~n41868 ;
  assign y20147 = ~n41869 ;
  assign y20148 = n41872 ;
  assign y20149 = ~n41879 ;
  assign y20150 = ~1'b0 ;
  assign y20151 = ~1'b0 ;
  assign y20152 = n17646 ;
  assign y20153 = ~n41881 ;
  assign y20154 = n41884 ;
  assign y20155 = n13248 ;
  assign y20156 = ~n41886 ;
  assign y20157 = ~1'b0 ;
  assign y20158 = ~1'b0 ;
  assign y20159 = n41888 ;
  assign y20160 = 1'b0 ;
  assign y20161 = n41889 ;
  assign y20162 = ~n6553 ;
  assign y20163 = ~1'b0 ;
  assign y20164 = ~n41890 ;
  assign y20165 = ~n41891 ;
  assign y20166 = ~n41892 ;
  assign y20167 = ~n41894 ;
  assign y20168 = n20362 ;
  assign y20169 = n41897 ;
  assign y20170 = n41900 ;
  assign y20171 = n41901 ;
  assign y20172 = ~n41904 ;
  assign y20173 = ~n41909 ;
  assign y20174 = ~1'b0 ;
  assign y20175 = n41911 ;
  assign y20176 = ~n41912 ;
  assign y20177 = ~n41914 ;
  assign y20178 = ~1'b0 ;
  assign y20179 = ~n41916 ;
  assign y20180 = ~n5942 ;
  assign y20181 = n41919 ;
  assign y20182 = n41926 ;
  assign y20183 = n37342 ;
  assign y20184 = ~n35342 ;
  assign y20185 = ~1'b0 ;
  assign y20186 = ~1'b0 ;
  assign y20187 = ~n41927 ;
  assign y20188 = ~n13911 ;
  assign y20189 = ~n41928 ;
  assign y20190 = n41929 ;
  assign y20191 = ~1'b0 ;
  assign y20192 = n41933 ;
  assign y20193 = n41935 ;
  assign y20194 = n41936 ;
  assign y20195 = n41940 ;
  assign y20196 = ~n12270 ;
  assign y20197 = n41946 ;
  assign y20198 = ~n41950 ;
  assign y20199 = n41951 ;
  assign y20200 = n41953 ;
  assign y20201 = n41956 ;
  assign y20202 = ~n41957 ;
  assign y20203 = n41958 ;
  assign y20204 = ~n41959 ;
  assign y20205 = ~1'b0 ;
  assign y20206 = ~n41961 ;
  assign y20207 = ~1'b0 ;
  assign y20208 = ~n41962 ;
  assign y20209 = n41963 ;
  assign y20210 = ~n41966 ;
  assign y20211 = ~1'b0 ;
  assign y20212 = n41968 ;
  assign y20213 = ~1'b0 ;
  assign y20214 = ~n41973 ;
  assign y20215 = ~n41974 ;
  assign y20216 = ~n41975 ;
  assign y20217 = ~n41981 ;
  assign y20218 = n41986 ;
  assign y20219 = n41987 ;
  assign y20220 = ~n41989 ;
  assign y20221 = ~n41991 ;
  assign y20222 = ~1'b0 ;
  assign y20223 = ~1'b0 ;
  assign y20224 = ~n41994 ;
  assign y20225 = ~1'b0 ;
  assign y20226 = ~n41995 ;
  assign y20227 = ~n39987 ;
  assign y20228 = ~n41997 ;
  assign y20229 = n42000 ;
  assign y20230 = n42004 ;
  assign y20231 = ~n42010 ;
  assign y20232 = ~n42015 ;
  assign y20233 = ~n31189 ;
  assign y20234 = n42017 ;
  assign y20235 = ~n42019 ;
  assign y20236 = ~n42021 ;
  assign y20237 = n42026 ;
  assign y20238 = ~n42027 ;
  assign y20239 = 1'b0 ;
  assign y20240 = n42028 ;
  assign y20241 = ~n42029 ;
  assign y20242 = n42033 ;
  assign y20243 = ~1'b0 ;
  assign y20244 = ~n42035 ;
  assign y20245 = ~1'b0 ;
  assign y20246 = n42037 ;
  assign y20247 = ~n42046 ;
  assign y20248 = ~n42048 ;
  assign y20249 = n42049 ;
  assign y20250 = ~n42050 ;
  assign y20251 = n42051 ;
  assign y20252 = ~n42053 ;
  assign y20253 = n37864 ;
  assign y20254 = 1'b0 ;
  assign y20255 = n42054 ;
  assign y20256 = ~n42056 ;
  assign y20257 = ~1'b0 ;
  assign y20258 = ~1'b0 ;
  assign y20259 = ~1'b0 ;
  assign y20260 = ~n42058 ;
  assign y20261 = ~n42060 ;
  assign y20262 = n42068 ;
  assign y20263 = n31592 ;
  assign y20264 = ~n42070 ;
  assign y20265 = ~1'b0 ;
  assign y20266 = n42078 ;
  assign y20267 = ~1'b0 ;
  assign y20268 = ~1'b0 ;
  assign y20269 = ~1'b0 ;
  assign y20270 = n42080 ;
  assign y20271 = n20989 ;
  assign y20272 = n42083 ;
  assign y20273 = n42086 ;
  assign y20274 = ~1'b0 ;
  assign y20275 = ~n42088 ;
  assign y20276 = ~1'b0 ;
  assign y20277 = n3355 ;
  assign y20278 = n42089 ;
  assign y20279 = n42090 ;
  assign y20280 = ~n9965 ;
  assign y20281 = n42096 ;
  assign y20282 = ~1'b0 ;
  assign y20283 = ~1'b0 ;
  assign y20284 = ~n42101 ;
  assign y20285 = n42103 ;
  assign y20286 = ~1'b0 ;
  assign y20287 = ~n42104 ;
  assign y20288 = n42107 ;
  assign y20289 = ~n42110 ;
  assign y20290 = ~n42116 ;
  assign y20291 = ~1'b0 ;
  assign y20292 = ~1'b0 ;
  assign y20293 = ~1'b0 ;
  assign y20294 = n42118 ;
  assign y20295 = ~n42119 ;
  assign y20296 = ~1'b0 ;
  assign y20297 = n42121 ;
  assign y20298 = ~1'b0 ;
  assign y20299 = ~n42122 ;
  assign y20300 = ~1'b0 ;
  assign y20301 = ~n42124 ;
  assign y20302 = ~n42126 ;
  assign y20303 = n42128 ;
  assign y20304 = n42129 ;
  assign y20305 = ~1'b0 ;
  assign y20306 = n42131 ;
  assign y20307 = 1'b0 ;
  assign y20308 = n42133 ;
  assign y20309 = ~n42135 ;
  assign y20310 = ~n42138 ;
  assign y20311 = ~1'b0 ;
  assign y20312 = ~n42143 ;
  assign y20313 = n42144 ;
  assign y20314 = ~1'b0 ;
  assign y20315 = n42154 ;
  assign y20316 = ~1'b0 ;
  assign y20317 = ~1'b0 ;
  assign y20318 = ~1'b0 ;
  assign y20319 = n42155 ;
  assign y20320 = ~n42159 ;
  assign y20321 = n42160 ;
  assign y20322 = ~n42163 ;
  assign y20323 = n42164 ;
  assign y20324 = ~1'b0 ;
  assign y20325 = ~1'b0 ;
  assign y20326 = ~1'b0 ;
  assign y20327 = ~1'b0 ;
  assign y20328 = n22277 ;
  assign y20329 = ~n34089 ;
  assign y20330 = ~1'b0 ;
  assign y20331 = ~n42165 ;
  assign y20332 = ~n42166 ;
  assign y20333 = ~1'b0 ;
  assign y20334 = n42170 ;
  assign y20335 = ~n42171 ;
  assign y20336 = ~1'b0 ;
  assign y20337 = ~1'b0 ;
  assign y20338 = n42174 ;
  assign y20339 = ~1'b0 ;
  assign y20340 = n42176 ;
  assign y20341 = ~n42181 ;
  assign y20342 = n42182 ;
  assign y20343 = ~n42184 ;
  assign y20344 = n42187 ;
  assign y20345 = ~1'b0 ;
  assign y20346 = n42188 ;
  assign y20347 = ~n42190 ;
  assign y20348 = ~n42193 ;
  assign y20349 = n30948 ;
  assign y20350 = n42199 ;
  assign y20351 = n42201 ;
  assign y20352 = ~1'b0 ;
  assign y20353 = n42203 ;
  assign y20354 = ~1'b0 ;
  assign y20355 = ~n42206 ;
  assign y20356 = n42207 ;
  assign y20357 = ~n42209 ;
  assign y20358 = n42211 ;
  assign y20359 = ~n42213 ;
  assign y20360 = ~n42214 ;
  assign y20361 = ~1'b0 ;
  assign y20362 = ~n42217 ;
  assign y20363 = ~n42218 ;
  assign y20364 = ~n42220 ;
  assign y20365 = n42222 ;
  assign y20366 = ~1'b0 ;
  assign y20367 = ~1'b0 ;
  assign y20368 = ~1'b0 ;
  assign y20369 = ~n33405 ;
  assign y20370 = n42230 ;
  assign y20371 = ~n42233 ;
  assign y20372 = ~n42235 ;
  assign y20373 = ~1'b0 ;
  assign y20374 = n42237 ;
  assign y20375 = ~1'b0 ;
  assign y20376 = ~n42240 ;
  assign y20377 = ~n42242 ;
  assign y20378 = n42247 ;
  assign y20379 = ~1'b0 ;
  assign y20380 = ~n42249 ;
  assign y20381 = ~n42252 ;
  assign y20382 = n42255 ;
  assign y20383 = ~1'b0 ;
  assign y20384 = n42256 ;
  assign y20385 = ~n36327 ;
  assign y20386 = ~n42260 ;
  assign y20387 = ~n42263 ;
  assign y20388 = ~1'b0 ;
  assign y20389 = ~n42266 ;
  assign y20390 = ~n42271 ;
  assign y20391 = ~n42272 ;
  assign y20392 = n42274 ;
  assign y20393 = ~n42275 ;
  assign y20394 = ~n42279 ;
  assign y20395 = ~1'b0 ;
  assign y20396 = n42284 ;
  assign y20397 = ~n42285 ;
  assign y20398 = ~1'b0 ;
  assign y20399 = n42286 ;
  assign y20400 = n42289 ;
  assign y20401 = n42295 ;
  assign y20402 = n42296 ;
  assign y20403 = ~1'b0 ;
  assign y20404 = ~1'b0 ;
  assign y20405 = ~1'b0 ;
  assign y20406 = n42297 ;
  assign y20407 = n23593 ;
  assign y20408 = n42300 ;
  assign y20409 = n42302 ;
  assign y20410 = ~1'b0 ;
  assign y20411 = ~n42303 ;
  assign y20412 = ~1'b0 ;
  assign y20413 = ~n17226 ;
  assign y20414 = n42306 ;
  assign y20415 = n42307 ;
  assign y20416 = n42309 ;
  assign y20417 = n42310 ;
  assign y20418 = ~n7863 ;
  assign y20419 = ~1'b0 ;
  assign y20420 = ~n42312 ;
  assign y20421 = n42314 ;
  assign y20422 = n42315 ;
  assign y20423 = ~1'b0 ;
  assign y20424 = ~n42316 ;
  assign y20425 = ~1'b0 ;
  assign y20426 = ~n42319 ;
  assign y20427 = 1'b0 ;
  assign y20428 = ~n42320 ;
  assign y20429 = n42325 ;
  assign y20430 = ~n42329 ;
  assign y20431 = n42330 ;
  assign y20432 = n42331 ;
  assign y20433 = ~n42333 ;
  assign y20434 = n19872 ;
  assign y20435 = ~n42340 ;
  assign y20436 = n17925 ;
  assign y20437 = n42342 ;
  assign y20438 = 1'b0 ;
  assign y20439 = ~n42343 ;
  assign y20440 = ~n42345 ;
  assign y20441 = n42349 ;
  assign y20442 = ~1'b0 ;
  assign y20443 = n42350 ;
  assign y20444 = n2229 ;
  assign y20445 = n42354 ;
  assign y20446 = ~n21691 ;
  assign y20447 = ~1'b0 ;
  assign y20448 = n42356 ;
  assign y20449 = ~1'b0 ;
  assign y20450 = ~1'b0 ;
  assign y20451 = ~n42358 ;
  assign y20452 = n42361 ;
  assign y20453 = ~n42362 ;
  assign y20454 = n42363 ;
  assign y20455 = ~n42364 ;
  assign y20456 = ~n42369 ;
  assign y20457 = n42375 ;
  assign y20458 = ~1'b0 ;
  assign y20459 = ~1'b0 ;
  assign y20460 = ~n42378 ;
  assign y20461 = ~1'b0 ;
  assign y20462 = n42379 ;
  assign y20463 = n42380 ;
  assign y20464 = n42382 ;
  assign y20465 = ~n42384 ;
  assign y20466 = ~n42386 ;
  assign y20467 = n42387 ;
  assign y20468 = ~n42389 ;
  assign y20469 = ~n42391 ;
  assign y20470 = ~n42394 ;
  assign y20471 = ~n42395 ;
  assign y20472 = n42396 ;
  assign y20473 = ~1'b0 ;
  assign y20474 = ~1'b0 ;
  assign y20475 = n42397 ;
  assign y20476 = n42398 ;
  assign y20477 = ~n42399 ;
  assign y20478 = ~1'b0 ;
  assign y20479 = n42400 ;
  assign y20480 = ~n42402 ;
  assign y20481 = ~n42406 ;
  assign y20482 = ~1'b0 ;
  assign y20483 = n42407 ;
  assign y20484 = ~1'b0 ;
  assign y20485 = ~1'b0 ;
  assign y20486 = ~n42409 ;
  assign y20487 = n42415 ;
  assign y20488 = ~1'b0 ;
  assign y20489 = ~n42417 ;
  assign y20490 = n42418 ;
  assign y20491 = ~1'b0 ;
  assign y20492 = ~n42419 ;
  assign y20493 = ~n42420 ;
  assign y20494 = n42421 ;
  assign y20495 = ~n42426 ;
  assign y20496 = n42427 ;
  assign y20497 = n42428 ;
  assign y20498 = ~n42435 ;
  assign y20499 = n42443 ;
  assign y20500 = ~1'b0 ;
  assign y20501 = n42447 ;
  assign y20502 = ~n42451 ;
  assign y20503 = ~n42452 ;
  assign y20504 = ~1'b0 ;
  assign y20505 = ~n42454 ;
  assign y20506 = n42455 ;
  assign y20507 = n42457 ;
  assign y20508 = ~1'b0 ;
  assign y20509 = ~n42463 ;
  assign y20510 = ~n42466 ;
  assign y20511 = ~n9332 ;
  assign y20512 = ~n42468 ;
  assign y20513 = ~n42473 ;
  assign y20514 = ~1'b0 ;
  assign y20515 = ~n42476 ;
  assign y20516 = n29413 ;
  assign y20517 = ~n42479 ;
  assign y20518 = ~1'b0 ;
  assign y20519 = n42481 ;
  assign y20520 = ~1'b0 ;
  assign y20521 = n19373 ;
  assign y20522 = ~1'b0 ;
  assign y20523 = ~1'b0 ;
  assign y20524 = ~1'b0 ;
  assign y20525 = n42483 ;
  assign y20526 = n42486 ;
  assign y20527 = ~1'b0 ;
  assign y20528 = ~1'b0 ;
  assign y20529 = 1'b0 ;
  assign y20530 = ~1'b0 ;
  assign y20531 = ~1'b0 ;
  assign y20532 = ~n42489 ;
  assign y20533 = ~1'b0 ;
  assign y20534 = ~n42490 ;
  assign y20535 = ~n42494 ;
  assign y20536 = ~n42495 ;
  assign y20537 = n42498 ;
  assign y20538 = n42499 ;
  assign y20539 = ~n42501 ;
  assign y20540 = n42502 ;
  assign y20541 = ~n42508 ;
  assign y20542 = n42509 ;
  assign y20543 = ~n42516 ;
  assign y20544 = n42517 ;
  assign y20545 = ~1'b0 ;
  assign y20546 = ~n42519 ;
  assign y20547 = n42524 ;
  assign y20548 = n42526 ;
  assign y20549 = ~n42531 ;
  assign y20550 = n42532 ;
  assign y20551 = n42538 ;
  assign y20552 = ~1'b0 ;
  assign y20553 = n42539 ;
  assign y20554 = ~1'b0 ;
  assign y20555 = ~1'b0 ;
  assign y20556 = ~n42543 ;
  assign y20557 = n42547 ;
  assign y20558 = ~1'b0 ;
  assign y20559 = ~1'b0 ;
  assign y20560 = ~n42550 ;
  assign y20561 = ~n42554 ;
  assign y20562 = ~n38421 ;
  assign y20563 = n42555 ;
  assign y20564 = n42559 ;
  assign y20565 = ~n42560 ;
  assign y20566 = ~n42561 ;
  assign y20567 = 1'b0 ;
  assign y20568 = ~n9132 ;
  assign y20569 = ~n42562 ;
  assign y20570 = n42563 ;
  assign y20571 = ~n42566 ;
  assign y20572 = ~n9365 ;
  assign y20573 = n42567 ;
  assign y20574 = ~n42568 ;
  assign y20575 = ~n42569 ;
  assign y20576 = ~n42570 ;
  assign y20577 = ~n42573 ;
  assign y20578 = n42575 ;
  assign y20579 = n42581 ;
  assign y20580 = n42582 ;
  assign y20581 = n42583 ;
  assign y20582 = ~1'b0 ;
  assign y20583 = ~1'b0 ;
  assign y20584 = n42584 ;
  assign y20585 = ~n42586 ;
  assign y20586 = ~n6409 ;
  assign y20587 = ~1'b0 ;
  assign y20588 = ~n1140 ;
  assign y20589 = ~1'b0 ;
  assign y20590 = ~1'b0 ;
  assign y20591 = n42590 ;
  assign y20592 = ~n42592 ;
  assign y20593 = n42593 ;
  assign y20594 = ~n15388 ;
  assign y20595 = n42594 ;
  assign y20596 = ~n42595 ;
  assign y20597 = ~1'b0 ;
  assign y20598 = ~1'b0 ;
  assign y20599 = n42600 ;
  assign y20600 = ~1'b0 ;
  assign y20601 = n20290 ;
  assign y20602 = ~n42604 ;
  assign y20603 = ~1'b0 ;
  assign y20604 = ~1'b0 ;
  assign y20605 = ~n42605 ;
  assign y20606 = ~1'b0 ;
  assign y20607 = ~n42607 ;
  assign y20608 = n30338 ;
  assign y20609 = ~n42611 ;
  assign y20610 = n42612 ;
  assign y20611 = ~n42614 ;
  assign y20612 = ~n42616 ;
  assign y20613 = n42618 ;
  assign y20614 = ~n42622 ;
  assign y20615 = ~n42626 ;
  assign y20616 = n42627 ;
  assign y20617 = n42630 ;
  assign y20618 = ~n42631 ;
  assign y20619 = 1'b0 ;
  assign y20620 = ~n42633 ;
  assign y20621 = ~n42635 ;
  assign y20622 = n42636 ;
  assign y20623 = ~n42637 ;
  assign y20624 = ~1'b0 ;
  assign y20625 = ~n42638 ;
  assign y20626 = n42640 ;
  assign y20627 = ~1'b0 ;
  assign y20628 = n42641 ;
  assign y20629 = ~1'b0 ;
  assign y20630 = ~n5010 ;
  assign y20631 = ~1'b0 ;
  assign y20632 = ~1'b0 ;
  assign y20633 = ~n42644 ;
  assign y20634 = ~n42645 ;
  assign y20635 = n42646 ;
  assign y20636 = n42648 ;
  assign y20637 = n42649 ;
  assign y20638 = n10950 ;
  assign y20639 = ~n42662 ;
  assign y20640 = ~1'b0 ;
  assign y20641 = n42666 ;
  assign y20642 = ~1'b0 ;
  assign y20643 = ~n42668 ;
  assign y20644 = ~n42670 ;
  assign y20645 = ~n42671 ;
  assign y20646 = n42673 ;
  assign y20647 = ~1'b0 ;
  assign y20648 = n42674 ;
  assign y20649 = ~n42675 ;
  assign y20650 = ~n42676 ;
  assign y20651 = ~n42679 ;
  assign y20652 = ~n42680 ;
  assign y20653 = ~1'b0 ;
  assign y20654 = n42681 ;
  assign y20655 = n42683 ;
  assign y20656 = ~1'b0 ;
  assign y20657 = n42685 ;
  assign y20658 = ~1'b0 ;
  assign y20659 = ~n42687 ;
  assign y20660 = n42691 ;
  assign y20661 = n42693 ;
  assign y20662 = ~1'b0 ;
  assign y20663 = ~1'b0 ;
  assign y20664 = ~n42695 ;
  assign y20665 = ~n42696 ;
  assign y20666 = n12608 ;
  assign y20667 = ~n42697 ;
  assign y20668 = ~n42699 ;
  assign y20669 = ~1'b0 ;
  assign y20670 = ~1'b0 ;
  assign y20671 = ~n11401 ;
  assign y20672 = ~1'b0 ;
  assign y20673 = ~n42705 ;
  assign y20674 = ~n42708 ;
  assign y20675 = ~n42712 ;
  assign y20676 = ~n42714 ;
  assign y20677 = ~n42720 ;
  assign y20678 = ~n42721 ;
  assign y20679 = ~n42723 ;
  assign y20680 = ~n42725 ;
  assign y20681 = ~n42727 ;
  assign y20682 = n42733 ;
  assign y20683 = ~n42734 ;
  assign y20684 = n42738 ;
  assign y20685 = n42743 ;
  assign y20686 = n42745 ;
  assign y20687 = ~1'b0 ;
  assign y20688 = 1'b0 ;
  assign y20689 = ~n6754 ;
  assign y20690 = n42751 ;
  assign y20691 = n42754 ;
  assign y20692 = ~1'b0 ;
  assign y20693 = n42758 ;
  assign y20694 = ~n42759 ;
  assign y20695 = ~n42761 ;
  assign y20696 = ~1'b0 ;
  assign y20697 = n42763 ;
  assign y20698 = ~n40659 ;
  assign y20699 = ~n42769 ;
  assign y20700 = ~n42771 ;
  assign y20701 = n42772 ;
  assign y20702 = n42774 ;
  assign y20703 = n42775 ;
  assign y20704 = n42780 ;
  assign y20705 = ~n42783 ;
  assign y20706 = n42792 ;
  assign y20707 = n42801 ;
  assign y20708 = n42802 ;
  assign y20709 = ~n42803 ;
  assign y20710 = ~n42807 ;
  assign y20711 = ~n42811 ;
  assign y20712 = ~n42812 ;
  assign y20713 = ~1'b0 ;
  assign y20714 = n42814 ;
  assign y20715 = ~n42819 ;
  assign y20716 = ~1'b0 ;
  assign y20717 = ~n3478 ;
  assign y20718 = ~n42823 ;
  assign y20719 = ~n42826 ;
  assign y20720 = ~n42828 ;
  assign y20721 = ~n42831 ;
  assign y20722 = n42833 ;
  assign y20723 = ~1'b0 ;
  assign y20724 = ~n42836 ;
  assign y20725 = n42840 ;
  assign y20726 = ~n42844 ;
  assign y20727 = ~1'b0 ;
  assign y20728 = n42845 ;
  assign y20729 = ~n42849 ;
  assign y20730 = ~n5741 ;
  assign y20731 = ~1'b0 ;
  assign y20732 = ~n27605 ;
  assign y20733 = n42853 ;
  assign y20734 = ~1'b0 ;
  assign y20735 = n42854 ;
  assign y20736 = ~1'b0 ;
  assign y20737 = ~n42859 ;
  assign y20738 = n42860 ;
  assign y20739 = ~n42861 ;
  assign y20740 = ~n42863 ;
  assign y20741 = ~1'b0 ;
  assign y20742 = ~n42869 ;
  assign y20743 = ~1'b0 ;
  assign y20744 = ~n42870 ;
  assign y20745 = ~n42871 ;
  assign y20746 = n42873 ;
  assign y20747 = n42874 ;
  assign y20748 = ~1'b0 ;
  assign y20749 = ~n42876 ;
  assign y20750 = n42882 ;
  assign y20751 = ~1'b0 ;
  assign y20752 = ~1'b0 ;
  assign y20753 = ~1'b0 ;
  assign y20754 = ~1'b0 ;
  assign y20755 = n42883 ;
  assign y20756 = ~n42884 ;
  assign y20757 = n42885 ;
  assign y20758 = ~1'b0 ;
  assign y20759 = ~1'b0 ;
  assign y20760 = ~1'b0 ;
  assign y20761 = ~n42890 ;
  assign y20762 = n42894 ;
  assign y20763 = n42895 ;
  assign y20764 = ~1'b0 ;
  assign y20765 = n42896 ;
  assign y20766 = ~n42899 ;
  assign y20767 = n42900 ;
  assign y20768 = ~1'b0 ;
  assign y20769 = n42902 ;
  assign y20770 = ~1'b0 ;
  assign y20771 = n42903 ;
  assign y20772 = n42904 ;
  assign y20773 = ~n42912 ;
  assign y20774 = ~1'b0 ;
  assign y20775 = ~n42914 ;
  assign y20776 = ~1'b0 ;
  assign y20777 = ~n17977 ;
  assign y20778 = ~n42915 ;
  assign y20779 = ~n42916 ;
  assign y20780 = ~n42918 ;
  assign y20781 = ~n42921 ;
  assign y20782 = n42922 ;
  assign y20783 = ~1'b0 ;
  assign y20784 = n42925 ;
  assign y20785 = n42931 ;
  assign y20786 = n42933 ;
  assign y20787 = ~1'b0 ;
  assign y20788 = ~1'b0 ;
  assign y20789 = ~1'b0 ;
  assign y20790 = ~n42934 ;
  assign y20791 = n42935 ;
  assign y20792 = n42936 ;
  assign y20793 = n42937 ;
  assign y20794 = ~1'b0 ;
  assign y20795 = 1'b0 ;
  assign y20796 = ~1'b0 ;
  assign y20797 = n42938 ;
  assign y20798 = 1'b0 ;
  assign y20799 = ~n42941 ;
  assign y20800 = n42948 ;
  assign y20801 = ~n42950 ;
  assign y20802 = ~n42952 ;
  assign y20803 = ~n42954 ;
  assign y20804 = ~n42956 ;
  assign y20805 = 1'b0 ;
  assign y20806 = 1'b0 ;
  assign y20807 = ~n42958 ;
  assign y20808 = n42959 ;
  assign y20809 = ~n42965 ;
  assign y20810 = n42969 ;
  assign y20811 = n42980 ;
  assign y20812 = ~1'b0 ;
  assign y20813 = ~1'b0 ;
  assign y20814 = n42986 ;
  assign y20815 = ~n42990 ;
  assign y20816 = ~n42992 ;
  assign y20817 = ~1'b0 ;
  assign y20818 = n42997 ;
  assign y20819 = n42999 ;
  assign y20820 = ~1'b0 ;
  assign y20821 = n12695 ;
  assign y20822 = n43000 ;
  assign y20823 = ~1'b0 ;
  assign y20824 = n43001 ;
  assign y20825 = n43006 ;
  assign y20826 = ~n43010 ;
  assign y20827 = ~1'b0 ;
  assign y20828 = 1'b0 ;
  assign y20829 = n43011 ;
  assign y20830 = ~1'b0 ;
  assign y20831 = ~1'b0 ;
  assign y20832 = ~n43013 ;
  assign y20833 = ~n43014 ;
  assign y20834 = ~n43016 ;
  assign y20835 = ~n23244 ;
  assign y20836 = n43017 ;
  assign y20837 = ~1'b0 ;
  assign y20838 = n43019 ;
  assign y20839 = n43022 ;
  assign y20840 = 1'b0 ;
  assign y20841 = n43025 ;
  assign y20842 = ~n43029 ;
  assign y20843 = ~n43031 ;
  assign y20844 = ~n43035 ;
  assign y20845 = ~1'b0 ;
  assign y20846 = ~1'b0 ;
  assign y20847 = ~n43036 ;
  assign y20848 = n43038 ;
  assign y20849 = n43039 ;
  assign y20850 = n43040 ;
  assign y20851 = ~n43045 ;
  assign y20852 = n43046 ;
  assign y20853 = ~n43047 ;
  assign y20854 = ~1'b0 ;
  assign y20855 = n43048 ;
  assign y20856 = n43052 ;
  assign y20857 = n43057 ;
  assign y20858 = n43060 ;
  assign y20859 = ~n43062 ;
  assign y20860 = n43070 ;
  assign y20861 = n43076 ;
  assign y20862 = ~n43078 ;
  assign y20863 = n43080 ;
  assign y20864 = ~n43082 ;
  assign y20865 = n43085 ;
  assign y20866 = ~n32989 ;
  assign y20867 = n43086 ;
  assign y20868 = n6175 ;
  assign y20869 = n43087 ;
  assign y20870 = ~1'b0 ;
  assign y20871 = n43094 ;
  assign y20872 = n43095 ;
  assign y20873 = ~n43096 ;
  assign y20874 = ~1'b0 ;
  assign y20875 = ~n43098 ;
  assign y20876 = n43102 ;
  assign y20877 = ~1'b0 ;
  assign y20878 = n43106 ;
  assign y20879 = ~n43108 ;
  assign y20880 = n43110 ;
  assign y20881 = ~n43113 ;
  assign y20882 = ~1'b0 ;
  assign y20883 = ~1'b0 ;
  assign y20884 = ~n43115 ;
  assign y20885 = ~n43118 ;
  assign y20886 = ~n43123 ;
  assign y20887 = ~n43124 ;
  assign y20888 = n43125 ;
  assign y20889 = ~n43126 ;
  assign y20890 = n43127 ;
  assign y20891 = ~1'b0 ;
  assign y20892 = n43128 ;
  assign y20893 = n43129 ;
  assign y20894 = ~n43131 ;
  assign y20895 = ~n43136 ;
  assign y20896 = n43138 ;
  assign y20897 = ~n43140 ;
  assign y20898 = ~1'b0 ;
  assign y20899 = n43141 ;
  assign y20900 = n43147 ;
  assign y20901 = ~n43150 ;
  assign y20902 = ~1'b0 ;
  assign y20903 = ~n43155 ;
  assign y20904 = n43157 ;
  assign y20905 = ~1'b0 ;
  assign y20906 = ~1'b0 ;
  assign y20907 = n43159 ;
  assign y20908 = ~n43160 ;
  assign y20909 = ~n43162 ;
  assign y20910 = n43164 ;
  assign y20911 = ~1'b0 ;
  assign y20912 = ~1'b0 ;
  assign y20913 = ~1'b0 ;
  assign y20914 = ~n43165 ;
  assign y20915 = n43170 ;
  assign y20916 = ~n11330 ;
  assign y20917 = ~1'b0 ;
  assign y20918 = ~n43180 ;
  assign y20919 = n6674 ;
  assign y20920 = ~n43181 ;
  assign y20921 = ~n43183 ;
  assign y20922 = n43185 ;
  assign y20923 = ~n6929 ;
  assign y20924 = ~n43186 ;
  assign y20925 = ~n3100 ;
  assign y20926 = n4211 ;
  assign y20927 = ~1'b0 ;
  assign y20928 = ~n43188 ;
  assign y20929 = ~n43189 ;
  assign y20930 = ~1'b0 ;
  assign y20931 = ~1'b0 ;
  assign y20932 = ~1'b0 ;
  assign y20933 = ~1'b0 ;
  assign y20934 = ~n43191 ;
  assign y20935 = ~n43192 ;
  assign y20936 = ~1'b0 ;
  assign y20937 = ~1'b0 ;
  assign y20938 = ~1'b0 ;
  assign y20939 = ~n5048 ;
  assign y20940 = n43197 ;
  assign y20941 = ~n43200 ;
  assign y20942 = ~n43201 ;
  assign y20943 = n43203 ;
  assign y20944 = n43211 ;
  assign y20945 = n43212 ;
  assign y20946 = ~1'b0 ;
  assign y20947 = ~1'b0 ;
  assign y20948 = n43214 ;
  assign y20949 = ~n43218 ;
  assign y20950 = ~n43220 ;
  assign y20951 = ~n43221 ;
  assign y20952 = ~1'b0 ;
  assign y20953 = ~n43222 ;
  assign y20954 = ~n43224 ;
  assign y20955 = ~n43227 ;
  assign y20956 = ~n43228 ;
  assign y20957 = ~n43231 ;
  assign y20958 = n43235 ;
  assign y20959 = n43242 ;
  assign y20960 = ~n43243 ;
  assign y20961 = n43244 ;
  assign y20962 = ~n43246 ;
  assign y20963 = n43248 ;
  assign y20964 = ~1'b0 ;
  assign y20965 = ~n43250 ;
  assign y20966 = ~n11065 ;
  assign y20967 = n43252 ;
  assign y20968 = ~1'b0 ;
  assign y20969 = ~n8115 ;
  assign y20970 = n43255 ;
  assign y20971 = n43256 ;
  assign y20972 = n43257 ;
  assign y20973 = n43258 ;
  assign y20974 = n43259 ;
  assign y20975 = ~1'b0 ;
  assign y20976 = n43263 ;
  assign y20977 = ~1'b0 ;
  assign y20978 = n43268 ;
  assign y20979 = ~1'b0 ;
  assign y20980 = ~1'b0 ;
  assign y20981 = ~n43270 ;
  assign y20982 = ~n43274 ;
  assign y20983 = ~n43279 ;
  assign y20984 = ~n37915 ;
  assign y20985 = ~n43283 ;
  assign y20986 = ~1'b0 ;
  assign y20987 = ~n43289 ;
  assign y20988 = ~n43294 ;
  assign y20989 = ~1'b0 ;
  assign y20990 = ~1'b0 ;
  assign y20991 = n43298 ;
  assign y20992 = n43299 ;
  assign y20993 = n43302 ;
  assign y20994 = ~n43308 ;
  assign y20995 = n43310 ;
  assign y20996 = ~n43314 ;
  assign y20997 = ~1'b0 ;
  assign y20998 = n43315 ;
  assign y20999 = n43317 ;
  assign y21000 = n43322 ;
  assign y21001 = ~n43327 ;
  assign y21002 = ~1'b0 ;
  assign y21003 = ~n43328 ;
  assign y21004 = ~n43329 ;
  assign y21005 = ~n43330 ;
  assign y21006 = ~1'b0 ;
  assign y21007 = ~1'b0 ;
  assign y21008 = n43331 ;
  assign y21009 = n43333 ;
  assign y21010 = ~n43337 ;
  assign y21011 = ~n33955 ;
  assign y21012 = n43342 ;
  assign y21013 = ~n43347 ;
  assign y21014 = ~1'b0 ;
  assign y21015 = ~1'b0 ;
  assign y21016 = n43348 ;
  assign y21017 = n43350 ;
  assign y21018 = ~1'b0 ;
  assign y21019 = n43352 ;
  assign y21020 = ~n43354 ;
  assign y21021 = n43359 ;
  assign y21022 = ~1'b0 ;
  assign y21023 = n43362 ;
  assign y21024 = ~1'b0 ;
  assign y21025 = n1019 ;
  assign y21026 = ~1'b0 ;
  assign y21027 = ~n43363 ;
  assign y21028 = ~n29073 ;
  assign y21029 = n43364 ;
  assign y21030 = ~n43367 ;
  assign y21031 = n43368 ;
  assign y21032 = n43370 ;
  assign y21033 = ~1'b0 ;
  assign y21034 = ~1'b0 ;
  assign y21035 = n22983 ;
  assign y21036 = ~n43373 ;
  assign y21037 = ~n43374 ;
  assign y21038 = n43375 ;
  assign y21039 = ~1'b0 ;
  assign y21040 = n43377 ;
  assign y21041 = n43378 ;
  assign y21042 = n43380 ;
  assign y21043 = ~1'b0 ;
  assign y21044 = ~1'b0 ;
  assign y21045 = n43387 ;
  assign y21046 = ~n43388 ;
  assign y21047 = ~n43389 ;
  assign y21048 = n43394 ;
  assign y21049 = ~1'b0 ;
  assign y21050 = ~1'b0 ;
  assign y21051 = n43396 ;
  assign y21052 = n43397 ;
  assign y21053 = ~n43398 ;
  assign y21054 = ~n43400 ;
  assign y21055 = ~n43403 ;
  assign y21056 = n43404 ;
  assign y21057 = ~n43407 ;
  assign y21058 = n43409 ;
  assign y21059 = ~1'b0 ;
  assign y21060 = ~1'b0 ;
  assign y21061 = ~n43415 ;
  assign y21062 = ~n43416 ;
  assign y21063 = ~n43421 ;
  assign y21064 = ~n43422 ;
  assign y21065 = ~n43423 ;
  assign y21066 = n43424 ;
  assign y21067 = ~1'b0 ;
  assign y21068 = ~1'b0 ;
  assign y21069 = ~n43426 ;
  assign y21070 = ~n43428 ;
  assign y21071 = ~n15627 ;
  assign y21072 = n43429 ;
  assign y21073 = ~n43432 ;
  assign y21074 = ~1'b0 ;
  assign y21075 = ~1'b0 ;
  assign y21076 = n43433 ;
  assign y21077 = n43434 ;
  assign y21078 = ~1'b0 ;
  assign y21079 = ~n43435 ;
  assign y21080 = ~n43440 ;
  assign y21081 = ~n43442 ;
  assign y21082 = n43448 ;
  assign y21083 = ~n43452 ;
  assign y21084 = ~n43457 ;
  assign y21085 = ~n43458 ;
  assign y21086 = ~1'b0 ;
  assign y21087 = ~n43462 ;
  assign y21088 = ~1'b0 ;
  assign y21089 = n43465 ;
  assign y21090 = n43466 ;
  assign y21091 = n11430 ;
  assign y21092 = n43468 ;
  assign y21093 = n43469 ;
  assign y21094 = ~n43471 ;
  assign y21095 = n43472 ;
  assign y21096 = ~1'b0 ;
  assign y21097 = n43474 ;
  assign y21098 = ~n43482 ;
  assign y21099 = n43484 ;
  assign y21100 = ~n43490 ;
  assign y21101 = n43492 ;
  assign y21102 = n43494 ;
  assign y21103 = n43495 ;
  assign y21104 = n43501 ;
  assign y21105 = n43505 ;
  assign y21106 = ~n43510 ;
  assign y21107 = ~n43513 ;
  assign y21108 = n43514 ;
  assign y21109 = n43521 ;
  assign y21110 = n43522 ;
  assign y21111 = ~1'b0 ;
  assign y21112 = ~n43526 ;
  assign y21113 = n43531 ;
  assign y21114 = ~n43532 ;
  assign y21115 = ~n43536 ;
  assign y21116 = ~n43543 ;
  assign y21117 = n21226 ;
  assign y21118 = ~n43547 ;
  assign y21119 = n43551 ;
  assign y21120 = ~n43553 ;
  assign y21121 = ~1'b0 ;
  assign y21122 = ~1'b0 ;
  assign y21123 = ~1'b0 ;
  assign y21124 = ~1'b0 ;
  assign y21125 = ~n43556 ;
  assign y21126 = ~n43558 ;
  assign y21127 = n43563 ;
  assign y21128 = n43566 ;
  assign y21129 = n43567 ;
  assign y21130 = ~1'b0 ;
  assign y21131 = 1'b0 ;
  assign y21132 = ~1'b0 ;
  assign y21133 = n43568 ;
  assign y21134 = n43574 ;
  assign y21135 = n43575 ;
  assign y21136 = ~1'b0 ;
  assign y21137 = n43579 ;
  assign y21138 = ~n43580 ;
  assign y21139 = ~n43583 ;
  assign y21140 = ~n20426 ;
  assign y21141 = ~n43584 ;
  assign y21142 = ~n43585 ;
  assign y21143 = ~1'b0 ;
  assign y21144 = n43586 ;
  assign y21145 = ~n43594 ;
  assign y21146 = ~n15566 ;
  assign y21147 = ~n43597 ;
  assign y21148 = n43600 ;
  assign y21149 = n43601 ;
  assign y21150 = n43603 ;
  assign y21151 = ~1'b0 ;
  assign y21152 = n10269 ;
  assign y21153 = n43604 ;
  assign y21154 = ~n43606 ;
  assign y21155 = ~1'b0 ;
  assign y21156 = n43610 ;
  assign y21157 = n43621 ;
  assign y21158 = ~n43622 ;
  assign y21159 = n16118 ;
  assign y21160 = ~n43627 ;
  assign y21161 = ~n43631 ;
  assign y21162 = n23304 ;
  assign y21163 = ~1'b0 ;
  assign y21164 = n43632 ;
  assign y21165 = ~n43635 ;
  assign y21166 = ~n43639 ;
  assign y21167 = n43643 ;
  assign y21168 = ~1'b0 ;
  assign y21169 = ~1'b0 ;
  assign y21170 = ~n43647 ;
  assign y21171 = n43650 ;
  assign y21172 = n43653 ;
  assign y21173 = ~1'b0 ;
  assign y21174 = ~n43655 ;
  assign y21175 = n43657 ;
  assign y21176 = n37483 ;
  assign y21177 = ~n43658 ;
  assign y21178 = n43662 ;
  assign y21179 = ~1'b0 ;
  assign y21180 = ~n43664 ;
  assign y21181 = ~1'b0 ;
  assign y21182 = n43669 ;
  assign y21183 = ~1'b0 ;
  assign y21184 = n43671 ;
  assign y21185 = ~n43672 ;
  assign y21186 = n43675 ;
  assign y21187 = ~n18793 ;
  assign y21188 = ~n43680 ;
  assign y21189 = n18485 ;
  assign y21190 = ~1'b0 ;
  assign y21191 = ~1'b0 ;
  assign y21192 = n36818 ;
  assign y21193 = ~n43681 ;
  assign y21194 = 1'b0 ;
  assign y21195 = ~n43682 ;
  assign y21196 = n43684 ;
  assign y21197 = n43685 ;
  assign y21198 = ~n43686 ;
  assign y21199 = ~n43689 ;
  assign y21200 = ~1'b0 ;
  assign y21201 = n43692 ;
  assign y21202 = ~n43693 ;
  assign y21203 = n43696 ;
  assign y21204 = ~1'b0 ;
  assign y21205 = n43700 ;
  assign y21206 = ~1'b0 ;
  assign y21207 = ~1'b0 ;
  assign y21208 = ~n43706 ;
  assign y21209 = 1'b0 ;
  assign y21210 = ~1'b0 ;
  assign y21211 = ~1'b0 ;
  assign y21212 = ~n43714 ;
  assign y21213 = ~n43717 ;
  assign y21214 = ~1'b0 ;
  assign y21215 = ~1'b0 ;
  assign y21216 = ~1'b0 ;
  assign y21217 = n43721 ;
  assign y21218 = ~n43722 ;
  assign y21219 = ~n43725 ;
  assign y21220 = ~1'b0 ;
  assign y21221 = ~1'b0 ;
  assign y21222 = n43726 ;
  assign y21223 = n43728 ;
  assign y21224 = 1'b0 ;
  assign y21225 = ~n43732 ;
  assign y21226 = n43733 ;
  assign y21227 = ~1'b0 ;
  assign y21228 = n2425 ;
  assign y21229 = ~1'b0 ;
  assign y21230 = ~1'b0 ;
  assign y21231 = ~1'b0 ;
  assign y21232 = ~n43736 ;
  assign y21233 = ~n43738 ;
  assign y21234 = ~1'b0 ;
  assign y21235 = n43741 ;
  assign y21236 = ~n43743 ;
  assign y21237 = ~n6369 ;
  assign y21238 = ~n43745 ;
  assign y21239 = n43747 ;
  assign y21240 = ~n43750 ;
  assign y21241 = ~n43752 ;
  assign y21242 = n43755 ;
  assign y21243 = n43758 ;
  assign y21244 = ~1'b0 ;
  assign y21245 = n43761 ;
  assign y21246 = n43762 ;
  assign y21247 = ~1'b0 ;
  assign y21248 = ~1'b0 ;
  assign y21249 = 1'b0 ;
  assign y21250 = n43764 ;
  assign y21251 = n32576 ;
  assign y21252 = ~1'b0 ;
  assign y21253 = ~1'b0 ;
  assign y21254 = n74 ;
  assign y21255 = ~n43766 ;
  assign y21256 = ~n43769 ;
  assign y21257 = ~n43771 ;
  assign y21258 = n43774 ;
  assign y21259 = ~n43775 ;
  assign y21260 = ~n43781 ;
  assign y21261 = ~1'b0 ;
  assign y21262 = ~n43783 ;
  assign y21263 = n43784 ;
  assign y21264 = ~1'b0 ;
  assign y21265 = n43787 ;
  assign y21266 = n43790 ;
  assign y21267 = ~n43791 ;
  assign y21268 = n43795 ;
  assign y21269 = ~n43797 ;
  assign y21270 = ~n43798 ;
  assign y21271 = n43802 ;
  assign y21272 = n13188 ;
  assign y21273 = ~1'b0 ;
  assign y21274 = ~n43803 ;
  assign y21275 = ~n43804 ;
  assign y21276 = ~n43806 ;
  assign y21277 = ~1'b0 ;
  assign y21278 = ~n43813 ;
  assign y21279 = ~1'b0 ;
  assign y21280 = n43814 ;
  assign y21281 = ~1'b0 ;
  assign y21282 = n43819 ;
  assign y21283 = n11138 ;
  assign y21284 = ~n43821 ;
  assign y21285 = ~n43826 ;
  assign y21286 = n43828 ;
  assign y21287 = ~1'b0 ;
  assign y21288 = 1'b0 ;
  assign y21289 = ~1'b0 ;
  assign y21290 = ~1'b0 ;
  assign y21291 = ~n43831 ;
  assign y21292 = n43832 ;
  assign y21293 = n43835 ;
  assign y21294 = ~1'b0 ;
  assign y21295 = ~n43839 ;
  assign y21296 = ~n43842 ;
  assign y21297 = ~n43846 ;
  assign y21298 = ~n43848 ;
  assign y21299 = ~n43849 ;
  assign y21300 = ~n43853 ;
  assign y21301 = ~n43856 ;
  assign y21302 = ~n43860 ;
  assign y21303 = n43861 ;
  assign y21304 = n43862 ;
  assign y21305 = n43864 ;
  assign y21306 = n43865 ;
  assign y21307 = ~1'b0 ;
  assign y21308 = ~1'b0 ;
  assign y21309 = ~n43868 ;
  assign y21310 = n43869 ;
  assign y21311 = ~1'b0 ;
  assign y21312 = ~n43870 ;
  assign y21313 = n43874 ;
  assign y21314 = n43876 ;
  assign y21315 = ~n43881 ;
  assign y21316 = ~n43883 ;
  assign y21317 = ~1'b0 ;
  assign y21318 = ~n43885 ;
  assign y21319 = ~n43887 ;
  assign y21320 = ~n43890 ;
  assign y21321 = n14460 ;
  assign y21322 = ~1'b0 ;
  assign y21323 = ~1'b0 ;
  assign y21324 = ~1'b0 ;
  assign y21325 = ~n30721 ;
  assign y21326 = n43891 ;
  assign y21327 = ~1'b0 ;
  assign y21328 = ~1'b0 ;
  assign y21329 = n43894 ;
  assign y21330 = n43901 ;
  assign y21331 = n43903 ;
  assign y21332 = n43908 ;
  assign y21333 = ~n43912 ;
  assign y21334 = n43914 ;
  assign y21335 = 1'b0 ;
  assign y21336 = ~n43916 ;
  assign y21337 = n43918 ;
  assign y21338 = ~n43281 ;
  assign y21339 = ~n43920 ;
  assign y21340 = ~n43923 ;
  assign y21341 = n43925 ;
  assign y21342 = 1'b0 ;
  assign y21343 = ~1'b0 ;
  assign y21344 = n43927 ;
  assign y21345 = ~n43929 ;
  assign y21346 = ~n43930 ;
  assign y21347 = ~1'b0 ;
  assign y21348 = n43932 ;
  assign y21349 = ~n43934 ;
  assign y21350 = n43935 ;
  assign y21351 = ~n43936 ;
  assign y21352 = ~n15311 ;
  assign y21353 = ~1'b0 ;
  assign y21354 = ~n43941 ;
  assign y21355 = ~1'b0 ;
  assign y21356 = ~1'b0 ;
  assign y21357 = n43945 ;
  assign y21358 = ~1'b0 ;
  assign y21359 = ~n43949 ;
  assign y21360 = ~n43950 ;
  assign y21361 = ~n43951 ;
  assign y21362 = n43953 ;
  assign y21363 = n43955 ;
  assign y21364 = ~n43956 ;
  assign y21365 = ~1'b0 ;
  assign y21366 = ~n43957 ;
  assign y21367 = n1875 ;
  assign y21368 = ~n43963 ;
  assign y21369 = ~n43965 ;
  assign y21370 = ~n43966 ;
  assign y21371 = ~n25648 ;
  assign y21372 = ~1'b0 ;
  assign y21373 = ~n43968 ;
  assign y21374 = ~n43970 ;
  assign y21375 = ~n43972 ;
  assign y21376 = ~n43976 ;
  assign y21377 = n43979 ;
  assign y21378 = ~n43980 ;
  assign y21379 = ~n43983 ;
  assign y21380 = ~n13421 ;
  assign y21381 = ~n43985 ;
  assign y21382 = ~1'b0 ;
  assign y21383 = 1'b0 ;
  assign y21384 = ~1'b0 ;
  assign y21385 = n43987 ;
  assign y21386 = n43990 ;
  assign y21387 = ~n43992 ;
  assign y21388 = ~n43993 ;
  assign y21389 = ~n43995 ;
  assign y21390 = n43998 ;
  assign y21391 = ~n44003 ;
  assign y21392 = n44004 ;
  assign y21393 = n44005 ;
  assign y21394 = ~n44006 ;
  assign y21395 = ~n44007 ;
  assign y21396 = n44008 ;
  assign y21397 = n44010 ;
  assign y21398 = ~1'b0 ;
  assign y21399 = ~n44012 ;
  assign y21400 = ~1'b0 ;
  assign y21401 = ~n44016 ;
  assign y21402 = ~n44018 ;
  assign y21403 = ~n44021 ;
  assign y21404 = n44022 ;
  assign y21405 = n44024 ;
  assign y21406 = n44027 ;
  assign y21407 = n44030 ;
  assign y21408 = ~1'b0 ;
  assign y21409 = ~1'b0 ;
  assign y21410 = n44031 ;
  assign y21411 = ~n44035 ;
  assign y21412 = ~n44037 ;
  assign y21413 = ~n44038 ;
  assign y21414 = ~n44040 ;
  assign y21415 = n44041 ;
  assign y21416 = n44051 ;
  assign y21417 = ~n44052 ;
  assign y21418 = n44053 ;
  assign y21419 = ~n44054 ;
  assign y21420 = n44055 ;
  assign y21421 = n44056 ;
  assign y21422 = ~n44059 ;
  assign y21423 = n44064 ;
  assign y21424 = n44066 ;
  assign y21425 = ~1'b0 ;
  assign y21426 = n44071 ;
  assign y21427 = n14375 ;
  assign y21428 = n44073 ;
  assign y21429 = ~1'b0 ;
  assign y21430 = ~n44078 ;
  assign y21431 = ~n44079 ;
  assign y21432 = n44086 ;
  assign y21433 = ~1'b0 ;
  assign y21434 = ~1'b0 ;
  assign y21435 = n44090 ;
  assign y21436 = n44096 ;
  assign y21437 = ~1'b0 ;
  assign y21438 = n44097 ;
  assign y21439 = ~n44099 ;
  assign y21440 = n44101 ;
  assign y21441 = n44105 ;
  assign y21442 = ~1'b0 ;
  assign y21443 = n44106 ;
  assign y21444 = ~n29154 ;
  assign y21445 = ~n44108 ;
  assign y21446 = ~n44110 ;
  assign y21447 = ~n44114 ;
  assign y21448 = ~n44121 ;
  assign y21449 = ~1'b0 ;
  assign y21450 = ~1'b0 ;
  assign y21451 = n44123 ;
  assign y21452 = ~n44125 ;
  assign y21453 = n44126 ;
  assign y21454 = ~1'b0 ;
  assign y21455 = ~n44129 ;
  assign y21456 = n44131 ;
  assign y21457 = ~n44132 ;
  assign y21458 = n44136 ;
  assign y21459 = ~1'b0 ;
  assign y21460 = ~1'b0 ;
  assign y21461 = ~n44139 ;
  assign y21462 = ~1'b0 ;
  assign y21463 = n44140 ;
  assign y21464 = n44141 ;
  assign y21465 = n44142 ;
  assign y21466 = ~n21429 ;
  assign y21467 = n44147 ;
  assign y21468 = n44150 ;
  assign y21469 = ~1'b0 ;
  assign y21470 = ~n44152 ;
  assign y21471 = n44157 ;
  assign y21472 = n44159 ;
  assign y21473 = ~1'b0 ;
  assign y21474 = ~n44161 ;
  assign y21475 = ~1'b0 ;
  assign y21476 = n44166 ;
  assign y21477 = n44167 ;
  assign y21478 = ~n44168 ;
  assign y21479 = n44171 ;
  assign y21480 = n44173 ;
  assign y21481 = ~n44181 ;
  assign y21482 = ~n44182 ;
  assign y21483 = ~n44184 ;
  assign y21484 = ~n44186 ;
  assign y21485 = n44187 ;
  assign y21486 = ~1'b0 ;
  assign y21487 = ~n44191 ;
  assign y21488 = ~n44195 ;
  assign y21489 = ~1'b0 ;
  assign y21490 = ~1'b0 ;
  assign y21491 = ~n44196 ;
  assign y21492 = ~1'b0 ;
  assign y21493 = ~n44201 ;
  assign y21494 = n44202 ;
  assign y21495 = ~n44206 ;
  assign y21496 = n44207 ;
  assign y21497 = ~n44209 ;
  assign y21498 = ~n44210 ;
  assign y21499 = n44211 ;
  assign y21500 = ~1'b0 ;
  assign y21501 = ~n44213 ;
  assign y21502 = n31634 ;
  assign y21503 = n41570 ;
  assign y21504 = n44216 ;
  assign y21505 = n44218 ;
  assign y21506 = ~1'b0 ;
  assign y21507 = ~n44220 ;
  assign y21508 = n2208 ;
  assign y21509 = 1'b0 ;
  assign y21510 = n44221 ;
  assign y21511 = n44222 ;
  assign y21512 = ~n44223 ;
  assign y21513 = n44224 ;
  assign y21514 = n44225 ;
  assign y21515 = n44230 ;
  assign y21516 = ~n44232 ;
  assign y21517 = ~1'b0 ;
  assign y21518 = ~1'b0 ;
  assign y21519 = ~1'b0 ;
  assign y21520 = n44235 ;
  assign y21521 = ~1'b0 ;
  assign y21522 = n44236 ;
  assign y21523 = ~n44239 ;
  assign y21524 = ~1'b0 ;
  assign y21525 = ~n44241 ;
  assign y21526 = ~n44243 ;
  assign y21527 = ~1'b0 ;
  assign y21528 = ~1'b0 ;
  assign y21529 = ~n44245 ;
  assign y21530 = n44246 ;
  assign y21531 = 1'b0 ;
  assign y21532 = n44249 ;
  assign y21533 = ~1'b0 ;
  assign y21534 = ~n44250 ;
  assign y21535 = n44253 ;
  assign y21536 = ~n44255 ;
  assign y21537 = ~n44256 ;
  assign y21538 = ~n9224 ;
  assign y21539 = ~n44258 ;
  assign y21540 = ~n44261 ;
  assign y21541 = ~n44263 ;
  assign y21542 = n44264 ;
  assign y21543 = ~1'b0 ;
  assign y21544 = n44266 ;
  assign y21545 = n44267 ;
  assign y21546 = n44270 ;
  assign y21547 = n44272 ;
  assign y21548 = n26566 ;
  assign y21549 = ~n44285 ;
  assign y21550 = n44289 ;
  assign y21551 = ~1'b0 ;
  assign y21552 = n44290 ;
  assign y21553 = ~1'b0 ;
  assign y21554 = ~1'b0 ;
  assign y21555 = ~1'b0 ;
  assign y21556 = n44291 ;
  assign y21557 = n44295 ;
  assign y21558 = n44299 ;
  assign y21559 = ~n44300 ;
  assign y21560 = n44301 ;
  assign y21561 = ~1'b0 ;
  assign y21562 = ~1'b0 ;
  assign y21563 = n44303 ;
  assign y21564 = ~n44305 ;
  assign y21565 = n44307 ;
  assign y21566 = n44310 ;
  assign y21567 = n44314 ;
  assign y21568 = n44316 ;
  assign y21569 = ~n13211 ;
  assign y21570 = ~1'b0 ;
  assign y21571 = n44321 ;
  assign y21572 = ~1'b0 ;
  assign y21573 = ~1'b0 ;
  assign y21574 = n44322 ;
  assign y21575 = ~n29995 ;
  assign y21576 = ~1'b0 ;
  assign y21577 = ~1'b0 ;
  assign y21578 = ~n44323 ;
  assign y21579 = ~1'b0 ;
  assign y21580 = ~1'b0 ;
  assign y21581 = ~n44330 ;
  assign y21582 = n44331 ;
  assign y21583 = ~n17441 ;
  assign y21584 = n44332 ;
  assign y21585 = ~n44335 ;
  assign y21586 = n44339 ;
  assign y21587 = ~1'b0 ;
  assign y21588 = n44343 ;
  assign y21589 = ~1'b0 ;
  assign y21590 = n44345 ;
  assign y21591 = ~n44349 ;
  assign y21592 = ~n44351 ;
  assign y21593 = ~1'b0 ;
  assign y21594 = ~1'b0 ;
  assign y21595 = ~n44356 ;
  assign y21596 = ~n44360 ;
  assign y21597 = n44365 ;
  assign y21598 = ~n44372 ;
  assign y21599 = ~n44374 ;
  assign y21600 = ~1'b0 ;
  assign y21601 = ~n44381 ;
  assign y21602 = ~n44383 ;
  assign y21603 = ~n44386 ;
  assign y21604 = n44396 ;
  assign y21605 = 1'b0 ;
  assign y21606 = n27136 ;
  assign y21607 = ~n44398 ;
  assign y21608 = n44402 ;
  assign y21609 = n21081 ;
  assign y21610 = n44404 ;
  assign y21611 = ~1'b0 ;
  assign y21612 = ~n44406 ;
  assign y21613 = n44409 ;
  assign y21614 = n7881 ;
  assign y21615 = ~1'b0 ;
  assign y21616 = ~n44414 ;
  assign y21617 = ~n44420 ;
  assign y21618 = ~1'b0 ;
  assign y21619 = n44425 ;
  assign y21620 = ~n44428 ;
  assign y21621 = ~n44431 ;
  assign y21622 = ~n44432 ;
  assign y21623 = ~1'b0 ;
  assign y21624 = n44435 ;
  assign y21625 = ~1'b0 ;
  assign y21626 = n44437 ;
  assign y21627 = n44440 ;
  assign y21628 = ~1'b0 ;
  assign y21629 = ~n44442 ;
  assign y21630 = ~n44444 ;
  assign y21631 = n44450 ;
  assign y21632 = ~n1465 ;
  assign y21633 = ~n206 ;
  assign y21634 = ~n44452 ;
  assign y21635 = n44455 ;
  assign y21636 = n44458 ;
  assign y21637 = ~n30369 ;
  assign y21638 = ~n44462 ;
  assign y21639 = ~n44463 ;
  assign y21640 = n44464 ;
  assign y21641 = n8950 ;
  assign y21642 = ~1'b0 ;
  assign y21643 = n44466 ;
  assign y21644 = ~n1172 ;
  assign y21645 = ~n44467 ;
  assign y21646 = n44468 ;
  assign y21647 = n44472 ;
  assign y21648 = n44473 ;
  assign y21649 = n44475 ;
  assign y21650 = n44477 ;
  assign y21651 = n44481 ;
  assign y21652 = ~n44485 ;
  assign y21653 = n44496 ;
  assign y21654 = ~n44500 ;
  assign y21655 = ~n44501 ;
  assign y21656 = n44504 ;
  assign y21657 = 1'b0 ;
  assign y21658 = n44506 ;
  assign y21659 = ~1'b0 ;
  assign y21660 = ~n44508 ;
  assign y21661 = ~n44510 ;
  assign y21662 = n44511 ;
  assign y21663 = ~n44513 ;
  assign y21664 = ~1'b0 ;
  assign y21665 = ~1'b0 ;
  assign y21666 = ~n44515 ;
  assign y21667 = ~1'b0 ;
  assign y21668 = n44516 ;
  assign y21669 = ~n44518 ;
  assign y21670 = n44519 ;
  assign y21671 = ~n44526 ;
  assign y21672 = ~n44528 ;
  assign y21673 = n39091 ;
  assign y21674 = n44530 ;
  assign y21675 = 1'b0 ;
  assign y21676 = n44532 ;
  assign y21677 = ~n44535 ;
  assign y21678 = ~n44536 ;
  assign y21679 = ~n44537 ;
  assign y21680 = ~n44538 ;
  assign y21681 = n44539 ;
  assign y21682 = n44540 ;
  assign y21683 = n44541 ;
  assign y21684 = ~1'b0 ;
  assign y21685 = n44543 ;
  assign y21686 = n8030 ;
  assign y21687 = ~n44544 ;
  assign y21688 = ~1'b0 ;
  assign y21689 = ~n2840 ;
  assign y21690 = n44546 ;
  assign y21691 = x4 ;
  assign y21692 = n44547 ;
  assign y21693 = n30991 ;
  assign y21694 = ~n44549 ;
  assign y21695 = ~1'b0 ;
  assign y21696 = n44550 ;
  assign y21697 = ~1'b0 ;
  assign y21698 = n44552 ;
  assign y21699 = ~1'b0 ;
  assign y21700 = ~n44553 ;
  assign y21701 = ~n44554 ;
  assign y21702 = ~n44556 ;
  assign y21703 = n44557 ;
  assign y21704 = ~n22094 ;
  assign y21705 = ~n44558 ;
  assign y21706 = ~1'b0 ;
  assign y21707 = ~1'b0 ;
  assign y21708 = n44560 ;
  assign y21709 = ~n44561 ;
  assign y21710 = n44564 ;
  assign y21711 = ~n44566 ;
  assign y21712 = n44570 ;
  assign y21713 = n44571 ;
  assign y21714 = n44574 ;
  assign y21715 = ~1'b0 ;
  assign y21716 = ~n44576 ;
  assign y21717 = ~1'b0 ;
  assign y21718 = ~1'b0 ;
  assign y21719 = ~n44578 ;
  assign y21720 = ~1'b0 ;
  assign y21721 = ~n44582 ;
  assign y21722 = n44586 ;
  assign y21723 = n37814 ;
  assign y21724 = ~1'b0 ;
  assign y21725 = n44589 ;
  assign y21726 = ~1'b0 ;
  assign y21727 = n44590 ;
  assign y21728 = ~n44591 ;
  assign y21729 = ~1'b0 ;
  assign y21730 = ~n44596 ;
  assign y21731 = ~1'b0 ;
  assign y21732 = ~n9975 ;
  assign y21733 = ~n44597 ;
  assign y21734 = ~n44600 ;
  assign y21735 = n44602 ;
  assign y21736 = 1'b0 ;
  assign y21737 = n44603 ;
  assign y21738 = n44605 ;
  assign y21739 = ~1'b0 ;
  assign y21740 = n44607 ;
  assign y21741 = n44611 ;
  assign y21742 = n44614 ;
  assign y21743 = n44615 ;
  assign y21744 = n10507 ;
  assign y21745 = ~n44619 ;
  assign y21746 = ~n44622 ;
  assign y21747 = ~1'b0 ;
  assign y21748 = ~n44626 ;
  assign y21749 = ~n44627 ;
  assign y21750 = ~n44631 ;
  assign y21751 = n44632 ;
  assign y21752 = ~n44635 ;
  assign y21753 = n44638 ;
  assign y21754 = n2581 ;
  assign y21755 = ~1'b0 ;
  assign y21756 = ~1'b0 ;
  assign y21757 = n44639 ;
  assign y21758 = ~n22142 ;
  assign y21759 = ~1'b0 ;
  assign y21760 = n44640 ;
  assign y21761 = ~n44641 ;
  assign y21762 = ~1'b0 ;
  assign y21763 = ~n44643 ;
  assign y21764 = n44644 ;
  assign y21765 = ~n44647 ;
  assign y21766 = ~n4044 ;
  assign y21767 = ~n44648 ;
  assign y21768 = ~1'b0 ;
  assign y21769 = n44650 ;
  assign y21770 = ~n44654 ;
  assign y21771 = ~n38341 ;
  assign y21772 = ~1'b0 ;
  assign y21773 = ~n44657 ;
  assign y21774 = n44663 ;
  assign y21775 = n44665 ;
  assign y21776 = n44669 ;
  assign y21777 = ~n44670 ;
  assign y21778 = ~n20648 ;
  assign y21779 = n44674 ;
  assign y21780 = ~n44675 ;
  assign y21781 = ~1'b0 ;
  assign y21782 = ~n9956 ;
  assign y21783 = ~n44677 ;
  assign y21784 = ~1'b0 ;
  assign y21785 = ~n44680 ;
  assign y21786 = ~n44682 ;
  assign y21787 = n44684 ;
  assign y21788 = n18504 ;
  assign y21789 = ~n44686 ;
  assign y21790 = n18669 ;
  assign y21791 = ~1'b0 ;
  assign y21792 = ~n44687 ;
  assign y21793 = ~n44691 ;
  assign y21794 = n44692 ;
  assign y21795 = ~n44694 ;
  assign y21796 = n44702 ;
  assign y21797 = n44703 ;
  assign y21798 = n44704 ;
  assign y21799 = n44706 ;
  assign y21800 = ~1'b0 ;
  assign y21801 = ~n44710 ;
  assign y21802 = ~n44712 ;
  assign y21803 = ~n9238 ;
  assign y21804 = ~1'b0 ;
  assign y21805 = n30995 ;
  assign y21806 = ~n44713 ;
  assign y21807 = n3523 ;
  assign y21808 = n44714 ;
  assign y21809 = ~1'b0 ;
  assign y21810 = ~n44717 ;
  assign y21811 = ~n44719 ;
  assign y21812 = ~1'b0 ;
  assign y21813 = ~n44720 ;
  assign y21814 = ~n44721 ;
  assign y21815 = ~1'b0 ;
  assign y21816 = ~1'b0 ;
  assign y21817 = ~n44722 ;
  assign y21818 = n44723 ;
  assign y21819 = n44727 ;
  assign y21820 = ~n44729 ;
  assign y21821 = ~1'b0 ;
  assign y21822 = ~1'b0 ;
  assign y21823 = ~1'b0 ;
  assign y21824 = ~1'b0 ;
  assign y21825 = ~1'b0 ;
  assign y21826 = ~n44731 ;
  assign y21827 = ~n44732 ;
  assign y21828 = n44736 ;
  assign y21829 = ~1'b0 ;
  assign y21830 = ~1'b0 ;
  assign y21831 = ~1'b0 ;
  assign y21832 = ~n44738 ;
  assign y21833 = ~n44739 ;
  assign y21834 = ~n44740 ;
  assign y21835 = n44744 ;
  assign y21836 = n44749 ;
  assign y21837 = n44752 ;
  assign y21838 = ~n44756 ;
  assign y21839 = ~n44760 ;
  assign y21840 = ~n44761 ;
  assign y21841 = ~n44762 ;
  assign y21842 = ~n44763 ;
  assign y21843 = ~1'b0 ;
  assign y21844 = ~n44764 ;
  assign y21845 = ~1'b0 ;
  assign y21846 = ~n44765 ;
  assign y21847 = n44766 ;
  assign y21848 = ~n44768 ;
  assign y21849 = n44769 ;
  assign y21850 = ~n44772 ;
  assign y21851 = n44773 ;
  assign y21852 = n44774 ;
  assign y21853 = n44776 ;
  assign y21854 = n44779 ;
  assign y21855 = n44781 ;
  assign y21856 = ~n44783 ;
  assign y21857 = ~n44785 ;
  assign y21858 = n44786 ;
  assign y21859 = ~n44792 ;
  assign y21860 = ~1'b0 ;
  assign y21861 = ~1'b0 ;
  assign y21862 = n44794 ;
  assign y21863 = ~n44797 ;
  assign y21864 = ~1'b0 ;
  assign y21865 = ~n44798 ;
  assign y21866 = ~1'b0 ;
  assign y21867 = ~n44800 ;
  assign y21868 = ~1'b0 ;
  assign y21869 = n44802 ;
  assign y21870 = ~n44805 ;
  assign y21871 = ~n27280 ;
  assign y21872 = ~n44806 ;
  assign y21873 = n3314 ;
  assign y21874 = n44809 ;
  assign y21875 = ~1'b0 ;
  assign y21876 = ~1'b0 ;
  assign y21877 = ~n44810 ;
  assign y21878 = ~n44815 ;
  assign y21879 = ~1'b0 ;
  assign y21880 = n44816 ;
  assign y21881 = n44818 ;
  assign y21882 = n44821 ;
  assign y21883 = ~1'b0 ;
  assign y21884 = ~1'b0 ;
  assign y21885 = n44824 ;
  assign y21886 = ~n44825 ;
  assign y21887 = ~n44828 ;
  assign y21888 = ~n44829 ;
  assign y21889 = n44832 ;
  assign y21890 = n44837 ;
  assign y21891 = n44840 ;
  assign y21892 = n43572 ;
  assign y21893 = n44841 ;
  assign y21894 = 1'b0 ;
  assign y21895 = ~1'b0 ;
  assign y21896 = ~1'b0 ;
  assign y21897 = ~n44842 ;
  assign y21898 = ~n44844 ;
  assign y21899 = n44847 ;
  assign y21900 = ~1'b0 ;
  assign y21901 = n44849 ;
  assign y21902 = ~1'b0 ;
  assign y21903 = ~1'b0 ;
  assign y21904 = ~n6167 ;
  assign y21905 = ~n44850 ;
  assign y21906 = n3306 ;
  assign y21907 = ~1'b0 ;
  assign y21908 = ~n44852 ;
  assign y21909 = ~1'b0 ;
  assign y21910 = ~n44854 ;
  assign y21911 = n44856 ;
  assign y21912 = ~n44859 ;
  assign y21913 = ~n44860 ;
  assign y21914 = ~1'b0 ;
  assign y21915 = ~1'b0 ;
  assign y21916 = ~1'b0 ;
  assign y21917 = ~n44863 ;
  assign y21918 = ~1'b0 ;
  assign y21919 = n130 ;
  assign y21920 = ~n44865 ;
  assign y21921 = ~n44866 ;
  assign y21922 = ~n44867 ;
  assign y21923 = n44868 ;
  assign y21924 = ~n44869 ;
  assign y21925 = ~n44871 ;
  assign y21926 = ~n44873 ;
  assign y21927 = ~1'b0 ;
  assign y21928 = ~1'b0 ;
  assign y21929 = ~n44874 ;
  assign y21930 = ~n44876 ;
  assign y21931 = ~n44878 ;
  assign y21932 = n44879 ;
  assign y21933 = n44886 ;
  assign y21934 = ~n44887 ;
  assign y21935 = n44889 ;
  assign y21936 = n44893 ;
  assign y21937 = ~n44896 ;
  assign y21938 = ~n44897 ;
  assign y21939 = ~n44905 ;
  assign y21940 = ~n44906 ;
  assign y21941 = n38608 ;
  assign y21942 = ~1'b0 ;
  assign y21943 = ~1'b0 ;
  assign y21944 = ~n44908 ;
  assign y21945 = ~n44911 ;
  assign y21946 = n44913 ;
  assign y21947 = ~n44916 ;
  assign y21948 = ~n12430 ;
  assign y21949 = n44917 ;
  assign y21950 = n44918 ;
  assign y21951 = n44921 ;
  assign y21952 = ~n44926 ;
  assign y21953 = n44928 ;
  assign y21954 = ~n28683 ;
  assign y21955 = ~1'b0 ;
  assign y21956 = n44933 ;
  assign y21957 = ~1'b0 ;
  assign y21958 = ~1'b0 ;
  assign y21959 = ~1'b0 ;
  assign y21960 = ~n44936 ;
  assign y21961 = ~1'b0 ;
  assign y21962 = ~n29303 ;
  assign y21963 = ~n44937 ;
  assign y21964 = ~n44942 ;
  assign y21965 = n44945 ;
  assign y21966 = ~n44947 ;
  assign y21967 = ~1'b0 ;
  assign y21968 = n44949 ;
  assign y21969 = n44950 ;
  assign y21970 = n44951 ;
  assign y21971 = n44952 ;
  assign y21972 = n44953 ;
  assign y21973 = ~1'b0 ;
  assign y21974 = ~n44955 ;
  assign y21975 = ~1'b0 ;
  assign y21976 = ~n44974 ;
  assign y21977 = ~n44980 ;
  assign y21978 = ~n44982 ;
  assign y21979 = ~1'b0 ;
  assign y21980 = ~n44983 ;
  assign y21981 = n44984 ;
  assign y21982 = n44985 ;
  assign y21983 = ~1'b0 ;
  assign y21984 = 1'b0 ;
  assign y21985 = ~n44986 ;
  assign y21986 = ~n44990 ;
  assign y21987 = n24908 ;
  assign y21988 = ~1'b0 ;
  assign y21989 = ~1'b0 ;
  assign y21990 = n44991 ;
  assign y21991 = n44994 ;
  assign y21992 = ~1'b0 ;
  assign y21993 = ~n44995 ;
  assign y21994 = n44996 ;
  assign y21995 = ~n45001 ;
  assign y21996 = ~1'b0 ;
  assign y21997 = n45002 ;
  assign y21998 = ~n45004 ;
  assign y21999 = ~n45008 ;
  assign y22000 = n45009 ;
  assign y22001 = ~1'b0 ;
  assign y22002 = ~1'b0 ;
  assign y22003 = n45012 ;
  assign y22004 = ~n45019 ;
  assign y22005 = ~n45020 ;
  assign y22006 = ~n45021 ;
  assign y22007 = ~n43365 ;
  assign y22008 = ~n45024 ;
  assign y22009 = ~1'b0 ;
  assign y22010 = ~1'b0 ;
  assign y22011 = ~n45025 ;
  assign y22012 = ~n45026 ;
  assign y22013 = ~1'b0 ;
  assign y22014 = ~n45027 ;
  assign y22015 = ~1'b0 ;
  assign y22016 = ~n45030 ;
  assign y22017 = ~n45033 ;
  assign y22018 = n45041 ;
  assign y22019 = n45042 ;
  assign y22020 = ~n45045 ;
  assign y22021 = ~n11346 ;
  assign y22022 = ~n45054 ;
  assign y22023 = n45056 ;
  assign y22024 = n45058 ;
  assign y22025 = n4336 ;
  assign y22026 = ~n45063 ;
  assign y22027 = ~n45067 ;
  assign y22028 = n45071 ;
  assign y22029 = n45076 ;
  assign y22030 = ~1'b0 ;
  assign y22031 = ~n45080 ;
  assign y22032 = n45083 ;
  assign y22033 = n45084 ;
  assign y22034 = ~n45086 ;
  assign y22035 = ~1'b0 ;
  assign y22036 = n45087 ;
  assign y22037 = ~1'b0 ;
  assign y22038 = ~1'b0 ;
  assign y22039 = n43886 ;
  assign y22040 = ~n45088 ;
  assign y22041 = ~1'b0 ;
  assign y22042 = ~1'b0 ;
  assign y22043 = ~1'b0 ;
  assign y22044 = n45092 ;
  assign y22045 = n45093 ;
  assign y22046 = n45097 ;
  assign y22047 = n45100 ;
  assign y22048 = n45103 ;
  assign y22049 = n45104 ;
  assign y22050 = ~n45107 ;
  assign y22051 = ~n45110 ;
  assign y22052 = n45114 ;
  assign y22053 = ~n45117 ;
  assign y22054 = ~1'b0 ;
  assign y22055 = ~n45123 ;
  assign y22056 = ~1'b0 ;
  assign y22057 = n45130 ;
  assign y22058 = ~1'b0 ;
  assign y22059 = n45132 ;
  assign y22060 = ~n45134 ;
  assign y22061 = ~n45137 ;
  assign y22062 = ~n45138 ;
  assign y22063 = n45139 ;
  assign y22064 = ~1'b0 ;
  assign y22065 = ~n45141 ;
  assign y22066 = n45145 ;
  assign y22067 = ~1'b0 ;
  assign y22068 = n12101 ;
  assign y22069 = n45147 ;
  assign y22070 = ~1'b0 ;
  assign y22071 = ~1'b0 ;
  assign y22072 = n45151 ;
  assign y22073 = n45152 ;
  assign y22074 = ~1'b0 ;
  assign y22075 = ~1'b0 ;
  assign y22076 = n45155 ;
  assign y22077 = ~1'b0 ;
  assign y22078 = n45157 ;
  assign y22079 = ~1'b0 ;
  assign y22080 = ~1'b0 ;
  assign y22081 = n45160 ;
  assign y22082 = n45162 ;
  assign y22083 = ~1'b0 ;
  assign y22084 = n45167 ;
  assign y22085 = n45170 ;
  assign y22086 = ~n45172 ;
  assign y22087 = ~1'b0 ;
  assign y22088 = ~n23023 ;
  assign y22089 = ~1'b0 ;
  assign y22090 = n45176 ;
  assign y22091 = n45177 ;
  assign y22092 = ~n45178 ;
  assign y22093 = n45180 ;
  assign y22094 = ~1'b0 ;
  assign y22095 = ~1'b0 ;
  assign y22096 = n45182 ;
  assign y22097 = n45183 ;
  assign y22098 = n45185 ;
  assign y22099 = n45187 ;
  assign y22100 = n45194 ;
  assign y22101 = ~n45200 ;
  assign y22102 = ~1'b0 ;
  assign y22103 = n45204 ;
  assign y22104 = ~1'b0 ;
  assign y22105 = n45205 ;
  assign y22106 = ~1'b0 ;
  assign y22107 = n45210 ;
  assign y22108 = n45212 ;
  assign y22109 = n45214 ;
  assign y22110 = ~n45216 ;
  assign y22111 = ~n45217 ;
  assign y22112 = ~n45218 ;
  assign y22113 = n45226 ;
  assign y22114 = n45229 ;
  assign y22115 = ~1'b0 ;
  assign y22116 = ~n45233 ;
  assign y22117 = n45237 ;
  assign y22118 = n45239 ;
  assign y22119 = ~n45240 ;
  assign y22120 = ~n45241 ;
  assign y22121 = ~n45242 ;
  assign y22122 = ~1'b0 ;
  assign y22123 = ~1'b0 ;
  assign y22124 = ~n45246 ;
  assign y22125 = ~n45247 ;
  assign y22126 = n45249 ;
  assign y22127 = ~1'b0 ;
  assign y22128 = ~n45254 ;
  assign y22129 = ~n45257 ;
  assign y22130 = n45258 ;
  assign y22131 = n45261 ;
  assign y22132 = n45264 ;
  assign y22133 = ~1'b0 ;
  assign y22134 = n45267 ;
  assign y22135 = ~n45268 ;
  assign y22136 = ~1'b0 ;
  assign y22137 = n45269 ;
  assign y22138 = ~1'b0 ;
  assign y22139 = ~1'b0 ;
  assign y22140 = ~1'b0 ;
  assign y22141 = ~n45278 ;
  assign y22142 = ~n45284 ;
  assign y22143 = ~n45285 ;
  assign y22144 = n45286 ;
  assign y22145 = n45287 ;
  assign y22146 = n45290 ;
  assign y22147 = n45293 ;
  assign y22148 = ~n45297 ;
  assign y22149 = n45298 ;
  assign y22150 = ~1'b0 ;
  assign y22151 = ~n45307 ;
  assign y22152 = ~n45309 ;
  assign y22153 = ~n45311 ;
  assign y22154 = ~n45314 ;
  assign y22155 = ~n45315 ;
  assign y22156 = n45318 ;
  assign y22157 = n45320 ;
  assign y22158 = ~1'b0 ;
  assign y22159 = ~n45322 ;
  assign y22160 = n45324 ;
  assign y22161 = ~n21431 ;
  assign y22162 = n45329 ;
  assign y22163 = ~1'b0 ;
  assign y22164 = ~n45332 ;
  assign y22165 = ~n45333 ;
  assign y22166 = ~n45335 ;
  assign y22167 = ~1'b0 ;
  assign y22168 = n45338 ;
  assign y22169 = n45339 ;
  assign y22170 = n45340 ;
  assign y22171 = n45344 ;
  assign y22172 = ~n45346 ;
  assign y22173 = n45348 ;
  assign y22174 = n45350 ;
  assign y22175 = ~1'b0 ;
  assign y22176 = n45352 ;
  assign y22177 = n45354 ;
  assign y22178 = n45357 ;
  assign y22179 = ~1'b0 ;
  assign y22180 = ~n45359 ;
  assign y22181 = n45360 ;
  assign y22182 = ~n45362 ;
  assign y22183 = ~n45363 ;
  assign y22184 = n45366 ;
  assign y22185 = ~1'b0 ;
  assign y22186 = ~1'b0 ;
  assign y22187 = ~n45368 ;
  assign y22188 = ~1'b0 ;
  assign y22189 = ~1'b0 ;
  assign y22190 = ~1'b0 ;
  assign y22191 = ~n45371 ;
  assign y22192 = n45372 ;
  assign y22193 = n45380 ;
  assign y22194 = n45387 ;
  assign y22195 = ~1'b0 ;
  assign y22196 = ~1'b0 ;
  assign y22197 = ~1'b0 ;
  assign y22198 = n45388 ;
  assign y22199 = n45390 ;
  assign y22200 = 1'b0 ;
  assign y22201 = n45391 ;
  assign y22202 = n45395 ;
  assign y22203 = n45397 ;
  assign y22204 = ~1'b0 ;
  assign y22205 = ~n45399 ;
  assign y22206 = n45400 ;
  assign y22207 = ~n45403 ;
  assign y22208 = ~n5531 ;
  assign y22209 = n13684 ;
  assign y22210 = ~1'b0 ;
  assign y22211 = ~1'b0 ;
  assign y22212 = ~n45405 ;
  assign y22213 = ~n45408 ;
  assign y22214 = ~n45409 ;
  assign y22215 = ~n45410 ;
  assign y22216 = n45415 ;
  assign y22217 = n45416 ;
  assign y22218 = n12696 ;
  assign y22219 = ~1'b0 ;
  assign y22220 = ~1'b0 ;
  assign y22221 = ~n45418 ;
  assign y22222 = ~n45421 ;
  assign y22223 = ~1'b0 ;
  assign y22224 = n45422 ;
  assign y22225 = n45425 ;
  assign y22226 = n45427 ;
  assign y22227 = n45432 ;
  assign y22228 = ~n45437 ;
  assign y22229 = ~n45438 ;
  assign y22230 = ~1'b0 ;
  assign y22231 = ~n45440 ;
  assign y22232 = ~n45443 ;
  assign y22233 = ~n45444 ;
  assign y22234 = ~n45445 ;
  assign y22235 = ~n35111 ;
  assign y22236 = ~1'b0 ;
  assign y22237 = n45447 ;
  assign y22238 = ~1'b0 ;
  assign y22239 = ~1'b0 ;
  assign y22240 = ~n45452 ;
  assign y22241 = ~n45459 ;
  assign y22242 = ~n45461 ;
  assign y22243 = ~1'b0 ;
  assign y22244 = n45464 ;
  assign y22245 = ~n45467 ;
  assign y22246 = n45469 ;
  assign y22247 = 1'b0 ;
  assign y22248 = ~1'b0 ;
  assign y22249 = n45471 ;
  assign y22250 = ~n45473 ;
  assign y22251 = n45474 ;
  assign y22252 = n45480 ;
  assign y22253 = ~1'b0 ;
  assign y22254 = ~1'b0 ;
  assign y22255 = ~1'b0 ;
  assign y22256 = ~1'b0 ;
  assign y22257 = ~1'b0 ;
  assign y22258 = ~n45484 ;
  assign y22259 = n30162 ;
  assign y22260 = n45488 ;
  assign y22261 = ~1'b0 ;
  assign y22262 = n45491 ;
  assign y22263 = ~n45493 ;
  assign y22264 = 1'b0 ;
  assign y22265 = ~1'b0 ;
  assign y22266 = ~1'b0 ;
  assign y22267 = ~n45498 ;
  assign y22268 = ~1'b0 ;
  assign y22269 = ~1'b0 ;
  assign y22270 = n45499 ;
  assign y22271 = ~n45502 ;
  assign y22272 = ~1'b0 ;
  assign y22273 = ~n45503 ;
  assign y22274 = ~1'b0 ;
  assign y22275 = n45504 ;
  assign y22276 = ~n45505 ;
  assign y22277 = ~n30753 ;
  assign y22278 = n45507 ;
  assign y22279 = n45508 ;
  assign y22280 = n45510 ;
  assign y22281 = 1'b0 ;
  assign y22282 = n45512 ;
  assign y22283 = ~1'b0 ;
  assign y22284 = ~n42443 ;
  assign y22285 = n45515 ;
  assign y22286 = ~n5654 ;
  assign y22287 = n45519 ;
  assign y22288 = n45523 ;
  assign y22289 = ~1'b0 ;
  assign y22290 = ~n45525 ;
  assign y22291 = ~n45526 ;
  assign y22292 = n45528 ;
  assign y22293 = ~1'b0 ;
  assign y22294 = ~n45529 ;
  assign y22295 = ~n45531 ;
  assign y22296 = n45532 ;
  assign y22297 = n45534 ;
  assign y22298 = n45535 ;
  assign y22299 = ~n45537 ;
  assign y22300 = n45539 ;
  assign y22301 = ~1'b0 ;
  assign y22302 = ~n45547 ;
  assign y22303 = n45551 ;
  assign y22304 = n45552 ;
  assign y22305 = ~1'b0 ;
  assign y22306 = ~n45554 ;
  assign y22307 = n45557 ;
  assign y22308 = n45562 ;
  assign y22309 = ~n45567 ;
  assign y22310 = ~1'b0 ;
  assign y22311 = ~n45572 ;
  assign y22312 = n45575 ;
  assign y22313 = ~1'b0 ;
  assign y22314 = ~n45578 ;
  assign y22315 = ~n45579 ;
  assign y22316 = n45580 ;
  assign y22317 = ~n45582 ;
  assign y22318 = ~n45584 ;
  assign y22319 = n45587 ;
  assign y22320 = ~n42985 ;
  assign y22321 = n45588 ;
  assign y22322 = ~n45589 ;
  assign y22323 = n13585 ;
  assign y22324 = ~1'b0 ;
  assign y22325 = 1'b0 ;
  assign y22326 = ~1'b0 ;
  assign y22327 = ~1'b0 ;
  assign y22328 = ~n45596 ;
  assign y22329 = n45597 ;
  assign y22330 = ~n17628 ;
  assign y22331 = ~n45598 ;
  assign y22332 = ~1'b0 ;
  assign y22333 = ~1'b0 ;
  assign y22334 = ~1'b0 ;
  assign y22335 = n45602 ;
  assign y22336 = ~n45603 ;
  assign y22337 = n45608 ;
  assign y22338 = n45613 ;
  assign y22339 = ~n45614 ;
  assign y22340 = n45617 ;
  assign y22341 = ~n45619 ;
  assign y22342 = n45620 ;
  assign y22343 = ~n45623 ;
  assign y22344 = ~n45624 ;
  assign y22345 = n45625 ;
  assign y22346 = ~n45628 ;
  assign y22347 = n45630 ;
  assign y22348 = ~n45632 ;
  assign y22349 = ~n45637 ;
  assign y22350 = n45638 ;
  assign y22351 = ~n45639 ;
  assign y22352 = n45642 ;
  assign y22353 = n9687 ;
  assign y22354 = ~n45644 ;
  assign y22355 = ~1'b0 ;
  assign y22356 = ~1'b0 ;
  assign y22357 = ~1'b0 ;
  assign y22358 = n45648 ;
  assign y22359 = ~n45650 ;
  assign y22360 = n45653 ;
  assign y22361 = ~n45654 ;
  assign y22362 = ~n45655 ;
  assign y22363 = ~1'b0 ;
  assign y22364 = n45658 ;
  assign y22365 = ~1'b0 ;
  assign y22366 = ~n45659 ;
  assign y22367 = n45663 ;
  assign y22368 = ~n45664 ;
  assign y22369 = ~n45669 ;
  assign y22370 = ~n45672 ;
  assign y22371 = ~1'b0 ;
  assign y22372 = ~n45674 ;
  assign y22373 = n45677 ;
  assign y22374 = n398 ;
  assign y22375 = n45680 ;
  assign y22376 = ~n45683 ;
  assign y22377 = ~n45689 ;
  assign y22378 = ~1'b0 ;
  assign y22379 = ~1'b0 ;
  assign y22380 = ~n45691 ;
  assign y22381 = ~1'b0 ;
  assign y22382 = n45692 ;
  assign y22383 = ~1'b0 ;
  assign y22384 = ~1'b0 ;
  assign y22385 = ~n45697 ;
  assign y22386 = ~n45699 ;
  assign y22387 = ~1'b0 ;
  assign y22388 = ~1'b0 ;
  assign y22389 = ~1'b0 ;
  assign y22390 = ~1'b0 ;
  assign y22391 = n45702 ;
  assign y22392 = ~n45703 ;
  assign y22393 = ~1'b0 ;
  assign y22394 = ~n45704 ;
  assign y22395 = n45705 ;
  assign y22396 = n45707 ;
  assign y22397 = ~n45709 ;
  assign y22398 = ~1'b0 ;
  assign y22399 = ~n45713 ;
  assign y22400 = ~n45720 ;
  assign y22401 = n45722 ;
  assign y22402 = ~n45725 ;
  assign y22403 = n45727 ;
  assign y22404 = n45729 ;
  assign y22405 = ~n45730 ;
  assign y22406 = ~n45732 ;
  assign y22407 = ~1'b0 ;
  assign y22408 = 1'b0 ;
  assign y22409 = ~n45733 ;
  assign y22410 = ~n12543 ;
  assign y22411 = ~1'b0 ;
  assign y22412 = ~n45740 ;
  assign y22413 = ~1'b0 ;
  assign y22414 = ~1'b0 ;
  assign y22415 = ~1'b0 ;
  assign y22416 = ~n45741 ;
  assign y22417 = ~n45743 ;
  assign y22418 = ~n45749 ;
  assign y22419 = ~n45755 ;
  assign y22420 = ~1'b0 ;
  assign y22421 = ~n45756 ;
  assign y22422 = n45757 ;
  assign y22423 = ~n45759 ;
  assign y22424 = n45761 ;
  assign y22425 = ~n45768 ;
  assign y22426 = ~1'b0 ;
  assign y22427 = n45769 ;
  assign y22428 = n45772 ;
  assign y22429 = ~1'b0 ;
  assign y22430 = ~1'b0 ;
  assign y22431 = ~1'b0 ;
  assign y22432 = ~n45774 ;
  assign y22433 = ~1'b0 ;
  assign y22434 = ~1'b0 ;
  assign y22435 = ~n27334 ;
  assign y22436 = ~1'b0 ;
  assign y22437 = 1'b0 ;
  assign y22438 = n45775 ;
  assign y22439 = n45776 ;
  assign y22440 = ~n45780 ;
  assign y22441 = ~n45784 ;
  assign y22442 = n45789 ;
  assign y22443 = n45799 ;
  assign y22444 = ~n11207 ;
  assign y22445 = ~n45804 ;
  assign y22446 = ~n45806 ;
  assign y22447 = ~1'b0 ;
  assign y22448 = ~n45811 ;
  assign y22449 = ~1'b0 ;
  assign y22450 = n7319 ;
  assign y22451 = n45812 ;
  assign y22452 = ~n17839 ;
  assign y22453 = n45817 ;
  assign y22454 = ~n45819 ;
  assign y22455 = ~n45820 ;
  assign y22456 = n45821 ;
  assign y22457 = ~1'b0 ;
  assign y22458 = ~1'b0 ;
  assign y22459 = n45823 ;
  assign y22460 = ~n45826 ;
  assign y22461 = ~n27433 ;
  assign y22462 = ~1'b0 ;
  assign y22463 = ~n45827 ;
  assign y22464 = n45830 ;
  assign y22465 = n45831 ;
  assign y22466 = ~1'b0 ;
  assign y22467 = ~1'b0 ;
  assign y22468 = ~1'b0 ;
  assign y22469 = ~n45834 ;
  assign y22470 = n45835 ;
  assign y22471 = n45836 ;
  assign y22472 = ~n45837 ;
  assign y22473 = n45839 ;
  assign y22474 = n45842 ;
  assign y22475 = ~n45843 ;
  assign y22476 = ~1'b0 ;
  assign y22477 = n45844 ;
  assign y22478 = n45849 ;
  assign y22479 = ~n18089 ;
  assign y22480 = n45851 ;
  assign y22481 = n45852 ;
  assign y22482 = n3824 ;
  assign y22483 = ~n45853 ;
  assign y22484 = n45856 ;
  assign y22485 = n45858 ;
  assign y22486 = n37994 ;
  assign y22487 = n45861 ;
  assign y22488 = ~n45862 ;
  assign y22489 = n45863 ;
  assign y22490 = n45865 ;
  assign y22491 = ~n27721 ;
  assign y22492 = ~1'b0 ;
  assign y22493 = ~n45866 ;
  assign y22494 = ~n45867 ;
  assign y22495 = ~n45868 ;
  assign y22496 = ~n45869 ;
  assign y22497 = n14204 ;
  assign y22498 = n45870 ;
  assign y22499 = ~n45874 ;
  assign y22500 = ~n45875 ;
  assign y22501 = ~1'b0 ;
  assign y22502 = n45876 ;
  assign y22503 = ~1'b0 ;
  assign y22504 = ~n45877 ;
  assign y22505 = ~n45878 ;
  assign y22506 = ~n45882 ;
  assign y22507 = n45884 ;
  assign y22508 = ~n45885 ;
  assign y22509 = n45886 ;
  assign y22510 = ~n45888 ;
  assign y22511 = ~1'b0 ;
  assign y22512 = ~n8777 ;
  assign y22513 = ~n45889 ;
  assign y22514 = ~1'b0 ;
  assign y22515 = n774 ;
  assign y22516 = n45890 ;
  assign y22517 = n45893 ;
  assign y22518 = ~1'b0 ;
  assign y22519 = n45895 ;
  assign y22520 = ~n45899 ;
  assign y22521 = ~1'b0 ;
  assign y22522 = n45901 ;
  assign y22523 = 1'b0 ;
  assign y22524 = ~n45903 ;
  assign y22525 = ~1'b0 ;
  assign y22526 = ~n45907 ;
  assign y22527 = ~1'b0 ;
  assign y22528 = n45908 ;
  assign y22529 = n45912 ;
  assign y22530 = n45913 ;
  assign y22531 = n45914 ;
  assign y22532 = ~n45918 ;
  assign y22533 = ~n45919 ;
  assign y22534 = ~n45928 ;
  assign y22535 = ~n45929 ;
  assign y22536 = ~n45933 ;
  assign y22537 = ~n45936 ;
  assign y22538 = ~n45940 ;
  assign y22539 = ~n45941 ;
  assign y22540 = ~n45942 ;
  assign y22541 = ~n45945 ;
  assign y22542 = n14145 ;
  assign y22543 = ~n45946 ;
  assign y22544 = ~1'b0 ;
  assign y22545 = ~1'b0 ;
  assign y22546 = n45947 ;
  assign y22547 = ~n45948 ;
  assign y22548 = 1'b0 ;
  assign y22549 = ~n45950 ;
  assign y22550 = ~1'b0 ;
  assign y22551 = n32108 ;
  assign y22552 = ~n45954 ;
  assign y22553 = n45957 ;
  assign y22554 = n45961 ;
  assign y22555 = n45964 ;
  assign y22556 = ~n45973 ;
  assign y22557 = ~n45978 ;
  assign y22558 = ~n45981 ;
  assign y22559 = ~n34610 ;
  assign y22560 = ~n45984 ;
  assign y22561 = ~1'b0 ;
  assign y22562 = ~n45985 ;
  assign y22563 = n45987 ;
  assign y22564 = n45995 ;
  assign y22565 = ~n45996 ;
  assign y22566 = ~n45999 ;
  assign y22567 = ~1'b0 ;
  assign y22568 = ~1'b0 ;
  assign y22569 = ~n46000 ;
  assign y22570 = ~1'b0 ;
  assign y22571 = n46001 ;
  assign y22572 = 1'b0 ;
  assign y22573 = n46002 ;
  assign y22574 = ~n46004 ;
  assign y22575 = ~n46011 ;
  assign y22576 = ~1'b0 ;
  assign y22577 = n46015 ;
  assign y22578 = n46021 ;
  assign y22579 = ~n46022 ;
  assign y22580 = ~n46028 ;
  assign y22581 = n46030 ;
  assign y22582 = ~1'b0 ;
  assign y22583 = ~1'b0 ;
  assign y22584 = ~1'b0 ;
  assign y22585 = n46032 ;
  assign y22586 = ~1'b0 ;
  assign y22587 = n46033 ;
  assign y22588 = n46037 ;
  assign y22589 = ~1'b0 ;
  assign y22590 = n46038 ;
  assign y22591 = ~n46040 ;
  assign y22592 = ~1'b0 ;
  assign y22593 = ~1'b0 ;
  assign y22594 = ~n46043 ;
  assign y22595 = n46047 ;
  assign y22596 = n46050 ;
  assign y22597 = ~n46051 ;
  assign y22598 = n46054 ;
  assign y22599 = n46056 ;
  assign y22600 = ~1'b0 ;
  assign y22601 = ~n28246 ;
  assign y22602 = ~n46060 ;
  assign y22603 = n12767 ;
  assign y22604 = n46062 ;
  assign y22605 = n46064 ;
  assign y22606 = ~n18967 ;
  assign y22607 = n10804 ;
  assign y22608 = ~1'b0 ;
  assign y22609 = ~n46068 ;
  assign y22610 = n46069 ;
  assign y22611 = ~n46070 ;
  assign y22612 = n46073 ;
  assign y22613 = n46074 ;
  assign y22614 = ~1'b0 ;
  assign y22615 = ~1'b0 ;
  assign y22616 = ~1'b0 ;
  assign y22617 = ~1'b0 ;
  assign y22618 = n46076 ;
  assign y22619 = n46078 ;
  assign y22620 = n46082 ;
  assign y22621 = ~1'b0 ;
  assign y22622 = ~1'b0 ;
  assign y22623 = ~1'b0 ;
  assign y22624 = n34491 ;
  assign y22625 = n46083 ;
  assign y22626 = ~n46086 ;
  assign y22627 = ~n46088 ;
  assign y22628 = ~n46094 ;
  assign y22629 = n5281 ;
  assign y22630 = ~1'b0 ;
  assign y22631 = ~1'b0 ;
  assign y22632 = ~n46095 ;
  assign y22633 = ~n46096 ;
  assign y22634 = n46098 ;
  assign y22635 = ~1'b0 ;
  assign y22636 = n46106 ;
  assign y22637 = ~n46110 ;
  assign y22638 = ~1'b0 ;
  assign y22639 = ~1'b0 ;
  assign y22640 = ~1'b0 ;
  assign y22641 = ~1'b0 ;
  assign y22642 = ~n46111 ;
  assign y22643 = ~1'b0 ;
  assign y22644 = n46112 ;
  assign y22645 = n46115 ;
  assign y22646 = ~n46116 ;
  assign y22647 = ~1'b0 ;
  assign y22648 = ~1'b0 ;
  assign y22649 = ~n46118 ;
  assign y22650 = ~1'b0 ;
  assign y22651 = ~1'b0 ;
  assign y22652 = ~n46119 ;
  assign y22653 = n46121 ;
  assign y22654 = ~n46122 ;
  assign y22655 = ~n46123 ;
  assign y22656 = ~1'b0 ;
  assign y22657 = ~1'b0 ;
  assign y22658 = ~n46125 ;
  assign y22659 = ~1'b0 ;
  assign y22660 = n46127 ;
  assign y22661 = n46128 ;
  assign y22662 = ~n46130 ;
  assign y22663 = n46133 ;
  assign y22664 = n46135 ;
  assign y22665 = ~1'b0 ;
  assign y22666 = n46136 ;
  assign y22667 = n46137 ;
  assign y22668 = ~n46138 ;
  assign y22669 = ~n18765 ;
  assign y22670 = ~n46142 ;
  assign y22671 = n46143 ;
  assign y22672 = ~n46144 ;
  assign y22673 = ~n46147 ;
  assign y22674 = ~n46148 ;
  assign y22675 = n46151 ;
  assign y22676 = ~1'b0 ;
  assign y22677 = ~n46159 ;
  assign y22678 = n46162 ;
  assign y22679 = n46166 ;
  assign y22680 = ~n46168 ;
  assign y22681 = ~n46171 ;
  assign y22682 = n46172 ;
  assign y22683 = ~n46174 ;
  assign y22684 = n15321 ;
  assign y22685 = ~n46176 ;
  assign y22686 = n46177 ;
  assign y22687 = ~1'b0 ;
  assign y22688 = ~n46178 ;
  assign y22689 = n46179 ;
  assign y22690 = ~n46181 ;
  assign y22691 = n46183 ;
  assign y22692 = n4706 ;
  assign y22693 = ~1'b0 ;
  assign y22694 = ~1'b0 ;
  assign y22695 = n46185 ;
  assign y22696 = ~n46201 ;
  assign y22697 = n46204 ;
  assign y22698 = ~1'b0 ;
  assign y22699 = ~1'b0 ;
  assign y22700 = ~1'b0 ;
  assign y22701 = ~n46205 ;
  assign y22702 = 1'b0 ;
  assign y22703 = n46210 ;
  assign y22704 = ~1'b0 ;
  assign y22705 = ~1'b0 ;
  assign y22706 = ~n46211 ;
  assign y22707 = n46212 ;
  assign y22708 = n46214 ;
  assign y22709 = ~n46218 ;
  assign y22710 = ~n46219 ;
  assign y22711 = n46221 ;
  assign y22712 = n46226 ;
  assign y22713 = n46227 ;
  assign y22714 = ~1'b0 ;
  assign y22715 = n46228 ;
  assign y22716 = ~n46231 ;
  assign y22717 = ~n46232 ;
  assign y22718 = ~1'b0 ;
  assign y22719 = n46234 ;
  assign y22720 = ~1'b0 ;
  assign y22721 = n46236 ;
  assign y22722 = ~n46237 ;
  assign y22723 = ~n46239 ;
  assign y22724 = n46241 ;
  assign y22725 = n46242 ;
  assign y22726 = n46246 ;
  assign y22727 = ~n46254 ;
  assign y22728 = ~1'b0 ;
  assign y22729 = ~1'b0 ;
  assign y22730 = n46256 ;
  assign y22731 = ~n46257 ;
  assign y22732 = n30251 ;
  assign y22733 = n8580 ;
  assign y22734 = ~n46259 ;
  assign y22735 = n46261 ;
  assign y22736 = ~1'b0 ;
  assign y22737 = n46264 ;
  assign y22738 = ~n46265 ;
  assign y22739 = ~n46267 ;
  assign y22740 = n46269 ;
  assign y22741 = ~n46272 ;
  assign y22742 = ~n46274 ;
  assign y22743 = ~n46276 ;
  assign y22744 = ~1'b0 ;
  assign y22745 = ~1'b0 ;
  assign y22746 = ~1'b0 ;
  assign y22747 = ~1'b0 ;
  assign y22748 = ~1'b0 ;
  assign y22749 = ~n46284 ;
  assign y22750 = ~n3187 ;
  assign y22751 = n46285 ;
  assign y22752 = ~1'b0 ;
  assign y22753 = ~n46287 ;
  assign y22754 = ~n46291 ;
  assign y22755 = n46292 ;
  assign y22756 = ~1'b0 ;
  assign y22757 = n46297 ;
  assign y22758 = n46299 ;
  assign y22759 = ~n46301 ;
  assign y22760 = ~n46304 ;
  assign y22761 = n8789 ;
  assign y22762 = ~n32919 ;
  assign y22763 = ~1'b0 ;
  assign y22764 = ~1'b0 ;
  assign y22765 = ~1'b0 ;
  assign y22766 = ~n46306 ;
  assign y22767 = ~n46313 ;
  assign y22768 = ~n46315 ;
  assign y22769 = n46321 ;
  assign y22770 = ~n46323 ;
  assign y22771 = ~n46329 ;
  assign y22772 = n46330 ;
  assign y22773 = ~1'b0 ;
  assign y22774 = n46331 ;
  assign y22775 = ~n46340 ;
  assign y22776 = n46343 ;
  assign y22777 = ~1'b0 ;
  assign y22778 = n46344 ;
  assign y22779 = n46350 ;
  assign y22780 = ~1'b0 ;
  assign y22781 = n27001 ;
  assign y22782 = n46352 ;
  assign y22783 = ~n46354 ;
  assign y22784 = n46356 ;
  assign y22785 = ~n46359 ;
  assign y22786 = n46365 ;
  assign y22787 = 1'b0 ;
  assign y22788 = n46366 ;
  assign y22789 = n46368 ;
  assign y22790 = ~n46370 ;
  assign y22791 = n46371 ;
  assign y22792 = n46378 ;
  assign y22793 = n46381 ;
  assign y22794 = ~n29982 ;
  assign y22795 = n46382 ;
  assign y22796 = ~1'b0 ;
  assign y22797 = ~n24951 ;
  assign y22798 = ~n46385 ;
  assign y22799 = ~n46387 ;
  assign y22800 = n27890 ;
  assign y22801 = n46390 ;
  assign y22802 = n30967 ;
  assign y22803 = n46391 ;
  assign y22804 = ~n46396 ;
  assign y22805 = ~n46397 ;
  assign y22806 = ~1'b0 ;
  assign y22807 = ~n46399 ;
  assign y22808 = n24446 ;
  assign y22809 = ~1'b0 ;
  assign y22810 = n46401 ;
  assign y22811 = n46406 ;
  assign y22812 = n46411 ;
  assign y22813 = ~n24408 ;
  assign y22814 = ~n27221 ;
  assign y22815 = ~n46413 ;
  assign y22816 = ~1'b0 ;
  assign y22817 = ~n46415 ;
  assign y22818 = n46416 ;
  assign y22819 = n46417 ;
  assign y22820 = ~n46420 ;
  assign y22821 = n46426 ;
  assign y22822 = ~1'b0 ;
  assign y22823 = ~n46428 ;
  assign y22824 = n46430 ;
  assign y22825 = ~1'b0 ;
  assign y22826 = ~n46435 ;
  assign y22827 = ~n46440 ;
  assign y22828 = n46443 ;
  assign y22829 = n46445 ;
  assign y22830 = ~n46447 ;
  assign y22831 = n46450 ;
  assign y22832 = ~n46453 ;
  assign y22833 = n46455 ;
  assign y22834 = ~n46458 ;
  assign y22835 = n2108 ;
  assign y22836 = ~1'b0 ;
  assign y22837 = ~1'b0 ;
  assign y22838 = ~n12715 ;
  assign y22839 = ~n46461 ;
  assign y22840 = ~n46465 ;
  assign y22841 = ~n46466 ;
  assign y22842 = n46468 ;
  assign y22843 = ~n46471 ;
  assign y22844 = n3614 ;
  assign y22845 = ~1'b0 ;
  assign y22846 = ~1'b0 ;
  assign y22847 = n46472 ;
  assign y22848 = ~n46473 ;
  assign y22849 = n46477 ;
  assign y22850 = n46478 ;
  assign y22851 = ~1'b0 ;
  assign y22852 = n46479 ;
  assign y22853 = n2674 ;
  assign y22854 = ~n46481 ;
  assign y22855 = n46483 ;
  assign y22856 = ~n46487 ;
  assign y22857 = n46490 ;
  assign y22858 = ~n46496 ;
  assign y22859 = 1'b0 ;
  assign y22860 = n46499 ;
  assign y22861 = ~n46500 ;
  assign y22862 = ~1'b0 ;
  assign y22863 = ~1'b0 ;
  assign y22864 = ~1'b0 ;
  assign y22865 = ~1'b0 ;
  assign y22866 = ~n46501 ;
  assign y22867 = ~n46506 ;
  assign y22868 = ~n46509 ;
  assign y22869 = ~1'b0 ;
  assign y22870 = ~n46513 ;
  assign y22871 = ~1'b0 ;
  assign y22872 = n30189 ;
  assign y22873 = ~1'b0 ;
  assign y22874 = n46515 ;
  assign y22875 = ~n46519 ;
  assign y22876 = n46520 ;
  assign y22877 = ~1'b0 ;
  assign y22878 = ~n46521 ;
  assign y22879 = ~1'b0 ;
  assign y22880 = n22900 ;
  assign y22881 = ~1'b0 ;
  assign y22882 = ~1'b0 ;
  assign y22883 = ~n46522 ;
  assign y22884 = ~n46525 ;
  assign y22885 = ~1'b0 ;
  assign y22886 = ~n46529 ;
  assign y22887 = ~n46530 ;
  assign y22888 = ~1'b0 ;
  assign y22889 = n46533 ;
  assign y22890 = ~n46539 ;
  assign y22891 = ~1'b0 ;
  assign y22892 = ~n46541 ;
  assign y22893 = n46542 ;
  assign y22894 = ~1'b0 ;
  assign y22895 = ~n46544 ;
  assign y22896 = n46550 ;
  assign y22897 = ~1'b0 ;
  assign y22898 = ~1'b0 ;
  assign y22899 = ~1'b0 ;
  assign y22900 = n46555 ;
  assign y22901 = ~n46556 ;
  assign y22902 = ~n46558 ;
  assign y22903 = ~n46560 ;
  assign y22904 = ~1'b0 ;
  assign y22905 = ~n46563 ;
  assign y22906 = ~n46569 ;
  assign y22907 = ~1'b0 ;
  assign y22908 = ~n46571 ;
  assign y22909 = ~n46573 ;
  assign y22910 = n46574 ;
  assign y22911 = n46575 ;
  assign y22912 = n46576 ;
  assign y22913 = n46579 ;
  assign y22914 = n46580 ;
  assign y22915 = ~1'b0 ;
  assign y22916 = n46583 ;
  assign y22917 = n46586 ;
  assign y22918 = ~n46595 ;
  assign y22919 = n46600 ;
  assign y22920 = ~1'b0 ;
  assign y22921 = n46602 ;
  assign y22922 = n46606 ;
  assign y22923 = 1'b0 ;
  assign y22924 = n46608 ;
  assign y22925 = ~n41681 ;
  assign y22926 = ~n46611 ;
  assign y22927 = ~1'b0 ;
  assign y22928 = ~n46612 ;
  assign y22929 = n46614 ;
  assign y22930 = ~1'b0 ;
  assign y22931 = ~1'b0 ;
  assign y22932 = 1'b0 ;
  assign y22933 = ~n46615 ;
  assign y22934 = ~n46617 ;
  assign y22935 = n46618 ;
  assign y22936 = ~1'b0 ;
  assign y22937 = n46620 ;
  assign y22938 = ~1'b0 ;
  assign y22939 = n46621 ;
  assign y22940 = ~n46629 ;
  assign y22941 = ~n46637 ;
  assign y22942 = ~n46639 ;
  assign y22943 = n46640 ;
  assign y22944 = n46642 ;
  assign y22945 = ~n46645 ;
  assign y22946 = ~n46648 ;
  assign y22947 = ~1'b0 ;
  assign y22948 = ~1'b0 ;
  assign y22949 = ~n46650 ;
  assign y22950 = ~n46652 ;
  assign y22951 = n46653 ;
  assign y22952 = ~n46654 ;
  assign y22953 = ~n46657 ;
  assign y22954 = ~n46659 ;
  assign y22955 = ~n46662 ;
  assign y22956 = n46666 ;
  assign y22957 = ~n46667 ;
  assign y22958 = n46669 ;
  assign y22959 = n46672 ;
  assign y22960 = ~n46674 ;
  assign y22961 = n46679 ;
  assign y22962 = ~n46680 ;
  assign y22963 = n46682 ;
  assign y22964 = n46685 ;
  assign y22965 = 1'b0 ;
  assign y22966 = n46687 ;
  assign y22967 = ~n46689 ;
  assign y22968 = ~n46690 ;
  assign y22969 = ~n46697 ;
  assign y22970 = n26253 ;
  assign y22971 = n46698 ;
  assign y22972 = ~n46699 ;
  assign y22973 = n46701 ;
  assign y22974 = ~n6433 ;
  assign y22975 = ~1'b0 ;
  assign y22976 = ~n46703 ;
  assign y22977 = ~n46707 ;
  assign y22978 = ~1'b0 ;
  assign y22979 = ~n4328 ;
  assign y22980 = n46710 ;
  assign y22981 = 1'b0 ;
  assign y22982 = n46712 ;
  assign y22983 = ~n46715 ;
  assign y22984 = 1'b0 ;
  assign y22985 = ~1'b0 ;
  assign y22986 = n46716 ;
  assign y22987 = n46720 ;
  assign y22988 = ~1'b0 ;
  assign y22989 = ~n46722 ;
  assign y22990 = n46726 ;
  assign y22991 = ~1'b0 ;
  assign y22992 = n46728 ;
  assign y22993 = ~n46729 ;
  assign y22994 = n46733 ;
  assign y22995 = n46735 ;
  assign y22996 = ~1'b0 ;
  assign y22997 = ~1'b0 ;
  assign y22998 = n46736 ;
  assign y22999 = ~n46741 ;
  assign y23000 = n46742 ;
  assign y23001 = n46744 ;
  assign y23002 = n30662 ;
  assign y23003 = n46749 ;
  assign y23004 = ~n46750 ;
  assign y23005 = ~n46752 ;
  assign y23006 = ~1'b0 ;
  assign y23007 = ~1'b0 ;
  assign y23008 = ~n46754 ;
  assign y23009 = n46758 ;
  assign y23010 = n46760 ;
  assign y23011 = ~n46762 ;
  assign y23012 = ~n46764 ;
  assign y23013 = n46767 ;
  assign y23014 = n46771 ;
  assign y23015 = n18469 ;
  assign y23016 = ~n46773 ;
  assign y23017 = ~n46775 ;
  assign y23018 = ~n46776 ;
  assign y23019 = ~n46777 ;
  assign y23020 = ~1'b0 ;
  assign y23021 = ~1'b0 ;
  assign y23022 = n46778 ;
  assign y23023 = ~1'b0 ;
  assign y23024 = ~1'b0 ;
  assign y23025 = ~n46780 ;
  assign y23026 = n46782 ;
  assign y23027 = ~n46783 ;
  assign y23028 = n46784 ;
  assign y23029 = ~n46788 ;
  assign y23030 = ~n38027 ;
  assign y23031 = n46790 ;
  assign y23032 = n46791 ;
  assign y23033 = n46793 ;
  assign y23034 = ~1'b0 ;
  assign y23035 = ~n46794 ;
  assign y23036 = n46798 ;
  assign y23037 = n46801 ;
  assign y23038 = n46802 ;
  assign y23039 = ~n46803 ;
  assign y23040 = ~1'b0 ;
  assign y23041 = ~n46804 ;
  assign y23042 = ~1'b0 ;
  assign y23043 = ~1'b0 ;
  assign y23044 = n46805 ;
  assign y23045 = ~1'b0 ;
  assign y23046 = n46809 ;
  assign y23047 = ~n46810 ;
  assign y23048 = ~1'b0 ;
  assign y23049 = n46816 ;
  assign y23050 = ~1'b0 ;
  assign y23051 = ~1'b0 ;
  assign y23052 = n46817 ;
  assign y23053 = n46819 ;
  assign y23054 = ~1'b0 ;
  assign y23055 = n46820 ;
  assign y23056 = n36998 ;
  assign y23057 = ~n46821 ;
  assign y23058 = n46822 ;
  assign y23059 = n46826 ;
  assign y23060 = n46829 ;
  assign y23061 = ~n46830 ;
  assign y23062 = ~1'b0 ;
  assign y23063 = ~1'b0 ;
  assign y23064 = ~1'b0 ;
  assign y23065 = ~1'b0 ;
  assign y23066 = ~1'b0 ;
  assign y23067 = n46833 ;
  assign y23068 = n46834 ;
  assign y23069 = ~n46838 ;
  assign y23070 = ~n46839 ;
  assign y23071 = n46841 ;
  assign y23072 = 1'b0 ;
  assign y23073 = ~n46845 ;
  assign y23074 = n46846 ;
  assign y23075 = ~n46847 ;
  assign y23076 = ~n46848 ;
  assign y23077 = ~n46849 ;
  assign y23078 = n46852 ;
  assign y23079 = n46853 ;
  assign y23080 = ~1'b0 ;
  assign y23081 = n46857 ;
  assign y23082 = n46858 ;
  assign y23083 = ~n46863 ;
  assign y23084 = n46864 ;
  assign y23085 = ~n19761 ;
  assign y23086 = n46865 ;
  assign y23087 = ~1'b0 ;
  assign y23088 = ~1'b0 ;
  assign y23089 = ~1'b0 ;
  assign y23090 = 1'b0 ;
  assign y23091 = ~n46875 ;
  assign y23092 = ~n46880 ;
  assign y23093 = ~n46885 ;
  assign y23094 = ~n46887 ;
  assign y23095 = ~n46889 ;
  assign y23096 = ~1'b0 ;
  assign y23097 = ~1'b0 ;
  assign y23098 = n46897 ;
  assign y23099 = ~1'b0 ;
  assign y23100 = ~1'b0 ;
  assign y23101 = n46898 ;
  assign y23102 = n31823 ;
  assign y23103 = ~1'b0 ;
  assign y23104 = n46902 ;
  assign y23105 = ~1'b0 ;
  assign y23106 = n46904 ;
  assign y23107 = ~n46913 ;
  assign y23108 = ~n46915 ;
  assign y23109 = n46917 ;
  assign y23110 = n46918 ;
  assign y23111 = ~n46921 ;
  assign y23112 = n46924 ;
  assign y23113 = n41188 ;
  assign y23114 = ~n46926 ;
  assign y23115 = n46930 ;
  assign y23116 = ~1'b0 ;
  assign y23117 = n46931 ;
  assign y23118 = ~n46933 ;
  assign y23119 = n46934 ;
  assign y23120 = ~n46935 ;
  assign y23121 = n46941 ;
  assign y23122 = ~1'b0 ;
  assign y23123 = ~1'b0 ;
  assign y23124 = ~1'b0 ;
  assign y23125 = n35081 ;
  assign y23126 = n46942 ;
  assign y23127 = n46944 ;
  assign y23128 = ~n45330 ;
  assign y23129 = n46946 ;
  assign y23130 = ~n46952 ;
  assign y23131 = n46953 ;
  assign y23132 = ~n21610 ;
  assign y23133 = ~n46955 ;
  assign y23134 = ~1'b0 ;
  assign y23135 = n46956 ;
  assign y23136 = ~n46957 ;
  assign y23137 = ~1'b0 ;
  assign y23138 = ~1'b0 ;
  assign y23139 = ~1'b0 ;
  assign y23140 = ~n46960 ;
  assign y23141 = n46961 ;
  assign y23142 = ~n46962 ;
  assign y23143 = ~n46966 ;
  assign y23144 = n46969 ;
  assign y23145 = n46978 ;
  assign y23146 = ~1'b0 ;
  assign y23147 = ~1'b0 ;
  assign y23148 = n46980 ;
  assign y23149 = ~n46981 ;
  assign y23150 = ~1'b0 ;
  assign y23151 = n46984 ;
  assign y23152 = ~n46985 ;
  assign y23153 = n46988 ;
  assign y23154 = ~n46989 ;
  assign y23155 = ~1'b0 ;
  assign y23156 = ~n46990 ;
  assign y23157 = ~1'b0 ;
  assign y23158 = ~1'b0 ;
  assign y23159 = n9070 ;
  assign y23160 = ~1'b0 ;
  assign y23161 = ~n21495 ;
  assign y23162 = n46991 ;
  assign y23163 = n46994 ;
  assign y23164 = n46995 ;
  assign y23165 = ~n46997 ;
  assign y23166 = n46998 ;
  assign y23167 = ~n46999 ;
  assign y23168 = n47002 ;
  assign y23169 = ~1'b0 ;
  assign y23170 = ~n47005 ;
  assign y23171 = ~1'b0 ;
  assign y23172 = n47006 ;
  assign y23173 = n26668 ;
  assign y23174 = n47008 ;
  assign y23175 = ~1'b0 ;
  assign y23176 = n47009 ;
  assign y23177 = ~n47012 ;
  assign y23178 = n47013 ;
  assign y23179 = ~n47014 ;
  assign y23180 = n47016 ;
  assign y23181 = ~n47020 ;
  assign y23182 = n47023 ;
  assign y23183 = n47024 ;
  assign y23184 = ~n47030 ;
  assign y23185 = ~n47032 ;
  assign y23186 = n47035 ;
  assign y23187 = ~n47040 ;
  assign y23188 = ~1'b0 ;
  assign y23189 = ~n47043 ;
  assign y23190 = ~n23793 ;
  assign y23191 = ~n47045 ;
  assign y23192 = ~n47046 ;
  assign y23193 = n47047 ;
  assign y23194 = ~1'b0 ;
  assign y23195 = ~n47051 ;
  assign y23196 = n47055 ;
  assign y23197 = n47056 ;
  assign y23198 = n13876 ;
  assign y23199 = ~n32532 ;
  assign y23200 = ~n21839 ;
  assign y23201 = ~n47058 ;
  assign y23202 = ~n47061 ;
  assign y23203 = n47067 ;
  assign y23204 = ~n47074 ;
  assign y23205 = ~n47076 ;
  assign y23206 = n47077 ;
  assign y23207 = n47078 ;
  assign y23208 = n47079 ;
  assign y23209 = ~n47081 ;
  assign y23210 = ~1'b0 ;
  assign y23211 = n47082 ;
  assign y23212 = ~n47084 ;
  assign y23213 = ~1'b0 ;
  assign y23214 = n47085 ;
  assign y23215 = n47086 ;
  assign y23216 = ~n47087 ;
  assign y23217 = ~n47090 ;
  assign y23218 = ~1'b0 ;
  assign y23219 = ~1'b0 ;
  assign y23220 = n47093 ;
  assign y23221 = n47096 ;
  assign y23222 = ~n26910 ;
  assign y23223 = ~n47097 ;
  assign y23224 = ~n47099 ;
  assign y23225 = n47103 ;
  assign y23226 = ~1'b0 ;
  assign y23227 = ~1'b0 ;
  assign y23228 = ~n34008 ;
  assign y23229 = 1'b0 ;
  assign y23230 = ~1'b0 ;
  assign y23231 = n47104 ;
  assign y23232 = n47105 ;
  assign y23233 = ~1'b0 ;
  assign y23234 = ~1'b0 ;
  assign y23235 = ~n47110 ;
  assign y23236 = ~n47111 ;
  assign y23237 = ~1'b0 ;
  assign y23238 = n47112 ;
  assign y23239 = ~n47115 ;
  assign y23240 = ~1'b0 ;
  assign y23241 = n47117 ;
  assign y23242 = ~n47120 ;
  assign y23243 = ~1'b0 ;
  assign y23244 = ~n47123 ;
  assign y23245 = ~n22661 ;
  assign y23246 = n47128 ;
  assign y23247 = ~n47129 ;
  assign y23248 = ~1'b0 ;
  assign y23249 = n47130 ;
  assign y23250 = ~1'b0 ;
  assign y23251 = ~n47133 ;
  assign y23252 = n47135 ;
  assign y23253 = n47136 ;
  assign y23254 = ~1'b0 ;
  assign y23255 = n47139 ;
  assign y23256 = ~n47141 ;
  assign y23257 = n47142 ;
  assign y23258 = ~1'b0 ;
  assign y23259 = ~1'b0 ;
  assign y23260 = ~1'b0 ;
  assign y23261 = n47143 ;
  assign y23262 = ~1'b0 ;
  assign y23263 = n47144 ;
  assign y23264 = n47145 ;
  assign y23265 = ~1'b0 ;
  assign y23266 = ~n47149 ;
  assign y23267 = ~n47151 ;
  assign y23268 = ~1'b0 ;
  assign y23269 = ~1'b0 ;
  assign y23270 = ~n43084 ;
  assign y23271 = ~1'b0 ;
  assign y23272 = ~1'b0 ;
  assign y23273 = ~n47153 ;
  assign y23274 = ~n47156 ;
  assign y23275 = n47163 ;
  assign y23276 = n47168 ;
  assign y23277 = 1'b0 ;
  assign y23278 = n47170 ;
  assign y23279 = n47173 ;
  assign y23280 = ~1'b0 ;
  assign y23281 = 1'b0 ;
  assign y23282 = n47175 ;
  assign y23283 = ~1'b0 ;
  assign y23284 = n47176 ;
  assign y23285 = n47181 ;
  assign y23286 = n47184 ;
  assign y23287 = n6681 ;
  assign y23288 = ~n47189 ;
  assign y23289 = ~n47192 ;
  assign y23290 = n47195 ;
  assign y23291 = ~1'b0 ;
  assign y23292 = n47196 ;
  assign y23293 = n47199 ;
  assign y23294 = 1'b0 ;
  assign y23295 = ~1'b0 ;
  assign y23296 = ~1'b0 ;
  assign y23297 = ~n47201 ;
  assign y23298 = n47204 ;
  assign y23299 = n47207 ;
  assign y23300 = n47209 ;
  assign y23301 = n47212 ;
  assign y23302 = n6437 ;
  assign y23303 = n47214 ;
  assign y23304 = n47216 ;
  assign y23305 = ~1'b0 ;
  assign y23306 = ~1'b0 ;
  assign y23307 = n47217 ;
  assign y23308 = n47222 ;
  assign y23309 = ~n47223 ;
  assign y23310 = 1'b0 ;
  assign y23311 = ~1'b0 ;
  assign y23312 = ~1'b0 ;
  assign y23313 = n47225 ;
  assign y23314 = ~1'b0 ;
  assign y23315 = ~1'b0 ;
  assign y23316 = ~n47227 ;
  assign y23317 = n47228 ;
  assign y23318 = ~1'b0 ;
  assign y23319 = ~n47230 ;
  assign y23320 = ~n47233 ;
  assign y23321 = ~n47237 ;
  assign y23322 = ~n47239 ;
  assign y23323 = n47240 ;
  assign y23324 = n47246 ;
  assign y23325 = n47253 ;
  assign y23326 = ~1'b0 ;
  assign y23327 = n47258 ;
  assign y23328 = ~n47259 ;
  assign y23329 = ~n47263 ;
  assign y23330 = ~n47264 ;
  assign y23331 = ~n47270 ;
  assign y23332 = n47275 ;
  assign y23333 = n47277 ;
  assign y23334 = n47281 ;
  assign y23335 = ~n7192 ;
  assign y23336 = ~n47283 ;
  assign y23337 = n47285 ;
  assign y23338 = ~n47287 ;
  assign y23339 = n47288 ;
  assign y23340 = ~1'b0 ;
  assign y23341 = ~n47290 ;
  assign y23342 = ~1'b0 ;
  assign y23343 = n47292 ;
  assign y23344 = ~n47297 ;
  assign y23345 = ~n47299 ;
  assign y23346 = ~n47302 ;
  assign y23347 = ~n47303 ;
  assign y23348 = ~n47305 ;
  assign y23349 = ~n36627 ;
  assign y23350 = ~1'b0 ;
  assign y23351 = ~n47309 ;
  assign y23352 = ~1'b0 ;
  assign y23353 = ~1'b0 ;
  assign y23354 = ~n47310 ;
  assign y23355 = ~n47311 ;
  assign y23356 = n47319 ;
  assign y23357 = ~1'b0 ;
  assign y23358 = ~n47321 ;
  assign y23359 = ~1'b0 ;
  assign y23360 = n47322 ;
  assign y23361 = ~n47324 ;
  assign y23362 = ~1'b0 ;
  assign y23363 = ~1'b0 ;
  assign y23364 = ~1'b0 ;
  assign y23365 = ~n47331 ;
  assign y23366 = ~1'b0 ;
  assign y23367 = ~n47334 ;
  assign y23368 = n47336 ;
  assign y23369 = ~n47340 ;
  assign y23370 = ~1'b0 ;
  assign y23371 = ~1'b0 ;
  assign y23372 = ~n47341 ;
  assign y23373 = ~n47344 ;
  assign y23374 = ~n7908 ;
  assign y23375 = n47345 ;
  assign y23376 = ~n47346 ;
  assign y23377 = ~1'b0 ;
  assign y23378 = n47351 ;
  assign y23379 = ~1'b0 ;
  assign y23380 = ~n31183 ;
  assign y23381 = n47354 ;
  assign y23382 = ~n47356 ;
  assign y23383 = n47357 ;
  assign y23384 = ~n47358 ;
  assign y23385 = ~n47360 ;
  assign y23386 = ~n47362 ;
  assign y23387 = ~n47364 ;
  assign y23388 = ~n47367 ;
  assign y23389 = ~1'b0 ;
  assign y23390 = ~1'b0 ;
  assign y23391 = ~1'b0 ;
  assign y23392 = ~n47372 ;
  assign y23393 = n47374 ;
  assign y23394 = n47375 ;
  assign y23395 = n47376 ;
  assign y23396 = n47384 ;
  assign y23397 = ~n47386 ;
  assign y23398 = ~n47388 ;
  assign y23399 = ~n47393 ;
  assign y23400 = n47394 ;
  assign y23401 = ~1'b0 ;
  assign y23402 = ~1'b0 ;
  assign y23403 = n47398 ;
  assign y23404 = n47399 ;
  assign y23405 = ~n47408 ;
  assign y23406 = ~n47409 ;
  assign y23407 = ~n47410 ;
  assign y23408 = ~n47411 ;
  assign y23409 = n47412 ;
  assign y23410 = ~1'b0 ;
  assign y23411 = n47415 ;
  assign y23412 = ~n732 ;
  assign y23413 = n22218 ;
  assign y23414 = n47417 ;
  assign y23415 = n47419 ;
  assign y23416 = ~1'b0 ;
  assign y23417 = n47421 ;
  assign y23418 = ~1'b0 ;
  assign y23419 = ~n47425 ;
  assign y23420 = ~n47429 ;
  assign y23421 = ~1'b0 ;
  assign y23422 = n28090 ;
  assign y23423 = n47432 ;
  assign y23424 = ~n47435 ;
  assign y23425 = n47436 ;
  assign y23426 = ~1'b0 ;
  assign y23427 = ~n26047 ;
  assign y23428 = ~1'b0 ;
  assign y23429 = ~n47438 ;
  assign y23430 = ~n47442 ;
  assign y23431 = n47445 ;
  assign y23432 = ~1'b0 ;
  assign y23433 = n47447 ;
  assign y23434 = ~1'b0 ;
  assign y23435 = n47449 ;
  assign y23436 = n47453 ;
  assign y23437 = ~1'b0 ;
  assign y23438 = ~n47455 ;
  assign y23439 = ~n47456 ;
  assign y23440 = n47458 ;
  assign y23441 = n47459 ;
  assign y23442 = ~1'b0 ;
  assign y23443 = ~n47460 ;
  assign y23444 = n25773 ;
  assign y23445 = ~n47463 ;
  assign y23446 = ~1'b0 ;
  assign y23447 = n47467 ;
  assign y23448 = ~n47471 ;
  assign y23449 = ~n47475 ;
  assign y23450 = n17893 ;
  assign y23451 = n47476 ;
  assign y23452 = n47478 ;
  assign y23453 = n47480 ;
  assign y23454 = ~n47483 ;
  assign y23455 = ~1'b0 ;
  assign y23456 = ~1'b0 ;
  assign y23457 = ~1'b0 ;
  assign y23458 = ~n47485 ;
  assign y23459 = n47492 ;
  assign y23460 = ~n47494 ;
  assign y23461 = n47496 ;
  assign y23462 = ~n2120 ;
  assign y23463 = ~n47500 ;
  assign y23464 = ~1'b0 ;
  assign y23465 = ~n47504 ;
  assign y23466 = ~1'b0 ;
  assign y23467 = n47506 ;
  assign y23468 = n47509 ;
  assign y23469 = n47510 ;
  assign y23470 = ~1'b0 ;
  assign y23471 = n47512 ;
  assign y23472 = ~n47514 ;
  assign y23473 = ~n47516 ;
  assign y23474 = n47517 ;
  assign y23475 = ~n47518 ;
  assign y23476 = ~n47521 ;
  assign y23477 = n47522 ;
  assign y23478 = ~n47524 ;
  assign y23479 = ~n47525 ;
  assign y23480 = ~1'b0 ;
  assign y23481 = ~n47528 ;
  assign y23482 = ~n47529 ;
  assign y23483 = n47530 ;
  assign y23484 = ~n36171 ;
  assign y23485 = n10374 ;
  assign y23486 = ~1'b0 ;
  assign y23487 = ~1'b0 ;
  assign y23488 = ~1'b0 ;
  assign y23489 = n47532 ;
  assign y23490 = ~n47533 ;
  assign y23491 = 1'b0 ;
  assign y23492 = n11912 ;
  assign y23493 = ~n47535 ;
  assign y23494 = n6790 ;
  assign y23495 = ~1'b0 ;
  assign y23496 = ~1'b0 ;
  assign y23497 = n47540 ;
  assign y23498 = ~1'b0 ;
  assign y23499 = ~n47541 ;
  assign y23500 = ~1'b0 ;
  assign y23501 = ~1'b0 ;
  assign y23502 = ~n47542 ;
  assign y23503 = n47545 ;
  assign y23504 = ~n47549 ;
  assign y23505 = ~n47551 ;
  assign y23506 = ~n47554 ;
  assign y23507 = ~1'b0 ;
  assign y23508 = ~n47557 ;
  assign y23509 = n47558 ;
  assign y23510 = n47560 ;
  assign y23511 = n10784 ;
  assign y23512 = n47562 ;
  assign y23513 = n47563 ;
  assign y23514 = n47565 ;
  assign y23515 = n47566 ;
  assign y23516 = ~1'b0 ;
  assign y23517 = n47568 ;
  assign y23518 = 1'b0 ;
  assign y23519 = ~n47569 ;
  assign y23520 = ~n47571 ;
  assign y23521 = n1320 ;
  assign y23522 = n47573 ;
  assign y23523 = ~n47574 ;
  assign y23524 = ~n47576 ;
  assign y23525 = n47578 ;
  assign y23526 = n47580 ;
  assign y23527 = n5262 ;
  assign y23528 = n119 ;
  assign y23529 = ~n47584 ;
  assign y23530 = ~n47586 ;
  assign y23531 = ~n47587 ;
  assign y23532 = ~n47588 ;
  assign y23533 = n47590 ;
  assign y23534 = ~1'b0 ;
  assign y23535 = n47595 ;
  assign y23536 = ~1'b0 ;
  assign y23537 = n47598 ;
  assign y23538 = ~n47601 ;
  assign y23539 = ~n47602 ;
  assign y23540 = n47603 ;
  assign y23541 = n16233 ;
  assign y23542 = n47605 ;
  assign y23543 = ~1'b0 ;
  assign y23544 = ~1'b0 ;
  assign y23545 = n24938 ;
  assign y23546 = ~1'b0 ;
  assign y23547 = ~n47607 ;
  assign y23548 = ~n47609 ;
  assign y23549 = ~n47613 ;
  assign y23550 = ~n47614 ;
  assign y23551 = n47615 ;
  assign y23552 = ~1'b0 ;
  assign y23553 = n47618 ;
  assign y23554 = n47621 ;
  assign y23555 = ~n47623 ;
  assign y23556 = ~n47627 ;
  assign y23557 = ~n47630 ;
  assign y23558 = n47631 ;
  assign y23559 = ~n18727 ;
  assign y23560 = n47633 ;
  assign y23561 = ~n47636 ;
  assign y23562 = ~1'b0 ;
  assign y23563 = ~n47637 ;
  assign y23564 = ~1'b0 ;
  assign y23565 = n47638 ;
  assign y23566 = n47642 ;
  assign y23567 = n47643 ;
  assign y23568 = ~n47644 ;
  assign y23569 = ~n47645 ;
  assign y23570 = ~n41499 ;
  assign y23571 = ~1'b0 ;
  assign y23572 = 1'b0 ;
  assign y23573 = ~n47648 ;
  assign y23574 = ~1'b0 ;
  assign y23575 = n47652 ;
  assign y23576 = ~n47653 ;
  assign y23577 = n47657 ;
  assign y23578 = ~n47661 ;
  assign y23579 = ~1'b0 ;
  assign y23580 = ~n47664 ;
  assign y23581 = n47666 ;
  assign y23582 = n47671 ;
  assign y23583 = ~1'b0 ;
  assign y23584 = ~1'b0 ;
  assign y23585 = ~1'b0 ;
  assign y23586 = n47673 ;
  assign y23587 = ~n47674 ;
  assign y23588 = n47675 ;
  assign y23589 = n47676 ;
  assign y23590 = 1'b0 ;
  assign y23591 = ~n47680 ;
  assign y23592 = ~n47683 ;
  assign y23593 = ~n47687 ;
  assign y23594 = ~n47693 ;
  assign y23595 = ~1'b0 ;
  assign y23596 = n47695 ;
  assign y23597 = ~n47698 ;
  assign y23598 = n47699 ;
  assign y23599 = n47702 ;
  assign y23600 = ~n11199 ;
  assign y23601 = ~n47706 ;
  assign y23602 = n47707 ;
  assign y23603 = ~n47709 ;
  assign y23604 = ~1'b0 ;
  assign y23605 = n47711 ;
  assign y23606 = n40115 ;
  assign y23607 = ~n47712 ;
  assign y23608 = n47713 ;
  assign y23609 = n47714 ;
  assign y23610 = ~1'b0 ;
  assign y23611 = n47717 ;
  assign y23612 = ~1'b0 ;
  assign y23613 = n47718 ;
  assign y23614 = n47719 ;
  assign y23615 = ~1'b0 ;
  assign y23616 = ~n47720 ;
  assign y23617 = n47721 ;
  assign y23618 = n47723 ;
  assign y23619 = 1'b0 ;
  assign y23620 = 1'b0 ;
  assign y23621 = ~1'b0 ;
  assign y23622 = ~1'b0 ;
  assign y23623 = n47725 ;
  assign y23624 = ~n47728 ;
  assign y23625 = ~n47731 ;
  assign y23626 = n47737 ;
  assign y23627 = ~1'b0 ;
  assign y23628 = ~1'b0 ;
  assign y23629 = ~n11783 ;
  assign y23630 = ~n47740 ;
  assign y23631 = n47743 ;
  assign y23632 = n47746 ;
  assign y23633 = ~n47748 ;
  assign y23634 = ~n47753 ;
  assign y23635 = n47756 ;
  assign y23636 = ~1'b0 ;
  assign y23637 = ~1'b0 ;
  assign y23638 = ~n47759 ;
  assign y23639 = n47768 ;
  assign y23640 = ~n47772 ;
  assign y23641 = n47774 ;
  assign y23642 = n47775 ;
  assign y23643 = ~n47778 ;
  assign y23644 = ~1'b0 ;
  assign y23645 = ~n47779 ;
  assign y23646 = ~1'b0 ;
  assign y23647 = n47782 ;
  assign y23648 = ~n47783 ;
  assign y23649 = n47784 ;
  assign y23650 = ~1'b0 ;
  assign y23651 = ~n47786 ;
  assign y23652 = ~n47789 ;
  assign y23653 = ~1'b0 ;
  assign y23654 = ~n47791 ;
  assign y23655 = n47792 ;
  assign y23656 = ~1'b0 ;
  assign y23657 = ~n47794 ;
  assign y23658 = n47795 ;
  assign y23659 = ~n47798 ;
  assign y23660 = n47805 ;
  assign y23661 = n47807 ;
  assign y23662 = ~1'b0 ;
  assign y23663 = n4769 ;
  assign y23664 = ~1'b0 ;
  assign y23665 = ~1'b0 ;
  assign y23666 = ~1'b0 ;
  assign y23667 = ~n47812 ;
  assign y23668 = ~n47815 ;
  assign y23669 = ~n47816 ;
  assign y23670 = n47821 ;
  assign y23671 = n47830 ;
  assign y23672 = n47832 ;
  assign y23673 = n47834 ;
  assign y23674 = ~n47836 ;
  assign y23675 = ~n47837 ;
  assign y23676 = ~n9275 ;
  assign y23677 = n47838 ;
  assign y23678 = ~n47842 ;
  assign y23679 = ~1'b0 ;
  assign y23680 = n47844 ;
  assign y23681 = ~1'b0 ;
  assign y23682 = n47848 ;
  assign y23683 = ~n47850 ;
  assign y23684 = n47854 ;
  assign y23685 = ~n47855 ;
  assign y23686 = ~n15336 ;
  assign y23687 = ~n47857 ;
  assign y23688 = ~1'b0 ;
  assign y23689 = ~n47860 ;
  assign y23690 = ~n47862 ;
  assign y23691 = n47865 ;
  assign y23692 = n26872 ;
  assign y23693 = ~n47867 ;
  assign y23694 = ~n47868 ;
  assign y23695 = n47870 ;
  assign y23696 = ~n47873 ;
  assign y23697 = ~1'b0 ;
  assign y23698 = n47874 ;
  assign y23699 = n23447 ;
  assign y23700 = ~n47878 ;
  assign y23701 = ~1'b0 ;
  assign y23702 = ~n47882 ;
  assign y23703 = ~1'b0 ;
  assign y23704 = ~n47883 ;
  assign y23705 = ~n47884 ;
  assign y23706 = ~n47885 ;
  assign y23707 = ~1'b0 ;
  assign y23708 = ~n47886 ;
  assign y23709 = ~1'b0 ;
  assign y23710 = n47887 ;
  assign y23711 = ~n47889 ;
  assign y23712 = n47893 ;
  assign y23713 = ~n47896 ;
  assign y23714 = n47897 ;
  assign y23715 = ~n47898 ;
  assign y23716 = ~1'b0 ;
  assign y23717 = n47899 ;
  assign y23718 = ~n47902 ;
  assign y23719 = ~1'b0 ;
  assign y23720 = ~n47903 ;
  assign y23721 = n47913 ;
  assign y23722 = ~n47915 ;
  assign y23723 = n47916 ;
  assign y23724 = ~1'b0 ;
  assign y23725 = ~n47918 ;
  assign y23726 = n47921 ;
  assign y23727 = ~n47924 ;
  assign y23728 = ~n47925 ;
  assign y23729 = ~n47926 ;
  assign y23730 = n47932 ;
  assign y23731 = ~n47935 ;
  assign y23732 = ~n47936 ;
  assign y23733 = ~n47942 ;
  assign y23734 = ~1'b0 ;
  assign y23735 = n9595 ;
  assign y23736 = ~n47945 ;
  assign y23737 = ~1'b0 ;
  assign y23738 = n47946 ;
  assign y23739 = ~n47947 ;
  assign y23740 = ~n47952 ;
  assign y23741 = n47953 ;
  assign y23742 = ~n2254 ;
  assign y23743 = n47954 ;
  assign y23744 = ~1'b0 ;
  assign y23745 = ~1'b0 ;
  assign y23746 = ~1'b0 ;
  assign y23747 = ~1'b0 ;
  assign y23748 = ~n47958 ;
  assign y23749 = n47965 ;
  assign y23750 = ~n47966 ;
  assign y23751 = n47967 ;
  assign y23752 = n47969 ;
  assign y23753 = ~n47970 ;
  assign y23754 = n47976 ;
  assign y23755 = ~n47978 ;
  assign y23756 = n47979 ;
  assign y23757 = ~1'b0 ;
  assign y23758 = n47980 ;
  assign y23759 = n47981 ;
  assign y23760 = n47984 ;
  assign y23761 = n47987 ;
  assign y23762 = ~n47988 ;
  assign y23763 = ~1'b0 ;
  assign y23764 = n47989 ;
  assign y23765 = ~1'b0 ;
  assign y23766 = n47991 ;
  assign y23767 = ~n47995 ;
  assign y23768 = ~1'b0 ;
  assign y23769 = n47996 ;
  assign y23770 = ~n47997 ;
  assign y23771 = ~n47998 ;
  assign y23772 = n47999 ;
  assign y23773 = n48001 ;
  assign y23774 = n48003 ;
  assign y23775 = ~n48004 ;
  assign y23776 = ~1'b0 ;
  assign y23777 = ~1'b0 ;
  assign y23778 = n48005 ;
  assign y23779 = ~n48006 ;
  assign y23780 = ~n48007 ;
  assign y23781 = ~n48011 ;
  assign y23782 = n48015 ;
  assign y23783 = n48016 ;
  assign y23784 = ~1'b0 ;
  assign y23785 = ~1'b0 ;
  assign y23786 = ~1'b0 ;
  assign y23787 = ~n48017 ;
  assign y23788 = ~1'b0 ;
  assign y23789 = ~n48019 ;
  assign y23790 = n48022 ;
  assign y23791 = n48023 ;
  assign y23792 = ~n48026 ;
  assign y23793 = ~n48028 ;
  assign y23794 = n48029 ;
  assign y23795 = ~n48030 ;
  assign y23796 = ~1'b0 ;
  assign y23797 = ~n48033 ;
  assign y23798 = n48034 ;
  assign y23799 = ~1'b0 ;
  assign y23800 = ~n48036 ;
  assign y23801 = ~n43767 ;
  assign y23802 = ~n48039 ;
  assign y23803 = n43515 ;
  assign y23804 = n48044 ;
  assign y23805 = ~1'b0 ;
  assign y23806 = ~1'b0 ;
  assign y23807 = n48046 ;
  assign y23808 = n48047 ;
  assign y23809 = ~1'b0 ;
  assign y23810 = ~n48048 ;
  assign y23811 = ~1'b0 ;
  assign y23812 = ~n48054 ;
  assign y23813 = n48060 ;
  assign y23814 = ~n48064 ;
  assign y23815 = n48068 ;
  assign y23816 = ~1'b0 ;
  assign y23817 = ~n48071 ;
  assign y23818 = n48072 ;
  assign y23819 = n48073 ;
  assign y23820 = n48074 ;
  assign y23821 = ~n48076 ;
  assign y23822 = ~1'b0 ;
  assign y23823 = ~n48078 ;
  assign y23824 = ~1'b0 ;
  assign y23825 = ~1'b0 ;
  assign y23826 = ~n48083 ;
  assign y23827 = ~n48085 ;
  assign y23828 = ~n48092 ;
  assign y23829 = ~1'b0 ;
  assign y23830 = ~n48093 ;
  assign y23831 = n48096 ;
  assign y23832 = n48097 ;
  assign y23833 = ~n35640 ;
  assign y23834 = n48099 ;
  assign y23835 = ~1'b0 ;
  assign y23836 = 1'b0 ;
  assign y23837 = n48102 ;
  assign y23838 = ~n48105 ;
  assign y23839 = n48106 ;
  assign y23840 = ~n48108 ;
  assign y23841 = ~1'b0 ;
  assign y23842 = ~1'b0 ;
  assign y23843 = ~n48113 ;
  assign y23844 = n28636 ;
  assign y23845 = ~1'b0 ;
  assign y23846 = ~n48114 ;
  assign y23847 = n48117 ;
  assign y23848 = ~n48119 ;
  assign y23849 = n48125 ;
  assign y23850 = ~n48126 ;
  assign y23851 = ~1'b0 ;
  assign y23852 = n48127 ;
  assign y23853 = ~n48129 ;
  assign y23854 = ~n48131 ;
  assign y23855 = ~1'b0 ;
  assign y23856 = n48134 ;
  assign y23857 = ~1'b0 ;
  assign y23858 = ~1'b0 ;
  assign y23859 = ~n48140 ;
  assign y23860 = n48147 ;
  assign y23861 = n48149 ;
  assign y23862 = n48155 ;
  assign y23863 = n48157 ;
  assign y23864 = n488 ;
  assign y23865 = ~1'b0 ;
  assign y23866 = ~n48158 ;
  assign y23867 = n48160 ;
  assign y23868 = ~n48161 ;
  assign y23869 = ~n48163 ;
  assign y23870 = n48165 ;
  assign y23871 = ~n48166 ;
  assign y23872 = ~n48172 ;
  assign y23873 = n48173 ;
  assign y23874 = ~1'b0 ;
  assign y23875 = n48174 ;
  assign y23876 = n48175 ;
  assign y23877 = ~n48176 ;
  assign y23878 = n48177 ;
  assign y23879 = ~n48179 ;
  assign y23880 = ~1'b0 ;
  assign y23881 = ~1'b0 ;
  assign y23882 = n48180 ;
  assign y23883 = n48181 ;
  assign y23884 = ~n48184 ;
  assign y23885 = ~1'b0 ;
  assign y23886 = ~n48192 ;
  assign y23887 = ~1'b0 ;
  assign y23888 = n48195 ;
  assign y23889 = n48197 ;
  assign y23890 = ~n48198 ;
  assign y23891 = n48200 ;
  assign y23892 = n48201 ;
  assign y23893 = n19150 ;
  assign y23894 = ~1'b0 ;
  assign y23895 = n48205 ;
  assign y23896 = n48206 ;
  assign y23897 = n48208 ;
  assign y23898 = ~n48211 ;
  assign y23899 = ~n48212 ;
  assign y23900 = n48214 ;
  assign y23901 = ~n48217 ;
  assign y23902 = ~n48219 ;
  assign y23903 = ~n36693 ;
  assign y23904 = n48220 ;
  assign y23905 = ~1'b0 ;
  assign y23906 = ~n48228 ;
  assign y23907 = ~n48229 ;
  assign y23908 = ~1'b0 ;
  assign y23909 = ~1'b0 ;
  assign y23910 = n48232 ;
  assign y23911 = ~n48233 ;
  assign y23912 = ~n48234 ;
  assign y23913 = n48236 ;
  assign y23914 = ~1'b0 ;
  assign y23915 = n18336 ;
  assign y23916 = n48237 ;
  assign y23917 = ~n48243 ;
  assign y23918 = ~1'b0 ;
  assign y23919 = ~1'b0 ;
  assign y23920 = ~n48244 ;
  assign y23921 = ~n13666 ;
  assign y23922 = n48247 ;
  assign y23923 = ~n48249 ;
  assign y23924 = ~1'b0 ;
  assign y23925 = ~n48250 ;
  assign y23926 = ~1'b0 ;
  assign y23927 = ~1'b0 ;
  assign y23928 = n48251 ;
  assign y23929 = n48253 ;
  assign y23930 = ~n48254 ;
  assign y23931 = ~n48255 ;
  assign y23932 = ~n48257 ;
  assign y23933 = ~1'b0 ;
  assign y23934 = ~1'b0 ;
  assign y23935 = ~n16815 ;
  assign y23936 = ~n48259 ;
  assign y23937 = n48262 ;
  assign y23938 = n48268 ;
  assign y23939 = ~1'b0 ;
  assign y23940 = ~n48270 ;
  assign y23941 = ~n48271 ;
  assign y23942 = ~n48273 ;
  assign y23943 = n48275 ;
  assign y23944 = n48279 ;
  assign y23945 = ~n48280 ;
  assign y23946 = n48282 ;
  assign y23947 = n18730 ;
  assign y23948 = ~1'b0 ;
  assign y23949 = ~n21443 ;
  assign y23950 = n48285 ;
  assign y23951 = n48289 ;
  assign y23952 = ~n48290 ;
  assign y23953 = ~n48296 ;
  assign y23954 = ~1'b0 ;
  assign y23955 = ~n43802 ;
  assign y23956 = ~n48298 ;
  assign y23957 = ~n48300 ;
  assign y23958 = ~n48301 ;
  assign y23959 = n48302 ;
  assign y23960 = ~n48303 ;
  assign y23961 = 1'b0 ;
  assign y23962 = ~1'b0 ;
  assign y23963 = n48304 ;
  assign y23964 = ~n48306 ;
  assign y23965 = n48308 ;
  assign y23966 = ~1'b0 ;
  assign y23967 = n48309 ;
  assign y23968 = ~n6105 ;
  assign y23969 = n48310 ;
  assign y23970 = ~1'b0 ;
  assign y23971 = ~1'b0 ;
  assign y23972 = n10821 ;
  assign y23973 = ~n48315 ;
  assign y23974 = ~1'b0 ;
  assign y23975 = ~n48318 ;
  assign y23976 = ~1'b0 ;
  assign y23977 = ~n48319 ;
  assign y23978 = n48321 ;
  assign y23979 = ~n48322 ;
  assign y23980 = ~1'b0 ;
  assign y23981 = ~n3797 ;
  assign y23982 = ~n48325 ;
  assign y23983 = ~1'b0 ;
  assign y23984 = ~1'b0 ;
  assign y23985 = n48331 ;
  assign y23986 = n48333 ;
  assign y23987 = n48334 ;
  assign y23988 = ~1'b0 ;
  assign y23989 = ~n48336 ;
  assign y23990 = n48338 ;
  assign y23991 = n48339 ;
  assign y23992 = n48341 ;
  assign y23993 = n48343 ;
  assign y23994 = n48345 ;
  assign y23995 = ~n48349 ;
  assign y23996 = ~n48350 ;
  assign y23997 = ~n38668 ;
  assign y23998 = n18280 ;
  assign y23999 = ~1'b0 ;
  assign y24000 = ~n23644 ;
  assign y24001 = n48356 ;
  assign y24002 = ~n48358 ;
  assign y24003 = ~n48361 ;
  assign y24004 = n48366 ;
  assign y24005 = ~n48368 ;
  assign y24006 = n48369 ;
  assign y24007 = ~1'b0 ;
  assign y24008 = n5078 ;
  assign y24009 = ~n48373 ;
  assign y24010 = n48374 ;
  assign y24011 = n48380 ;
  assign y24012 = ~n48381 ;
  assign y24013 = n48382 ;
  assign y24014 = n48385 ;
  assign y24015 = ~n48386 ;
  assign y24016 = n48389 ;
  assign y24017 = ~n48391 ;
  assign y24018 = ~n48394 ;
  assign y24019 = ~n48399 ;
  assign y24020 = ~1'b0 ;
  assign y24021 = ~1'b0 ;
  assign y24022 = ~1'b0 ;
  assign y24023 = n48400 ;
  assign y24024 = ~n48401 ;
  assign y24025 = n48403 ;
  assign y24026 = ~n48406 ;
  assign y24027 = ~1'b0 ;
  assign y24028 = n48408 ;
  assign y24029 = ~n48411 ;
  assign y24030 = ~1'b0 ;
  assign y24031 = ~1'b0 ;
  assign y24032 = n48412 ;
  assign y24033 = n48413 ;
  assign y24034 = ~n48414 ;
  assign y24035 = ~n48415 ;
  assign y24036 = n48417 ;
  assign y24037 = ~n48421 ;
  assign y24038 = ~1'b0 ;
  assign y24039 = ~1'b0 ;
  assign y24040 = ~n48422 ;
  assign y24041 = n48424 ;
  assign y24042 = ~n48426 ;
  assign y24043 = ~n48427 ;
  assign y24044 = n48429 ;
  assign y24045 = n48431 ;
  assign y24046 = ~1'b0 ;
  assign y24047 = ~n48436 ;
  assign y24048 = ~n41534 ;
  assign y24049 = ~n48437 ;
  assign y24050 = n48439 ;
  assign y24051 = n48443 ;
  assign y24052 = ~n48444 ;
  assign y24053 = ~n48446 ;
  assign y24054 = ~1'b0 ;
  assign y24055 = n48449 ;
  assign y24056 = ~n48450 ;
  assign y24057 = n48451 ;
  assign y24058 = n48452 ;
  assign y24059 = n48453 ;
  assign y24060 = ~n48454 ;
  assign y24061 = n48456 ;
  assign y24062 = ~n48457 ;
  assign y24063 = ~1'b0 ;
  assign y24064 = ~1'b0 ;
  assign y24065 = n2064 ;
  assign y24066 = ~1'b0 ;
  assign y24067 = ~n48460 ;
  assign y24068 = ~1'b0 ;
  assign y24069 = ~n48462 ;
  assign y24070 = ~n48466 ;
  assign y24071 = ~n48469 ;
  assign y24072 = ~n48473 ;
  assign y24073 = ~1'b0 ;
  assign y24074 = ~n48474 ;
  assign y24075 = ~1'b0 ;
  assign y24076 = ~n48477 ;
  assign y24077 = n48480 ;
  assign y24078 = n48483 ;
  assign y24079 = n48484 ;
  assign y24080 = n48486 ;
  assign y24081 = ~n48487 ;
  assign y24082 = n48489 ;
  assign y24083 = ~n48490 ;
  assign y24084 = n48492 ;
  assign y24085 = n48494 ;
  assign y24086 = n48496 ;
  assign y24087 = n48498 ;
  assign y24088 = n48500 ;
  assign y24089 = ~n48502 ;
  assign y24090 = ~n48504 ;
  assign y24091 = n48505 ;
  assign y24092 = n48506 ;
  assign y24093 = ~1'b0 ;
  assign y24094 = ~n48508 ;
  assign y24095 = ~1'b0 ;
  assign y24096 = n48510 ;
  assign y24097 = ~n48511 ;
  assign y24098 = n48513 ;
  assign y24099 = n9045 ;
  assign y24100 = ~n48514 ;
  assign y24101 = n48520 ;
  assign y24102 = n48525 ;
  assign y24103 = ~1'b0 ;
  assign y24104 = ~1'b0 ;
  assign y24105 = n48526 ;
  assign y24106 = ~n48527 ;
  assign y24107 = ~n48528 ;
  assign y24108 = n48530 ;
  assign y24109 = n4617 ;
  assign y24110 = ~n48531 ;
  assign y24111 = ~n48535 ;
  assign y24112 = ~n48536 ;
  assign y24113 = ~n48537 ;
  assign y24114 = n48538 ;
  assign y24115 = ~1'b0 ;
  assign y24116 = ~n48541 ;
  assign y24117 = n48545 ;
  assign y24118 = n48546 ;
  assign y24119 = ~n48549 ;
  assign y24120 = ~n48553 ;
  assign y24121 = ~n48555 ;
  assign y24122 = n48556 ;
  assign y24123 = n48558 ;
  assign y24124 = 1'b0 ;
  assign y24125 = ~1'b0 ;
  assign y24126 = n48559 ;
  assign y24127 = ~n48561 ;
  assign y24128 = ~1'b0 ;
  assign y24129 = ~n48563 ;
  assign y24130 = n48567 ;
  assign y24131 = ~1'b0 ;
  assign y24132 = ~n48571 ;
  assign y24133 = n48574 ;
  assign y24134 = ~n48575 ;
  assign y24135 = ~n48578 ;
  assign y24136 = ~n48581 ;
  assign y24137 = n48582 ;
  assign y24138 = ~n48585 ;
  assign y24139 = n48591 ;
  assign y24140 = ~n48594 ;
  assign y24141 = ~1'b0 ;
  assign y24142 = n48595 ;
  assign y24143 = n48597 ;
  assign y24144 = ~1'b0 ;
  assign y24145 = n48600 ;
  assign y24146 = ~n48601 ;
  assign y24147 = ~n48604 ;
  assign y24148 = ~1'b0 ;
  assign y24149 = ~n48606 ;
  assign y24150 = n48609 ;
  assign y24151 = ~n48616 ;
  assign y24152 = ~n48617 ;
  assign y24153 = n48620 ;
  assign y24154 = n48621 ;
  assign y24155 = n48624 ;
  assign y24156 = 1'b0 ;
  assign y24157 = n48629 ;
  assign y24158 = ~n48631 ;
  assign y24159 = 1'b0 ;
  assign y24160 = ~1'b0 ;
  assign y24161 = ~n48637 ;
  assign y24162 = n48640 ;
  assign y24163 = n48645 ;
  assign y24164 = n48332 ;
  assign y24165 = ~1'b0 ;
  assign y24166 = ~n48647 ;
  assign y24167 = ~n48648 ;
  assign y24168 = ~1'b0 ;
  assign y24169 = ~1'b0 ;
  assign y24170 = ~n48650 ;
  assign y24171 = ~n48652 ;
  assign y24172 = ~n6875 ;
  assign y24173 = ~n48653 ;
  assign y24174 = ~n48654 ;
  assign y24175 = n48658 ;
  assign y24176 = ~1'b0 ;
  assign y24177 = ~1'b0 ;
  assign y24178 = n48660 ;
  assign y24179 = ~n24268 ;
  assign y24180 = ~n48663 ;
  assign y24181 = ~n48664 ;
  assign y24182 = ~1'b0 ;
  assign y24183 = ~1'b0 ;
  assign y24184 = ~n48667 ;
  assign y24185 = ~n48671 ;
  assign y24186 = n48673 ;
  assign y24187 = 1'b0 ;
  assign y24188 = ~n48675 ;
  assign y24189 = ~1'b0 ;
  assign y24190 = ~n48677 ;
  assign y24191 = n48680 ;
  assign y24192 = ~1'b0 ;
  assign y24193 = n48682 ;
  assign y24194 = n48685 ;
  assign y24195 = ~n48686 ;
  assign y24196 = ~n48689 ;
  assign y24197 = n48690 ;
  assign y24198 = ~1'b0 ;
  assign y24199 = n48693 ;
  assign y24200 = ~1'b0 ;
  assign y24201 = ~n48696 ;
  assign y24202 = n48698 ;
  assign y24203 = ~n48700 ;
  assign y24204 = n48706 ;
  assign y24205 = ~n48710 ;
  assign y24206 = ~n48712 ;
  assign y24207 = ~1'b0 ;
  assign y24208 = ~n42243 ;
  assign y24209 = ~1'b0 ;
  assign y24210 = n48714 ;
  assign y24211 = n48718 ;
  assign y24212 = ~n48720 ;
  assign y24213 = n48724 ;
  assign y24214 = n48726 ;
  assign y24215 = ~n48727 ;
  assign y24216 = ~1'b0 ;
  assign y24217 = ~1'b0 ;
  assign y24218 = 1'b0 ;
  assign y24219 = n48728 ;
  assign y24220 = n48731 ;
  assign y24221 = ~n2170 ;
  assign y24222 = ~n48734 ;
  assign y24223 = ~1'b0 ;
  assign y24224 = n48737 ;
  assign y24225 = ~n48739 ;
  assign y24226 = n48743 ;
  assign y24227 = ~1'b0 ;
  assign y24228 = ~n48744 ;
  assign y24229 = n48746 ;
  assign y24230 = ~n48748 ;
  assign y24231 = n48751 ;
  assign y24232 = ~n48753 ;
  assign y24233 = n48754 ;
  assign y24234 = n48755 ;
  assign y24235 = ~n48759 ;
  assign y24236 = ~1'b0 ;
  assign y24237 = 1'b0 ;
  assign y24238 = ~1'b0 ;
  assign y24239 = n48764 ;
  assign y24240 = ~n48765 ;
  assign y24241 = ~1'b0 ;
  assign y24242 = ~n14973 ;
  assign y24243 = ~n48771 ;
  assign y24244 = ~1'b0 ;
  assign y24245 = ~1'b0 ;
  assign y24246 = ~n48775 ;
  assign y24247 = ~n48779 ;
  assign y24248 = ~n30060 ;
  assign y24249 = ~1'b0 ;
  assign y24250 = ~n48780 ;
  assign y24251 = ~1'b0 ;
  assign y24252 = n48782 ;
  assign y24253 = n48785 ;
  assign y24254 = n48790 ;
  assign y24255 = ~n48794 ;
  assign y24256 = ~n48795 ;
  assign y24257 = n48798 ;
  assign y24258 = ~1'b0 ;
  assign y24259 = ~n48799 ;
  assign y24260 = n48800 ;
  assign y24261 = ~1'b0 ;
  assign y24262 = n23113 ;
  assign y24263 = ~n48803 ;
  assign y24264 = ~1'b0 ;
  assign y24265 = ~1'b0 ;
  assign y24266 = n48804 ;
  assign y24267 = n48805 ;
  assign y24268 = ~1'b0 ;
  assign y24269 = ~n48806 ;
  assign y24270 = ~n48808 ;
  assign y24271 = ~1'b0 ;
  assign y24272 = ~n48810 ;
  assign y24273 = n48811 ;
  assign y24274 = ~n48813 ;
  assign y24275 = ~1'b0 ;
  assign y24276 = ~1'b0 ;
  assign y24277 = ~n48817 ;
  assign y24278 = n48818 ;
  assign y24279 = 1'b0 ;
  assign y24280 = 1'b0 ;
  assign y24281 = ~n48819 ;
  assign y24282 = ~1'b0 ;
  assign y24283 = n48820 ;
  assign y24284 = n48826 ;
  assign y24285 = n48827 ;
  assign y24286 = n48829 ;
  assign y24287 = ~1'b0 ;
  assign y24288 = n48836 ;
  assign y24289 = ~n48840 ;
  assign y24290 = n48841 ;
  assign y24291 = ~n48847 ;
  assign y24292 = ~n48851 ;
  assign y24293 = n48852 ;
  assign y24294 = n48854 ;
  assign y24295 = n48856 ;
  assign y24296 = n33946 ;
  assign y24297 = ~n48862 ;
  assign y24298 = ~1'b0 ;
  assign y24299 = ~n48871 ;
  assign y24300 = ~n48875 ;
  assign y24301 = n40264 ;
  assign y24302 = ~1'b0 ;
  assign y24303 = ~n48877 ;
  assign y24304 = ~n48883 ;
  assign y24305 = ~1'b0 ;
  assign y24306 = ~n48884 ;
  assign y24307 = n48887 ;
  assign y24308 = n48889 ;
  assign y24309 = ~n48892 ;
  assign y24310 = n48895 ;
  assign y24311 = ~1'b0 ;
  assign y24312 = n31009 ;
  assign y24313 = ~1'b0 ;
  assign y24314 = ~1'b0 ;
  assign y24315 = n7356 ;
  assign y24316 = n48896 ;
  assign y24317 = ~n48897 ;
  assign y24318 = n48900 ;
  assign y24319 = ~1'b0 ;
  assign y24320 = n48903 ;
  assign y24321 = n48906 ;
  assign y24322 = ~1'b0 ;
  assign y24323 = n48908 ;
  assign y24324 = ~n48912 ;
  assign y24325 = n48914 ;
  assign y24326 = ~n48916 ;
  assign y24327 = ~n48917 ;
  assign y24328 = ~n48920 ;
  assign y24329 = ~n48923 ;
  assign y24330 = ~1'b0 ;
  assign y24331 = n48929 ;
  assign y24332 = n48931 ;
  assign y24333 = ~n48932 ;
  assign y24334 = ~n48933 ;
  assign y24335 = ~n48936 ;
  assign y24336 = n36113 ;
  assign y24337 = n48938 ;
  assign y24338 = n48939 ;
  assign y24339 = ~n48940 ;
  assign y24340 = ~1'b0 ;
  assign y24341 = ~1'b0 ;
  assign y24342 = n48945 ;
  assign y24343 = ~n48950 ;
  assign y24344 = n48951 ;
  assign y24345 = ~n48954 ;
  assign y24346 = n48958 ;
  assign y24347 = ~1'b0 ;
  assign y24348 = ~1'b0 ;
  assign y24349 = n25341 ;
  assign y24350 = ~n48961 ;
  assign y24351 = ~n48963 ;
  assign y24352 = ~n48966 ;
  assign y24353 = ~n48970 ;
  assign y24354 = ~n48971 ;
  assign y24355 = ~1'b0 ;
  assign y24356 = n48972 ;
  assign y24357 = n48976 ;
  assign y24358 = ~1'b0 ;
  assign y24359 = ~n48977 ;
  assign y24360 = n48980 ;
  assign y24361 = ~n48982 ;
  assign y24362 = n48983 ;
  assign y24363 = ~n48984 ;
  assign y24364 = n48987 ;
  assign y24365 = n29903 ;
  assign y24366 = n48989 ;
  assign y24367 = n48991 ;
  assign y24368 = ~1'b0 ;
  assign y24369 = ~n48993 ;
  assign y24370 = n48994 ;
  assign y24371 = ~1'b0 ;
  assign y24372 = ~1'b0 ;
  assign y24373 = n48996 ;
  assign y24374 = ~n49002 ;
  assign y24375 = ~n49003 ;
  assign y24376 = ~n49006 ;
  assign y24377 = ~1'b0 ;
  assign y24378 = ~n28410 ;
  assign y24379 = ~1'b0 ;
  assign y24380 = n49009 ;
  assign y24381 = ~n49010 ;
  assign y24382 = n49011 ;
  assign y24383 = ~1'b0 ;
  assign y24384 = n49015 ;
  assign y24385 = ~n49018 ;
  assign y24386 = ~1'b0 ;
  assign y24387 = ~n49021 ;
  assign y24388 = n49027 ;
  assign y24389 = ~n49028 ;
  assign y24390 = n49030 ;
  assign y24391 = n49031 ;
  assign y24392 = ~n49033 ;
  assign y24393 = ~n49034 ;
  assign y24394 = ~n49035 ;
  assign y24395 = ~n49038 ;
  assign y24396 = ~1'b0 ;
  assign y24397 = n49041 ;
  assign y24398 = n26391 ;
  assign y24399 = ~1'b0 ;
  assign y24400 = n49042 ;
  assign y24401 = ~n49044 ;
  assign y24402 = n49048 ;
  assign y24403 = ~1'b0 ;
  assign y24404 = ~1'b0 ;
  assign y24405 = n49049 ;
  assign y24406 = n49051 ;
  assign y24407 = ~1'b0 ;
  assign y24408 = ~n49054 ;
  assign y24409 = n49056 ;
  assign y24410 = ~n49059 ;
  assign y24411 = ~n49061 ;
  assign y24412 = n49062 ;
  assign y24413 = ~n49067 ;
  assign y24414 = ~n49069 ;
  assign y24415 = ~n49071 ;
  assign y24416 = ~n49072 ;
  assign y24417 = ~n17079 ;
  assign y24418 = n49073 ;
  assign y24419 = n49074 ;
  assign y24420 = ~1'b0 ;
  assign y24421 = n49076 ;
  assign y24422 = n23442 ;
  assign y24423 = ~1'b0 ;
  assign y24424 = ~n49077 ;
  assign y24425 = n49078 ;
  assign y24426 = n49082 ;
  assign y24427 = ~1'b0 ;
  assign y24428 = n49089 ;
  assign y24429 = ~n49090 ;
  assign y24430 = ~1'b0 ;
  assign y24431 = n49093 ;
  assign y24432 = ~n49095 ;
  assign y24433 = ~1'b0 ;
  assign y24434 = ~n49096 ;
  assign y24435 = ~n49099 ;
  assign y24436 = ~n49103 ;
  assign y24437 = n49104 ;
  assign y24438 = ~1'b0 ;
  assign y24439 = ~n49106 ;
  assign y24440 = ~1'b0 ;
  assign y24441 = ~n49111 ;
  assign y24442 = n49113 ;
  assign y24443 = 1'b0 ;
  assign y24444 = ~1'b0 ;
  assign y24445 = ~n49114 ;
  assign y24446 = ~n49115 ;
  assign y24447 = ~n49116 ;
  assign y24448 = n49120 ;
  assign y24449 = ~n29478 ;
  assign y24450 = ~1'b0 ;
  assign y24451 = ~n49122 ;
  assign y24452 = n49123 ;
  assign y24453 = ~1'b0 ;
  assign y24454 = ~n49126 ;
  assign y24455 = n13067 ;
  assign y24456 = n49132 ;
  assign y24457 = ~n49136 ;
  assign y24458 = ~1'b0 ;
  assign y24459 = ~n49137 ;
  assign y24460 = ~1'b0 ;
  assign y24461 = n33166 ;
  assign y24462 = ~n49138 ;
  assign y24463 = ~n49143 ;
  assign y24464 = ~n49146 ;
  assign y24465 = ~1'b0 ;
  assign y24466 = n49148 ;
  assign y24467 = ~n49149 ;
  assign y24468 = ~n49150 ;
  assign y24469 = ~n49153 ;
  assign y24470 = n33304 ;
  assign y24471 = n49154 ;
  assign y24472 = ~1'b0 ;
  assign y24473 = ~1'b0 ;
  assign y24474 = ~n49156 ;
  assign y24475 = ~n49158 ;
  assign y24476 = n49161 ;
  assign y24477 = ~n49165 ;
  assign y24478 = n49168 ;
  assign y24479 = n15065 ;
  assign y24480 = ~n49169 ;
  assign y24481 = n49175 ;
  assign y24482 = ~1'b0 ;
  assign y24483 = ~1'b0 ;
  assign y24484 = ~1'b0 ;
  assign y24485 = ~1'b0 ;
  assign y24486 = ~n49181 ;
  assign y24487 = ~n49183 ;
  assign y24488 = ~1'b0 ;
  assign y24489 = n49185 ;
  assign y24490 = n49187 ;
  assign y24491 = n49188 ;
  assign y24492 = n49190 ;
  assign y24493 = ~1'b0 ;
  assign y24494 = ~1'b0 ;
  assign y24495 = ~1'b0 ;
  assign y24496 = n49192 ;
  assign y24497 = ~1'b0 ;
  assign y24498 = ~n49194 ;
  assign y24499 = n49197 ;
  assign y24500 = ~1'b0 ;
  assign y24501 = ~n49199 ;
  assign y24502 = ~n49202 ;
  assign y24503 = ~n46216 ;
  assign y24504 = ~n49206 ;
  assign y24505 = n49208 ;
  assign y24506 = ~1'b0 ;
  assign y24507 = n49210 ;
  assign y24508 = ~n49211 ;
  assign y24509 = n49212 ;
  assign y24510 = n49213 ;
  assign y24511 = 1'b0 ;
  assign y24512 = ~n49214 ;
  assign y24513 = n49215 ;
  assign y24514 = ~1'b0 ;
  assign y24515 = ~n49216 ;
  assign y24516 = n2701 ;
  assign y24517 = ~1'b0 ;
  assign y24518 = ~n49217 ;
  assign y24519 = ~1'b0 ;
  assign y24520 = ~n49218 ;
  assign y24521 = n49221 ;
  assign y24522 = ~n49222 ;
  assign y24523 = ~n49229 ;
  assign y24524 = ~1'b0 ;
  assign y24525 = ~n49232 ;
  assign y24526 = n49234 ;
  assign y24527 = n49236 ;
  assign y24528 = ~n49238 ;
  assign y24529 = ~n49243 ;
  assign y24530 = ~n12929 ;
  assign y24531 = ~n49246 ;
  assign y24532 = n49248 ;
  assign y24533 = ~n49251 ;
  assign y24534 = n49252 ;
  assign y24535 = n49253 ;
  assign y24536 = ~n49258 ;
  assign y24537 = n49260 ;
  assign y24538 = ~n49262 ;
  assign y24539 = ~n49263 ;
  assign y24540 = ~1'b0 ;
  assign y24541 = ~n49264 ;
  assign y24542 = ~n49266 ;
  assign y24543 = ~n49269 ;
  assign y24544 = n49272 ;
  assign y24545 = n49273 ;
  assign y24546 = ~n49276 ;
  assign y24547 = ~n49278 ;
  assign y24548 = n49280 ;
  assign y24549 = ~1'b0 ;
  assign y24550 = ~n49282 ;
  assign y24551 = ~n49284 ;
  assign y24552 = n49286 ;
  assign y24553 = n49287 ;
  assign y24554 = ~n49291 ;
  assign y24555 = n49292 ;
  assign y24556 = ~n49294 ;
  assign y24557 = n49298 ;
  assign y24558 = ~1'b0 ;
  assign y24559 = ~n49299 ;
  assign y24560 = n49300 ;
  assign y24561 = ~n49301 ;
  assign y24562 = ~n49303 ;
  assign y24563 = ~n49305 ;
  assign y24564 = ~1'b0 ;
  assign y24565 = n49307 ;
  assign y24566 = n49309 ;
  assign y24567 = ~1'b0 ;
  assign y24568 = ~n49312 ;
  assign y24569 = ~n49318 ;
  assign y24570 = ~1'b0 ;
  assign y24571 = 1'b0 ;
  assign y24572 = ~n49321 ;
  assign y24573 = ~n49323 ;
  assign y24574 = n49325 ;
  assign y24575 = ~1'b0 ;
  assign y24576 = ~1'b0 ;
  assign y24577 = ~n49327 ;
  assign y24578 = ~n49329 ;
  assign y24579 = n49332 ;
  assign y24580 = ~n49339 ;
  assign y24581 = ~n49341 ;
  assign y24582 = n49342 ;
  assign y24583 = n49344 ;
  assign y24584 = ~1'b0 ;
  assign y24585 = ~1'b0 ;
  assign y24586 = n49348 ;
  assign y24587 = ~n49350 ;
  assign y24588 = ~n49354 ;
  assign y24589 = ~1'b0 ;
  assign y24590 = n49356 ;
  assign y24591 = n49358 ;
  assign y24592 = ~n49359 ;
  assign y24593 = 1'b0 ;
  assign y24594 = ~1'b0 ;
  assign y24595 = n49363 ;
  assign y24596 = n49365 ;
  assign y24597 = ~n49366 ;
  assign y24598 = n49368 ;
  assign y24599 = n49369 ;
  assign y24600 = n30974 ;
  assign y24601 = ~n49370 ;
  assign y24602 = n49371 ;
  assign y24603 = n49372 ;
  assign y24604 = 1'b0 ;
  assign y24605 = n49381 ;
  assign y24606 = ~n49382 ;
  assign y24607 = ~1'b0 ;
  assign y24608 = n49383 ;
  assign y24609 = n49385 ;
  assign y24610 = ~n49392 ;
  assign y24611 = ~1'b0 ;
  assign y24612 = ~n1768 ;
  assign y24613 = n49397 ;
  assign y24614 = ~1'b0 ;
  assign y24615 = ~n49400 ;
  assign y24616 = ~n9528 ;
  assign y24617 = n49401 ;
  assign y24618 = n49405 ;
  assign y24619 = ~1'b0 ;
  assign y24620 = ~n49409 ;
  assign y24621 = ~1'b0 ;
  assign y24622 = n49411 ;
  assign y24623 = n49412 ;
  assign y24624 = 1'b0 ;
  assign y24625 = 1'b0 ;
  assign y24626 = n49413 ;
  assign y24627 = n49414 ;
  assign y24628 = ~1'b0 ;
  assign y24629 = n49417 ;
  assign y24630 = n49418 ;
  assign y24631 = ~n49419 ;
  assign y24632 = n49422 ;
  assign y24633 = ~n49425 ;
  assign y24634 = n49426 ;
  assign y24635 = ~n49428 ;
  assign y24636 = n49433 ;
  assign y24637 = ~n49434 ;
  assign y24638 = ~1'b0 ;
  assign y24639 = ~n49438 ;
  assign y24640 = ~n49440 ;
  assign y24641 = ~n49442 ;
  assign y24642 = ~1'b0 ;
  assign y24643 = n49444 ;
  assign y24644 = ~n49445 ;
  assign y24645 = ~n49446 ;
  assign y24646 = ~n49449 ;
  assign y24647 = ~1'b0 ;
  assign y24648 = n49450 ;
  assign y24649 = ~1'b0 ;
  assign y24650 = ~1'b0 ;
  assign y24651 = ~1'b0 ;
  assign y24652 = ~1'b0 ;
  assign y24653 = ~n49451 ;
  assign y24654 = n49454 ;
  assign y24655 = ~n49458 ;
  assign y24656 = ~n49459 ;
  assign y24657 = n49463 ;
  assign y24658 = ~n49465 ;
  assign y24659 = n49469 ;
  assign y24660 = n49472 ;
  assign y24661 = n49474 ;
  assign y24662 = ~n49475 ;
  assign y24663 = ~n27432 ;
  assign y24664 = ~n49477 ;
  assign y24665 = n49481 ;
  assign y24666 = ~n49487 ;
  assign y24667 = n49489 ;
  assign y24668 = ~n49490 ;
  assign y24669 = n49494 ;
  assign y24670 = ~n49495 ;
  assign y24671 = ~n49498 ;
  assign y24672 = ~n6101 ;
  assign y24673 = n39479 ;
  assign y24674 = n49501 ;
  assign y24675 = ~n49503 ;
  assign y24676 = ~1'b0 ;
  assign y24677 = n46989 ;
  assign y24678 = n49506 ;
  assign y24679 = ~1'b0 ;
  assign y24680 = ~n49508 ;
  assign y24681 = n49515 ;
  assign y24682 = ~n49520 ;
  assign y24683 = ~1'b0 ;
  assign y24684 = ~n49523 ;
  assign y24685 = ~n49526 ;
  assign y24686 = n49527 ;
  assign y24687 = ~n49529 ;
  assign y24688 = ~1'b0 ;
  assign y24689 = n49535 ;
  assign y24690 = ~1'b0 ;
  assign y24691 = ~n49536 ;
  assign y24692 = n49538 ;
  assign y24693 = ~n49539 ;
  assign y24694 = n49541 ;
  assign y24695 = ~1'b0 ;
  assign y24696 = n49544 ;
  assign y24697 = ~1'b0 ;
  assign y24698 = 1'b0 ;
  assign y24699 = n49547 ;
  assign y24700 = ~n49549 ;
  assign y24701 = ~n49550 ;
  assign y24702 = n16907 ;
  assign y24703 = ~1'b0 ;
  assign y24704 = n49552 ;
  assign y24705 = ~1'b0 ;
  assign y24706 = ~1'b0 ;
  assign y24707 = n49553 ;
  assign y24708 = ~1'b0 ;
  assign y24709 = ~n49555 ;
  assign y24710 = n49556 ;
  assign y24711 = ~n49557 ;
  assign y24712 = ~1'b0 ;
  assign y24713 = ~1'b0 ;
  assign y24714 = ~1'b0 ;
  assign y24715 = ~n6569 ;
  assign y24716 = n49560 ;
  assign y24717 = ~n49562 ;
  assign y24718 = n49565 ;
  assign y24719 = ~n49566 ;
  assign y24720 = n49567 ;
  assign y24721 = ~n49569 ;
  assign y24722 = n24781 ;
  assign y24723 = n49570 ;
  assign y24724 = ~n49571 ;
  assign y24725 = 1'b0 ;
  assign y24726 = n49574 ;
  assign y24727 = ~n49575 ;
  assign y24728 = ~n49584 ;
  assign y24729 = ~n7902 ;
  assign y24730 = n49586 ;
  assign y24731 = ~1'b0 ;
  assign y24732 = n49588 ;
  assign y24733 = n49596 ;
  assign y24734 = ~n49600 ;
  assign y24735 = ~n49604 ;
  assign y24736 = ~n49605 ;
  assign y24737 = n49609 ;
  assign y24738 = ~n49614 ;
  assign y24739 = ~n49615 ;
  assign y24740 = ~n49621 ;
  assign y24741 = ~1'b0 ;
  assign y24742 = ~1'b0 ;
  assign y24743 = ~n49622 ;
  assign y24744 = ~1'b0 ;
  assign y24745 = ~1'b0 ;
  assign y24746 = ~n49623 ;
  assign y24747 = n49624 ;
  assign y24748 = ~1'b0 ;
  assign y24749 = ~1'b0 ;
  assign y24750 = n49625 ;
  assign y24751 = n49630 ;
  assign y24752 = n7944 ;
  assign y24753 = n49631 ;
  assign y24754 = 1'b0 ;
  assign y24755 = n49634 ;
  assign y24756 = n49636 ;
  assign y24757 = ~n49639 ;
  assign y24758 = ~n49641 ;
  assign y24759 = ~n49644 ;
  assign y24760 = ~1'b0 ;
  assign y24761 = n49646 ;
  assign y24762 = 1'b0 ;
  assign y24763 = n49648 ;
  assign y24764 = ~n5287 ;
  assign y24765 = n49649 ;
  assign y24766 = ~n49652 ;
  assign y24767 = ~n49658 ;
  assign y24768 = n49662 ;
  assign y24769 = ~n49666 ;
  assign y24770 = ~n49669 ;
  assign y24771 = ~n49674 ;
  assign y24772 = n49675 ;
  assign y24773 = n49678 ;
  assign y24774 = ~n39299 ;
  assign y24775 = ~n49680 ;
  assign y24776 = n49682 ;
  assign y24777 = ~n49683 ;
  assign y24778 = ~n49684 ;
  assign y24779 = n49688 ;
  assign y24780 = ~1'b0 ;
  assign y24781 = ~n49690 ;
  assign y24782 = ~1'b0 ;
  assign y24783 = ~1'b0 ;
  assign y24784 = ~1'b0 ;
  assign y24785 = ~n49691 ;
  assign y24786 = n49693 ;
  assign y24787 = ~n49698 ;
  assign y24788 = ~1'b0 ;
  assign y24789 = ~n49700 ;
  assign y24790 = n49702 ;
  assign y24791 = ~n49704 ;
  assign y24792 = n49706 ;
  assign y24793 = ~1'b0 ;
  assign y24794 = n49712 ;
  assign y24795 = n49713 ;
  assign y24796 = ~n49714 ;
  assign y24797 = n49723 ;
  assign y24798 = ~1'b0 ;
  assign y24799 = ~n49729 ;
  assign y24800 = n49733 ;
  assign y24801 = ~n49739 ;
  assign y24802 = n49741 ;
  assign y24803 = ~n49743 ;
  assign y24804 = ~n49748 ;
  assign y24805 = n49752 ;
  assign y24806 = n49754 ;
  assign y24807 = n49756 ;
  assign y24808 = ~n49757 ;
  assign y24809 = ~n49761 ;
  assign y24810 = ~n49763 ;
  assign y24811 = ~n49766 ;
  assign y24812 = n49770 ;
  assign y24813 = ~n49773 ;
  assign y24814 = ~n49780 ;
  assign y24815 = ~n49781 ;
  assign y24816 = ~n49782 ;
  assign y24817 = n49785 ;
  assign y24818 = n49786 ;
  assign y24819 = ~1'b0 ;
  assign y24820 = ~n49787 ;
  assign y24821 = ~1'b0 ;
  assign y24822 = n5594 ;
  assign y24823 = n49788 ;
  assign y24824 = ~1'b0 ;
  assign y24825 = ~n49793 ;
  assign y24826 = ~n49795 ;
  assign y24827 = n49796 ;
  assign y24828 = ~n49800 ;
  assign y24829 = ~n49801 ;
  assign y24830 = ~1'b0 ;
  assign y24831 = ~n49802 ;
  assign y24832 = ~1'b0 ;
  assign y24833 = n49803 ;
  assign y24834 = n49805 ;
  assign y24835 = ~n49806 ;
  assign y24836 = ~n49811 ;
  assign y24837 = 1'b0 ;
  assign y24838 = ~n49814 ;
  assign y24839 = 1'b0 ;
  assign y24840 = n49816 ;
  assign y24841 = ~n49817 ;
  assign y24842 = ~n49819 ;
  assign y24843 = ~1'b0 ;
  assign y24844 = n49821 ;
  assign y24845 = 1'b0 ;
  assign y24846 = n49825 ;
  assign y24847 = n49827 ;
  assign y24848 = ~1'b0 ;
  assign y24849 = n49833 ;
  assign y24850 = ~1'b0 ;
  assign y24851 = n49835 ;
  assign y24852 = ~n49848 ;
  assign y24853 = ~n24149 ;
  assign y24854 = ~1'b0 ;
  assign y24855 = ~n22796 ;
  assign y24856 = ~1'b0 ;
  assign y24857 = ~n49852 ;
  assign y24858 = ~1'b0 ;
  assign y24859 = ~1'b0 ;
  assign y24860 = ~1'b0 ;
  assign y24861 = ~1'b0 ;
  assign y24862 = ~n49853 ;
  assign y24863 = ~n49856 ;
  assign y24864 = n49861 ;
  assign y24865 = ~n2179 ;
  assign y24866 = ~1'b0 ;
  assign y24867 = ~1'b0 ;
  assign y24868 = ~n49863 ;
  assign y24869 = n49864 ;
  assign y24870 = n49868 ;
  assign y24871 = ~1'b0 ;
  assign y24872 = ~1'b0 ;
  assign y24873 = n49869 ;
  assign y24874 = n49870 ;
  assign y24875 = n49871 ;
  assign y24876 = ~1'b0 ;
  assign y24877 = ~n49872 ;
  assign y24878 = ~1'b0 ;
  assign y24879 = n49874 ;
  assign y24880 = ~n49875 ;
  assign y24881 = 1'b0 ;
  assign y24882 = ~n49878 ;
  assign y24883 = ~1'b0 ;
  assign y24884 = n49881 ;
  assign y24885 = ~1'b0 ;
  assign y24886 = ~n49886 ;
  assign y24887 = n49888 ;
  assign y24888 = ~1'b0 ;
  assign y24889 = n49890 ;
  assign y24890 = ~n6820 ;
  assign y24891 = ~1'b0 ;
  assign y24892 = ~1'b0 ;
  assign y24893 = ~n49891 ;
  assign y24894 = ~n49895 ;
  assign y24895 = n49900 ;
  assign y24896 = n49901 ;
  assign y24897 = 1'b0 ;
  assign y24898 = n12867 ;
  assign y24899 = ~n49902 ;
  assign y24900 = ~1'b0 ;
  assign y24901 = n49903 ;
  assign y24902 = ~n49908 ;
  assign y24903 = n49909 ;
  assign y24904 = n49910 ;
  assign y24905 = n49913 ;
  assign y24906 = ~1'b0 ;
  assign y24907 = n49914 ;
  assign y24908 = ~1'b0 ;
  assign y24909 = ~1'b0 ;
  assign y24910 = ~1'b0 ;
  assign y24911 = n49916 ;
  assign y24912 = ~n49920 ;
  assign y24913 = ~n49923 ;
  assign y24914 = n49925 ;
  assign y24915 = ~1'b0 ;
  assign y24916 = 1'b0 ;
  assign y24917 = n49929 ;
  assign y24918 = ~n49931 ;
  assign y24919 = ~1'b0 ;
  assign y24920 = ~n49935 ;
  assign y24921 = n49940 ;
  assign y24922 = ~1'b0 ;
  assign y24923 = n49943 ;
  assign y24924 = ~n49944 ;
  assign y24925 = n49945 ;
  assign y24926 = ~1'b0 ;
  assign y24927 = ~1'b0 ;
  assign y24928 = n49946 ;
  assign y24929 = ~1'b0 ;
  assign y24930 = ~n49947 ;
  assign y24931 = ~1'b0 ;
  assign y24932 = n49952 ;
  assign y24933 = ~n49953 ;
  assign y24934 = ~n49956 ;
  assign y24935 = ~1'b0 ;
  assign y24936 = ~n49957 ;
  assign y24937 = ~n49960 ;
  assign y24938 = ~1'b0 ;
  assign y24939 = ~1'b0 ;
  assign y24940 = ~1'b0 ;
  assign y24941 = ~1'b0 ;
  assign y24942 = n49962 ;
  assign y24943 = ~n49965 ;
  assign y24944 = ~n49966 ;
  assign y24945 = n49968 ;
  assign y24946 = ~1'b0 ;
  assign y24947 = ~n49969 ;
  assign y24948 = n49971 ;
  assign y24949 = ~n49973 ;
  assign y24950 = ~n33628 ;
  assign y24951 = n12860 ;
  assign y24952 = ~n49974 ;
  assign y24953 = n49975 ;
  assign y24954 = ~n49976 ;
  assign y24955 = n12185 ;
  assign y24956 = ~1'b0 ;
  assign y24957 = n49980 ;
  assign y24958 = ~n49986 ;
  assign y24959 = n49991 ;
  assign y24960 = ~n49992 ;
  assign y24961 = n49997 ;
  assign y24962 = n49999 ;
  assign y24963 = ~n50000 ;
  assign y24964 = ~n50002 ;
  assign y24965 = ~1'b0 ;
  assign y24966 = ~n50004 ;
  assign y24967 = ~n50005 ;
  assign y24968 = ~1'b0 ;
  assign y24969 = ~1'b0 ;
  assign y24970 = ~1'b0 ;
  assign y24971 = ~n50011 ;
  assign y24972 = n50012 ;
  assign y24973 = ~n50013 ;
  assign y24974 = ~1'b0 ;
  assign y24975 = 1'b0 ;
  assign y24976 = ~n50014 ;
  assign y24977 = ~n50015 ;
  assign y24978 = n50016 ;
  assign y24979 = n50017 ;
  assign y24980 = ~1'b0 ;
  assign y24981 = ~n50019 ;
  assign y24982 = n50020 ;
  assign y24983 = n50022 ;
  assign y24984 = n50023 ;
  assign y24985 = ~n4214 ;
  assign y24986 = n50028 ;
  assign y24987 = n46563 ;
  assign y24988 = ~1'b0 ;
  assign y24989 = ~1'b0 ;
  assign y24990 = ~n50029 ;
  assign y24991 = ~n50030 ;
  assign y24992 = n50031 ;
  assign y24993 = n50034 ;
  assign y24994 = n5561 ;
  assign y24995 = n50036 ;
  assign y24996 = n50037 ;
  assign y24997 = ~1'b0 ;
  assign y24998 = n50039 ;
  assign y24999 = ~n2083 ;
  assign y25000 = n50046 ;
  assign y25001 = ~n50048 ;
  assign y25002 = ~1'b0 ;
  assign y25003 = n50050 ;
  assign y25004 = n50051 ;
  assign y25005 = ~1'b0 ;
  assign y25006 = n50052 ;
  assign y25007 = n50054 ;
  assign y25008 = ~1'b0 ;
  assign y25009 = ~n49118 ;
  assign y25010 = n25265 ;
  assign y25011 = n50055 ;
  assign y25012 = ~n50056 ;
  assign y25013 = ~n50057 ;
  assign y25014 = ~n50058 ;
  assign y25015 = ~n50062 ;
  assign y25016 = ~1'b0 ;
  assign y25017 = ~n50063 ;
  assign y25018 = ~1'b0 ;
  assign y25019 = n50064 ;
  assign y25020 = ~n50067 ;
  assign y25021 = n50071 ;
  assign y25022 = ~n50072 ;
  assign y25023 = ~1'b0 ;
  assign y25024 = ~1'b0 ;
  assign y25025 = n50074 ;
  assign y25026 = ~n50076 ;
  assign y25027 = ~n50081 ;
  assign y25028 = n50083 ;
  assign y25029 = ~n9275 ;
  assign y25030 = n50084 ;
  assign y25031 = ~n50085 ;
  assign y25032 = ~n50086 ;
  assign y25033 = n50089 ;
  assign y25034 = ~n50091 ;
  assign y25035 = n50092 ;
  assign y25036 = ~n50095 ;
  assign y25037 = ~1'b0 ;
  assign y25038 = n50098 ;
  assign y25039 = n50102 ;
  assign y25040 = ~n50103 ;
  assign y25041 = ~1'b0 ;
  assign y25042 = ~1'b0 ;
  assign y25043 = ~n50107 ;
  assign y25044 = ~1'b0 ;
  assign y25045 = ~1'b0 ;
  assign y25046 = n50108 ;
  assign y25047 = n50110 ;
  assign y25048 = ~1'b0 ;
  assign y25049 = n50111 ;
  assign y25050 = n50112 ;
  assign y25051 = n50116 ;
  assign y25052 = ~n50119 ;
  assign y25053 = ~1'b0 ;
  assign y25054 = ~1'b0 ;
  assign y25055 = n50120 ;
  assign y25056 = n50121 ;
  assign y25057 = ~n50122 ;
  assign y25058 = n50123 ;
  assign y25059 = ~n50126 ;
  assign y25060 = ~n50132 ;
  assign y25061 = ~1'b0 ;
  assign y25062 = ~1'b0 ;
  assign y25063 = ~n50135 ;
  assign y25064 = ~n50136 ;
  assign y25065 = ~n50137 ;
  assign y25066 = ~n50139 ;
  assign y25067 = n50140 ;
  assign y25068 = n50143 ;
  assign y25069 = n50144 ;
  assign y25070 = n50145 ;
  assign y25071 = ~n50146 ;
  assign y25072 = ~n50148 ;
  assign y25073 = ~n50153 ;
  assign y25074 = ~n50158 ;
  assign y25075 = ~n50162 ;
  assign y25076 = ~n50170 ;
  assign y25077 = ~1'b0 ;
  assign y25078 = ~1'b0 ;
  assign y25079 = n50171 ;
  assign y25080 = ~n50174 ;
  assign y25081 = ~n50177 ;
  assign y25082 = n50180 ;
  assign y25083 = ~1'b0 ;
  assign y25084 = ~1'b0 ;
  assign y25085 = ~n50182 ;
  assign y25086 = n50184 ;
  assign y25087 = ~n50187 ;
  assign y25088 = n50191 ;
  assign y25089 = n50193 ;
  assign y25090 = n50197 ;
  assign y25091 = ~n50200 ;
  assign y25092 = ~n50207 ;
  assign y25093 = ~n50211 ;
  assign y25094 = ~1'b0 ;
  assign y25095 = ~n50213 ;
  assign y25096 = ~n50214 ;
  assign y25097 = ~1'b0 ;
  assign y25098 = n50216 ;
  assign y25099 = ~n50218 ;
  assign y25100 = n50219 ;
  assign y25101 = ~1'b0 ;
  assign y25102 = ~1'b0 ;
  assign y25103 = n50221 ;
  assign y25104 = ~n50222 ;
  assign y25105 = ~n50226 ;
  assign y25106 = n50227 ;
  assign y25107 = ~1'b0 ;
  assign y25108 = ~n50229 ;
  assign y25109 = ~n50232 ;
  assign y25110 = n50236 ;
  assign y25111 = ~n6767 ;
  assign y25112 = n3792 ;
  assign y25113 = ~1'b0 ;
  assign y25114 = ~n50238 ;
  assign y25115 = ~1'b0 ;
  assign y25116 = n50239 ;
  assign y25117 = ~n50240 ;
  assign y25118 = ~n50242 ;
  assign y25119 = ~1'b0 ;
  assign y25120 = ~1'b0 ;
  assign y25121 = ~n50243 ;
  assign y25122 = ~n50245 ;
  assign y25123 = n50247 ;
  assign y25124 = ~n50252 ;
  assign y25125 = ~n50253 ;
  assign y25126 = ~n50258 ;
  assign y25127 = ~n50260 ;
  assign y25128 = n50262 ;
  assign y25129 = n34157 ;
  assign y25130 = ~n50264 ;
  assign y25131 = ~1'b0 ;
  assign y25132 = ~1'b0 ;
  assign y25133 = ~1'b0 ;
  assign y25134 = ~1'b0 ;
  assign y25135 = n50265 ;
  assign y25136 = n50266 ;
  assign y25137 = ~1'b0 ;
  assign y25138 = ~n18236 ;
  assign y25139 = ~1'b0 ;
  assign y25140 = ~n50272 ;
  assign y25141 = ~n50274 ;
  assign y25142 = ~n50278 ;
  assign y25143 = ~1'b0 ;
  assign y25144 = n50279 ;
  assign y25145 = ~1'b0 ;
  assign y25146 = n50283 ;
  assign y25147 = n50285 ;
  assign y25148 = ~n50289 ;
  assign y25149 = ~n16771 ;
  assign y25150 = ~1'b0 ;
  assign y25151 = ~n50292 ;
  assign y25152 = ~n50295 ;
  assign y25153 = n50298 ;
  assign y25154 = n50299 ;
  assign y25155 = ~n50300 ;
  assign y25156 = ~1'b0 ;
  assign y25157 = n50302 ;
  assign y25158 = ~n1105 ;
  assign y25159 = ~1'b0 ;
  assign y25160 = ~n22562 ;
  assign y25161 = ~n50304 ;
  assign y25162 = n50305 ;
  assign y25163 = n50306 ;
  assign y25164 = n50308 ;
  assign y25165 = n50314 ;
  assign y25166 = n50316 ;
  assign y25167 = n50317 ;
  assign y25168 = ~n50319 ;
  assign y25169 = n50325 ;
  assign y25170 = ~n50326 ;
  assign y25171 = ~n11998 ;
  assign y25172 = n50328 ;
  assign y25173 = ~n5303 ;
  assign y25174 = ~n50333 ;
  assign y25175 = n50335 ;
  assign y25176 = ~n50337 ;
  assign y25177 = ~n50339 ;
  assign y25178 = n50341 ;
  assign y25179 = ~1'b0 ;
  assign y25180 = n50342 ;
  assign y25181 = ~n9281 ;
  assign y25182 = ~n50352 ;
  assign y25183 = ~1'b0 ;
  assign y25184 = ~n50355 ;
  assign y25185 = n50364 ;
  assign y25186 = n50366 ;
  assign y25187 = ~n50371 ;
  assign y25188 = ~n50373 ;
  assign y25189 = ~n50375 ;
  assign y25190 = ~n50376 ;
  assign y25191 = ~1'b0 ;
  assign y25192 = ~1'b0 ;
  assign y25193 = ~1'b0 ;
  assign y25194 = ~n50381 ;
  assign y25195 = n50382 ;
  assign y25196 = n50387 ;
  assign y25197 = n50390 ;
  assign y25198 = ~n50391 ;
  assign y25199 = ~1'b0 ;
  assign y25200 = ~n50394 ;
  assign y25201 = ~n50397 ;
  assign y25202 = 1'b0 ;
  assign y25203 = ~1'b0 ;
  assign y25204 = ~1'b0 ;
  assign y25205 = n50401 ;
  assign y25206 = ~n50405 ;
  assign y25207 = ~n50407 ;
  assign y25208 = ~n50408 ;
  assign y25209 = n50412 ;
  assign y25210 = ~n50414 ;
  assign y25211 = n50416 ;
  assign y25212 = n50417 ;
  assign y25213 = ~n50418 ;
  assign y25214 = ~1'b0 ;
  assign y25215 = ~1'b0 ;
  assign y25216 = n50420 ;
  assign y25217 = n50425 ;
  assign y25218 = ~n50426 ;
  assign y25219 = n50427 ;
  assign y25220 = n50429 ;
  assign y25221 = ~1'b0 ;
  assign y25222 = ~n50434 ;
  assign y25223 = n17830 ;
  assign y25224 = ~1'b0 ;
  assign y25225 = ~1'b0 ;
  assign y25226 = n50438 ;
  assign y25227 = ~1'b0 ;
  assign y25228 = ~1'b0 ;
  assign y25229 = ~1'b0 ;
  assign y25230 = ~1'b0 ;
  assign y25231 = ~1'b0 ;
  assign y25232 = ~n20964 ;
  assign y25233 = n50440 ;
  assign y25234 = n50442 ;
  assign y25235 = n50443 ;
  assign y25236 = ~n50450 ;
  assign y25237 = n38357 ;
  assign y25238 = ~n50453 ;
  assign y25239 = n50455 ;
  assign y25240 = ~1'b0 ;
  assign y25241 = ~n50457 ;
  assign y25242 = ~n50463 ;
  assign y25243 = n50464 ;
  assign y25244 = ~n50465 ;
  assign y25245 = n50467 ;
  assign y25246 = n50469 ;
  assign y25247 = n50470 ;
  assign y25248 = n50471 ;
  assign y25249 = ~n50473 ;
  assign y25250 = ~1'b0 ;
  assign y25251 = n50474 ;
  assign y25252 = ~1'b0 ;
  assign y25253 = ~1'b0 ;
  assign y25254 = n50476 ;
  assign y25255 = ~1'b0 ;
  assign y25256 = ~n50479 ;
  assign y25257 = n50482 ;
  assign y25258 = ~1'b0 ;
  assign y25259 = n50486 ;
  assign y25260 = ~1'b0 ;
  assign y25261 = n50488 ;
  assign y25262 = ~1'b0 ;
  assign y25263 = ~1'b0 ;
  assign y25264 = ~n50490 ;
  assign y25265 = ~1'b0 ;
  assign y25266 = n50491 ;
  assign y25267 = ~n50496 ;
  assign y25268 = ~1'b0 ;
  assign y25269 = ~n50500 ;
  assign y25270 = ~n50503 ;
  assign y25271 = n43904 ;
  assign y25272 = ~n50504 ;
  assign y25273 = ~n37685 ;
  assign y25274 = n50508 ;
  assign y25275 = ~n50509 ;
  assign y25276 = ~n50511 ;
  assign y25277 = ~n50516 ;
  assign y25278 = ~1'b0 ;
  assign y25279 = ~1'b0 ;
  assign y25280 = ~n50518 ;
  assign y25281 = n50522 ;
  assign y25282 = n50524 ;
  assign y25283 = ~1'b0 ;
  assign y25284 = ~1'b0 ;
  assign y25285 = ~n50526 ;
  assign y25286 = n50529 ;
  assign y25287 = n50532 ;
  assign y25288 = n50533 ;
  assign y25289 = n50537 ;
  assign y25290 = ~n50538 ;
  assign y25291 = ~n50539 ;
  assign y25292 = 1'b0 ;
  assign y25293 = n34753 ;
  assign y25294 = ~n50540 ;
  assign y25295 = n50541 ;
  assign y25296 = n50542 ;
  assign y25297 = ~n50545 ;
  assign y25298 = ~1'b0 ;
  assign y25299 = n50547 ;
  assign y25300 = ~1'b0 ;
  assign y25301 = ~1'b0 ;
  assign y25302 = n50548 ;
  assign y25303 = ~n4694 ;
  assign y25304 = n50553 ;
  assign y25305 = n50556 ;
  assign y25306 = n50557 ;
  assign y25307 = n50559 ;
  assign y25308 = n50561 ;
  assign y25309 = n50562 ;
  assign y25310 = ~n50564 ;
  assign y25311 = ~n50565 ;
  assign y25312 = ~n50566 ;
  assign y25313 = n50569 ;
  assign y25314 = n50572 ;
  assign y25315 = n4126 ;
  assign y25316 = ~n50574 ;
  assign y25317 = n50578 ;
  assign y25318 = n50579 ;
  assign y25319 = ~1'b0 ;
  assign y25320 = ~n50582 ;
  assign y25321 = ~n50584 ;
  assign y25322 = n50588 ;
  assign y25323 = n50589 ;
  assign y25324 = ~1'b0 ;
  assign y25325 = ~n50591 ;
  assign y25326 = ~n50594 ;
  assign y25327 = ~n50595 ;
  assign y25328 = ~n50600 ;
  assign y25329 = n50605 ;
  assign y25330 = ~n50606 ;
  assign y25331 = ~n50608 ;
  assign y25332 = ~n50611 ;
  assign y25333 = n50612 ;
  assign y25334 = 1'b0 ;
  assign y25335 = ~1'b0 ;
  assign y25336 = 1'b0 ;
  assign y25337 = n50614 ;
  assign y25338 = n50617 ;
  assign y25339 = ~n50619 ;
  assign y25340 = ~1'b0 ;
  assign y25341 = n50621 ;
  assign y25342 = ~1'b0 ;
  assign y25343 = n50624 ;
  assign y25344 = ~n50626 ;
  assign y25345 = ~1'b0 ;
  assign y25346 = n50628 ;
  assign y25347 = ~n50629 ;
  assign y25348 = ~n50631 ;
  assign y25349 = ~1'b0 ;
  assign y25350 = n18726 ;
  assign y25351 = ~n50632 ;
  assign y25352 = ~1'b0 ;
  assign y25353 = ~n50633 ;
  assign y25354 = ~n50637 ;
  assign y25355 = n50641 ;
  assign y25356 = n50642 ;
  assign y25357 = ~n50643 ;
  assign y25358 = ~1'b0 ;
  assign y25359 = ~1'b0 ;
  assign y25360 = ~1'b0 ;
  assign y25361 = ~n50645 ;
  assign y25362 = n50648 ;
  assign y25363 = n50665 ;
  assign y25364 = ~n50666 ;
  assign y25365 = ~n50669 ;
  assign y25366 = ~n50674 ;
  assign y25367 = n50675 ;
  assign y25368 = n50680 ;
  assign y25369 = 1'b0 ;
  assign y25370 = ~n37673 ;
  assign y25371 = n50681 ;
  assign y25372 = n50682 ;
  assign y25373 = ~n50683 ;
  assign y25374 = ~n50684 ;
  assign y25375 = ~n50687 ;
  assign y25376 = ~1'b0 ;
  assign y25377 = ~n50688 ;
  assign y25378 = ~n50689 ;
  assign y25379 = ~n50692 ;
  assign y25380 = ~1'b0 ;
  assign y25381 = ~n50693 ;
  assign y25382 = ~n50695 ;
  assign y25383 = ~n50699 ;
  assign y25384 = n50700 ;
  assign y25385 = ~n50703 ;
  assign y25386 = ~n50705 ;
  assign y25387 = n50708 ;
  assign y25388 = ~n50711 ;
  assign y25389 = n50712 ;
  assign y25390 = ~n50713 ;
  assign y25391 = ~n50714 ;
  assign y25392 = n50716 ;
  assign y25393 = n50718 ;
  assign y25394 = ~n50721 ;
  assign y25395 = ~n50722 ;
  assign y25396 = ~n50725 ;
  assign y25397 = ~n50727 ;
  assign y25398 = n50729 ;
  assign y25399 = ~n50731 ;
  assign y25400 = n50732 ;
  assign y25401 = n50734 ;
  assign y25402 = ~1'b0 ;
  assign y25403 = ~n50736 ;
  assign y25404 = ~1'b0 ;
  assign y25405 = n50738 ;
  assign y25406 = n50739 ;
  assign y25407 = ~n50740 ;
  assign y25408 = n50741 ;
  assign y25409 = 1'b0 ;
  assign y25410 = ~n50744 ;
  assign y25411 = n50746 ;
  assign y25412 = n50748 ;
  assign y25413 = ~n50753 ;
  assign y25414 = ~n50755 ;
  assign y25415 = ~n50756 ;
  assign y25416 = n50757 ;
  assign y25417 = n50758 ;
  assign y25418 = n50759 ;
  assign y25419 = n50761 ;
  assign y25420 = ~n50765 ;
  assign y25421 = ~1'b0 ;
  assign y25422 = ~n50768 ;
  assign y25423 = ~n50771 ;
  assign y25424 = ~1'b0 ;
  assign y25425 = ~n50772 ;
  assign y25426 = n50780 ;
  assign y25427 = ~1'b0 ;
  assign y25428 = ~1'b0 ;
  assign y25429 = ~1'b0 ;
  assign y25430 = ~1'b0 ;
  assign y25431 = ~n50782 ;
  assign y25432 = ~1'b0 ;
  assign y25433 = n50785 ;
  assign y25434 = n50786 ;
  assign y25435 = ~n50787 ;
  assign y25436 = n50788 ;
  assign y25437 = ~1'b0 ;
  assign y25438 = n50791 ;
  assign y25439 = n50792 ;
  assign y25440 = ~n50793 ;
  assign y25441 = ~1'b0 ;
  assign y25442 = n50794 ;
  assign y25443 = n50796 ;
  assign y25444 = ~1'b0 ;
  assign y25445 = ~n31249 ;
  assign y25446 = n50798 ;
  assign y25447 = ~n50799 ;
  assign y25448 = ~1'b0 ;
  assign y25449 = ~n50803 ;
  assign y25450 = ~n50804 ;
  assign y25451 = ~n50806 ;
  assign y25452 = n4974 ;
  assign y25453 = ~1'b0 ;
  assign y25454 = ~n50808 ;
  assign y25455 = ~n50809 ;
  assign y25456 = ~n50812 ;
  assign y25457 = ~n50813 ;
  assign y25458 = ~n20830 ;
  assign y25459 = ~n50814 ;
  assign y25460 = n50818 ;
  assign y25461 = ~1'b0 ;
  assign y25462 = n50819 ;
  assign y25463 = n50820 ;
  assign y25464 = ~n50822 ;
  assign y25465 = n50824 ;
  assign y25466 = ~n50826 ;
  assign y25467 = n50829 ;
  assign y25468 = ~1'b0 ;
  assign y25469 = n50830 ;
  assign y25470 = n50834 ;
  assign y25471 = n1447 ;
  assign y25472 = ~1'b0 ;
  assign y25473 = n50837 ;
  assign y25474 = ~n50841 ;
  assign y25475 = ~n50842 ;
  assign y25476 = n50844 ;
  assign y25477 = ~n50845 ;
  assign y25478 = ~n50849 ;
  assign y25479 = ~n50853 ;
  assign y25480 = n50854 ;
  assign y25481 = ~1'b0 ;
  assign y25482 = ~1'b0 ;
  assign y25483 = ~1'b0 ;
  assign y25484 = ~n38051 ;
  assign y25485 = n50856 ;
  assign y25486 = ~n50857 ;
  assign y25487 = ~1'b0 ;
  assign y25488 = 1'b0 ;
  assign y25489 = ~1'b0 ;
  assign y25490 = ~1'b0 ;
  assign y25491 = ~1'b0 ;
  assign y25492 = n50860 ;
  assign y25493 = n50861 ;
  assign y25494 = n50863 ;
  assign y25495 = n50864 ;
  assign y25496 = ~n50865 ;
  assign y25497 = n50868 ;
  assign y25498 = ~n50869 ;
  assign y25499 = n19515 ;
  assign y25500 = ~n50870 ;
  assign y25501 = ~n50873 ;
  assign y25502 = ~1'b0 ;
  assign y25503 = ~n50876 ;
  assign y25504 = ~n50878 ;
  assign y25505 = ~1'b0 ;
  assign y25506 = ~1'b0 ;
  assign y25507 = ~n50879 ;
  assign y25508 = ~1'b0 ;
  assign y25509 = ~1'b0 ;
  assign y25510 = ~n50881 ;
  assign y25511 = n50882 ;
  assign y25512 = ~n40930 ;
  assign y25513 = ~n50883 ;
  assign y25514 = ~n50891 ;
  assign y25515 = n50894 ;
  assign y25516 = n50896 ;
  assign y25517 = ~1'b0 ;
  assign y25518 = 1'b0 ;
  assign y25519 = ~n41748 ;
  assign y25520 = ~1'b0 ;
  assign y25521 = ~n50897 ;
  assign y25522 = ~1'b0 ;
  assign y25523 = ~n50902 ;
  assign y25524 = ~n38522 ;
  assign y25525 = ~n50906 ;
  assign y25526 = ~n1668 ;
  assign y25527 = ~n50908 ;
  assign y25528 = n50909 ;
  assign y25529 = n48 ;
  assign y25530 = ~1'b0 ;
  assign y25531 = ~1'b0 ;
  assign y25532 = ~n50910 ;
  assign y25533 = n4884 ;
  assign y25534 = ~1'b0 ;
  assign y25535 = ~1'b0 ;
  assign y25536 = ~n50912 ;
  assign y25537 = ~1'b0 ;
  assign y25538 = 1'b0 ;
  assign y25539 = ~1'b0 ;
  assign y25540 = ~1'b0 ;
  assign y25541 = ~1'b0 ;
  assign y25542 = n50916 ;
  assign y25543 = n50918 ;
  assign y25544 = ~n50922 ;
  assign y25545 = ~n50926 ;
  assign y25546 = n50928 ;
  assign y25547 = ~n50930 ;
  assign y25548 = ~1'b0 ;
  assign y25549 = ~n50932 ;
  assign y25550 = n50933 ;
  assign y25551 = ~n37549 ;
  assign y25552 = ~n50935 ;
  assign y25553 = ~n50936 ;
  assign y25554 = ~n50937 ;
  assign y25555 = ~n50941 ;
  assign y25556 = ~1'b0 ;
  assign y25557 = ~n24161 ;
  assign y25558 = ~1'b0 ;
  assign y25559 = ~1'b0 ;
  assign y25560 = n50943 ;
  assign y25561 = 1'b0 ;
  assign y25562 = n50946 ;
  assign y25563 = n50947 ;
  assign y25564 = ~n50954 ;
  assign y25565 = ~1'b0 ;
  assign y25566 = ~n50958 ;
  assign y25567 = ~1'b0 ;
  assign y25568 = ~1'b0 ;
  assign y25569 = ~n50960 ;
  assign y25570 = n50961 ;
  assign y25571 = n50965 ;
  assign y25572 = ~n50966 ;
  assign y25573 = n50967 ;
  assign y25574 = ~n50969 ;
  assign y25575 = ~1'b0 ;
  assign y25576 = n50971 ;
  assign y25577 = n10903 ;
  assign y25578 = ~n50973 ;
  assign y25579 = n50980 ;
  assign y25580 = n50982 ;
  assign y25581 = ~n50983 ;
  assign y25582 = ~n50984 ;
  assign y25583 = ~n50987 ;
  assign y25584 = ~n50988 ;
  assign y25585 = ~n50989 ;
  assign y25586 = n50991 ;
  assign y25587 = ~n51004 ;
  assign y25588 = ~n51009 ;
  assign y25589 = n51016 ;
  assign y25590 = ~n51017 ;
  assign y25591 = ~1'b0 ;
  assign y25592 = ~1'b0 ;
  assign y25593 = n51018 ;
  assign y25594 = ~n6305 ;
  assign y25595 = ~n51019 ;
  assign y25596 = ~n51020 ;
  assign y25597 = ~1'b0 ;
  assign y25598 = n2441 ;
  assign y25599 = n51025 ;
  assign y25600 = ~n42771 ;
  assign y25601 = ~n51026 ;
  assign y25602 = n51027 ;
  assign y25603 = ~1'b0 ;
  assign y25604 = ~1'b0 ;
  assign y25605 = ~1'b0 ;
  assign y25606 = ~n14433 ;
  assign y25607 = ~1'b0 ;
  assign y25608 = 1'b0 ;
  assign y25609 = n51030 ;
  assign y25610 = n51034 ;
  assign y25611 = n51035 ;
  assign y25612 = n51036 ;
  assign y25613 = n51037 ;
  assign y25614 = ~n51042 ;
  assign y25615 = ~1'b0 ;
  assign y25616 = n51043 ;
  assign y25617 = ~n51045 ;
  assign y25618 = n51048 ;
  assign y25619 = ~n51050 ;
  assign y25620 = n51055 ;
  assign y25621 = ~1'b0 ;
  assign y25622 = ~1'b0 ;
  assign y25623 = ~n51059 ;
  assign y25624 = ~1'b0 ;
  assign y25625 = ~n51061 ;
  assign y25626 = ~n51063 ;
  assign y25627 = ~1'b0 ;
  assign y25628 = ~n51064 ;
  assign y25629 = n10975 ;
  assign y25630 = ~1'b0 ;
  assign y25631 = ~1'b0 ;
  assign y25632 = ~n36771 ;
  assign y25633 = ~n51066 ;
  assign y25634 = n51069 ;
  assign y25635 = n51072 ;
  assign y25636 = ~n51075 ;
  assign y25637 = n51076 ;
  assign y25638 = ~n51079 ;
  assign y25639 = n51081 ;
  assign y25640 = ~1'b0 ;
  assign y25641 = ~n51083 ;
  assign y25642 = ~n51084 ;
  assign y25643 = ~1'b0 ;
  assign y25644 = n51088 ;
  assign y25645 = n51090 ;
  assign y25646 = n51092 ;
  assign y25647 = ~1'b0 ;
  assign y25648 = ~1'b0 ;
  assign y25649 = ~n51095 ;
  assign y25650 = ~n51098 ;
  assign y25651 = ~n51099 ;
  assign y25652 = ~n51102 ;
  assign y25653 = n51105 ;
  assign y25654 = n51109 ;
  assign y25655 = ~n51110 ;
  assign y25656 = ~n51112 ;
  assign y25657 = ~1'b0 ;
  assign y25658 = ~1'b0 ;
  assign y25659 = ~1'b0 ;
  assign y25660 = ~n51113 ;
  assign y25661 = ~1'b0 ;
  assign y25662 = ~n51114 ;
  assign y25663 = ~n51122 ;
  assign y25664 = ~n4867 ;
  assign y25665 = n51123 ;
  assign y25666 = ~n51125 ;
  assign y25667 = ~1'b0 ;
  assign y25668 = ~1'b0 ;
  assign y25669 = ~n51127 ;
  assign y25670 = ~1'b0 ;
  assign y25671 = ~n51129 ;
  assign y25672 = ~n51131 ;
  assign y25673 = ~n51141 ;
  assign y25674 = n51144 ;
  assign y25675 = ~n51145 ;
  assign y25676 = 1'b0 ;
  assign y25677 = ~n51147 ;
  assign y25678 = n51150 ;
  assign y25679 = n32 ;
  assign y25680 = ~1'b0 ;
  assign y25681 = ~1'b0 ;
  assign y25682 = ~1'b0 ;
  assign y25683 = ~n51153 ;
  assign y25684 = n51155 ;
  assign y25685 = ~n51157 ;
  assign y25686 = n51160 ;
  assign y25687 = ~1'b0 ;
  assign y25688 = n51165 ;
  assign y25689 = n3782 ;
  assign y25690 = n51168 ;
  assign y25691 = ~1'b0 ;
  assign y25692 = n51170 ;
  assign y25693 = ~1'b0 ;
  assign y25694 = n51171 ;
  assign y25695 = ~1'b0 ;
  assign y25696 = ~1'b0 ;
  assign y25697 = ~1'b0 ;
  assign y25698 = ~n51173 ;
  assign y25699 = ~n51174 ;
  assign y25700 = ~1'b0 ;
  assign y25701 = ~n51182 ;
  assign y25702 = n51186 ;
  assign y25703 = n51188 ;
  assign y25704 = ~n51191 ;
  assign y25705 = ~n51196 ;
  assign y25706 = n51198 ;
  assign y25707 = ~1'b0 ;
  assign y25708 = ~n51199 ;
  assign y25709 = ~1'b0 ;
  assign y25710 = n51203 ;
  assign y25711 = ~n51205 ;
  assign y25712 = ~n51206 ;
  assign y25713 = ~n51207 ;
  assign y25714 = ~n51209 ;
  assign y25715 = ~n51212 ;
  assign y25716 = ~1'b0 ;
  assign y25717 = ~n51214 ;
  assign y25718 = n14858 ;
  assign y25719 = n51215 ;
  assign y25720 = n51217 ;
  assign y25721 = ~1'b0 ;
  assign y25722 = n51220 ;
  assign y25723 = n35687 ;
  assign y25724 = ~1'b0 ;
  assign y25725 = ~n51224 ;
  assign y25726 = n51225 ;
  assign y25727 = n51227 ;
  assign y25728 = ~n51231 ;
  assign y25729 = ~1'b0 ;
  assign y25730 = ~n51235 ;
  assign y25731 = n51238 ;
  assign y25732 = ~n51241 ;
  assign y25733 = n51245 ;
  assign y25734 = n51248 ;
  assign y25735 = ~1'b0 ;
  assign y25736 = ~n51249 ;
  assign y25737 = n51250 ;
  assign y25738 = ~n51253 ;
  assign y25739 = ~n51254 ;
  assign y25740 = n51259 ;
  assign y25741 = ~n51262 ;
  assign y25742 = ~1'b0 ;
  assign y25743 = ~n51263 ;
  assign y25744 = ~n51267 ;
  assign y25745 = ~n51270 ;
  assign y25746 = ~1'b0 ;
  assign y25747 = n51272 ;
  assign y25748 = ~n51274 ;
  assign y25749 = n51275 ;
  assign y25750 = ~n51277 ;
  assign y25751 = ~1'b0 ;
  assign y25752 = ~1'b0 ;
  assign y25753 = ~1'b0 ;
  assign y25754 = n51279 ;
  assign y25755 = ~1'b0 ;
  assign y25756 = n51281 ;
  assign y25757 = ~n51283 ;
  assign y25758 = n51286 ;
  assign y25759 = ~n51287 ;
  assign y25760 = ~1'b0 ;
  assign y25761 = n51288 ;
  assign y25762 = ~n51290 ;
  assign y25763 = ~1'b0 ;
  assign y25764 = ~1'b0 ;
  assign y25765 = ~1'b0 ;
  assign y25766 = n51291 ;
  assign y25767 = n51296 ;
  assign y25768 = n51299 ;
  assign y25769 = ~n50493 ;
  assign y25770 = 1'b0 ;
  assign y25771 = ~1'b0 ;
  assign y25772 = ~n51300 ;
  assign y25773 = ~1'b0 ;
  assign y25774 = ~n51301 ;
  assign y25775 = ~n51303 ;
  assign y25776 = n51305 ;
  assign y25777 = ~n51310 ;
  assign y25778 = ~1'b0 ;
  assign y25779 = ~n51312 ;
  assign y25780 = ~1'b0 ;
  assign y25781 = ~n51313 ;
  assign y25782 = n51314 ;
  assign y25783 = ~n51317 ;
  assign y25784 = ~n51319 ;
  assign y25785 = n51320 ;
  assign y25786 = ~1'b0 ;
  assign y25787 = n51323 ;
  assign y25788 = n12200 ;
  assign y25789 = ~1'b0 ;
  assign y25790 = ~1'b0 ;
  assign y25791 = ~1'b0 ;
  assign y25792 = ~n51325 ;
  assign y25793 = ~n51327 ;
  assign y25794 = ~1'b0 ;
  assign y25795 = ~n51330 ;
  assign y25796 = ~n51332 ;
  assign y25797 = n51337 ;
  assign y25798 = n51338 ;
  assign y25799 = n51340 ;
  assign y25800 = ~1'b0 ;
  assign y25801 = ~1'b0 ;
  assign y25802 = n51343 ;
  assign y25803 = n51346 ;
  assign y25804 = ~n51347 ;
  assign y25805 = ~n51349 ;
  assign y25806 = ~1'b0 ;
  assign y25807 = ~n51350 ;
  assign y25808 = ~n51352 ;
  assign y25809 = ~1'b0 ;
  assign y25810 = ~n51355 ;
  assign y25811 = n51359 ;
  assign y25812 = n51362 ;
  assign y25813 = ~n51363 ;
  assign y25814 = n51367 ;
  assign y25815 = n25391 ;
  assign y25816 = ~n51368 ;
  assign y25817 = n51373 ;
  assign y25818 = ~n31050 ;
  assign y25819 = ~n51377 ;
  assign y25820 = n17599 ;
  assign y25821 = ~1'b0 ;
  assign y25822 = ~1'b0 ;
  assign y25823 = n35496 ;
  assign y25824 = n51378 ;
  assign y25825 = ~n51380 ;
  assign y25826 = ~1'b0 ;
  assign y25827 = ~n51381 ;
  assign y25828 = ~1'b0 ;
  assign y25829 = ~n51387 ;
  assign y25830 = ~1'b0 ;
  assign y25831 = ~n51391 ;
  assign y25832 = n51393 ;
  assign y25833 = ~n51396 ;
  assign y25834 = n51402 ;
  assign y25835 = ~1'b0 ;
  assign y25836 = n51406 ;
  assign y25837 = n51410 ;
  assign y25838 = n51411 ;
  assign y25839 = n51417 ;
  assign y25840 = ~1'b0 ;
  assign y25841 = ~n51421 ;
  assign y25842 = n51424 ;
  assign y25843 = n51425 ;
  assign y25844 = ~1'b0 ;
  assign y25845 = ~1'b0 ;
  assign y25846 = ~1'b0 ;
  assign y25847 = n51426 ;
  assign y25848 = ~1'b0 ;
  assign y25849 = n51430 ;
  assign y25850 = n51432 ;
  assign y25851 = ~n51433 ;
  assign y25852 = 1'b0 ;
  assign y25853 = ~n51437 ;
  assign y25854 = ~n51438 ;
  assign y25855 = n9437 ;
  assign y25856 = n51442 ;
  assign y25857 = ~1'b0 ;
  assign y25858 = ~1'b0 ;
  assign y25859 = ~n51445 ;
  assign y25860 = n51449 ;
  assign y25861 = ~1'b0 ;
  assign y25862 = ~1'b0 ;
  assign y25863 = n51450 ;
  assign y25864 = ~n51451 ;
  assign y25865 = n2606 ;
  assign y25866 = n51452 ;
  assign y25867 = ~n51453 ;
  assign y25868 = n51455 ;
  assign y25869 = ~1'b0 ;
  assign y25870 = ~n51460 ;
  assign y25871 = n10228 ;
  assign y25872 = ~n27691 ;
  assign y25873 = ~n51462 ;
  assign y25874 = ~1'b0 ;
  assign y25875 = ~n51466 ;
  assign y25876 = ~n51468 ;
  assign y25877 = 1'b0 ;
  assign y25878 = ~n51470 ;
  assign y25879 = n51473 ;
  assign y25880 = n51474 ;
  assign y25881 = ~n51475 ;
  assign y25882 = ~n51476 ;
  assign y25883 = ~1'b0 ;
  assign y25884 = ~n51479 ;
  assign y25885 = n51480 ;
  assign y25886 = 1'b0 ;
  assign y25887 = n51483 ;
  assign y25888 = ~1'b0 ;
  assign y25889 = ~n51484 ;
  assign y25890 = n51487 ;
  assign y25891 = ~n51488 ;
  assign y25892 = ~n51490 ;
  assign y25893 = n51491 ;
  assign y25894 = ~1'b0 ;
  assign y25895 = ~n51493 ;
  assign y25896 = ~1'b0 ;
  assign y25897 = ~1'b0 ;
  assign y25898 = ~n51494 ;
  assign y25899 = n51495 ;
  assign y25900 = 1'b0 ;
  assign y25901 = n51498 ;
  assign y25902 = ~n51500 ;
  assign y25903 = ~n51501 ;
  assign y25904 = ~n51502 ;
  assign y25905 = n51503 ;
  assign y25906 = ~1'b0 ;
  assign y25907 = ~n51506 ;
  assign y25908 = ~1'b0 ;
  assign y25909 = ~1'b0 ;
  assign y25910 = ~n51507 ;
  assign y25911 = ~1'b0 ;
  assign y25912 = n12754 ;
  assign y25913 = n51508 ;
  assign y25914 = ~1'b0 ;
  assign y25915 = ~n51510 ;
  assign y25916 = n51511 ;
  assign y25917 = ~1'b0 ;
  assign y25918 = ~1'b0 ;
  assign y25919 = ~1'b0 ;
  assign y25920 = n3013 ;
  assign y25921 = ~n51515 ;
  assign y25922 = ~n51516 ;
  assign y25923 = ~n51519 ;
  assign y25924 = n51520 ;
  assign y25925 = n51521 ;
  assign y25926 = ~1'b0 ;
  assign y25927 = n51523 ;
  assign y25928 = ~n51527 ;
  assign y25929 = ~1'b0 ;
  assign y25930 = ~n51528 ;
  assign y25931 = ~1'b0 ;
  assign y25932 = ~n10068 ;
  assign y25933 = n51532 ;
  assign y25934 = n51535 ;
  assign y25935 = ~n7380 ;
  assign y25936 = n42835 ;
  assign y25937 = n51538 ;
  assign y25938 = n51544 ;
  assign y25939 = ~1'b0 ;
  assign y25940 = ~1'b0 ;
  assign y25941 = n51546 ;
  assign y25942 = ~n51547 ;
  assign y25943 = n51551 ;
  assign y25944 = n51552 ;
  assign y25945 = ~1'b0 ;
  assign y25946 = n51553 ;
  assign y25947 = n51554 ;
  assign y25948 = ~n51558 ;
  assign y25949 = ~n51561 ;
  assign y25950 = n51562 ;
  assign y25951 = ~n51571 ;
  assign y25952 = ~1'b0 ;
  assign y25953 = n51573 ;
  assign y25954 = n51579 ;
  assign y25955 = ~1'b0 ;
  assign y25956 = ~1'b0 ;
  assign y25957 = n51582 ;
  assign y25958 = n51586 ;
  assign y25959 = n51588 ;
  assign y25960 = n51590 ;
  assign y25961 = ~n51593 ;
  assign y25962 = ~n51597 ;
  assign y25963 = ~n51599 ;
  assign y25964 = n51601 ;
  assign y25965 = ~1'b0 ;
  assign y25966 = ~n51603 ;
  assign y25967 = ~1'b0 ;
  assign y25968 = n51608 ;
  assign y25969 = ~n51611 ;
  assign y25970 = ~n51617 ;
  assign y25971 = n51620 ;
  assign y25972 = n51621 ;
  assign y25973 = n51622 ;
  assign y25974 = ~n51623 ;
  assign y25975 = ~1'b0 ;
  assign y25976 = ~n51624 ;
  assign y25977 = n51626 ;
  assign y25978 = ~n51628 ;
  assign y25979 = n51631 ;
  assign y25980 = n51632 ;
  assign y25981 = n51634 ;
  assign y25982 = ~1'b0 ;
  assign y25983 = n51635 ;
  assign y25984 = n51637 ;
  assign y25985 = ~n51638 ;
  assign y25986 = n51639 ;
  assign y25987 = n51644 ;
  assign y25988 = n51646 ;
  assign y25989 = ~1'b0 ;
  assign y25990 = n51647 ;
  assign y25991 = ~n51650 ;
  assign y25992 = n51651 ;
  assign y25993 = ~1'b0 ;
  assign y25994 = ~n51653 ;
  assign y25995 = ~1'b0 ;
  assign y25996 = ~1'b0 ;
  assign y25997 = ~n51656 ;
  assign y25998 = ~n51659 ;
  assign y25999 = ~n51662 ;
  assign y26000 = ~n51664 ;
  assign y26001 = ~1'b0 ;
  assign y26002 = ~n51665 ;
  assign y26003 = ~n51666 ;
  assign y26004 = ~n51667 ;
  assign y26005 = ~1'b0 ;
  assign y26006 = ~1'b0 ;
  assign y26007 = ~1'b0 ;
  assign y26008 = ~1'b0 ;
  assign y26009 = n51669 ;
  assign y26010 = n51673 ;
  assign y26011 = ~1'b0 ;
  assign y26012 = ~1'b0 ;
  assign y26013 = ~n51676 ;
  assign y26014 = ~n51678 ;
  assign y26015 = ~n51683 ;
  assign y26016 = ~1'b0 ;
  assign y26017 = n11304 ;
  assign y26018 = ~1'b0 ;
  assign y26019 = ~1'b0 ;
  assign y26020 = ~n51684 ;
  assign y26021 = n51686 ;
  assign y26022 = n51688 ;
  assign y26023 = n51689 ;
  assign y26024 = ~n51693 ;
  assign y26025 = ~n51694 ;
  assign y26026 = ~n51696 ;
  assign y26027 = ~1'b0 ;
  assign y26028 = n51698 ;
  assign y26029 = ~1'b0 ;
  assign y26030 = ~n43564 ;
  assign y26031 = ~n51699 ;
  assign y26032 = ~1'b0 ;
  assign y26033 = ~n51702 ;
  assign y26034 = ~1'b0 ;
  assign y26035 = ~n51703 ;
  assign y26036 = ~n51705 ;
  assign y26037 = ~n51707 ;
  assign y26038 = n51709 ;
  assign y26039 = n51717 ;
  assign y26040 = ~1'b0 ;
  assign y26041 = ~n51721 ;
  assign y26042 = n51728 ;
  assign y26043 = ~n51738 ;
  assign y26044 = ~n51741 ;
  assign y26045 = ~1'b0 ;
  assign y26046 = ~n51742 ;
  assign y26047 = n51743 ;
  assign y26048 = n51747 ;
  assign y26049 = n51748 ;
  assign y26050 = ~n51749 ;
  assign y26051 = n51752 ;
  assign y26052 = n51754 ;
  assign y26053 = n51759 ;
  assign y26054 = ~n51761 ;
  assign y26055 = 1'b0 ;
  assign y26056 = ~n51762 ;
  assign y26057 = n51763 ;
  assign y26058 = ~n51765 ;
  assign y26059 = ~n5372 ;
  assign y26060 = n51766 ;
  assign y26061 = ~n51767 ;
  assign y26062 = ~n51771 ;
  assign y26063 = n9517 ;
  assign y26064 = n51774 ;
  assign y26065 = ~n51776 ;
  assign y26066 = ~1'b0 ;
  assign y26067 = n51779 ;
  assign y26068 = n51782 ;
  assign y26069 = ~n51783 ;
  assign y26070 = ~n51784 ;
  assign y26071 = ~n51785 ;
  assign y26072 = n51787 ;
  assign y26073 = n51788 ;
  assign y26074 = ~n51790 ;
  assign y26075 = n51794 ;
  assign y26076 = ~n51796 ;
  assign y26077 = ~1'b0 ;
  assign y26078 = n51797 ;
  assign y26079 = ~1'b0 ;
  assign y26080 = n51800 ;
  assign y26081 = ~n32888 ;
  assign y26082 = ~n51801 ;
  assign y26083 = n51802 ;
  assign y26084 = ~1'b0 ;
  assign y26085 = ~1'b0 ;
  assign y26086 = ~1'b0 ;
  assign y26087 = ~1'b0 ;
  assign y26088 = ~1'b0 ;
  assign y26089 = 1'b0 ;
  assign y26090 = ~n51803 ;
  assign y26091 = ~1'b0 ;
  assign y26092 = ~n51804 ;
  assign y26093 = ~n51808 ;
  assign y26094 = n51809 ;
  assign y26095 = ~1'b0 ;
  assign y26096 = ~1'b0 ;
  assign y26097 = ~1'b0 ;
  assign y26098 = ~n51811 ;
  assign y26099 = ~1'b0 ;
  assign y26100 = n51813 ;
  assign y26101 = ~n51816 ;
  assign y26102 = ~n51817 ;
  assign y26103 = ~n51820 ;
  assign y26104 = n15708 ;
  assign y26105 = n51825 ;
  assign y26106 = n51828 ;
  assign y26107 = ~n51831 ;
  assign y26108 = ~n51832 ;
  assign y26109 = n51833 ;
  assign y26110 = n51835 ;
  assign y26111 = n51837 ;
  assign y26112 = n51842 ;
  assign y26113 = ~n45963 ;
  assign y26114 = n34041 ;
  assign y26115 = ~n51847 ;
  assign y26116 = ~n51848 ;
  assign y26117 = ~1'b0 ;
  assign y26118 = ~1'b0 ;
  assign y26119 = ~1'b0 ;
  assign y26120 = ~n51849 ;
  assign y26121 = n51850 ;
  assign y26122 = ~n51853 ;
  assign y26123 = n51858 ;
  assign y26124 = ~1'b0 ;
  assign y26125 = ~n51864 ;
  assign y26126 = n51866 ;
  assign y26127 = ~n51868 ;
  assign y26128 = n51871 ;
  assign y26129 = n51873 ;
  assign y26130 = n24896 ;
  assign y26131 = ~1'b0 ;
  assign y26132 = ~n51875 ;
  assign y26133 = ~n51880 ;
  assign y26134 = ~n51681 ;
  assign y26135 = ~n51882 ;
  assign y26136 = n15396 ;
  assign y26137 = ~n51886 ;
  assign y26138 = n511 ;
  assign y26139 = ~1'b0 ;
  assign y26140 = n51887 ;
  assign y26141 = ~1'b0 ;
  assign y26142 = n46282 ;
  assign y26143 = ~n51888 ;
  assign y26144 = n51889 ;
  assign y26145 = ~1'b0 ;
  assign y26146 = n51890 ;
  assign y26147 = ~n51892 ;
  assign y26148 = n51896 ;
  assign y26149 = ~n51898 ;
  assign y26150 = n51900 ;
  assign y26151 = ~1'b0 ;
  assign y26152 = ~n51903 ;
  assign y26153 = ~n51326 ;
  assign y26154 = n51905 ;
  assign y26155 = n51906 ;
  assign y26156 = ~n51907 ;
  assign y26157 = ~1'b0 ;
  assign y26158 = ~n28817 ;
  assign y26159 = ~1'b0 ;
  assign y26160 = n51917 ;
  assign y26161 = ~n50347 ;
  assign y26162 = ~n51920 ;
  assign y26163 = n5051 ;
  assign y26164 = ~n51924 ;
  assign y26165 = ~1'b0 ;
  assign y26166 = n51927 ;
  assign y26167 = ~n51930 ;
  assign y26168 = n51937 ;
  assign y26169 = n51941 ;
  assign y26170 = ~n51948 ;
  assign y26171 = ~n51950 ;
  assign y26172 = n51951 ;
  assign y26173 = n51952 ;
  assign y26174 = ~n51954 ;
  assign y26175 = n51956 ;
  assign y26176 = n51958 ;
  assign y26177 = ~1'b0 ;
  assign y26178 = 1'b0 ;
  assign y26179 = n51959 ;
  assign y26180 = ~n51964 ;
  assign y26181 = ~1'b0 ;
  assign y26182 = ~n51965 ;
  assign y26183 = ~1'b0 ;
  assign y26184 = ~n51967 ;
  assign y26185 = ~1'b0 ;
  assign y26186 = ~n51973 ;
  assign y26187 = n51975 ;
  assign y26188 = ~1'b0 ;
  assign y26189 = ~n51979 ;
  assign y26190 = ~n51983 ;
  assign y26191 = ~n51985 ;
  assign y26192 = n51988 ;
  assign y26193 = ~1'b0 ;
  assign y26194 = n51990 ;
  assign y26195 = ~1'b0 ;
  assign y26196 = n51991 ;
  assign y26197 = n51992 ;
  assign y26198 = n3255 ;
  assign y26199 = n51993 ;
  assign y26200 = ~1'b0 ;
  assign y26201 = ~n51994 ;
  assign y26202 = ~1'b0 ;
  assign y26203 = ~1'b0 ;
  assign y26204 = ~1'b0 ;
  assign y26205 = n22645 ;
  assign y26206 = ~n51996 ;
  assign y26207 = ~n51998 ;
  assign y26208 = ~n52004 ;
  assign y26209 = ~n52007 ;
  assign y26210 = n52008 ;
  assign y26211 = n31449 ;
  assign y26212 = ~n52010 ;
  assign y26213 = n52013 ;
  assign y26214 = ~n52018 ;
  assign y26215 = ~1'b0 ;
  assign y26216 = ~1'b0 ;
  assign y26217 = ~1'b0 ;
  assign y26218 = n52019 ;
  assign y26219 = n52020 ;
  assign y26220 = n52022 ;
  assign y26221 = ~1'b0 ;
  assign y26222 = ~n52025 ;
  assign y26223 = n52026 ;
  assign y26224 = ~1'b0 ;
  assign y26225 = n52028 ;
  assign y26226 = ~n52030 ;
  assign y26227 = ~n52031 ;
  assign y26228 = ~n52032 ;
  assign y26229 = n52033 ;
  assign y26230 = n52044 ;
  assign y26231 = n52046 ;
  assign y26232 = ~n52048 ;
  assign y26233 = ~n52054 ;
  assign y26234 = ~1'b0 ;
  assign y26235 = n52057 ;
  assign y26236 = ~n52059 ;
  assign y26237 = n52060 ;
  assign y26238 = ~n52062 ;
  assign y26239 = 1'b0 ;
  assign y26240 = ~n52064 ;
  assign y26241 = n52066 ;
  assign y26242 = ~n52068 ;
  assign y26243 = ~1'b0 ;
  assign y26244 = 1'b0 ;
  assign y26245 = n17830 ;
  assign y26246 = n52069 ;
  assign y26247 = ~n52070 ;
  assign y26248 = ~n10771 ;
  assign y26249 = n52072 ;
  assign y26250 = ~1'b0 ;
  assign y26251 = n52073 ;
  assign y26252 = n52074 ;
  assign y26253 = ~n52077 ;
  assign y26254 = ~n52078 ;
  assign y26255 = ~n52079 ;
  assign y26256 = ~n52080 ;
  assign y26257 = ~n52083 ;
  assign y26258 = ~n52085 ;
  assign y26259 = n52086 ;
  assign y26260 = ~n52088 ;
  assign y26261 = n52089 ;
  assign y26262 = ~n14411 ;
  assign y26263 = n52093 ;
  assign y26264 = ~1'b0 ;
  assign y26265 = ~n52094 ;
  assign y26266 = ~n52098 ;
  assign y26267 = ~n52101 ;
  assign y26268 = ~n52103 ;
  assign y26269 = ~n52109 ;
  assign y26270 = n52111 ;
  assign y26271 = n52112 ;
  assign y26272 = ~1'b0 ;
  assign y26273 = ~n52116 ;
  assign y26274 = n52120 ;
  assign y26275 = ~1'b0 ;
  assign y26276 = n52122 ;
  assign y26277 = ~n52123 ;
  assign y26278 = ~n52125 ;
  assign y26279 = ~1'b0 ;
  assign y26280 = n52128 ;
  assign y26281 = ~1'b0 ;
  assign y26282 = ~1'b0 ;
  assign y26283 = n52129 ;
  assign y26284 = n52132 ;
  assign y26285 = n52136 ;
  assign y26286 = ~1'b0 ;
  assign y26287 = ~n52137 ;
  assign y26288 = ~n52138 ;
  assign y26289 = n52142 ;
  assign y26290 = ~1'b0 ;
  assign y26291 = ~n52146 ;
  assign y26292 = ~n52148 ;
  assign y26293 = ~1'b0 ;
  assign y26294 = ~n52149 ;
  assign y26295 = n52151 ;
  assign y26296 = ~1'b0 ;
  assign y26297 = ~n52153 ;
  assign y26298 = ~n52154 ;
  assign y26299 = ~n52155 ;
  assign y26300 = ~n52157 ;
  assign y26301 = ~1'b0 ;
  assign y26302 = ~n52159 ;
  assign y26303 = ~n52162 ;
  assign y26304 = ~1'b0 ;
  assign y26305 = n52164 ;
  assign y26306 = n52169 ;
  assign y26307 = n52170 ;
  assign y26308 = n52172 ;
  assign y26309 = n52173 ;
  assign y26310 = n52175 ;
  assign y26311 = n52179 ;
  assign y26312 = n25301 ;
  assign y26313 = n52180 ;
  assign y26314 = n52181 ;
  assign y26315 = ~1'b0 ;
  assign y26316 = 1'b0 ;
  assign y26317 = ~1'b0 ;
  assign y26318 = ~n3751 ;
  assign y26319 = ~n52184 ;
  assign y26320 = n30164 ;
  assign y26321 = n52186 ;
  assign y26322 = ~1'b0 ;
  assign y26323 = n52187 ;
  assign y26324 = n52189 ;
  assign y26325 = n52191 ;
  assign y26326 = ~n52196 ;
  assign y26327 = ~n52199 ;
  assign y26328 = ~n52202 ;
  assign y26329 = ~n52204 ;
  assign y26330 = n52207 ;
  assign y26331 = ~1'b0 ;
  assign y26332 = n52209 ;
  assign y26333 = ~1'b0 ;
  assign y26334 = ~1'b0 ;
  assign y26335 = ~n52211 ;
  assign y26336 = ~n52216 ;
  assign y26337 = n52218 ;
  assign y26338 = ~n52221 ;
  assign y26339 = n52228 ;
  assign y26340 = n52230 ;
  assign y26341 = ~n52232 ;
  assign y26342 = ~n52234 ;
  assign y26343 = ~1'b0 ;
  assign y26344 = ~1'b0 ;
  assign y26345 = ~n52236 ;
  assign y26346 = ~1'b0 ;
  assign y26347 = n52238 ;
  assign y26348 = ~n52240 ;
  assign y26349 = n52242 ;
  assign y26350 = n52244 ;
  assign y26351 = n52246 ;
  assign y26352 = ~1'b0 ;
  assign y26353 = n52250 ;
  assign y26354 = ~n52253 ;
  assign y26355 = ~1'b0 ;
  assign y26356 = ~1'b0 ;
  assign y26357 = ~1'b0 ;
  assign y26358 = n52261 ;
  assign y26359 = ~n52264 ;
  assign y26360 = ~n52266 ;
  assign y26361 = n52270 ;
  assign y26362 = ~n52272 ;
  assign y26363 = ~n52273 ;
  assign y26364 = ~n52275 ;
  assign y26365 = ~n52280 ;
  assign y26366 = n52283 ;
  assign y26367 = ~1'b0 ;
  assign y26368 = ~n52285 ;
  assign y26369 = n52288 ;
  assign y26370 = ~n52289 ;
  assign y26371 = ~n52294 ;
  assign y26372 = n52295 ;
  assign y26373 = ~1'b0 ;
  assign y26374 = 1'b0 ;
  assign y26375 = n52297 ;
  assign y26376 = ~1'b0 ;
  assign y26377 = n52298 ;
  assign y26378 = ~1'b0 ;
  assign y26379 = n12249 ;
  assign y26380 = ~n52301 ;
  assign y26381 = n52302 ;
  assign y26382 = n52304 ;
  assign y26383 = ~n52307 ;
  assign y26384 = n52309 ;
  assign y26385 = ~n52313 ;
  assign y26386 = n52314 ;
  assign y26387 = n52318 ;
  assign y26388 = ~n52320 ;
  assign y26389 = n52323 ;
  assign y26390 = ~1'b0 ;
  assign y26391 = n52324 ;
  assign y26392 = 1'b0 ;
  assign y26393 = ~n52325 ;
  assign y26394 = ~1'b0 ;
  assign y26395 = ~n52326 ;
  assign y26396 = ~n52329 ;
  assign y26397 = ~n52331 ;
  assign y26398 = ~n52333 ;
  assign y26399 = ~n52334 ;
  assign y26400 = ~n52336 ;
  assign y26401 = n12955 ;
  assign y26402 = ~1'b0 ;
  assign y26403 = ~n52340 ;
  assign y26404 = ~1'b0 ;
  assign y26405 = ~n42212 ;
  assign y26406 = ~1'b0 ;
  assign y26407 = ~1'b0 ;
  assign y26408 = ~n52343 ;
  assign y26409 = ~n52344 ;
  assign y26410 = ~n52345 ;
  assign y26411 = ~n52347 ;
  assign y26412 = ~1'b0 ;
  assign y26413 = ~1'b0 ;
  assign y26414 = n52348 ;
  assign y26415 = n52351 ;
  assign y26416 = ~n52352 ;
  assign y26417 = ~n52355 ;
  assign y26418 = ~1'b0 ;
  assign y26419 = n52356 ;
  assign y26420 = ~n52363 ;
  assign y26421 = ~1'b0 ;
  assign y26422 = ~1'b0 ;
  assign y26423 = ~1'b0 ;
  assign y26424 = 1'b0 ;
  assign y26425 = ~1'b0 ;
  assign y26426 = ~1'b0 ;
  assign y26427 = ~1'b0 ;
  assign y26428 = n25283 ;
  assign y26429 = ~n52366 ;
  assign y26430 = ~n52374 ;
  assign y26431 = n52376 ;
  assign y26432 = ~1'b0 ;
  assign y26433 = ~n52378 ;
  assign y26434 = n52381 ;
  assign y26435 = ~1'b0 ;
  assign y26436 = ~1'b0 ;
  assign y26437 = n52383 ;
  assign y26438 = ~n52384 ;
  assign y26439 = n52386 ;
  assign y26440 = n52389 ;
  assign y26441 = ~n52394 ;
  assign y26442 = n52398 ;
  assign y26443 = ~1'b0 ;
  assign y26444 = ~n52401 ;
  assign y26445 = ~n52402 ;
  assign y26446 = ~1'b0 ;
  assign y26447 = n52405 ;
  assign y26448 = ~1'b0 ;
  assign y26449 = ~1'b0 ;
  assign y26450 = n52407 ;
  assign y26451 = n52412 ;
  assign y26452 = ~n52414 ;
  assign y26453 = n52415 ;
  assign y26454 = ~n52418 ;
  assign y26455 = ~1'b0 ;
  assign y26456 = n52419 ;
  assign y26457 = n52420 ;
  assign y26458 = ~n52421 ;
  assign y26459 = n1171 ;
  assign y26460 = ~1'b0 ;
  assign y26461 = n52422 ;
  assign y26462 = ~n52425 ;
  assign y26463 = ~n52427 ;
  assign y26464 = ~n52429 ;
  assign y26465 = ~n52432 ;
  assign y26466 = n52436 ;
  assign y26467 = n52440 ;
  assign y26468 = 1'b0 ;
  assign y26469 = n52442 ;
  assign y26470 = ~1'b0 ;
  assign y26471 = ~n20564 ;
  assign y26472 = ~n52443 ;
  assign y26473 = ~n52447 ;
  assign y26474 = n52448 ;
  assign y26475 = ~n52449 ;
  assign y26476 = ~1'b0 ;
  assign y26477 = ~n52451 ;
  assign y26478 = n52452 ;
  assign y26479 = ~n52454 ;
  assign y26480 = ~1'b0 ;
  assign y26481 = ~1'b0 ;
  assign y26482 = n52455 ;
  assign y26483 = n52457 ;
  assign y26484 = ~n52458 ;
  assign y26485 = ~1'b0 ;
  assign y26486 = ~1'b0 ;
  assign y26487 = n52462 ;
  assign y26488 = ~1'b0 ;
  assign y26489 = n52463 ;
  assign y26490 = n16825 ;
  assign y26491 = n52464 ;
  assign y26492 = ~n52466 ;
  assign y26493 = n52467 ;
  assign y26494 = ~n52470 ;
  assign y26495 = ~n52471 ;
  assign y26496 = ~1'b0 ;
  assign y26497 = n52474 ;
  assign y26498 = n52475 ;
  assign y26499 = ~1'b0 ;
  assign y26500 = ~n708 ;
  assign y26501 = n52476 ;
  assign y26502 = ~n52477 ;
  assign y26503 = ~n52478 ;
  assign y26504 = ~n52480 ;
  assign y26505 = n52487 ;
  assign y26506 = ~1'b0 ;
  assign y26507 = n52490 ;
  assign y26508 = ~1'b0 ;
  assign y26509 = ~n52493 ;
  assign y26510 = ~1'b0 ;
  assign y26511 = ~n52494 ;
  assign y26512 = ~1'b0 ;
  assign y26513 = n52495 ;
  assign y26514 = ~n3255 ;
  assign y26515 = ~1'b0 ;
  assign y26516 = n52498 ;
  assign y26517 = ~n52500 ;
  assign y26518 = ~1'b0 ;
  assign y26519 = n52504 ;
  assign y26520 = ~1'b0 ;
  assign y26521 = ~1'b0 ;
  assign y26522 = n52508 ;
  assign y26523 = n52509 ;
  assign y26524 = ~n52510 ;
  assign y26525 = ~n52513 ;
  assign y26526 = ~n52514 ;
  assign y26527 = n52517 ;
  assign y26528 = ~1'b0 ;
  assign y26529 = n52523 ;
  assign y26530 = n52524 ;
  assign y26531 = ~1'b0 ;
  assign y26532 = n52527 ;
  assign y26533 = n22596 ;
  assign y26534 = ~n52528 ;
  assign y26535 = ~1'b0 ;
  assign y26536 = ~n52530 ;
  assign y26537 = 1'b0 ;
  assign y26538 = ~n52541 ;
  assign y26539 = ~n52542 ;
  assign y26540 = 1'b0 ;
  assign y26541 = ~n52543 ;
  assign y26542 = n42434 ;
  assign y26543 = ~n52547 ;
  assign y26544 = n52548 ;
  assign y26545 = ~n52549 ;
  assign y26546 = ~n52551 ;
  assign y26547 = n52552 ;
  assign y26548 = ~n52554 ;
  assign y26549 = ~n18851 ;
  assign y26550 = ~1'b0 ;
  assign y26551 = ~n52556 ;
  assign y26552 = n52558 ;
  assign y26553 = ~1'b0 ;
  assign y26554 = n52559 ;
  assign y26555 = ~1'b0 ;
  assign y26556 = ~1'b0 ;
  assign y26557 = ~1'b0 ;
  assign y26558 = ~n52562 ;
  assign y26559 = n52568 ;
  assign y26560 = ~n52571 ;
  assign y26561 = n52573 ;
  assign y26562 = ~n52575 ;
  assign y26563 = ~1'b0 ;
  assign y26564 = n52577 ;
  assign y26565 = n52580 ;
  assign y26566 = ~1'b0 ;
  assign y26567 = ~n52584 ;
  assign y26568 = ~1'b0 ;
  assign y26569 = n52589 ;
  assign y26570 = ~n52595 ;
  assign y26571 = n52604 ;
  assign y26572 = ~n52608 ;
  assign y26573 = n32079 ;
  assign y26574 = ~n52612 ;
  assign y26575 = ~n52614 ;
  assign y26576 = ~n52616 ;
  assign y26577 = ~n52617 ;
  assign y26578 = ~n41310 ;
  assign y26579 = ~1'b0 ;
  assign y26580 = ~n11947 ;
  assign y26581 = n52619 ;
  assign y26582 = n52620 ;
  assign y26583 = n52621 ;
  assign y26584 = ~n52625 ;
  assign y26585 = ~n4803 ;
  assign y26586 = n52629 ;
  assign y26587 = n52631 ;
  assign y26588 = n52633 ;
  assign y26589 = ~1'b0 ;
  assign y26590 = ~n52634 ;
  assign y26591 = ~n52640 ;
  assign y26592 = ~1'b0 ;
  assign y26593 = n52642 ;
  assign y26594 = n52649 ;
  assign y26595 = n14114 ;
  assign y26596 = ~1'b0 ;
  assign y26597 = ~n52651 ;
  assign y26598 = ~1'b0 ;
  assign y26599 = ~n52655 ;
  assign y26600 = ~n52656 ;
  assign y26601 = ~n52657 ;
  assign y26602 = n52662 ;
  assign y26603 = n52667 ;
  assign y26604 = ~n52668 ;
  assign y26605 = ~n52670 ;
  assign y26606 = n52672 ;
  assign y26607 = ~1'b0 ;
  assign y26608 = n52675 ;
  assign y26609 = n52677 ;
  assign y26610 = n52679 ;
  assign y26611 = ~n52684 ;
  assign y26612 = n52686 ;
  assign y26613 = ~n52688 ;
  assign y26614 = ~n52689 ;
  assign y26615 = ~1'b0 ;
  assign y26616 = ~n52691 ;
  assign y26617 = ~n52696 ;
  assign y26618 = ~n52699 ;
  assign y26619 = n2992 ;
  assign y26620 = 1'b0 ;
  assign y26621 = ~1'b0 ;
  assign y26622 = ~1'b0 ;
  assign y26623 = n52700 ;
  assign y26624 = ~n52704 ;
  assign y26625 = ~n52705 ;
  assign y26626 = n27266 ;
  assign y26627 = ~1'b0 ;
  assign y26628 = ~n52709 ;
  assign y26629 = n52711 ;
  assign y26630 = n52712 ;
  assign y26631 = ~n52713 ;
  assign y26632 = n52714 ;
  assign y26633 = ~n52715 ;
  assign y26634 = n52716 ;
  assign y26635 = ~n52718 ;
  assign y26636 = ~1'b0 ;
  assign y26637 = ~n52720 ;
  assign y26638 = ~n52723 ;
  assign y26639 = ~n4511 ;
  assign y26640 = n52728 ;
  assign y26641 = n52732 ;
  assign y26642 = ~n52737 ;
  assign y26643 = ~n24820 ;
  assign y26644 = n52740 ;
  assign y26645 = ~n52743 ;
  assign y26646 = n52745 ;
  assign y26647 = n52747 ;
  assign y26648 = ~n52750 ;
  assign y26649 = n52754 ;
  assign y26650 = ~n52756 ;
  assign y26651 = ~n52757 ;
  assign y26652 = n52760 ;
  assign y26653 = ~n52762 ;
  assign y26654 = n52765 ;
  assign y26655 = n52768 ;
  assign y26656 = n52769 ;
  assign y26657 = ~1'b0 ;
  assign y26658 = n52771 ;
  assign y26659 = ~n52773 ;
  assign y26660 = ~n52777 ;
  assign y26661 = n52785 ;
  assign y26662 = ~1'b0 ;
  assign y26663 = ~1'b0 ;
  assign y26664 = ~1'b0 ;
  assign y26665 = n52789 ;
  assign y26666 = ~1'b0 ;
  assign y26667 = ~1'b0 ;
  assign y26668 = n52790 ;
  assign y26669 = ~n52791 ;
  assign y26670 = ~n52792 ;
  assign y26671 = ~n52793 ;
  assign y26672 = ~1'b0 ;
  assign y26673 = ~n52795 ;
  assign y26674 = n52797 ;
  assign y26675 = n52798 ;
  assign y26676 = n52799 ;
  assign y26677 = ~n52805 ;
  assign y26678 = ~n52806 ;
  assign y26679 = ~n52809 ;
  assign y26680 = ~n52810 ;
  assign y26681 = ~n52812 ;
  assign y26682 = ~n52813 ;
  assign y26683 = ~n52816 ;
  assign y26684 = ~n52818 ;
  assign y26685 = ~n52820 ;
  assign y26686 = n52822 ;
  assign y26687 = n52828 ;
  assign y26688 = ~n52829 ;
  assign y26689 = ~n52832 ;
  assign y26690 = n1204 ;
  assign y26691 = n52834 ;
  assign y26692 = ~n52837 ;
  assign y26693 = ~n52838 ;
  assign y26694 = n52842 ;
  assign y26695 = ~1'b0 ;
  assign y26696 = n52844 ;
  assign y26697 = n49901 ;
  assign y26698 = n52848 ;
  assign y26699 = n52852 ;
  assign y26700 = n52857 ;
  assign y26701 = ~n43085 ;
  assign y26702 = ~n52858 ;
  assign y26703 = n52860 ;
  assign y26704 = n52862 ;
  assign y26705 = ~1'b0 ;
  assign y26706 = n52863 ;
  assign y26707 = ~n52867 ;
  assign y26708 = ~n52871 ;
  assign y26709 = n52872 ;
  assign y26710 = n52874 ;
  assign y26711 = ~1'b0 ;
  assign y26712 = ~1'b0 ;
  assign y26713 = ~1'b0 ;
  assign y26714 = ~n19652 ;
  assign y26715 = ~1'b0 ;
  assign y26716 = n52875 ;
  assign y26717 = n52877 ;
  assign y26718 = ~1'b0 ;
  assign y26719 = n37523 ;
  assign y26720 = ~n52879 ;
  assign y26721 = n52883 ;
  assign y26722 = ~n52885 ;
  assign y26723 = ~1'b0 ;
  assign y26724 = ~n52887 ;
  assign y26725 = ~1'b0 ;
  assign y26726 = ~1'b0 ;
  assign y26727 = ~1'b0 ;
  assign y26728 = ~n52888 ;
  assign y26729 = ~n52889 ;
  assign y26730 = ~n52890 ;
  assign y26731 = ~n52894 ;
  assign y26732 = n52895 ;
  assign y26733 = ~n52897 ;
  assign y26734 = ~1'b0 ;
  assign y26735 = n52902 ;
  assign y26736 = ~1'b0 ;
  assign y26737 = n52903 ;
  assign y26738 = n52906 ;
  assign y26739 = ~n52907 ;
  assign y26740 = ~n52908 ;
  assign y26741 = 1'b0 ;
  assign y26742 = ~n52910 ;
  assign y26743 = ~1'b0 ;
  assign y26744 = n52911 ;
  assign y26745 = n52914 ;
  assign y26746 = ~n52916 ;
  assign y26747 = n52917 ;
  assign y26748 = n52918 ;
  assign y26749 = ~1'b0 ;
  assign y26750 = ~n52919 ;
  assign y26751 = ~n52920 ;
  assign y26752 = ~1'b0 ;
  assign y26753 = ~n52921 ;
  assign y26754 = n52922 ;
  assign y26755 = ~n52924 ;
  assign y26756 = ~n52927 ;
  assign y26757 = n52928 ;
  assign y26758 = n52929 ;
  assign y26759 = n52933 ;
  assign y26760 = n52934 ;
  assign y26761 = n27699 ;
  assign y26762 = ~n52940 ;
  assign y26763 = n52942 ;
  assign y26764 = ~1'b0 ;
  assign y26765 = n52945 ;
  assign y26766 = ~n52950 ;
  assign y26767 = ~1'b0 ;
  assign y26768 = n52953 ;
  assign y26769 = ~1'b0 ;
  assign y26770 = ~n52954 ;
  assign y26771 = ~n52955 ;
  assign y26772 = ~1'b0 ;
  assign y26773 = n52958 ;
  assign y26774 = ~1'b0 ;
  assign y26775 = ~1'b0 ;
  assign y26776 = ~1'b0 ;
  assign y26777 = ~n52960 ;
  assign y26778 = ~1'b0 ;
  assign y26779 = ~n52962 ;
  assign y26780 = n52965 ;
  assign y26781 = n7464 ;
  assign y26782 = n52966 ;
  assign y26783 = n52969 ;
  assign y26784 = ~n52970 ;
  assign y26785 = ~n52979 ;
  assign y26786 = ~n52985 ;
  assign y26787 = ~n52992 ;
  assign y26788 = n52993 ;
  assign y26789 = n52996 ;
  assign y26790 = ~1'b0 ;
  assign y26791 = n52998 ;
  assign y26792 = n53002 ;
  assign y26793 = ~n53009 ;
  assign y26794 = n53017 ;
  assign y26795 = ~1'b0 ;
  assign y26796 = 1'b0 ;
  assign y26797 = ~n53019 ;
  assign y26798 = ~1'b0 ;
  assign y26799 = n53020 ;
  assign y26800 = n53021 ;
  assign y26801 = ~n53023 ;
  assign y26802 = ~n53024 ;
  assign y26803 = ~n53025 ;
  assign y26804 = ~n53030 ;
  assign y26805 = n53031 ;
  assign y26806 = ~n53033 ;
  assign y26807 = ~1'b0 ;
  assign y26808 = ~1'b0 ;
  assign y26809 = n53037 ;
  assign y26810 = ~1'b0 ;
  assign y26811 = ~n53039 ;
  assign y26812 = ~n53040 ;
  assign y26813 = n53044 ;
  assign y26814 = ~n53046 ;
  assign y26815 = n53050 ;
  assign y26816 = ~1'b0 ;
  assign y26817 = ~n53053 ;
  assign y26818 = ~n53055 ;
  assign y26819 = ~1'b0 ;
  assign y26820 = ~n53060 ;
  assign y26821 = n53065 ;
  assign y26822 = n53066 ;
  assign y26823 = ~1'b0 ;
  assign y26824 = ~1'b0 ;
  assign y26825 = ~n27996 ;
  assign y26826 = ~1'b0 ;
  assign y26827 = ~1'b0 ;
  assign y26828 = ~1'b0 ;
  assign y26829 = ~n53069 ;
  assign y26830 = ~1'b0 ;
  assign y26831 = ~1'b0 ;
  assign y26832 = n53073 ;
  assign y26833 = ~n53074 ;
  assign y26834 = ~1'b0 ;
  assign y26835 = n53080 ;
  assign y26836 = n14179 ;
  assign y26837 = ~n48433 ;
  assign y26838 = n53081 ;
  assign y26839 = ~n53083 ;
  assign y26840 = ~1'b0 ;
  assign y26841 = n1840 ;
  assign y26842 = ~1'b0 ;
  assign y26843 = ~n53086 ;
  assign y26844 = ~1'b0 ;
  assign y26845 = ~n53087 ;
  assign y26846 = n53088 ;
  assign y26847 = n53092 ;
  assign y26848 = n53094 ;
  assign y26849 = n53095 ;
  assign y26850 = ~1'b0 ;
  assign y26851 = ~n53100 ;
  assign y26852 = n53103 ;
  assign y26853 = n53104 ;
  assign y26854 = n53105 ;
  assign y26855 = n36054 ;
  assign y26856 = ~n53109 ;
  assign y26857 = ~n53111 ;
  assign y26858 = ~n53115 ;
  assign y26859 = ~1'b0 ;
  assign y26860 = ~n53120 ;
  assign y26861 = n53122 ;
  assign y26862 = ~n2628 ;
  assign y26863 = n53123 ;
  assign y26864 = n53125 ;
  assign y26865 = n53127 ;
  assign y26866 = ~1'b0 ;
  assign y26867 = ~1'b0 ;
  assign y26868 = ~1'b0 ;
  assign y26869 = n53128 ;
  assign y26870 = ~n53130 ;
  assign y26871 = ~1'b0 ;
  assign y26872 = ~1'b0 ;
  assign y26873 = ~n53132 ;
  assign y26874 = n53141 ;
  assign y26875 = ~n9317 ;
  assign y26876 = ~1'b0 ;
  assign y26877 = n19254 ;
  assign y26878 = n53144 ;
  assign y26879 = ~1'b0 ;
  assign y26880 = ~n53145 ;
  assign y26881 = ~n53146 ;
  assign y26882 = ~n53148 ;
  assign y26883 = ~n53153 ;
  assign y26884 = ~n53154 ;
  assign y26885 = n53158 ;
  assign y26886 = n53160 ;
  assign y26887 = ~1'b0 ;
  assign y26888 = ~n53161 ;
  assign y26889 = ~n53166 ;
  assign y26890 = n53171 ;
  assign y26891 = ~n53175 ;
  assign y26892 = ~n53180 ;
  assign y26893 = ~1'b0 ;
  assign y26894 = ~n53185 ;
  assign y26895 = n15646 ;
  assign y26896 = ~n53198 ;
  assign y26897 = ~1'b0 ;
  assign y26898 = ~1'b0 ;
  assign y26899 = n53202 ;
  assign y26900 = ~n25952 ;
  assign y26901 = n14812 ;
  assign y26902 = 1'b0 ;
  assign y26903 = ~n53204 ;
  assign y26904 = n53208 ;
  assign y26905 = ~n53210 ;
  assign y26906 = n53212 ;
  assign y26907 = ~1'b0 ;
  assign y26908 = ~n53214 ;
  assign y26909 = ~n53215 ;
  assign y26910 = ~1'b0 ;
  assign y26911 = n53216 ;
  assign y26912 = ~n53217 ;
  assign y26913 = n52325 ;
  assign y26914 = ~n53221 ;
  assign y26915 = ~n53224 ;
  assign y26916 = n53225 ;
  assign y26917 = n53226 ;
  assign y26918 = ~n53227 ;
  assign y26919 = ~n53228 ;
  assign y26920 = ~1'b0 ;
  assign y26921 = ~1'b0 ;
  assign y26922 = n53231 ;
  assign y26923 = ~1'b0 ;
  assign y26924 = n53236 ;
  assign y26925 = ~n53237 ;
  assign y26926 = ~n53238 ;
  assign y26927 = n53239 ;
  assign y26928 = ~1'b0 ;
  assign y26929 = n3435 ;
  assign y26930 = ~n53241 ;
  assign y26931 = ~n53242 ;
  assign y26932 = ~n53243 ;
  assign y26933 = ~1'b0 ;
  assign y26934 = ~n53246 ;
  assign y26935 = n53247 ;
  assign y26936 = ~n28139 ;
  assign y26937 = ~n53248 ;
  assign y26938 = n53252 ;
  assign y26939 = n53253 ;
  assign y26940 = ~1'b0 ;
  assign y26941 = ~n53259 ;
  assign y26942 = ~1'b0 ;
  assign y26943 = n53261 ;
  assign y26944 = n53263 ;
  assign y26945 = n53265 ;
  assign y26946 = ~n53266 ;
  assign y26947 = ~n53267 ;
  assign y26948 = n53274 ;
  assign y26949 = ~1'b0 ;
  assign y26950 = n26064 ;
  assign y26951 = ~1'b0 ;
  assign y26952 = ~n53275 ;
  assign y26953 = ~1'b0 ;
  assign y26954 = 1'b0 ;
  assign y26955 = ~n53277 ;
  assign y26956 = ~n53285 ;
  assign y26957 = n53287 ;
  assign y26958 = n53289 ;
  assign y26959 = n53292 ;
  assign y26960 = n53297 ;
  assign y26961 = ~n53303 ;
  assign y26962 = 1'b0 ;
  assign y26963 = ~1'b0 ;
  assign y26964 = ~n53305 ;
  assign y26965 = n53306 ;
  assign y26966 = n53309 ;
  assign y26967 = ~n12275 ;
  assign y26968 = ~n53312 ;
  assign y26969 = ~n53318 ;
  assign y26970 = n53321 ;
  assign y26971 = ~1'b0 ;
  assign y26972 = n53327 ;
  assign y26973 = ~1'b0 ;
  assign y26974 = n53332 ;
  assign y26975 = ~n53333 ;
  assign y26976 = ~1'b0 ;
  assign y26977 = n53334 ;
  assign y26978 = ~n53336 ;
  assign y26979 = n53341 ;
  assign y26980 = ~1'b0 ;
  assign y26981 = ~n53345 ;
  assign y26982 = n53347 ;
  assign y26983 = ~1'b0 ;
  assign y26984 = n53351 ;
  assign y26985 = n53354 ;
  assign y26986 = ~n53357 ;
  assign y26987 = n53358 ;
  assign y26988 = n53360 ;
  assign y26989 = ~n7089 ;
  assign y26990 = ~1'b0 ;
  assign y26991 = ~n21391 ;
  assign y26992 = ~n53364 ;
  assign y26993 = ~1'b0 ;
  assign y26994 = n53365 ;
  assign y26995 = ~n17597 ;
  assign y26996 = n53367 ;
  assign y26997 = n53369 ;
  assign y26998 = n39576 ;
  assign y26999 = n53370 ;
  assign y27000 = ~1'b0 ;
  assign y27001 = ~n53372 ;
  assign y27002 = ~n53376 ;
  assign y27003 = n53379 ;
  assign y27004 = n53384 ;
  assign y27005 = n53386 ;
  assign y27006 = ~n53387 ;
  assign y27007 = ~1'b0 ;
  assign y27008 = ~n53388 ;
  assign y27009 = n53389 ;
  assign y27010 = ~n53390 ;
  assign y27011 = n40579 ;
  assign y27012 = n38172 ;
  assign y27013 = ~n53391 ;
  assign y27014 = n53392 ;
  assign y27015 = n53393 ;
  assign y27016 = n53395 ;
  assign y27017 = ~1'b0 ;
  assign y27018 = ~n53396 ;
  assign y27019 = ~n53399 ;
  assign y27020 = ~n53402 ;
  assign y27021 = ~n53409 ;
  assign y27022 = ~1'b0 ;
  assign y27023 = ~1'b0 ;
  assign y27024 = ~n53410 ;
  assign y27025 = n53412 ;
  assign y27026 = ~1'b0 ;
  assign y27027 = ~n7974 ;
  assign y27028 = n11109 ;
  assign y27029 = ~1'b0 ;
  assign y27030 = ~n53413 ;
  assign y27031 = n53414 ;
  assign y27032 = ~n53416 ;
  assign y27033 = n53418 ;
  assign y27034 = ~1'b0 ;
  assign y27035 = ~1'b0 ;
  assign y27036 = n53419 ;
  assign y27037 = n53420 ;
  assign y27038 = 1'b0 ;
  assign y27039 = ~1'b0 ;
  assign y27040 = n53421 ;
  assign y27041 = n53422 ;
  assign y27042 = n53423 ;
  assign y27043 = ~n53425 ;
  assign y27044 = ~n53427 ;
  assign y27045 = n53429 ;
  assign y27046 = ~1'b0 ;
  assign y27047 = n53431 ;
  assign y27048 = ~n5147 ;
  assign y27049 = ~1'b0 ;
  assign y27050 = n53433 ;
  assign y27051 = n53435 ;
  assign y27052 = ~n53438 ;
  assign y27053 = ~n53440 ;
  assign y27054 = ~n53442 ;
  assign y27055 = n17936 ;
  assign y27056 = ~n22336 ;
  assign y27057 = ~1'b0 ;
  assign y27058 = ~1'b0 ;
  assign y27059 = ~n53445 ;
  assign y27060 = n53451 ;
  assign y27061 = 1'b0 ;
  assign y27062 = n53456 ;
  assign y27063 = ~n53457 ;
  assign y27064 = n53462 ;
  assign y27065 = ~n53465 ;
  assign y27066 = n53467 ;
  assign y27067 = ~n13153 ;
  assign y27068 = n53470 ;
  assign y27069 = ~n53475 ;
  assign y27070 = n53477 ;
  assign y27071 = 1'b0 ;
  assign y27072 = n53478 ;
  assign y27073 = ~n53482 ;
  assign y27074 = ~n53486 ;
  assign y27075 = ~n53491 ;
  assign y27076 = ~n53493 ;
  assign y27077 = ~n53496 ;
  assign y27078 = ~n53497 ;
  assign y27079 = ~1'b0 ;
  assign y27080 = ~n53498 ;
  assign y27081 = n53500 ;
  assign y27082 = n53503 ;
  assign y27083 = ~1'b0 ;
  assign y27084 = ~n53504 ;
  assign y27085 = n53505 ;
  assign y27086 = ~n53508 ;
  assign y27087 = ~1'b0 ;
  assign y27088 = ~n53510 ;
  assign y27089 = n53515 ;
  assign y27090 = ~1'b0 ;
  assign y27091 = n53516 ;
  assign y27092 = n53518 ;
  assign y27093 = ~1'b0 ;
  assign y27094 = n53519 ;
  assign y27095 = ~n53523 ;
  assign y27096 = n53527 ;
  assign y27097 = ~n53528 ;
  assign y27098 = ~n53533 ;
  assign y27099 = n53534 ;
  assign y27100 = n53537 ;
  assign y27101 = n53542 ;
  assign y27102 = ~1'b0 ;
  assign y27103 = n33946 ;
  assign y27104 = ~n53544 ;
  assign y27105 = ~n53550 ;
  assign y27106 = ~n53552 ;
  assign y27107 = ~1'b0 ;
  assign y27108 = ~n53553 ;
  assign y27109 = ~n53555 ;
  assign y27110 = ~n53560 ;
  assign y27111 = ~1'b0 ;
  assign y27112 = ~n53564 ;
  assign y27113 = n53565 ;
  assign y27114 = n53566 ;
  assign y27115 = n53568 ;
  assign y27116 = n53575 ;
  assign y27117 = ~n53576 ;
  assign y27118 = ~1'b0 ;
  assign y27119 = ~1'b0 ;
  assign y27120 = ~n53578 ;
  assign y27121 = ~1'b0 ;
  assign y27122 = ~n53583 ;
  assign y27123 = ~n53584 ;
  assign y27124 = n53587 ;
  assign y27125 = n53588 ;
  assign y27126 = ~n53590 ;
  assign y27127 = ~n53593 ;
  assign y27128 = ~n53594 ;
  assign y27129 = ~n53596 ;
  assign y27130 = n53598 ;
  assign y27131 = ~n53600 ;
  assign y27132 = ~1'b0 ;
  assign y27133 = 1'b0 ;
  assign y27134 = ~n3574 ;
  assign y27135 = ~1'b0 ;
  assign y27136 = n53605 ;
  assign y27137 = ~n53606 ;
  assign y27138 = ~n53608 ;
  assign y27139 = n53610 ;
  assign y27140 = ~1'b0 ;
  assign y27141 = n53611 ;
  assign y27142 = n53612 ;
  assign y27143 = ~n53614 ;
  assign y27144 = ~1'b0 ;
  assign y27145 = n53616 ;
  assign y27146 = ~n53618 ;
  assign y27147 = n14926 ;
  assign y27148 = n53619 ;
  assign y27149 = n53621 ;
  assign y27150 = ~n24923 ;
  assign y27151 = n53623 ;
  assign y27152 = ~n53625 ;
  assign y27153 = ~n53627 ;
  assign y27154 = n53631 ;
  assign y27155 = ~1'b0 ;
  assign y27156 = ~n53633 ;
  assign y27157 = n53635 ;
  assign y27158 = n53636 ;
  assign y27159 = ~n53640 ;
  assign y27160 = ~n22084 ;
  assign y27161 = ~n53643 ;
  assign y27162 = n53644 ;
  assign y27163 = ~n53650 ;
  assign y27164 = n53653 ;
  assign y27165 = ~1'b0 ;
  assign y27166 = ~1'b0 ;
  assign y27167 = n53658 ;
  assign y27168 = n53662 ;
  assign y27169 = ~n53665 ;
  assign y27170 = ~n53667 ;
  assign y27171 = ~n53669 ;
  assign y27172 = ~1'b0 ;
  assign y27173 = n53670 ;
  assign y27174 = n53671 ;
  assign y27175 = n53673 ;
  assign y27176 = ~n53675 ;
  assign y27177 = n53676 ;
  assign y27178 = n53678 ;
  assign y27179 = n53679 ;
  assign y27180 = ~1'b0 ;
  assign y27181 = ~1'b0 ;
  assign y27182 = ~1'b0 ;
  assign y27183 = ~n53685 ;
  assign y27184 = n53688 ;
  assign y27185 = ~1'b0 ;
  assign y27186 = ~1'b0 ;
  assign y27187 = ~n53690 ;
  assign y27188 = ~n53691 ;
  assign y27189 = ~n53693 ;
  assign y27190 = ~n6161 ;
  assign y27191 = ~n53694 ;
  assign y27192 = n53696 ;
  assign y27193 = ~1'b0 ;
  assign y27194 = n53699 ;
  assign y27195 = ~1'b0 ;
  assign y27196 = ~n53701 ;
  assign y27197 = ~n53703 ;
  assign y27198 = ~1'b0 ;
  assign y27199 = n53704 ;
  assign y27200 = n53709 ;
  assign y27201 = n53710 ;
  assign y27202 = ~1'b0 ;
  assign y27203 = n53711 ;
  assign y27204 = ~n53714 ;
  assign y27205 = ~n53715 ;
  assign y27206 = n53719 ;
  assign y27207 = ~n53720 ;
  assign y27208 = n53722 ;
  assign y27209 = ~1'b0 ;
  assign y27210 = ~n53725 ;
  assign y27211 = ~n53727 ;
  assign y27212 = ~n53728 ;
  assign y27213 = ~1'b0 ;
  assign y27214 = ~1'b0 ;
  assign y27215 = n53730 ;
  assign y27216 = ~n47543 ;
  assign y27217 = ~1'b0 ;
  assign y27218 = n53731 ;
  assign y27219 = ~n53733 ;
  assign y27220 = ~1'b0 ;
  assign y27221 = ~n53734 ;
  assign y27222 = n53735 ;
  assign y27223 = ~n53740 ;
  assign y27224 = ~n53742 ;
  assign y27225 = ~1'b0 ;
  assign y27226 = ~n53746 ;
  assign y27227 = n53747 ;
  assign y27228 = n53751 ;
  assign y27229 = ~n53754 ;
  assign y27230 = n53757 ;
  assign y27231 = ~n53760 ;
  assign y27232 = ~n53762 ;
  assign y27233 = n53764 ;
  assign y27234 = n53765 ;
  assign y27235 = n45171 ;
  assign y27236 = ~n53768 ;
  assign y27237 = ~n53769 ;
  assign y27238 = ~n53770 ;
  assign y27239 = ~n53774 ;
  assign y27240 = ~n53778 ;
  assign y27241 = n53783 ;
  assign y27242 = n53784 ;
  assign y27243 = n53786 ;
  assign y27244 = ~n53796 ;
  assign y27245 = ~1'b0 ;
  assign y27246 = n53798 ;
  assign y27247 = ~n10180 ;
  assign y27248 = n53803 ;
  assign y27249 = n4761 ;
  assign y27250 = ~n53806 ;
  assign y27251 = ~1'b0 ;
  assign y27252 = ~n53809 ;
  assign y27253 = n9165 ;
  assign y27254 = ~n4086 ;
  assign y27255 = ~n53811 ;
  assign y27256 = n53813 ;
  assign y27257 = ~1'b0 ;
  assign y27258 = ~1'b0 ;
  assign y27259 = ~n53815 ;
  assign y27260 = ~n53816 ;
  assign y27261 = ~1'b0 ;
  assign y27262 = ~1'b0 ;
  assign y27263 = n15555 ;
  assign y27264 = ~n5218 ;
  assign y27265 = ~n53817 ;
  assign y27266 = ~n53821 ;
  assign y27267 = n53823 ;
  assign y27268 = ~n53825 ;
  assign y27269 = n53827 ;
  assign y27270 = n53832 ;
  assign y27271 = ~1'b0 ;
  assign y27272 = n53833 ;
  assign y27273 = n53834 ;
  assign y27274 = n53836 ;
  assign y27275 = ~n53837 ;
  assign y27276 = ~n53839 ;
  assign y27277 = ~1'b0 ;
  assign y27278 = ~1'b0 ;
  assign y27279 = n53840 ;
  assign y27280 = n53843 ;
  assign y27281 = ~1'b0 ;
  assign y27282 = ~1'b0 ;
  assign y27283 = n53844 ;
  assign y27284 = n53846 ;
  assign y27285 = ~n7841 ;
  assign y27286 = ~n53848 ;
  assign y27287 = ~n53850 ;
  assign y27288 = n53853 ;
  assign y27289 = ~1'b0 ;
  assign y27290 = ~1'b0 ;
  assign y27291 = n53854 ;
  assign y27292 = ~n18679 ;
  assign y27293 = n30631 ;
  assign y27294 = n53855 ;
  assign y27295 = n53856 ;
  assign y27296 = n53857 ;
  assign y27297 = ~n53859 ;
  assign y27298 = 1'b0 ;
  assign y27299 = n53861 ;
  assign y27300 = ~1'b0 ;
  assign y27301 = ~1'b0 ;
  assign y27302 = ~n53864 ;
  assign y27303 = ~n53868 ;
  assign y27304 = ~1'b0 ;
  assign y27305 = n53869 ;
  assign y27306 = ~n53870 ;
  assign y27307 = ~n45362 ;
  assign y27308 = ~1'b0 ;
  assign y27309 = ~1'b0 ;
  assign y27310 = ~n53872 ;
  assign y27311 = ~1'b0 ;
  assign y27312 = ~1'b0 ;
  assign y27313 = ~1'b0 ;
  assign y27314 = ~n53874 ;
  assign y27315 = n53877 ;
  assign y27316 = ~n53878 ;
  assign y27317 = ~n53879 ;
  assign y27318 = ~1'b0 ;
  assign y27319 = ~n53881 ;
  assign y27320 = ~n53882 ;
  assign y27321 = ~n53884 ;
  assign y27322 = n53885 ;
  assign y27323 = ~1'b0 ;
  assign y27324 = ~n53887 ;
  assign y27325 = n23825 ;
  assign y27326 = ~n53889 ;
  assign y27327 = n53893 ;
  assign y27328 = n53894 ;
  assign y27329 = ~1'b0 ;
  assign y27330 = n53898 ;
  assign y27331 = ~1'b0 ;
  assign y27332 = n53901 ;
  assign y27333 = ~n53903 ;
  assign y27334 = n53905 ;
  assign y27335 = ~1'b0 ;
  assign y27336 = ~n53908 ;
  assign y27337 = ~n53909 ;
  assign y27338 = ~n53911 ;
  assign y27339 = n1334 ;
  assign y27340 = ~1'b0 ;
  assign y27341 = ~n6846 ;
  assign y27342 = ~1'b0 ;
  assign y27343 = ~1'b0 ;
  assign y27344 = ~1'b0 ;
  assign y27345 = ~n53913 ;
  assign y27346 = n53916 ;
  assign y27347 = n53917 ;
  assign y27348 = n53919 ;
  assign y27349 = ~n53920 ;
  assign y27350 = ~1'b0 ;
  assign y27351 = n53927 ;
  assign y27352 = ~n53932 ;
  assign y27353 = n53934 ;
  assign y27354 = ~1'b0 ;
  assign y27355 = ~1'b0 ;
  assign y27356 = n53936 ;
  assign y27357 = ~n53939 ;
  assign y27358 = n53940 ;
  assign y27359 = n53946 ;
  assign y27360 = ~1'b0 ;
  assign y27361 = ~n53950 ;
  assign y27362 = ~n53954 ;
  assign y27363 = ~n53955 ;
  assign y27364 = ~n53956 ;
  assign y27365 = n53959 ;
  assign y27366 = ~n53961 ;
  assign y27367 = ~1'b0 ;
  assign y27368 = ~n53967 ;
  assign y27369 = ~n53970 ;
  assign y27370 = ~n53974 ;
  assign y27371 = ~n2382 ;
  assign y27372 = ~n53975 ;
  assign y27373 = ~n53976 ;
  assign y27374 = ~1'b0 ;
  assign y27375 = ~n53980 ;
  assign y27376 = ~n53982 ;
  assign y27377 = ~1'b0 ;
  assign y27378 = n2484 ;
  assign y27379 = ~n53983 ;
  assign y27380 = ~n53985 ;
  assign y27381 = n53990 ;
  assign y27382 = ~1'b0 ;
  assign y27383 = n53991 ;
  assign y27384 = n53993 ;
  assign y27385 = ~1'b0 ;
  assign y27386 = ~1'b0 ;
  assign y27387 = ~n53994 ;
  assign y27388 = ~n27623 ;
  assign y27389 = ~n54001 ;
  assign y27390 = ~n54005 ;
  assign y27391 = n54009 ;
  assign y27392 = ~n54010 ;
  assign y27393 = ~1'b0 ;
  assign y27394 = n54011 ;
  assign y27395 = ~n54013 ;
  assign y27396 = n54014 ;
  assign y27397 = n54016 ;
  assign y27398 = ~1'b0 ;
  assign y27399 = ~n54017 ;
  assign y27400 = ~1'b0 ;
  assign y27401 = n54019 ;
  assign y27402 = ~n54023 ;
  assign y27403 = n54027 ;
  assign y27404 = ~n54030 ;
  assign y27405 = n54031 ;
  assign y27406 = n54033 ;
  assign y27407 = n54034 ;
  assign y27408 = ~1'b0 ;
  assign y27409 = ~1'b0 ;
  assign y27410 = ~n54037 ;
  assign y27411 = n54038 ;
  assign y27412 = ~1'b0 ;
  assign y27413 = n54043 ;
  assign y27414 = n54044 ;
  assign y27415 = ~n54047 ;
  assign y27416 = ~n54048 ;
  assign y27417 = ~1'b0 ;
  assign y27418 = ~1'b0 ;
  assign y27419 = n54054 ;
  assign y27420 = ~n54059 ;
  assign y27421 = ~n54060 ;
  assign y27422 = ~1'b0 ;
  assign y27423 = n54061 ;
  assign y27424 = ~n54065 ;
  assign y27425 = n54066 ;
  assign y27426 = ~1'b0 ;
  assign y27427 = ~1'b0 ;
  assign y27428 = ~1'b0 ;
  assign y27429 = ~n13282 ;
  assign y27430 = ~n859 ;
  assign y27431 = ~n54068 ;
  assign y27432 = n54070 ;
  assign y27433 = n54072 ;
  assign y27434 = ~1'b0 ;
  assign y27435 = ~1'b0 ;
  assign y27436 = n54073 ;
  assign y27437 = n54075 ;
  assign y27438 = n54076 ;
  assign y27439 = ~1'b0 ;
  assign y27440 = ~n54078 ;
  assign y27441 = ~n54079 ;
  assign y27442 = ~n54081 ;
  assign y27443 = ~n54082 ;
  assign y27444 = n18024 ;
  assign y27445 = n54086 ;
  assign y27446 = n54088 ;
  assign y27447 = ~1'b0 ;
  assign y27448 = n4005 ;
  assign y27449 = n54089 ;
  assign y27450 = n54091 ;
  assign y27451 = ~n54096 ;
  assign y27452 = n54099 ;
  assign y27453 = n17224 ;
  assign y27454 = ~n54111 ;
  assign y27455 = ~n54112 ;
  assign y27456 = n54113 ;
  assign y27457 = n54114 ;
  assign y27458 = ~1'b0 ;
  assign y27459 = n54115 ;
  assign y27460 = n54117 ;
  assign y27461 = ~n54121 ;
  assign y27462 = ~n54125 ;
  assign y27463 = n54128 ;
  assign y27464 = n54132 ;
  assign y27465 = 1'b0 ;
  assign y27466 = ~n54134 ;
  assign y27467 = ~1'b0 ;
  assign y27468 = n54137 ;
  assign y27469 = ~1'b0 ;
  assign y27470 = ~n54139 ;
  assign y27471 = n54141 ;
  assign y27472 = ~n54144 ;
  assign y27473 = ~n42346 ;
  assign y27474 = n54147 ;
  assign y27475 = 1'b0 ;
  assign y27476 = n45845 ;
  assign y27477 = ~n54149 ;
  assign y27478 = ~1'b0 ;
  assign y27479 = ~1'b0 ;
  assign y27480 = ~1'b0 ;
  assign y27481 = ~n54154 ;
  assign y27482 = ~1'b0 ;
  assign y27483 = n54155 ;
  assign y27484 = n54159 ;
  assign y27485 = ~n54160 ;
  assign y27486 = ~1'b0 ;
  assign y27487 = ~1'b0 ;
  assign y27488 = 1'b0 ;
  assign y27489 = n31130 ;
  assign y27490 = n54161 ;
  assign y27491 = n54162 ;
  assign y27492 = ~n54164 ;
  assign y27493 = n54166 ;
  assign y27494 = ~n54168 ;
  assign y27495 = ~n54170 ;
  assign y27496 = ~n54174 ;
  assign y27497 = n54177 ;
  assign y27498 = ~n54180 ;
  assign y27499 = n54183 ;
  assign y27500 = ~n54186 ;
  assign y27501 = n54191 ;
  assign y27502 = ~n54194 ;
  assign y27503 = ~1'b0 ;
  assign y27504 = n54195 ;
  assign y27505 = n54196 ;
  assign y27506 = ~n54197 ;
  assign y27507 = ~n54199 ;
  assign y27508 = ~1'b0 ;
  assign y27509 = ~n54201 ;
  assign y27510 = ~1'b0 ;
  assign y27511 = ~1'b0 ;
  assign y27512 = ~n54203 ;
  assign y27513 = ~n54205 ;
  assign y27514 = ~n54206 ;
  assign y27515 = ~n54211 ;
  assign y27516 = ~n54212 ;
  assign y27517 = n54214 ;
  assign y27518 = ~n26979 ;
  assign y27519 = n54216 ;
  assign y27520 = n54218 ;
  assign y27521 = n54222 ;
  assign y27522 = n54224 ;
  assign y27523 = ~n54225 ;
  assign y27524 = ~n54226 ;
  assign y27525 = ~n12422 ;
  assign y27526 = n54228 ;
  assign y27527 = n5160 ;
  assign y27528 = n54232 ;
  assign y27529 = ~n54234 ;
  assign y27530 = ~n54236 ;
  assign y27531 = n25797 ;
  assign y27532 = ~1'b0 ;
  assign y27533 = ~1'b0 ;
  assign y27534 = n54238 ;
  assign y27535 = ~1'b0 ;
  assign y27536 = n54240 ;
  assign y27537 = ~n54242 ;
  assign y27538 = ~n54243 ;
  assign y27539 = n54248 ;
  assign y27540 = n54252 ;
  assign y27541 = n16023 ;
  assign y27542 = n54254 ;
  assign y27543 = n54256 ;
  assign y27544 = ~1'b0 ;
  assign y27545 = ~n54257 ;
  assign y27546 = n54261 ;
  assign y27547 = ~n10339 ;
  assign y27548 = 1'b0 ;
  assign y27549 = n54262 ;
  assign y27550 = n54263 ;
  assign y27551 = ~1'b0 ;
  assign y27552 = ~1'b0 ;
  assign y27553 = ~1'b0 ;
  assign y27554 = ~1'b0 ;
  assign y27555 = n50365 ;
  assign y27556 = ~1'b0 ;
  assign y27557 = n15085 ;
  assign y27558 = n54264 ;
  assign y27559 = n7188 ;
  assign y27560 = n54266 ;
  assign y27561 = n39588 ;
  assign y27562 = n54268 ;
  assign y27563 = ~n54269 ;
  assign y27564 = ~n54271 ;
  assign y27565 = ~n54274 ;
  assign y27566 = ~n54275 ;
  assign y27567 = n54280 ;
  assign y27568 = ~n54282 ;
  assign y27569 = n54284 ;
  assign y27570 = n54285 ;
  assign y27571 = n54286 ;
  assign y27572 = ~1'b0 ;
  assign y27573 = ~n54289 ;
  assign y27574 = ~1'b0 ;
  assign y27575 = n54295 ;
  assign y27576 = ~1'b0 ;
  assign y27577 = ~1'b0 ;
  assign y27578 = ~1'b0 ;
  assign y27579 = ~n28974 ;
  assign y27580 = ~n54298 ;
  assign y27581 = ~n54299 ;
  assign y27582 = n54300 ;
  assign y27583 = ~n54304 ;
  assign y27584 = ~1'b0 ;
  assign y27585 = ~1'b0 ;
  assign y27586 = n54305 ;
  assign y27587 = ~n19071 ;
  assign y27588 = n54306 ;
  assign y27589 = n48464 ;
  assign y27590 = n54307 ;
  assign y27591 = ~n54309 ;
  assign y27592 = ~1'b0 ;
  assign y27593 = ~n45845 ;
  assign y27594 = ~1'b0 ;
  assign y27595 = ~1'b0 ;
  assign y27596 = ~n54312 ;
  assign y27597 = n54314 ;
  assign y27598 = n54315 ;
  assign y27599 = n54319 ;
  assign y27600 = n54321 ;
  assign y27601 = ~n54328 ;
  assign y27602 = n51566 ;
  assign y27603 = n54329 ;
  assign y27604 = ~n54330 ;
  assign y27605 = ~1'b0 ;
  assign y27606 = ~1'b0 ;
  assign y27607 = 1'b0 ;
  assign y27608 = ~n54332 ;
  assign y27609 = n54335 ;
  assign y27610 = 1'b0 ;
  assign y27611 = n54336 ;
  assign y27612 = ~n54337 ;
  assign y27613 = ~n54340 ;
  assign y27614 = n54342 ;
  assign y27615 = ~n54343 ;
  assign y27616 = ~n54351 ;
  assign y27617 = ~n54353 ;
  assign y27618 = n54354 ;
  assign y27619 = n54355 ;
  assign y27620 = n54359 ;
  assign y27621 = ~n54360 ;
  assign y27622 = ~n54361 ;
  assign y27623 = n54362 ;
  assign y27624 = ~n54363 ;
  assign y27625 = 1'b0 ;
  assign y27626 = 1'b0 ;
  assign y27627 = ~1'b0 ;
  assign y27628 = 1'b0 ;
  assign y27629 = ~n54366 ;
  assign y27630 = ~1'b0 ;
  assign y27631 = ~1'b0 ;
  assign y27632 = ~n54367 ;
  assign y27633 = ~n54371 ;
  assign y27634 = ~n54372 ;
  assign y27635 = n15900 ;
  assign y27636 = ~1'b0 ;
  assign y27637 = n54374 ;
  assign y27638 = ~n54376 ;
  assign y27639 = n54379 ;
  assign y27640 = n54382 ;
  assign y27641 = n54384 ;
  assign y27642 = ~1'b0 ;
  assign y27643 = ~n54385 ;
  assign y27644 = ~n13350 ;
  assign y27645 = n54386 ;
  assign y27646 = n46363 ;
  assign y27647 = ~1'b0 ;
  assign y27648 = ~n54387 ;
  assign y27649 = ~n54389 ;
  assign y27650 = n54391 ;
  assign y27651 = ~n54393 ;
  assign y27652 = n51603 ;
  assign y27653 = ~n54394 ;
  assign y27654 = ~n54395 ;
  assign y27655 = ~n54397 ;
  assign y27656 = ~1'b0 ;
  assign y27657 = n54402 ;
  assign y27658 = ~n54406 ;
  assign y27659 = n54407 ;
  assign y27660 = ~n54410 ;
  assign y27661 = ~1'b0 ;
  assign y27662 = ~1'b0 ;
  assign y27663 = n54411 ;
  assign y27664 = n54412 ;
  assign y27665 = n54413 ;
  assign y27666 = ~n54414 ;
  assign y27667 = 1'b0 ;
  assign y27668 = ~n54415 ;
  assign y27669 = ~n54416 ;
  assign y27670 = ~1'b0 ;
  assign y27671 = ~1'b0 ;
  assign y27672 = n54418 ;
  assign y27673 = ~n54420 ;
  assign y27674 = ~1'b0 ;
  assign y27675 = n54421 ;
  assign y27676 = ~n54427 ;
  assign y27677 = n54428 ;
  assign y27678 = ~1'b0 ;
  assign y27679 = ~1'b0 ;
  assign y27680 = n54430 ;
  assign y27681 = ~1'b0 ;
  assign y27682 = ~1'b0 ;
  assign y27683 = ~1'b0 ;
  assign y27684 = ~1'b0 ;
  assign y27685 = n54432 ;
  assign y27686 = n54433 ;
  assign y27687 = ~n54435 ;
  assign y27688 = ~n5675 ;
  assign y27689 = ~n10308 ;
  assign y27690 = ~1'b0 ;
  assign y27691 = n54436 ;
  assign y27692 = ~n54437 ;
  assign y27693 = ~1'b0 ;
  assign y27694 = ~1'b0 ;
  assign y27695 = ~1'b0 ;
  assign y27696 = ~n54438 ;
  assign y27697 = ~n54441 ;
  assign y27698 = ~n54447 ;
  assign y27699 = ~n49030 ;
  assign y27700 = ~1'b0 ;
  assign y27701 = ~n54449 ;
  assign y27702 = n54451 ;
  assign y27703 = ~n39001 ;
  assign y27704 = 1'b0 ;
  assign y27705 = n54452 ;
  assign y27706 = ~1'b0 ;
  assign y27707 = ~n54458 ;
  assign y27708 = ~n54459 ;
  assign y27709 = n54466 ;
  assign y27710 = ~1'b0 ;
  assign y27711 = n54467 ;
  assign y27712 = ~1'b0 ;
  assign y27713 = ~1'b0 ;
  assign y27714 = n54468 ;
  assign y27715 = ~1'b0 ;
  assign y27716 = ~n54470 ;
  assign y27717 = n54471 ;
  assign y27718 = n54472 ;
  assign y27719 = ~1'b0 ;
  assign y27720 = ~1'b0 ;
  assign y27721 = ~n54475 ;
  assign y27722 = n54476 ;
  assign y27723 = n46924 ;
  assign y27724 = ~n54477 ;
  assign y27725 = 1'b0 ;
  assign y27726 = ~1'b0 ;
  assign y27727 = n54479 ;
  assign y27728 = n54483 ;
  assign y27729 = ~n54484 ;
  assign y27730 = ~n54487 ;
  assign y27731 = 1'b0 ;
  assign y27732 = n8881 ;
  assign y27733 = n54489 ;
  assign y27734 = ~n54491 ;
  assign y27735 = ~1'b0 ;
  assign y27736 = ~1'b0 ;
  assign y27737 = n54492 ;
  assign y27738 = ~n54494 ;
  assign y27739 = ~n54495 ;
  assign y27740 = ~n46442 ;
  assign y27741 = ~n54497 ;
  assign y27742 = ~1'b0 ;
  assign y27743 = ~n54499 ;
  assign y27744 = ~1'b0 ;
  assign y27745 = n27600 ;
  assign y27746 = ~n54500 ;
  assign y27747 = ~n54501 ;
  assign y27748 = ~1'b0 ;
  assign y27749 = ~n40932 ;
  assign y27750 = ~1'b0 ;
  assign y27751 = n54503 ;
  assign y27752 = ~1'b0 ;
  assign y27753 = n54505 ;
  assign y27754 = n54507 ;
  assign y27755 = ~n54508 ;
  assign y27756 = ~1'b0 ;
  assign y27757 = n54509 ;
  assign y27758 = ~1'b0 ;
  assign y27759 = ~n54510 ;
  assign y27760 = n54523 ;
  assign y27761 = n771 ;
  assign y27762 = ~n54524 ;
  assign y27763 = ~n54528 ;
  assign y27764 = n54530 ;
  assign y27765 = n54531 ;
  assign y27766 = ~1'b0 ;
  assign y27767 = n54533 ;
  assign y27768 = ~n54535 ;
  assign y27769 = n2070 ;
  assign y27770 = ~1'b0 ;
  assign y27771 = n54536 ;
  assign y27772 = ~n54540 ;
  assign y27773 = ~n54541 ;
  assign y27774 = ~1'b0 ;
  assign y27775 = ~1'b0 ;
  assign y27776 = ~1'b0 ;
  assign y27777 = n54542 ;
  assign y27778 = n54543 ;
  assign y27779 = ~n54546 ;
  assign y27780 = ~1'b0 ;
  assign y27781 = n31468 ;
  assign y27782 = n54547 ;
  assign y27783 = ~1'b0 ;
  assign y27784 = ~1'b0 ;
  assign y27785 = ~n54550 ;
  assign y27786 = n54551 ;
  assign y27787 = 1'b0 ;
  assign y27788 = n54552 ;
  assign y27789 = n54553 ;
  assign y27790 = ~n54554 ;
  assign y27791 = n3926 ;
  assign y27792 = n54557 ;
  assign y27793 = n54559 ;
  assign y27794 = ~n54561 ;
  assign y27795 = ~n54562 ;
  assign y27796 = ~n54569 ;
  assign y27797 = n54570 ;
  assign y27798 = n54572 ;
  assign y27799 = n54573 ;
  assign y27800 = 1'b0 ;
  assign y27801 = ~n4083 ;
  assign y27802 = ~n54574 ;
  assign y27803 = ~n54575 ;
  assign y27804 = n54576 ;
  assign y27805 = n54579 ;
  assign y27806 = ~n23669 ;
  assign y27807 = n54583 ;
  assign y27808 = ~n20128 ;
  assign y27809 = ~n54584 ;
  assign y27810 = ~1'b0 ;
  assign y27811 = n54588 ;
  assign y27812 = ~n54592 ;
  assign y27813 = n54594 ;
  assign y27814 = ~n54599 ;
  assign y27815 = n54601 ;
  assign y27816 = ~1'b0 ;
  assign y27817 = ~1'b0 ;
  assign y27818 = n54604 ;
  assign y27819 = ~1'b0 ;
  assign y27820 = ~1'b0 ;
  assign y27821 = n54605 ;
  assign y27822 = ~1'b0 ;
  assign y27823 = ~1'b0 ;
  assign y27824 = ~n53686 ;
  assign y27825 = ~n54608 ;
  assign y27826 = n54613 ;
  assign y27827 = n54615 ;
  assign y27828 = ~1'b0 ;
  assign y27829 = ~1'b0 ;
  assign y27830 = ~n54617 ;
  assign y27831 = ~1'b0 ;
  assign y27832 = ~1'b0 ;
  assign y27833 = n54618 ;
  assign y27834 = n54622 ;
  assign y27835 = n34521 ;
  assign y27836 = ~n54623 ;
  assign y27837 = n54626 ;
  assign y27838 = ~n54633 ;
  assign y27839 = n54637 ;
  assign y27840 = ~1'b0 ;
  assign y27841 = n54639 ;
  assign y27842 = ~1'b0 ;
  assign y27843 = n54641 ;
  assign y27844 = ~n54642 ;
  assign y27845 = ~1'b0 ;
  assign y27846 = n54644 ;
  assign y27847 = 1'b0 ;
  assign y27848 = n38587 ;
  assign y27849 = ~1'b0 ;
  assign y27850 = n54645 ;
  assign y27851 = ~1'b0 ;
  assign y27852 = ~n54648 ;
  assign y27853 = n6638 ;
  assign y27854 = n54650 ;
  assign y27855 = ~n54652 ;
  assign y27856 = n54655 ;
  assign y27857 = n54656 ;
  assign y27858 = ~1'b0 ;
  assign y27859 = ~n54657 ;
  assign y27860 = n54662 ;
  assign y27861 = ~1'b0 ;
  assign y27862 = ~n5643 ;
  assign y27863 = n54663 ;
  assign y27864 = n54666 ;
  assign y27865 = ~1'b0 ;
  assign y27866 = ~n54667 ;
  assign y27867 = n29389 ;
  assign y27868 = n16670 ;
  assign y27869 = n54668 ;
  assign y27870 = ~n54671 ;
  assign y27871 = ~1'b0 ;
  assign y27872 = ~n54672 ;
  assign y27873 = ~n54674 ;
  assign y27874 = ~n54676 ;
  assign y27875 = ~n54682 ;
  assign y27876 = n54683 ;
  assign y27877 = ~1'b0 ;
  assign y27878 = ~1'b0 ;
  assign y27879 = n54685 ;
  assign y27880 = ~n1415 ;
  assign y27881 = n54688 ;
  assign y27882 = n54690 ;
  assign y27883 = ~n54691 ;
  assign y27884 = ~n54694 ;
  assign y27885 = ~1'b0 ;
  assign y27886 = ~n53757 ;
  assign y27887 = n54695 ;
  assign y27888 = ~n54696 ;
  assign y27889 = ~n54697 ;
  assign y27890 = n54699 ;
  assign y27891 = ~n54700 ;
  assign y27892 = n54703 ;
  assign y27893 = ~n54705 ;
  assign y27894 = ~1'b0 ;
  assign y27895 = ~n54712 ;
  assign y27896 = 1'b0 ;
  assign y27897 = ~n54493 ;
  assign y27898 = ~n54713 ;
  assign y27899 = ~n54715 ;
  assign y27900 = n54718 ;
  assign y27901 = ~n54719 ;
  assign y27902 = ~1'b0 ;
  assign y27903 = n54723 ;
  assign y27904 = ~1'b0 ;
  assign y27905 = ~1'b0 ;
  assign y27906 = n54724 ;
  assign y27907 = ~1'b0 ;
  assign y27908 = n54735 ;
  assign y27909 = n54738 ;
  assign y27910 = n54741 ;
  assign y27911 = n54747 ;
  assign y27912 = ~n54749 ;
  assign y27913 = ~1'b0 ;
  assign y27914 = ~1'b0 ;
  assign y27915 = ~n54750 ;
  assign y27916 = ~1'b0 ;
  assign y27917 = ~1'b0 ;
  assign y27918 = ~1'b0 ;
  assign y27919 = n54752 ;
  assign y27920 = n54755 ;
  assign y27921 = ~n54757 ;
  assign y27922 = ~n54758 ;
  assign y27923 = ~n54759 ;
  assign y27924 = n54761 ;
  assign y27925 = n54763 ;
  assign y27926 = ~1'b0 ;
  assign y27927 = n54765 ;
  assign y27928 = n54767 ;
  assign y27929 = ~n54768 ;
  assign y27930 = ~1'b0 ;
  assign y27931 = n54769 ;
  assign y27932 = n54773 ;
  assign y27933 = ~n54775 ;
  assign y27934 = n54778 ;
  assign y27935 = ~n54783 ;
  assign y27936 = n14925 ;
  assign y27937 = ~n20230 ;
  assign y27938 = ~1'b0 ;
  assign y27939 = ~n54784 ;
  assign y27940 = ~1'b0 ;
  assign y27941 = ~1'b0 ;
  assign y27942 = ~n54785 ;
  assign y27943 = ~1'b0 ;
  assign y27944 = ~n54786 ;
  assign y27945 = ~1'b0 ;
  assign y27946 = n54790 ;
  assign y27947 = n54791 ;
  assign y27948 = ~1'b0 ;
  assign y27949 = ~1'b0 ;
  assign y27950 = n54797 ;
  assign y27951 = ~n54800 ;
  assign y27952 = n54807 ;
  assign y27953 = n54808 ;
  assign y27954 = ~n54810 ;
  assign y27955 = ~n54814 ;
  assign y27956 = ~n54818 ;
  assign y27957 = ~n54820 ;
  assign y27958 = ~n54827 ;
  assign y27959 = ~n54828 ;
  assign y27960 = n54832 ;
  assign y27961 = ~n54835 ;
  assign y27962 = ~1'b0 ;
  assign y27963 = ~n5106 ;
  assign y27964 = n54837 ;
  assign y27965 = ~n54839 ;
  assign y27966 = ~n54841 ;
  assign y27967 = ~1'b0 ;
  assign y27968 = ~1'b0 ;
  assign y27969 = ~1'b0 ;
  assign y27970 = ~n54842 ;
  assign y27971 = n54844 ;
  assign y27972 = ~n54847 ;
  assign y27973 = n54848 ;
  assign y27974 = ~n54852 ;
  assign y27975 = ~n54856 ;
  assign y27976 = ~n4264 ;
  assign y27977 = n54858 ;
  assign y27978 = n54859 ;
  assign y27979 = n54862 ;
  assign y27980 = ~n54867 ;
  assign y27981 = ~1'b0 ;
  assign y27982 = ~1'b0 ;
  assign y27983 = ~1'b0 ;
  assign y27984 = ~n54870 ;
  assign y27985 = ~1'b0 ;
  assign y27986 = n54872 ;
  assign y27987 = n54874 ;
  assign y27988 = ~n54877 ;
  assign y27989 = ~n54883 ;
  assign y27990 = n54884 ;
  assign y27991 = x3 ;
  assign y27992 = n54890 ;
  assign y27993 = ~1'b0 ;
  assign y27994 = ~n54894 ;
  assign y27995 = ~n54895 ;
  assign y27996 = ~n54897 ;
  assign y27997 = ~n54898 ;
  assign y27998 = n54901 ;
  assign y27999 = n54902 ;
  assign y28000 = ~1'b0 ;
  assign y28001 = n54903 ;
  assign y28002 = n54904 ;
  assign y28003 = n20745 ;
  assign y28004 = ~1'b0 ;
  assign y28005 = n54906 ;
  assign y28006 = ~n54908 ;
  assign y28007 = n54910 ;
  assign y28008 = n54911 ;
  assign y28009 = ~n54914 ;
  assign y28010 = n54916 ;
  assign y28011 = ~n54920 ;
  assign y28012 = ~1'b0 ;
  assign y28013 = n54923 ;
  assign y28014 = ~n54928 ;
  assign y28015 = n54929 ;
  assign y28016 = n54933 ;
  assign y28017 = ~1'b0 ;
  assign y28018 = n54936 ;
  assign y28019 = ~n54937 ;
  assign y28020 = n38856 ;
  assign y28021 = n54938 ;
  assign y28022 = n54941 ;
  assign y28023 = ~1'b0 ;
  assign y28024 = n54945 ;
  assign y28025 = n54948 ;
  assign y28026 = ~1'b0 ;
  assign y28027 = ~1'b0 ;
  assign y28028 = n54950 ;
  assign y28029 = n54952 ;
  assign y28030 = n54953 ;
  assign y28031 = n54957 ;
  assign y28032 = ~n54958 ;
  assign y28033 = ~1'b0 ;
  assign y28034 = ~n54960 ;
  assign y28035 = ~n54963 ;
  assign y28036 = 1'b0 ;
  assign y28037 = n54965 ;
  assign y28038 = ~n54966 ;
  assign y28039 = ~n54968 ;
  assign y28040 = ~n54969 ;
  assign y28041 = ~n54970 ;
  assign y28042 = ~n54972 ;
  assign y28043 = ~1'b0 ;
  assign y28044 = n54973 ;
  assign y28045 = n54975 ;
  assign y28046 = ~n54979 ;
  assign y28047 = n54981 ;
  assign y28048 = ~1'b0 ;
  assign y28049 = ~n54983 ;
  assign y28050 = ~n54985 ;
  assign y28051 = n54986 ;
  assign y28052 = ~n54988 ;
  assign y28053 = ~n54990 ;
  assign y28054 = n54996 ;
  assign y28055 = ~1'b0 ;
  assign y28056 = n54998 ;
  assign y28057 = n55002 ;
  assign y28058 = ~n55004 ;
  assign y28059 = ~1'b0 ;
  assign y28060 = ~n55006 ;
  assign y28061 = ~n55009 ;
  assign y28062 = n55014 ;
  assign y28063 = ~1'b0 ;
  assign y28064 = ~1'b0 ;
  assign y28065 = ~1'b0 ;
  assign y28066 = n55016 ;
  assign y28067 = ~n55018 ;
  assign y28068 = n55021 ;
  assign y28069 = ~n55022 ;
  assign y28070 = n55024 ;
  assign y28071 = n55028 ;
  assign y28072 = ~1'b0 ;
  assign y28073 = 1'b0 ;
  assign y28074 = n55030 ;
  assign y28075 = ~n55033 ;
  assign y28076 = ~n55039 ;
  assign y28077 = ~n55040 ;
  assign y28078 = n55044 ;
  assign y28079 = ~1'b0 ;
  assign y28080 = ~n27156 ;
  assign y28081 = ~n55047 ;
  assign y28082 = ~1'b0 ;
  assign y28083 = n55049 ;
  assign y28084 = n55050 ;
  assign y28085 = ~n55054 ;
  assign y28086 = ~n55056 ;
  assign y28087 = ~1'b0 ;
  assign y28088 = ~n55058 ;
  assign y28089 = n55060 ;
  assign y28090 = n55061 ;
  assign y28091 = ~1'b0 ;
  assign y28092 = ~n55066 ;
  assign y28093 = ~n55067 ;
  assign y28094 = n55068 ;
  assign y28095 = ~n55073 ;
  assign y28096 = n55075 ;
  assign y28097 = n55077 ;
  assign y28098 = ~1'b0 ;
  assign y28099 = n55037 ;
  assign y28100 = ~n55078 ;
  assign y28101 = n55081 ;
  assign y28102 = ~1'b0 ;
  assign y28103 = n55082 ;
  assign y28104 = ~1'b0 ;
  assign y28105 = ~n55083 ;
  assign y28106 = n55084 ;
  assign y28107 = ~1'b0 ;
  assign y28108 = ~n55086 ;
  assign y28109 = ~1'b0 ;
  assign y28110 = n55088 ;
  assign y28111 = ~1'b0 ;
  assign y28112 = ~1'b0 ;
  assign y28113 = n55090 ;
  assign y28114 = ~n55094 ;
  assign y28115 = ~n43959 ;
  assign y28116 = ~n55096 ;
  assign y28117 = n55097 ;
  assign y28118 = ~1'b0 ;
  assign y28119 = ~1'b0 ;
  assign y28120 = ~1'b0 ;
  assign y28121 = ~n55098 ;
  assign y28122 = n55100 ;
  assign y28123 = ~n55101 ;
  assign y28124 = n55102 ;
  assign y28125 = n55103 ;
  assign y28126 = n55104 ;
  assign y28127 = ~1'b0 ;
  assign y28128 = n55107 ;
  assign y28129 = ~n55112 ;
  assign y28130 = ~n55114 ;
  assign y28131 = n55116 ;
  assign y28132 = ~n12146 ;
  assign y28133 = n48232 ;
  assign y28134 = ~n55125 ;
  assign y28135 = ~n30831 ;
  assign y28136 = n55127 ;
  assign y28137 = n55129 ;
  assign y28138 = ~n55130 ;
  assign y28139 = ~1'b0 ;
  assign y28140 = 1'b0 ;
  assign y28141 = ~n55132 ;
  assign y28142 = ~n55136 ;
  assign y28143 = ~n55137 ;
  assign y28144 = n55140 ;
  assign y28145 = ~n55141 ;
  assign y28146 = ~n55145 ;
  assign y28147 = ~n6374 ;
  assign y28148 = ~n55147 ;
  assign y28149 = n55148 ;
  assign y28150 = ~1'b0 ;
  assign y28151 = ~n37292 ;
  assign y28152 = n55150 ;
  assign y28153 = ~n55152 ;
  assign y28154 = n55154 ;
  assign y28155 = ~n55155 ;
  assign y28156 = n55157 ;
  assign y28157 = ~1'b0 ;
  assign y28158 = 1'b0 ;
  assign y28159 = n55158 ;
  assign y28160 = ~n55160 ;
  assign y28161 = ~n55161 ;
  assign y28162 = n55162 ;
  assign y28163 = ~1'b0 ;
  assign y28164 = n55164 ;
  assign y28165 = ~1'b0 ;
  assign y28166 = n55166 ;
  assign y28167 = ~1'b0 ;
  assign y28168 = ~n55167 ;
  assign y28169 = ~n55168 ;
  assign y28170 = ~n55169 ;
  assign y28171 = n55171 ;
  assign y28172 = ~1'b0 ;
  assign y28173 = n55173 ;
  assign y28174 = ~n55176 ;
  assign y28175 = ~1'b0 ;
  assign y28176 = ~n55178 ;
  assign y28177 = ~1'b0 ;
  assign y28178 = n55181 ;
  assign y28179 = n55185 ;
  assign y28180 = n13062 ;
  assign y28181 = ~n55186 ;
  assign y28182 = ~n55190 ;
  assign y28183 = ~n55192 ;
  assign y28184 = ~n25884 ;
  assign y28185 = ~1'b0 ;
  assign y28186 = ~1'b0 ;
  assign y28187 = n55193 ;
  assign y28188 = n7944 ;
  assign y28189 = ~1'b0 ;
  assign y28190 = n55194 ;
  assign y28191 = n55197 ;
  assign y28192 = n55198 ;
  assign y28193 = n55199 ;
  assign y28194 = 1'b0 ;
  assign y28195 = ~n55200 ;
  assign y28196 = ~n99 ;
  assign y28197 = ~n55202 ;
  assign y28198 = ~1'b0 ;
  assign y28199 = n55204 ;
  assign y28200 = ~n55209 ;
  assign y28201 = n55212 ;
  assign y28202 = ~n1412 ;
  assign y28203 = n55222 ;
  assign y28204 = ~n55223 ;
  assign y28205 = ~n55227 ;
  assign y28206 = ~n55229 ;
  assign y28207 = ~n55231 ;
  assign y28208 = ~n55234 ;
  assign y28209 = n55236 ;
  assign y28210 = ~1'b0 ;
  assign y28211 = ~1'b0 ;
  assign y28212 = ~1'b0 ;
  assign y28213 = n54156 ;
  assign y28214 = ~n55237 ;
  assign y28215 = ~n55238 ;
  assign y28216 = ~n55241 ;
  assign y28217 = n17737 ;
  assign y28218 = n55242 ;
  assign y28219 = n55243 ;
  assign y28220 = ~1'b0 ;
  assign y28221 = ~1'b0 ;
  assign y28222 = n55245 ;
  assign y28223 = n55246 ;
  assign y28224 = n55247 ;
  assign y28225 = ~n55251 ;
  assign y28226 = ~n55254 ;
  assign y28227 = ~1'b0 ;
  assign y28228 = ~1'b0 ;
  assign y28229 = n11696 ;
  assign y28230 = ~1'b0 ;
  assign y28231 = n55256 ;
  assign y28232 = ~1'b0 ;
  assign y28233 = ~n55257 ;
  assign y28234 = ~1'b0 ;
  assign y28235 = ~n55258 ;
  assign y28236 = ~n55259 ;
  assign y28237 = ~n55271 ;
  assign y28238 = n55273 ;
  assign y28239 = ~1'b0 ;
  assign y28240 = ~n55280 ;
  assign y28241 = ~1'b0 ;
  assign y28242 = ~1'b0 ;
  assign y28243 = n55283 ;
  assign y28244 = ~1'b0 ;
  assign y28245 = n55286 ;
  assign y28246 = n55287 ;
  assign y28247 = n55288 ;
  assign y28248 = n55290 ;
  assign y28249 = n55293 ;
  assign y28250 = ~1'b0 ;
  assign y28251 = 1'b0 ;
  assign y28252 = ~1'b0 ;
  assign y28253 = ~n55294 ;
  assign y28254 = 1'b0 ;
  assign y28255 = ~1'b0 ;
  assign y28256 = ~n55295 ;
  assign y28257 = ~n27956 ;
  assign y28258 = n55298 ;
  assign y28259 = n55300 ;
  assign y28260 = ~1'b0 ;
  assign y28261 = ~n55304 ;
  assign y28262 = n55306 ;
  assign y28263 = ~1'b0 ;
  assign y28264 = ~n18743 ;
  assign y28265 = n21843 ;
  assign y28266 = ~n55309 ;
  assign y28267 = ~1'b0 ;
  assign y28268 = n55310 ;
  assign y28269 = ~1'b0 ;
  assign y28270 = n55313 ;
  assign y28271 = n55315 ;
  assign y28272 = ~n55318 ;
  assign y28273 = ~1'b0 ;
  assign y28274 = n55319 ;
  assign y28275 = n55320 ;
  assign y28276 = ~1'b0 ;
  assign y28277 = ~n55324 ;
  assign y28278 = ~1'b0 ;
  assign y28279 = n55325 ;
  assign y28280 = ~n55327 ;
  assign y28281 = ~n55329 ;
  assign y28282 = ~1'b0 ;
  assign y28283 = n55334 ;
  assign y28284 = n55335 ;
  assign y28285 = ~n55342 ;
  assign y28286 = n55344 ;
  assign y28287 = n55347 ;
  assign y28288 = ~n32358 ;
  assign y28289 = ~1'b0 ;
  assign y28290 = n55349 ;
  assign y28291 = ~n55350 ;
  assign y28292 = ~n55351 ;
  assign y28293 = ~n55352 ;
  assign y28294 = n55354 ;
  assign y28295 = ~1'b0 ;
  assign y28296 = ~n55358 ;
  assign y28297 = ~n55362 ;
  assign y28298 = ~n55363 ;
  assign y28299 = ~1'b0 ;
  assign y28300 = ~1'b0 ;
  assign y28301 = ~n55367 ;
  assign y28302 = ~n55369 ;
  assign y28303 = n55371 ;
  assign y28304 = ~n43259 ;
  assign y28305 = n1109 ;
  assign y28306 = ~n55373 ;
  assign y28307 = n55376 ;
  assign y28308 = n55377 ;
  assign y28309 = ~n55379 ;
  assign y28310 = ~1'b0 ;
  assign y28311 = ~1'b0 ;
  assign y28312 = n55380 ;
  assign y28313 = ~n55381 ;
  assign y28314 = n55384 ;
  assign y28315 = n55385 ;
  assign y28316 = ~n55387 ;
  assign y28317 = ~n55392 ;
  assign y28318 = ~n55394 ;
  assign y28319 = ~1'b0 ;
  assign y28320 = n55397 ;
  assign y28321 = n55399 ;
  assign y28322 = n55402 ;
  assign y28323 = ~n55403 ;
  assign y28324 = ~n55404 ;
  assign y28325 = ~n55405 ;
  assign y28326 = ~1'b0 ;
  assign y28327 = ~n55413 ;
  assign y28328 = ~1'b0 ;
  assign y28329 = n55417 ;
  assign y28330 = ~n55420 ;
  assign y28331 = ~1'b0 ;
  assign y28332 = ~n55422 ;
  assign y28333 = ~n55424 ;
  assign y28334 = ~1'b0 ;
  assign y28335 = ~n55425 ;
  assign y28336 = ~n55426 ;
  assign y28337 = ~n55428 ;
  assign y28338 = ~n55430 ;
  assign y28339 = ~n55433 ;
  assign y28340 = ~1'b0 ;
  assign y28341 = ~n55435 ;
  assign y28342 = ~n55437 ;
  assign y28343 = n55438 ;
  assign y28344 = ~n17401 ;
  assign y28345 = ~n55439 ;
  assign y28346 = ~n55443 ;
  assign y28347 = ~n55444 ;
  assign y28348 = ~n55449 ;
  assign y28349 = ~n55451 ;
  assign y28350 = ~1'b0 ;
  assign y28351 = ~1'b0 ;
  assign y28352 = n55454 ;
  assign y28353 = ~n55459 ;
  assign y28354 = ~1'b0 ;
  assign y28355 = n55460 ;
  assign y28356 = n55461 ;
  assign y28357 = ~n55462 ;
  assign y28358 = n55463 ;
  assign y28359 = ~1'b0 ;
  assign y28360 = ~n55465 ;
  assign y28361 = 1'b0 ;
  assign y28362 = ~n55468 ;
  assign y28363 = ~n1602 ;
  assign y28364 = n55469 ;
  assign y28365 = n55471 ;
  assign y28366 = ~1'b0 ;
  assign y28367 = n55475 ;
  assign y28368 = 1'b0 ;
  assign y28369 = n55484 ;
  assign y28370 = n55485 ;
  assign y28371 = ~1'b0 ;
  assign y28372 = n21495 ;
  assign y28373 = ~n55487 ;
  assign y28374 = ~1'b0 ;
  assign y28375 = n55490 ;
  assign y28376 = n55492 ;
  assign y28377 = n55493 ;
  assign y28378 = 1'b0 ;
  assign y28379 = ~1'b0 ;
  assign y28380 = ~n55494 ;
  assign y28381 = ~1'b0 ;
  assign y28382 = ~1'b0 ;
  assign y28383 = ~1'b0 ;
  assign y28384 = n55497 ;
  assign y28385 = ~n55500 ;
  assign y28386 = ~1'b0 ;
  assign y28387 = ~1'b0 ;
  assign y28388 = n55501 ;
  assign y28389 = n18662 ;
  assign y28390 = n55507 ;
  assign y28391 = n55511 ;
  assign y28392 = ~n16798 ;
  assign y28393 = ~n39867 ;
  assign y28394 = n55515 ;
  assign y28395 = ~1'b0 ;
  assign y28396 = ~1'b0 ;
  assign y28397 = ~n55519 ;
  assign y28398 = ~n16947 ;
  assign y28399 = ~n55520 ;
  assign y28400 = ~n55527 ;
  assign y28401 = n55528 ;
  assign y28402 = 1'b0 ;
  assign y28403 = ~1'b0 ;
  assign y28404 = ~n55530 ;
  assign y28405 = ~1'b0 ;
  assign y28406 = ~1'b0 ;
  assign y28407 = ~n55531 ;
  assign y28408 = n55534 ;
  assign y28409 = ~n55538 ;
  assign y28410 = ~1'b0 ;
  assign y28411 = n55539 ;
  assign y28412 = ~1'b0 ;
  assign y28413 = ~n55541 ;
  assign y28414 = ~1'b0 ;
  assign y28415 = n55543 ;
  assign y28416 = ~1'b0 ;
  assign y28417 = ~1'b0 ;
  assign y28418 = ~n55544 ;
  assign y28419 = ~n13011 ;
  assign y28420 = n55545 ;
  assign y28421 = n55546 ;
  assign y28422 = ~n55550 ;
  assign y28423 = ~n55553 ;
  assign y28424 = ~n55554 ;
  assign y28425 = ~n55556 ;
  assign y28426 = n55563 ;
  assign y28427 = ~n55567 ;
  assign y28428 = ~1'b0 ;
  assign y28429 = ~n55573 ;
  assign y28430 = ~1'b0 ;
  assign y28431 = ~1'b0 ;
  assign y28432 = n35086 ;
  assign y28433 = n55575 ;
  assign y28434 = n55576 ;
  assign y28435 = n55578 ;
  assign y28436 = ~n55579 ;
  assign y28437 = ~1'b0 ;
  assign y28438 = ~1'b0 ;
  assign y28439 = ~1'b0 ;
  assign y28440 = ~n55580 ;
  assign y28441 = n55581 ;
  assign y28442 = ~n55582 ;
  assign y28443 = ~1'b0 ;
  assign y28444 = n55586 ;
  assign y28445 = n55587 ;
  assign y28446 = ~n55588 ;
  assign y28447 = ~1'b0 ;
  assign y28448 = ~1'b0 ;
  assign y28449 = ~1'b0 ;
  assign y28450 = ~n55589 ;
  assign y28451 = n55591 ;
  assign y28452 = n55594 ;
  assign y28453 = n55598 ;
  assign y28454 = ~1'b0 ;
  assign y28455 = ~n55600 ;
  assign y28456 = ~n55602 ;
  assign y28457 = n55603 ;
  assign y28458 = n55605 ;
  assign y28459 = n55608 ;
  assign y28460 = n55609 ;
  assign y28461 = n55611 ;
  assign y28462 = ~1'b0 ;
  assign y28463 = n55618 ;
  assign y28464 = ~n55619 ;
  assign y28465 = ~n55620 ;
  assign y28466 = ~n55624 ;
  assign y28467 = ~n55625 ;
  assign y28468 = n55628 ;
  assign y28469 = ~1'b0 ;
  assign y28470 = ~1'b0 ;
  assign y28471 = ~n28929 ;
  assign y28472 = ~n55629 ;
  assign y28473 = n55631 ;
  assign y28474 = ~1'b0 ;
  assign y28475 = ~n55633 ;
  assign y28476 = n55634 ;
  assign y28477 = n55636 ;
  assign y28478 = ~n55637 ;
  assign y28479 = ~n55643 ;
  assign y28480 = n55645 ;
  assign y28481 = n55646 ;
  assign y28482 = ~1'b0 ;
  assign y28483 = ~1'b0 ;
  assign y28484 = n55647 ;
  assign y28485 = ~n55649 ;
  assign y28486 = ~1'b0 ;
  assign y28487 = ~1'b0 ;
  assign y28488 = n55650 ;
  assign y28489 = n55654 ;
  assign y28490 = n53997 ;
  assign y28491 = ~n3575 ;
  assign y28492 = n55656 ;
  assign y28493 = n55659 ;
  assign y28494 = ~1'b0 ;
  assign y28495 = ~n55663 ;
  assign y28496 = n55665 ;
  assign y28497 = ~1'b0 ;
  assign y28498 = ~n55667 ;
  assign y28499 = ~n55668 ;
  assign y28500 = ~n55669 ;
  assign y28501 = ~n55674 ;
  assign y28502 = ~n55676 ;
  assign y28503 = ~n55677 ;
  assign y28504 = ~n55680 ;
  assign y28505 = ~1'b0 ;
  assign y28506 = n55683 ;
  assign y28507 = ~1'b0 ;
  assign y28508 = ~n55684 ;
  assign y28509 = ~n55686 ;
  assign y28510 = ~n55687 ;
  assign y28511 = ~n55688 ;
  assign y28512 = ~n55690 ;
  assign y28513 = n25668 ;
  assign y28514 = ~1'b0 ;
  assign y28515 = ~1'b0 ;
  assign y28516 = ~1'b0 ;
  assign y28517 = ~n55692 ;
  assign y28518 = ~n55693 ;
  assign y28519 = 1'b0 ;
  assign y28520 = ~n55694 ;
  assign y28521 = ~n16738 ;
  assign y28522 = n55696 ;
  assign y28523 = ~n55698 ;
  assign y28524 = ~1'b0 ;
  assign y28525 = ~1'b0 ;
  assign y28526 = ~n55700 ;
  assign y28527 = ~1'b0 ;
  assign y28528 = n55702 ;
  assign y28529 = n55704 ;
  assign y28530 = n55705 ;
  assign y28531 = n55706 ;
  assign y28532 = ~1'b0 ;
  assign y28533 = n55713 ;
  assign y28534 = ~n55718 ;
  assign y28535 = ~1'b0 ;
  assign y28536 = n55720 ;
  assign y28537 = ~n55723 ;
  assign y28538 = ~n55725 ;
  assign y28539 = ~n55726 ;
  assign y28540 = ~1'b0 ;
  assign y28541 = ~n55727 ;
  assign y28542 = ~n55730 ;
  assign y28543 = ~n55731 ;
  assign y28544 = ~n55732 ;
  assign y28545 = n24264 ;
  assign y28546 = n55733 ;
  assign y28547 = n55735 ;
  assign y28548 = ~1'b0 ;
  assign y28549 = ~n55737 ;
  assign y28550 = ~n55738 ;
  assign y28551 = ~1'b0 ;
  assign y28552 = ~n55741 ;
  assign y28553 = n55745 ;
  assign y28554 = ~n55746 ;
  assign y28555 = n55747 ;
  assign y28556 = ~n55748 ;
  assign y28557 = ~1'b0 ;
  assign y28558 = n55750 ;
  assign y28559 = ~n55752 ;
  assign y28560 = ~n55753 ;
  assign y28561 = ~1'b0 ;
  assign y28562 = n55754 ;
  assign y28563 = n55755 ;
  assign y28564 = n55756 ;
  assign y28565 = ~n55757 ;
  assign y28566 = n55759 ;
  assign y28567 = ~n55761 ;
  assign y28568 = n55762 ;
  assign y28569 = ~1'b0 ;
  assign y28570 = ~n55765 ;
  assign y28571 = ~1'b0 ;
  assign y28572 = n55768 ;
  assign y28573 = ~n55779 ;
  assign y28574 = ~n48133 ;
  assign y28575 = ~n55780 ;
  assign y28576 = n55783 ;
  assign y28577 = ~1'b0 ;
  assign y28578 = ~1'b0 ;
  assign y28579 = n55787 ;
  assign y28580 = ~1'b0 ;
  assign y28581 = n55791 ;
  assign y28582 = n55795 ;
  assign y28583 = ~1'b0 ;
  assign y28584 = n30927 ;
  assign y28585 = ~n55796 ;
  assign y28586 = ~n55798 ;
  assign y28587 = n55800 ;
  assign y28588 = ~n55805 ;
  assign y28589 = ~n9586 ;
  assign y28590 = n55806 ;
  assign y28591 = ~n55809 ;
  assign y28592 = n55812 ;
  assign y28593 = ~1'b0 ;
  assign y28594 = ~n55816 ;
  assign y28595 = n55817 ;
  assign y28596 = ~n55819 ;
  assign y28597 = ~n55820 ;
  assign y28598 = ~1'b0 ;
  assign y28599 = n55822 ;
  assign y28600 = ~1'b0 ;
  assign y28601 = ~1'b0 ;
  assign y28602 = ~1'b0 ;
  assign y28603 = 1'b0 ;
  assign y28604 = ~1'b0 ;
  assign y28605 = n55823 ;
  assign y28606 = n55827 ;
  assign y28607 = n55829 ;
  assign y28608 = n55837 ;
  assign y28609 = ~n55838 ;
  assign y28610 = ~n55847 ;
  assign y28611 = ~n55848 ;
  assign y28612 = ~1'b0 ;
  assign y28613 = ~1'b0 ;
  assign y28614 = ~1'b0 ;
  assign y28615 = n55850 ;
  assign y28616 = ~1'b0 ;
  assign y28617 = ~1'b0 ;
  assign y28618 = n55851 ;
  assign y28619 = ~n55852 ;
  assign y28620 = ~n55853 ;
  assign y28621 = ~n55854 ;
  assign y28622 = ~n55855 ;
  assign y28623 = ~n55856 ;
  assign y28624 = n55860 ;
  assign y28625 = ~n51503 ;
  assign y28626 = n55861 ;
  assign y28627 = ~1'b0 ;
  assign y28628 = ~n55864 ;
  assign y28629 = ~n55865 ;
  assign y28630 = ~n55866 ;
  assign y28631 = n55868 ;
  assign y28632 = ~n55871 ;
  assign y28633 = ~n55874 ;
  assign y28634 = ~1'b0 ;
  assign y28635 = n55877 ;
  assign y28636 = ~1'b0 ;
  assign y28637 = ~n55879 ;
  assign y28638 = n55881 ;
  assign y28639 = ~n55883 ;
  assign y28640 = ~n55884 ;
  assign y28641 = ~n55886 ;
  assign y28642 = ~n55889 ;
  assign y28643 = ~1'b0 ;
  assign y28644 = ~1'b0 ;
  assign y28645 = n55893 ;
  assign y28646 = ~1'b0 ;
  assign y28647 = ~n55894 ;
  assign y28648 = 1'b0 ;
  assign y28649 = ~n55899 ;
  assign y28650 = ~n55901 ;
  assign y28651 = n55902 ;
  assign y28652 = n55903 ;
  assign y28653 = n53906 ;
  assign y28654 = ~n55906 ;
  assign y28655 = ~n55908 ;
  assign y28656 = ~n55911 ;
  assign y28657 = ~n55914 ;
  assign y28658 = ~1'b0 ;
  assign y28659 = ~n55916 ;
  assign y28660 = ~n55926 ;
  assign y28661 = ~1'b0 ;
  assign y28662 = n55927 ;
  assign y28663 = n55930 ;
  assign y28664 = ~n55931 ;
  assign y28665 = ~1'b0 ;
  assign y28666 = n55933 ;
  assign y28667 = ~n55934 ;
  assign y28668 = n55935 ;
  assign y28669 = ~1'b0 ;
  assign y28670 = ~1'b0 ;
  assign y28671 = n55937 ;
  assign y28672 = ~1'b0 ;
  assign y28673 = n55939 ;
  assign y28674 = ~n55940 ;
  assign y28675 = 1'b0 ;
  assign y28676 = ~1'b0 ;
  assign y28677 = ~n55941 ;
  assign y28678 = n55942 ;
  assign y28679 = n55945 ;
  assign y28680 = n55948 ;
  assign y28681 = n55952 ;
  assign y28682 = n55953 ;
  assign y28683 = ~1'b0 ;
  assign y28684 = ~n55955 ;
  assign y28685 = n55956 ;
  assign y28686 = n55957 ;
  assign y28687 = n55959 ;
  assign y28688 = n55960 ;
  assign y28689 = ~n55962 ;
  assign y28690 = n55963 ;
  assign y28691 = ~n55965 ;
  assign y28692 = ~1'b0 ;
  assign y28693 = ~n55968 ;
  assign y28694 = n55970 ;
  assign y28695 = n55973 ;
  assign y28696 = ~n55974 ;
  assign y28697 = n55976 ;
  assign y28698 = ~n55982 ;
  assign y28699 = ~n55983 ;
  assign y28700 = ~n55986 ;
  assign y28701 = n55988 ;
  assign y28702 = ~n55990 ;
  assign y28703 = n55996 ;
  assign y28704 = n38205 ;
  assign y28705 = n56003 ;
  assign y28706 = ~n56006 ;
  assign y28707 = n56007 ;
  assign y28708 = ~n56012 ;
  assign y28709 = ~1'b0 ;
  assign y28710 = ~n56013 ;
  assign y28711 = ~n48235 ;
  assign y28712 = n56017 ;
  assign y28713 = ~1'b0 ;
  assign y28714 = ~n56021 ;
  assign y28715 = 1'b0 ;
  assign y28716 = ~n56023 ;
  assign y28717 = ~n56024 ;
  assign y28718 = ~n56029 ;
  assign y28719 = ~n56031 ;
  assign y28720 = ~n56032 ;
  assign y28721 = n56033 ;
  assign y28722 = ~n17243 ;
  assign y28723 = n56035 ;
  assign y28724 = ~n56036 ;
  assign y28725 = ~n56037 ;
  assign y28726 = ~1'b0 ;
  assign y28727 = ~n56038 ;
  assign y28728 = ~n1818 ;
  assign y28729 = ~n56039 ;
  assign y28730 = ~n56045 ;
  assign y28731 = ~n56046 ;
  assign y28732 = n56048 ;
  assign y28733 = ~1'b0 ;
  assign y28734 = ~n56050 ;
  assign y28735 = ~n39456 ;
  assign y28736 = ~n35198 ;
  assign y28737 = ~1'b0 ;
  assign y28738 = ~n56051 ;
  assign y28739 = ~n56053 ;
  assign y28740 = ~n56054 ;
  assign y28741 = n40025 ;
  assign y28742 = ~n56056 ;
  assign y28743 = ~n56058 ;
  assign y28744 = ~1'b0 ;
  assign y28745 = ~1'b0 ;
  assign y28746 = ~1'b0 ;
  assign y28747 = ~1'b0 ;
  assign y28748 = n56059 ;
  assign y28749 = ~1'b0 ;
  assign y28750 = ~n56064 ;
  assign y28751 = ~n56069 ;
  assign y28752 = ~n56072 ;
  assign y28753 = ~1'b0 ;
  assign y28754 = ~1'b0 ;
  assign y28755 = ~n56074 ;
  assign y28756 = n56075 ;
  assign y28757 = n56077 ;
  assign y28758 = n56081 ;
  assign y28759 = ~1'b0 ;
  assign y28760 = ~1'b0 ;
  assign y28761 = n56082 ;
  assign y28762 = n56086 ;
  assign y28763 = 1'b0 ;
  assign y28764 = n56087 ;
  assign y28765 = ~1'b0 ;
  assign y28766 = n56088 ;
  assign y28767 = ~n56089 ;
  assign y28768 = ~1'b0 ;
  assign y28769 = n56091 ;
  assign y28770 = ~n56095 ;
  assign y28771 = ~1'b0 ;
  assign y28772 = ~n56099 ;
  assign y28773 = ~n56100 ;
  assign y28774 = ~n56103 ;
  assign y28775 = ~n56104 ;
  assign y28776 = ~1'b0 ;
endmodule
